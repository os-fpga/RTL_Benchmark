library ieee;
use ieee.std_logic_1164.all;

entity top is
 port(opcode: in std_logic_vector(4 downto 0);
      op_ext: in std_logic_vector(1 downto 0);
      sel_reg_dst, sel_alu_opB: out std_logic_vector(1 downto 0);
      alu_op: out std_logic_vector(2 downto 0);
      alu_op_ext: out std_logic_vector(3 downto 0);
      halt, reg_write, sel_pc_opA, sel_pc_opB, beqz, bnez, bgez, bltz, jump, Cin, invA, invB, sign, mem_write, sel_wb: out std_logic);
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173: std_logic;

begin

w0 <= opcode(0) and not opcode(1);
w1 <= opcode(3) and opcode(4);
w2 <= w0 and w1;
w3 <= opcode(1) and opcode(3);
w4 <= opcode(4) and w3;
w5 <= not w2 and not w4;
w6 <= not opcode(2) and not w5;
w7 <= not opcode(1) and opcode(3);
w8 <= opcode(4) and w7;
w9 <= not opcode(3) and not opcode(4);
w10 <= not w1 and not w9;
w11 <= opcode(1) and not w10;
w12 <= not w8 and not w11;
w13 <= opcode(2) and not w12;
w14 <= not w6 and not w13;
w15 <= not opcode(0) and not w1;
w16 <= not opcode(0) and not w15;
w17 <= not opcode(1) and not w16;
w18 <= not opcode(3) and not w9;
w19 <= opcode(1) and not w18;
w20 <= not w17 and not w19;
w21 <= not opcode(2) and not w20;
w22 <= not opcode(3) and opcode(4);
w23 <= not opcode(3) and not w22;
w24 <= opcode(1) and not w23;
w25 <= opcode(1) and not w24;
w26 <= opcode(2) and not w25;
w27 <= not w21 and not w26;
w28 <= not opcode(0) and not w10;
w29 <= opcode(3) and not w1;
w30 <= opcode(0) and not w29;
w31 <= not w28 and not w30;
w32 <= opcode(1) and not w31;
w33 <= not w17 and not w32;
w34 <= not opcode(2) and not w33;
w35 <= not opcode(2) and not w34;
w36 <= not opcode(0) and not opcode(3);
w37 <= not w22 and w36;
w38 <= opcode(0) and not w10;
w39 <= not w37 and not w38;
w40 <= not opcode(1) and not w39;
w41 <= not w19 and not w40;
w42 <= not opcode(2) and not w41;
w43 <= opcode(2) and not w18;
w44 <= not w42 and not w43;
w45 <= not opcode(0) and opcode(3);
w46 <= opcode(4) and op_ext(0);
w47 <= w45 and w46;
w48 <= opcode(3) and not op_ext(1);
w49 <= not w1 and w48;
w50 <= opcode(3) and not op_ext(0);
w51 <= not w1 and w50;
w52 <= opcode(3) and op_ext(0);
w53 <= not w51 and not w52;
w54 <= op_ext(1) and not w53;
w55 <= not w49 and not w54;
w56 <= opcode(0) and not w55;
w57 <= not w47 and not w56;
w58 <= opcode(1) and not w57;
w59 <= not opcode(2) and not w58;
w60 <= opcode(0) and not w18;
w61 <= opcode(0) and not w60;
w62 <= opcode(2) and not w61;
w63 <= not w59 and not w62;
w64 <= opcode(3) and op_ext(1);
w65 <= not w49 and not w64;
w66 <= opcode(1) and not w65;
w67 <= not opcode(2) and not w66;
w68 <= opcode(1) and not w19;
w69 <= opcode(2) and not w68;
w70 <= not w67 and not w69;
w71 <= not opcode(1) and not w1;
w72 <= not w9 and w71;
w73 <= not w9 and w15;
w74 <= opcode(0) and not w23;
w75 <= not w73 and not w74;
w76 <= opcode(1) and not w75;
w77 <= not w72 and not w76;
w78 <= not opcode(2) and not w77;
w79 <= opcode(2) and opcode(3);
w80 <= opcode(4) and w79;
w81 <= not w78 and not w80;
w82 <= not opcode(1) and not opcode(2);
w83 <= not w17 and w82;
w84 <= opcode(1) and not w39;
w85 <= not w2 and not w84;
w86 <= opcode(2) and not w85;
w87 <= not w83 and not w86;
w88 <= not opcode(0) and not w18;
w89 <= not opcode(0) and not w88;
w90 <= opcode(1) and not w89;
w91 <= opcode(1) and not opcode(2);
w92 <= not w90 and w91;
w93 <= opcode(1) and opcode(2);
w94 <= not w10 and w93;
w95 <= not w92 and not w94;
w96 <= not w71 and not w90;
w97 <= not opcode(2) and not w96;
w98 <= not w26 and not w97;
w99 <= not w45 and not w74;
w100 <= opcode(1) and not w99;
w101 <= not opcode(2) and not w72;
w102 <= not w100 and w101;
w103 <= not w43 and not w102;
w104 <= not opcode(0) and not w23;
w105 <= not opcode(0) and not w104;
w106 <= not opcode(1) and not w105;
w107 <= not opcode(1) and not w106;
w108 <= not opcode(2) and not w107;
w109 <= not opcode(2) and not w108;
w110 <= not opcode(1) and not w99;
w111 <= not w24 and not w110;
w112 <= not opcode(2) and not w111;
w113 <= not opcode(1) and opcode(4);
w114 <= opcode(1) and not w29;
w115 <= not w113 and not w114;
w116 <= opcode(2) and not w115;
w117 <= not w112 and not w116;
w118 <= opcode(0) and not w74;
w119 <= opcode(2) and not w118;
w120 <= opcode(2) and not w119;
w121 <= opcode(2) and not w105;
w122 <= opcode(2) and not w121;
w123 <= not opcode(0) and not w29;
w124 <= not opcode(0) and not w123;
w125 <= not opcode(1) and not w124;
w126 <= not opcode(1) and not w125;
w127 <= opcode(2) and not w126;
w128 <= opcode(2) and not w127;
w129 <= opcode(0) and not w30;
w130 <= not opcode(1) and not w129;
w131 <= not opcode(1) and not w130;
w132 <= opcode(2) and not w131;
w133 <= opcode(2) and not w132;
w134 <= opcode(1) and not w129;
w135 <= opcode(1) and not w134;
w136 <= opcode(2) and not w135;
w137 <= opcode(2) and not w136;
w138 <= opcode(1) and not w124;
w139 <= opcode(1) and not w138;
w140 <= opcode(2) and not w139;
w141 <= opcode(2) and not w140;
w142 <= opcode(2) and not w23;
w143 <= opcode(2) and not w142;
w144 <= opcode(0) and opcode(1);
w145 <= not w53 and w144;
w146 <= w0 and not w30;
w147 <= not opcode(2) and not w146;
w148 <= not w145 and w147;
w149 <= opcode(1) and not w16;
w150 <= not w71 and not w149;
w151 <= opcode(2) and not w150;
w152 <= not w148 and not w151;
w153 <= op_ext(0) and w1;
w154 <= not op_ext(1) and not w153;
w155 <= not op_ext(1) and not w154;
w156 <= opcode(0) and not w155;
w157 <= opcode(0) and not w156;
w158 <= opcode(1) and not w157;
w159 <= not w130 and not w158;
w160 <= not opcode(2) and not w159;
w161 <= not opcode(2) and not w160;
w162 <= not w55 and w144;
w163 <= not opcode(2) and not w162;
w164 <= not w151 and not w163;
w165 <= not opcode(1) and not w89;
w166 <= opcode(1) and not w61;
w167 <= not w165 and not w166;
w168 <= not opcode(2) and not w167;
w169 <= not opcode(2) and not w168;
w170 <= not opcode(1) and not w61;
w171 <= not opcode(1) and not w170;
w172 <= not opcode(2) and not w171;
w173 <= not opcode(2) and not w172;
one <= '1';
sel_reg_dst(0) <= not w14;-- level 6
sel_reg_dst(1) <= w27;-- level 7
sel_alu_opB(0) <= w35;-- level 8
sel_alu_opB(1) <= w44;-- level 8
alu_op(0) <= w63;-- level 10
alu_op(1) <= w70;-- level 6
alu_op(2) <= not w81;-- level 8
alu_op_ext(0) <= not w87;-- level 8
alu_op_ext(1) <= not w95;-- level 7
alu_op_ext(2) <= w98;-- level 8
alu_op_ext(3) <= w103;-- level 7
halt <= w109;-- level 8
reg_write <= not w117;-- level 8
sel_pc_opA <= w120;-- level 6
sel_pc_opB <= w122;-- level 6
beqz <= w128;-- level 8
bnez <= w133;-- level 8
bgez <= w137;-- level 8
bltz <= w141;-- level 8
jump <= w143;-- level 4
Cin <= w152;-- level 7
invA <= w161;-- level 10
invB <= w164;-- level 8
sign <= one;-- level 0
mem_write <= w169;-- level 8
sel_wb <= w173;-- level 8
end Behavioral;