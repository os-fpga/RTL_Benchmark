// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: data_input_sequencer.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2016-04-18-EP on Sat Apr 27 13:59:59 2019
//=============================================================================
// Description: Sequencer for data_input
//=============================================================================

`ifndef DATA_INPUT_SEQUENCER_SV
`define DATA_INPUT_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(input_tx) data_input_sequencer_t;


`endif // DATA_INPUT_SEQUENCER_SV

