module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] ,
    \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] ,
    \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] ,
    \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ;
  output \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] ,
    \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] ,
    \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] ,
    \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24] ;
  wire n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
    n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
    n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
    n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
    n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
    n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
    n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
    n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
    n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
    n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
    n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
    n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
    n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
    n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
    n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
    n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
    n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
    n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
    n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
    n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
    n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
    n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
    n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
    n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
    n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
    n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
    n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
    n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
    n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
    n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
    n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
    n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
    n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
    n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
    n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
    n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
    n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
    n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
    n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
    n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
    n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
    n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
    n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
    n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
    n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
    n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
    n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
    n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
    n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
    n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
    n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
    n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
    n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
    n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
    n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
    n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
    n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
    n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
    n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
    n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
    n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
    n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
    n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
    n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
    n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
    n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
    n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
    n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
    n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
    n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
    n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
    n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
    n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
    n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
    n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
    n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
    n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
    n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
    n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
    n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
    n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
    n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
    n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
    n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
    n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
    n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
    n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
    n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
    n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
    n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
    n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
    n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
    n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
    n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
    n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
    n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
    n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
    n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
    n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
    n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
    n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
    n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
    n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
    n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
    n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
    n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
    n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
    n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
    n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
    n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
    n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
    n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
    n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
    n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
    n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
    n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
    n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
    n4277, n4278, n4279, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
    n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
    n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
    n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
    n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
    n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
    n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
    n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
    n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
    n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
    n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
    n4388, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
    n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
    n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
    n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
    n4499, n4500, n4501, n4502, n4503, n4505, n4506, n4507, n4508, n4509,
    n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
    n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
    n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
    n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
    n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
    n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
    n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
    n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
    n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
    n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
    n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
    n4711, n4712, n4713, n4714, n4715, n4717, n4718, n4719, n4720, n4721,
    n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
    n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
    n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
    n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
    n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
    n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
    n4812, n4813, n4814, n4815, n4817, n4818, n4819, n4820, n4821, n4822,
    n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
    n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
    n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
    n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
    n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898, n4900, n4901, n4902, n4903,
    n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
    n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
    n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
    n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
    n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
    n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
    n4984, n4985, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
    n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
    n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
    n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
    n5045, n5046, n5047, n5048, n5049, n5051, n5052, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
    n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
    n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
    n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
    n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
    n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
    n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
    n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
    n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
    n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
    n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
    n5238, n5239, n5240, n5241, n5242, n5244, n5245, n5246, n5247, n5248,
    n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
    n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
    n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5295, n5296, n5297, n5298, n5299,
    n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
    n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
    n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
    n5330, n5331, n5332, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
    n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
    n5351, n5352, n5353, n5354, n5356, n5357, n5358, n5359, n5360, n5361,
    n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
    n5372, n5373, n5374, n5375, n5376, n5377, n5379, n5380, n5381, n5382,
    n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
    n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5401, n5402, n5403,
    n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
    n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5424,
    n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
    n5435, n5436, n5437, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5451, n5452, n5453, n5454, n5455, n5456,
    n5457, n5458, n5459, n5461, n5462, n5463, n5464;
  assign n50 = \a[21]  & \a[22] ;
  assign n51 = ~\a[1]  & ~\a[2] ;
  assign n52 = ~\a[0]  & n51;
  assign n53 = ~\a[3]  & n52;
  assign n54 = ~\a[4]  & n53;
  assign n55 = ~\a[5]  & n54;
  assign n56 = ~\a[6]  & n55;
  assign n57 = ~\a[7]  & n56;
  assign n58 = ~\a[8]  & n57;
  assign n59 = ~\a[9]  & n58;
  assign n60 = ~\a[10]  & n59;
  assign n61 = ~\a[11]  & n60;
  assign n62 = ~\a[12]  & n61;
  assign n63 = ~\a[13]  & n62;
  assign n64 = ~\a[14]  & n63;
  assign n65 = ~\a[15]  & n64;
  assign n66 = ~\a[16]  & n65;
  assign n67 = ~\a[17]  & n66;
  assign n68 = ~\a[18]  & n67;
  assign n69 = ~\a[19]  & n68;
  assign n70 = ~\a[20]  & n69;
  assign n71 = ~\a[21]  & n70;
  assign n72 = \a[21]  & ~n70;
  assign n73 = ~n71 & ~n72;
  assign n74 = ~\a[22]  & n73;
  assign n75 = ~n50 & ~n74;
  assign n76 = \a[20]  & \a[22] ;
  assign n77 = \a[20]  & ~n69;
  assign n78 = ~n70 & ~n77;
  assign n79 = ~\a[22]  & n78;
  assign n80 = ~n76 & ~n79;
  assign n81 = n75 & n80;
  assign n82 = \a[15]  & \a[22] ;
  assign n83 = ~\a[22]  & ~n65;
  assign n84 = \a[15]  & ~n64;
  assign n85 = n83 & ~n84;
  assign n86 = ~n82 & ~n85;
  assign n87 = n81 & n86;
  assign n88 = ~\a[22]  & ~n68;
  assign n89 = \a[19]  & ~n88;
  assign n90 = ~\a[19]  & n88;
  assign n91 = ~n89 & ~n90;
  assign n92 = \a[18]  & \a[22] ;
  assign n93 = \a[18]  & ~n67;
  assign n94 = n88 & ~n93;
  assign n95 = ~n92 & ~n94;
  assign n96 = ~n91 & ~n95;
  assign n97 = ~\a[22]  & ~n66;
  assign n98 = \a[17]  & ~n97;
  assign n99 = ~\a[17]  & n97;
  assign n100 = ~n98 & ~n99;
  assign n101 = \a[16]  & ~n83;
  assign n102 = ~\a[16]  & n83;
  assign n103 = ~n101 & ~n102;
  assign n104 = ~n100 & n103;
  assign n105 = n96 & n104;
  assign n106 = n87 & n105;
  assign n107 = n100 & n103;
  assign n108 = n96 & n107;
  assign n109 = n75 & ~n80;
  assign n110 = n86 & n109;
  assign n111 = n108 & n110;
  assign n112 = ~n91 & n95;
  assign n113 = n107 & n112;
  assign n114 = n110 & n113;
  assign n115 = ~n86 & n109;
  assign n116 = n91 & ~n95;
  assign n117 = n107 & n116;
  assign n118 = n115 & n117;
  assign n119 = ~n75 & n80;
  assign n120 = ~n86 & n119;
  assign n121 = n100 & ~n103;
  assign n122 = n112 & n121;
  assign n123 = n120 & n122;
  assign n124 = ~n75 & ~n80;
  assign n125 = ~n86 & n124;
  assign n126 = n104 & n112;
  assign n127 = n125 & n126;
  assign n128 = n86 & n124;
  assign n129 = n105 & n128;
  assign n130 = n81 & ~n86;
  assign n131 = n104 & n116;
  assign n132 = n130 & n131;
  assign n133 = n105 & n120;
  assign n134 = n122 & n125;
  assign n135 = ~n100 & ~n103;
  assign n136 = n116 & n135;
  assign n137 = n125 & n136;
  assign n138 = n128 & n136;
  assign n139 = n122 & n128;
  assign n140 = n128 & n131;
  assign n141 = ~n139 & ~n140;
  assign n142 = n105 & n110;
  assign n143 = n96 & n121;
  assign n144 = n128 & n143;
  assign n145 = ~n142 & ~n144;
  assign n146 = n105 & n115;
  assign n147 = n116 & n121;
  assign n148 = n110 & n147;
  assign n149 = ~n146 & ~n148;
  assign n150 = n126 & n128;
  assign n151 = n112 & n135;
  assign n152 = n128 & n151;
  assign n153 = ~n150 & ~n152;
  assign n154 = n130 & n136;
  assign n155 = n105 & n125;
  assign n156 = ~n154 & ~n155;
  assign n157 = n153 & n156;
  assign n158 = n149 & n157;
  assign n159 = n145 & n158;
  assign n160 = n141 & n159;
  assign n161 = ~n138 & n160;
  assign n162 = ~n137 & n161;
  assign n163 = ~n134 & n162;
  assign n164 = ~n133 & n163;
  assign n165 = ~n132 & n164;
  assign n166 = n110 & n143;
  assign n167 = n120 & n151;
  assign n168 = n87 & n151;
  assign n169 = n115 & n122;
  assign n170 = n91 & n95;
  assign n171 = n107 & n170;
  assign n172 = n115 & n171;
  assign n173 = n86 & n119;
  assign n174 = n151 & n173;
  assign n175 = n108 & n125;
  assign n176 = n125 & n143;
  assign n177 = n117 & n173;
  assign n178 = n108 & n128;
  assign n179 = ~n177 & ~n178;
  assign n180 = ~n176 & n179;
  assign n181 = ~n175 & n180;
  assign n182 = ~n174 & n181;
  assign n183 = ~n172 & n182;
  assign n184 = ~n169 & n183;
  assign n185 = ~n168 & n184;
  assign n186 = n108 & n120;
  assign n187 = n135 & n170;
  assign n188 = n128 & n187;
  assign n189 = ~n186 & ~n188;
  assign n190 = n110 & n151;
  assign n191 = n117 & n120;
  assign n192 = n120 & n126;
  assign n193 = n121 & n170;
  assign n194 = n125 & n193;
  assign n195 = n96 & n135;
  assign n196 = n128 & n195;
  assign n197 = ~n194 & ~n196;
  assign n198 = ~n192 & n197;
  assign n199 = ~n191 & n198;
  assign n200 = ~n190 & n199;
  assign n201 = n189 & n200;
  assign n202 = n185 & n201;
  assign n203 = ~n167 & n202;
  assign n204 = ~n166 & n203;
  assign n205 = n104 & n170;
  assign n206 = n115 & n205;
  assign n207 = n120 & n131;
  assign n208 = n128 & n147;
  assign n209 = ~n207 & ~n208;
  assign n210 = ~n206 & n209;
  assign n211 = n130 & n147;
  assign n212 = n115 & n195;
  assign n213 = n171 & n173;
  assign n214 = n125 & n171;
  assign n215 = n117 & n130;
  assign n216 = n110 & n126;
  assign n217 = n120 & n147;
  assign n218 = n108 & n173;
  assign n219 = n125 & n187;
  assign n220 = n125 & n131;
  assign n221 = n125 & n147;
  assign n222 = n128 & n193;
  assign n223 = n122 & n130;
  assign n224 = n115 & n126;
  assign n225 = n120 & n143;
  assign n226 = n105 & n173;
  assign n227 = n125 & n151;
  assign n228 = n113 & n125;
  assign n229 = ~n227 & ~n228;
  assign n230 = ~n226 & n229;
  assign n231 = ~n225 & n230;
  assign n232 = ~n224 & n231;
  assign n233 = ~n223 & n232;
  assign n234 = n115 & n187;
  assign n235 = n105 & n130;
  assign n236 = ~n234 & ~n235;
  assign n237 = n130 & n187;
  assign n238 = n130 & n205;
  assign n239 = ~n237 & ~n238;
  assign n240 = n236 & n239;
  assign n241 = n233 & n240;
  assign n242 = ~n222 & n241;
  assign n243 = ~n221 & n242;
  assign n244 = ~n220 & n243;
  assign n245 = ~n219 & n244;
  assign n246 = ~n218 & n245;
  assign n247 = ~n217 & n246;
  assign n248 = ~n216 & n247;
  assign n249 = ~n215 & n248;
  assign n250 = ~n214 & n249;
  assign n251 = ~n213 & n250;
  assign n252 = ~n212 & n251;
  assign n253 = ~n211 & n252;
  assign n254 = n173 & n193;
  assign n255 = n120 & n195;
  assign n256 = ~n254 & ~n255;
  assign n257 = n113 & n173;
  assign n258 = n87 & n193;
  assign n259 = ~n257 & ~n258;
  assign n260 = n256 & n259;
  assign n261 = n253 & n260;
  assign n262 = n210 & n261;
  assign n263 = n204 & n262;
  assign n264 = n165 & n263;
  assign n265 = ~n129 & n264;
  assign n266 = ~n127 & n265;
  assign n267 = ~n123 & n266;
  assign n268 = ~n118 & n267;
  assign n269 = ~n114 & n268;
  assign n270 = ~n111 & n269;
  assign n271 = ~n106 & n270;
  assign n272 = ~\a[22]  & ~n54;
  assign n273 = \a[5]  & ~n272;
  assign n274 = ~\a[5]  & n272;
  assign n275 = ~n273 & ~n274;
  assign n276 = \a[4]  & \a[22] ;
  assign n277 = \a[4]  & ~n53;
  assign n278 = n272 & ~n277;
  assign n279 = ~n276 & ~n278;
  assign n280 = n275 & ~n279;
  assign n281 = ~n275 & n279;
  assign n282 = ~n280 & ~n281;
  assign n283 = ~\a[22]  & ~n52;
  assign n284 = \a[3]  & ~n283;
  assign n285 = ~\a[3]  & n283;
  assign n286 = ~n284 & ~n285;
  assign n287 = \a[2]  & \a[22] ;
  assign n288 = ~\a[0]  & ~\a[1] ;
  assign n289 = \a[2]  & ~n288;
  assign n290 = n283 & ~n289;
  assign n291 = ~n287 & ~n290;
  assign n292 = n286 & ~n291;
  assign n293 = ~n286 & n291;
  assign n294 = ~n292 & ~n293;
  assign n295 = n282 & ~n294;
  assign n296 = n130 & n151;
  assign n297 = n108 & n115;
  assign n298 = n113 & n115;
  assign n299 = n122 & n173;
  assign n300 = n120 & n205;
  assign n301 = ~n211 & ~n300;
  assign n302 = n115 & n131;
  assign n303 = ~n111 & ~n302;
  assign n304 = n179 & n303;
  assign n305 = n301 & n304;
  assign n306 = ~n137 & n305;
  assign n307 = ~n299 & n306;
  assign n308 = ~n191 & n307;
  assign n309 = ~n298 & n308;
  assign n310 = ~n297 & n309;
  assign n311 = ~n296 & n310;
  assign n312 = n173 & n195;
  assign n313 = n120 & n136;
  assign n314 = ~n221 & ~n313;
  assign n315 = n110 & n187;
  assign n316 = ~n114 & ~n315;
  assign n317 = n125 & n205;
  assign n318 = ~n129 & ~n317;
  assign n319 = ~n207 & n318;
  assign n320 = n316 & n319;
  assign n321 = n314 & n320;
  assign n322 = ~n312 & n321;
  assign n323 = ~n212 & n322;
  assign n324 = n87 & n171;
  assign n325 = ~n123 & ~n324;
  assign n326 = n87 & n147;
  assign n327 = n136 & n173;
  assign n328 = n128 & n205;
  assign n329 = n147 & n173;
  assign n330 = ~n328 & ~n329;
  assign n331 = ~n255 & n330;
  assign n332 = ~n327 & n331;
  assign n333 = ~n168 & n332;
  assign n334 = ~n326 & n333;
  assign n335 = n110 & n193;
  assign n336 = n113 & n120;
  assign n337 = n113 & n128;
  assign n338 = ~n188 & ~n337;
  assign n339 = ~n175 & n338;
  assign n340 = ~n336 & n339;
  assign n341 = ~n335 & n340;
  assign n342 = n108 & n130;
  assign n343 = n173 & n187;
  assign n344 = ~n342 & ~n343;
  assign n345 = n130 & n171;
  assign n346 = ~n150 & ~n345;
  assign n347 = n110 & n195;
  assign n348 = n131 & n173;
  assign n349 = ~n347 & ~n348;
  assign n350 = n126 & n173;
  assign n351 = n87 & n113;
  assign n352 = ~n192 & ~n226;
  assign n353 = ~n351 & n352;
  assign n354 = ~n217 & n353;
  assign n355 = ~n216 & n354;
  assign n356 = n110 & n171;
  assign n357 = n110 & n136;
  assign n358 = n110 & n205;
  assign n359 = n110 & n117;
  assign n360 = n120 & n187;
  assign n361 = n115 & n147;
  assign n362 = ~n360 & ~n361;
  assign n363 = ~n359 & n362;
  assign n364 = ~n358 & n363;
  assign n365 = ~n357 & n364;
  assign n366 = ~n356 & n365;
  assign n367 = n87 & n195;
  assign n368 = n87 & n126;
  assign n369 = ~n127 & ~n368;
  assign n370 = n173 & n205;
  assign n371 = n369 & ~n370;
  assign n372 = ~n367 & n371;
  assign n373 = ~n106 & ~n215;
  assign n374 = n372 & n373;
  assign n375 = n366 & n374;
  assign n376 = n355 & n375;
  assign n377 = ~n174 & n376;
  assign n378 = ~n133 & n377;
  assign n379 = ~n146 & n378;
  assign n380 = ~n223 & n379;
  assign n381 = n156 & n380;
  assign n382 = ~n350 & n381;
  assign n383 = n349 & n382;
  assign n384 = n346 & n383;
  assign n385 = n259 & n384;
  assign n386 = n344 & n385;
  assign n387 = n341 & n386;
  assign n388 = n334 & n387;
  assign n389 = n325 & n388;
  assign n390 = n323 & n389;
  assign n391 = n311 & n390;
  assign n392 = ~n208 & n391;
  assign n393 = ~n134 & n392;
  assign n394 = n125 & n195;
  assign n395 = ~n192 & ~n350;
  assign n396 = ~n174 & ~n337;
  assign n397 = ~n207 & ~n327;
  assign n398 = n396 & n397;
  assign n399 = n314 & n398;
  assign n400 = n141 & n399;
  assign n401 = ~n208 & n400;
  assign n402 = ~n228 & n401;
  assign n403 = n395 & n402;
  assign n404 = ~n167 & n403;
  assign n405 = n117 & n125;
  assign n406 = ~n137 & ~n257;
  assign n407 = ~n336 & n406;
  assign n408 = n117 & n128;
  assign n409 = ~n138 & ~n408;
  assign n410 = ~n220 & n409;
  assign n411 = ~n299 & n410;
  assign n412 = n407 & n411;
  assign n413 = ~n405 & n412;
  assign n414 = ~n123 & n413;
  assign n415 = n128 & n171;
  assign n416 = ~n255 & ~n415;
  assign n417 = n143 & n173;
  assign n418 = n153 & n189;
  assign n419 = ~n127 & n418;
  assign n420 = ~n219 & n419;
  assign n421 = ~n225 & n420;
  assign n422 = ~n417 & n421;
  assign n423 = ~n218 & n422;
  assign n424 = n416 & n423;
  assign n425 = n414 & n424;
  assign n426 = ~n222 & n425;
  assign n427 = ~n144 & n426;
  assign n428 = ~n129 & n427;
  assign n429 = ~n176 & n428;
  assign n430 = ~n214 & n429;
  assign n431 = ~n134 & n430;
  assign n432 = ~n155 & ~n194;
  assign n433 = ~n178 & ~n227;
  assign n434 = ~n175 & n433;
  assign n435 = ~n312 & n434;
  assign n436 = ~n226 & n435;
  assign n437 = ~n133 & n436;
  assign n438 = n432 & n437;
  assign n439 = n431 & n438;
  assign n440 = n404 & n439;
  assign n441 = ~n328 & n440;
  assign n442 = ~n196 & n441;
  assign n443 = ~n317 & n442;
  assign n444 = ~n394 & n443;
  assign n445 = n87 & n122;
  assign n446 = n120 & n171;
  assign n447 = n115 & n151;
  assign n448 = ~n190 & ~n447;
  assign n449 = n115 & n143;
  assign n450 = ~n297 & ~n449;
  assign n451 = ~n166 & n450;
  assign n452 = n448 & n451;
  assign n453 = ~n146 & n452;
  assign n454 = ~n254 & ~n343;
  assign n455 = ~n224 & n454;
  assign n456 = ~n212 & n455;
  assign n457 = ~n142 & n456;
  assign n458 = n120 & n193;
  assign n459 = ~n300 & ~n458;
  assign n460 = ~n360 & ~n370;
  assign n461 = n349 & n460;
  assign n462 = n459 & n461;
  assign n463 = n457 & n462;
  assign n464 = n453 & n463;
  assign n465 = ~n213 & n464;
  assign n466 = ~n446 & n465;
  assign n467 = ~n111 & n466;
  assign n468 = n113 & n130;
  assign n469 = n126 & n130;
  assign n470 = n87 & n108;
  assign n471 = n130 & n195;
  assign n472 = n87 & n143;
  assign n473 = ~n177 & ~n329;
  assign n474 = ~n235 & ~n356;
  assign n475 = ~n191 & ~n217;
  assign n476 = ~n172 & n475;
  assign n477 = n130 & n143;
  assign n478 = ~n342 & ~n477;
  assign n479 = n476 & n478;
  assign n480 = n474 & n479;
  assign n481 = n473 & n480;
  assign n482 = ~n106 & n481;
  assign n483 = ~n367 & n482;
  assign n484 = ~n472 & n483;
  assign n485 = ~n471 & n484;
  assign n486 = ~n470 & n485;
  assign n487 = ~n168 & n486;
  assign n488 = ~n296 & n487;
  assign n489 = ~n469 & n488;
  assign n490 = ~n468 & n489;
  assign n491 = n467 & n490;
  assign n492 = ~n368 & n491;
  assign n493 = ~n445 & n492;
  assign n494 = ~n223 & n493;
  assign n495 = n115 & n193;
  assign n496 = ~n118 & ~n335;
  assign n497 = ~n495 & n496;
  assign n498 = ~n358 & n497;
  assign n499 = ~n315 & n498;
  assign n500 = ~n234 & n499;
  assign n501 = ~n206 & n500;
  assign n502 = ~n359 & n501;
  assign n503 = n110 & n122;
  assign n504 = n115 & n136;
  assign n505 = ~n216 & ~n504;
  assign n506 = n110 & n131;
  assign n507 = ~n357 & ~n361;
  assign n508 = ~n506 & n507;
  assign n509 = n505 & n508;
  assign n510 = ~n302 & n509;
  assign n511 = ~n298 & n510;
  assign n512 = ~n169 & n511;
  assign n513 = ~n114 & n512;
  assign n514 = ~n503 & n513;
  assign n515 = n467 & n514;
  assign n516 = n475 & n515;
  assign n517 = n473 & n516;
  assign n518 = n502 & n517;
  assign n519 = ~n148 & n518;
  assign n520 = ~n494 & ~n519;
  assign n521 = \a[14]  & \a[22] ;
  assign n522 = \a[14]  & ~n63;
  assign n523 = ~n64 & ~n522;
  assign n524 = ~\a[22]  & n523;
  assign n525 = ~n521 & ~n524;
  assign n526 = ~\a[22]  & ~n62;
  assign n527 = \a[13]  & ~n526;
  assign n528 = ~\a[13]  & n526;
  assign n529 = ~n527 & ~n528;
  assign n530 = ~n525 & n529;
  assign n531 = n525 & ~n529;
  assign n532 = ~n530 & ~n531;
  assign n533 = n520 & n532;
  assign n534 = ~n520 & ~n532;
  assign n535 = ~n533 & ~n534;
  assign n536 = ~n444 & n535;
  assign n537 = n494 & ~n519;
  assign n538 = ~n494 & n519;
  assign n539 = ~n537 & ~n538;
  assign n540 = n494 & n519;
  assign n541 = n444 & ~n540;
  assign n542 = n539 & ~n541;
  assign n543 = ~n525 & n542;
  assign n544 = ~n444 & ~n520;
  assign n545 = ~n539 & ~n544;
  assign n546 = n525 & ~n544;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~n543 & n547;
  assign n549 = ~n444 & ~n529;
  assign n550 = n548 & ~n549;
  assign n551 = ~n548 & n549;
  assign n552 = n87 & n136;
  assign n553 = n87 & n205;
  assign n554 = n87 & n131;
  assign n555 = ~n238 & ~n554;
  assign n556 = ~n208 & n555;
  assign n557 = ~n221 & n556;
  assign n558 = ~n367 & n557;
  assign n559 = ~n225 & ~n417;
  assign n560 = ~n296 & n559;
  assign n561 = ~n234 & ~n471;
  assign n562 = ~n237 & n561;
  assign n563 = ~n227 & ~n394;
  assign n564 = ~n127 & n563;
  assign n565 = n562 & n564;
  assign n566 = n560 & n565;
  assign n567 = n558 & n566;
  assign n568 = n185 & n567;
  assign n569 = ~n129 & n568;
  assign n570 = ~n348 & n569;
  assign n571 = ~n553 & n570;
  assign n572 = ~n167 & ~n220;
  assign n573 = ~n191 & n572;
  assign n574 = ~n337 & n573;
  assign n575 = ~n360 & n574;
  assign n576 = ~n212 & n575;
  assign n577 = ~n470 & n576;
  assign n578 = ~n118 & ~n196;
  assign n579 = ~n114 & n578;
  assign n580 = ~n503 & n579;
  assign n581 = ~n469 & n580;
  assign n582 = ~n218 & ~n343;
  assign n583 = ~n329 & n582;
  assign n584 = ~n449 & n583;
  assign n585 = ~n298 & ~n347;
  assign n586 = ~n356 & n585;
  assign n587 = n165 & ~n228;
  assign n588 = ~n359 & n587;
  assign n589 = n87 & n187;
  assign n590 = ~n186 & ~n589;
  assign n591 = n588 & n590;
  assign n592 = n586 & n591;
  assign n593 = n584 & n592;
  assign n594 = n581 & n593;
  assign n595 = n577 & n594;
  assign n596 = n571 & n595;
  assign n597 = n355 & n596;
  assign n598 = ~n552 & n597;
  assign n599 = n87 & n117;
  assign n600 = n141 & n373;
  assign n601 = ~n220 & n600;
  assign n602 = ~n134 & n601;
  assign n603 = ~n172 & n602;
  assign n604 = ~n298 & n603;
  assign n605 = ~n506 & n604;
  assign n606 = ~n554 & n605;
  assign n607 = ~n222 & ~n337;
  assign n608 = ~n114 & n607;
  assign n609 = ~n317 & ~n405;
  assign n610 = n474 & n609;
  assign n611 = ~n227 & n610;
  assign n612 = ~n348 & n611;
  assign n613 = ~n329 & n612;
  assign n614 = ~n154 & n613;
  assign n615 = n153 & n432;
  assign n616 = n505 & n615;
  assign n617 = n614 & n616;
  assign n618 = ~n408 & n617;
  assign n619 = ~n188 & n618;
  assign n620 = ~n129 & n619;
  assign n621 = ~n217 & n620;
  assign n622 = ~n357 & n621;
  assign n623 = ~n326 & n622;
  assign n624 = ~n394 & n623;
  assign n625 = ~n351 & n624;
  assign n626 = ~n208 & ~n214;
  assign n627 = ~n137 & n626;
  assign n628 = ~n169 & n627;
  assign n629 = n625 & n628;
  assign n630 = n344 & n629;
  assign n631 = n608 & n630;
  assign n632 = n606 & n631;
  assign n633 = ~n191 & n632;
  assign n634 = ~n446 & n633;
  assign n635 = ~n599 & n634;
  assign n636 = ~n211 & n635;
  assign n637 = ~n312 & ~n415;
  assign n638 = ~n176 & ~n503;
  assign n639 = n637 & n638;
  assign n640 = ~n196 & n639;
  assign n641 = ~n175 & n640;
  assign n642 = ~n300 & n641;
  assign n643 = ~n302 & n642;
  assign n644 = ~n213 & ~n472;
  assign n645 = ~n138 & ~n228;
  assign n646 = ~n477 & n645;
  assign n647 = ~n127 & ~n328;
  assign n648 = ~n370 & n647;
  assign n649 = n256 & n648;
  assign n650 = ~n144 & n649;
  assign n651 = ~n221 & n650;
  assign n652 = ~n471 & n651;
  assign n653 = ~n132 & n652;
  assign n654 = ~n219 & n653;
  assign n655 = ~n458 & n654;
  assign n656 = n179 & n655;
  assign n657 = n646 & n656;
  assign n658 = n644 & n657;
  assign n659 = n643 & n658;
  assign n660 = n636 & n659;
  assign n661 = n362 & n660;
  assign n662 = ~n552 & n661;
  assign n663 = ~n367 & n662;
  assign n664 = ~n598 & ~n663;
  assign n665 = ~n494 & ~n664;
  assign n666 = ~\a[22]  & ~n60;
  assign n667 = \a[11]  & ~n666;
  assign n668 = ~\a[11]  & n666;
  assign n669 = ~n667 & ~n668;
  assign n670 = ~n444 & ~n669;
  assign n671 = ~n665 & n670;
  assign n672 = n665 & ~n670;
  assign n673 = ~n671 & ~n672;
  assign n674 = \a[12]  & \a[22] ;
  assign n675 = \a[12]  & ~n61;
  assign n676 = n526 & ~n675;
  assign n677 = ~n674 & ~n676;
  assign n678 = ~n444 & ~n677;
  assign n679 = n673 & n678;
  assign n680 = ~n671 & ~n679;
  assign n681 = ~n550 & ~n680;
  assign n682 = ~n551 & n681;
  assign n683 = ~n550 & ~n682;
  assign n684 = ~n539 & ~n541;
  assign n685 = ~n525 & n684;
  assign n686 = n525 & n545;
  assign n687 = n539 & ~n544;
  assign n688 = n529 & n687;
  assign n689 = ~n529 & n542;
  assign n690 = ~n688 & ~n689;
  assign n691 = ~n686 & n690;
  assign n692 = ~n685 & n691;
  assign n693 = n598 & ~n663;
  assign n694 = ~n598 & n663;
  assign n695 = ~n693 & ~n694;
  assign n696 = n598 & n663;
  assign n697 = n494 & ~n696;
  assign n698 = n695 & ~n697;
  assign n699 = ~n525 & n698;
  assign n700 = ~n665 & ~n695;
  assign n701 = n525 & ~n665;
  assign n702 = ~n700 & ~n701;
  assign n703 = ~n699 & n702;
  assign n704 = ~n670 & n703;
  assign n705 = ~n529 & n684;
  assign n706 = n529 & n545;
  assign n707 = n677 & n687;
  assign n708 = n542 & ~n677;
  assign n709 = ~n707 & ~n708;
  assign n710 = ~n706 & n709;
  assign n711 = ~n705 & n710;
  assign n712 = n670 & ~n703;
  assign n713 = ~n704 & ~n712;
  assign n714 = n711 & n713;
  assign n715 = ~n704 & ~n714;
  assign n716 = n692 & ~n715;
  assign n717 = ~n692 & n715;
  assign n718 = ~n716 & ~n717;
  assign n719 = ~n673 & ~n678;
  assign n720 = ~n679 & ~n719;
  assign n721 = n718 & n720;
  assign n722 = ~n716 & ~n721;
  assign n723 = ~n680 & ~n682;
  assign n724 = ~n551 & n683;
  assign n725 = ~n723 & ~n724;
  assign n726 = ~n722 & n725;
  assign n727 = n722 & ~n725;
  assign n728 = ~n726 & ~n727;
  assign n729 = ~n222 & ~n415;
  assign n730 = ~n219 & n729;
  assign n731 = ~n359 & n730;
  assign n732 = ~n166 & n731;
  assign n733 = ~n470 & n732;
  assign n734 = ~n368 & n733;
  assign n735 = ~n345 & n734;
  assign n736 = n130 & n193;
  assign n737 = ~n123 & ~n167;
  assign n738 = ~n216 & n737;
  assign n739 = ~n736 & n738;
  assign n740 = ~n337 & ~n495;
  assign n741 = ~n503 & n740;
  assign n742 = ~n506 & n741;
  assign n743 = ~n351 & n742;
  assign n744 = ~n235 & n743;
  assign n745 = n476 & n744;
  assign n746 = n739 & n745;
  assign n747 = ~n139 & n746;
  assign n748 = ~n504 & n747;
  assign n749 = ~n297 & n748;
  assign n750 = ~n206 & n749;
  assign n751 = ~n106 & n750;
  assign n752 = ~n238 & n751;
  assign n753 = ~n132 & ~n298;
  assign n754 = ~n348 & n645;
  assign n755 = ~n350 & n754;
  assign n756 = ~n218 & n755;
  assign n757 = ~n148 & n756;
  assign n758 = ~n177 & ~n211;
  assign n759 = ~n215 & n758;
  assign n760 = ~n212 & ~n472;
  assign n761 = n759 & n760;
  assign n762 = n757 & n761;
  assign n763 = n753 & n762;
  assign n764 = ~n188 & n763;
  assign n765 = ~n257 & n764;
  assign n766 = ~n142 & n765;
  assign n767 = ~n552 & n766;
  assign n768 = ~n445 & n767;
  assign n769 = ~n137 & ~n313;
  assign n770 = ~n447 & n769;
  assign n771 = ~n315 & n770;
  assign n772 = ~n168 & n771;
  assign n773 = ~n471 & n772;
  assign n774 = ~n214 & ~n405;
  assign n775 = ~n302 & n774;
  assign n776 = ~n254 & ~n300;
  assign n777 = ~n225 & n776;
  assign n778 = n775 & n777;
  assign n779 = n773 & n778;
  assign n780 = n768 & n779;
  assign n781 = n752 & n780;
  assign n782 = n735 & n781;
  assign n783 = ~n408 & n782;
  assign n784 = ~n226 & n783;
  assign n785 = ~n133 & n784;
  assign n786 = ~n237 & n785;
  assign n787 = ~n166 & ~n226;
  assign n788 = ~n237 & n787;
  assign n789 = ~n477 & n788;
  assign n790 = ~n169 & ~n186;
  assign n791 = ~n347 & n790;
  assign n792 = ~n223 & n791;
  assign n793 = ~n111 & ~n176;
  assign n794 = ~n470 & n793;
  assign n795 = ~n134 & ~n178;
  assign n796 = ~n212 & n795;
  assign n797 = n794 & n796;
  assign n798 = n648 & n797;
  assign n799 = n792 & n798;
  assign n800 = ~n219 & n799;
  assign n801 = ~n350 & n800;
  assign n802 = ~n417 & n801;
  assign n803 = ~n133 & n802;
  assign n804 = ~n315 & n803;
  assign n805 = ~n106 & n804;
  assign n806 = ~n225 & ~n299;
  assign n807 = ~n123 & ~n175;
  assign n808 = ~n144 & ~n336;
  assign n809 = ~n458 & ~n589;
  assign n810 = n301 & n809;
  assign n811 = n149 & n810;
  assign n812 = ~n258 & n811;
  assign n813 = ~n368 & n812;
  assign n814 = ~n297 & n813;
  assign n815 = ~n206 & n814;
  assign n816 = n625 & n815;
  assign n817 = n808 & n816;
  assign n818 = n807 & n817;
  assign n819 = n806 & n818;
  assign n820 = n805 & n819;
  assign n821 = n789 & n820;
  assign n822 = ~n172 & n821;
  assign n823 = n578 & n822;
  assign n824 = ~n358 & n823;
  assign n825 = ~n736 & n824;
  assign n826 = ~n296 & n825;
  assign n827 = ~n786 & ~n826;
  assign n828 = ~n598 & ~n827;
  assign n829 = ~\a[22]  & ~n58;
  assign n830 = \a[9]  & ~n829;
  assign n831 = ~\a[9]  & n829;
  assign n832 = ~n830 & ~n831;
  assign n833 = ~n444 & ~n832;
  assign n834 = ~n828 & n833;
  assign n835 = n828 & ~n833;
  assign n836 = ~n834 & ~n835;
  assign n837 = \a[10]  & \a[22] ;
  assign n838 = \a[10]  & ~n59;
  assign n839 = n666 & ~n838;
  assign n840 = ~n837 & ~n839;
  assign n841 = ~n444 & ~n840;
  assign n842 = n836 & n841;
  assign n843 = ~n834 & ~n842;
  assign n844 = ~n695 & ~n697;
  assign n845 = ~n525 & n844;
  assign n846 = n525 & n700;
  assign n847 = ~n665 & n695;
  assign n848 = n529 & n847;
  assign n849 = ~n529 & n698;
  assign n850 = ~n848 & ~n849;
  assign n851 = ~n846 & n850;
  assign n852 = ~n845 & n851;
  assign n853 = ~n677 & n684;
  assign n854 = n545 & n677;
  assign n855 = n669 & n687;
  assign n856 = n542 & ~n669;
  assign n857 = ~n855 & ~n856;
  assign n858 = ~n854 & n857;
  assign n859 = ~n853 & n858;
  assign n860 = n852 & n859;
  assign n861 = n786 & ~n826;
  assign n862 = ~n786 & n826;
  assign n863 = ~n861 & ~n862;
  assign n864 = n786 & n826;
  assign n865 = n598 & ~n864;
  assign n866 = n863 & ~n865;
  assign n867 = ~n525 & n866;
  assign n868 = ~n828 & ~n863;
  assign n869 = n525 & ~n828;
  assign n870 = ~n868 & ~n869;
  assign n871 = ~n867 & n870;
  assign n872 = ~n833 & n871;
  assign n873 = ~n529 & n844;
  assign n874 = n529 & n700;
  assign n875 = n677 & n847;
  assign n876 = ~n677 & n698;
  assign n877 = ~n875 & ~n876;
  assign n878 = ~n874 & n877;
  assign n879 = ~n873 & n878;
  assign n880 = n833 & ~n871;
  assign n881 = ~n872 & ~n880;
  assign n882 = n879 & n881;
  assign n883 = ~n872 & ~n882;
  assign n884 = ~n852 & ~n859;
  assign n885 = ~n860 & ~n884;
  assign n886 = ~n883 & n885;
  assign n887 = ~n860 & ~n886;
  assign n888 = ~n843 & ~n887;
  assign n889 = ~n843 & ~n888;
  assign n890 = ~n887 & ~n888;
  assign n891 = ~n889 & ~n890;
  assign n892 = ~n711 & ~n713;
  assign n893 = ~n714 & ~n892;
  assign n894 = ~n891 & n893;
  assign n895 = ~n888 & ~n894;
  assign n896 = ~n718 & ~n720;
  assign n897 = ~n721 & ~n896;
  assign n898 = ~n895 & n897;
  assign n899 = ~n669 & n684;
  assign n900 = n545 & n669;
  assign n901 = n687 & n840;
  assign n902 = n542 & ~n840;
  assign n903 = ~n901 & ~n902;
  assign n904 = ~n900 & n903;
  assign n905 = ~n899 & n904;
  assign n906 = ~n166 & ~n446;
  assign n907 = n145 & n906;
  assign n908 = ~n552 & n907;
  assign n909 = ~n238 & n908;
  assign n910 = ~n296 & n909;
  assign n911 = ~n174 & ~n470;
  assign n912 = ~n222 & n911;
  assign n913 = ~n350 & n912;
  assign n914 = ~n345 & n913;
  assign n915 = n303 & n914;
  assign n916 = n323 & n915;
  assign n917 = n910 & n916;
  assign n918 = ~n152 & n917;
  assign n919 = ~n196 & n918;
  assign n920 = ~n186 & n919;
  assign n921 = ~n504 & n920;
  assign n922 = ~n495 & n921;
  assign n923 = ~n154 & n922;
  assign n924 = ~n370 & ~n468;
  assign n925 = ~n347 & n924;
  assign n926 = ~n445 & n925;
  assign n927 = ~n127 & n407;
  assign n928 = ~n216 & n927;
  assign n929 = ~n589 & n928;
  assign n930 = ~n367 & n929;
  assign n931 = ~n139 & ~n327;
  assign n932 = n562 & n638;
  assign n933 = n931 & n932;
  assign n934 = n930 & n933;
  assign n935 = n926 & n934;
  assign n936 = ~n219 & n935;
  assign n937 = ~n299 & n936;
  assign n938 = ~n148 & n937;
  assign n939 = ~n177 & ~n214;
  assign n940 = ~n218 & n939;
  assign n941 = ~n192 & n940;
  assign n942 = ~n133 & n941;
  assign n943 = ~n736 & n942;
  assign n944 = ~n342 & n943;
  assign n945 = ~n190 & ~n394;
  assign n946 = ~n235 & n945;
  assign n947 = ~n155 & ~n405;
  assign n948 = ~n351 & n947;
  assign n949 = n496 & n573;
  assign n950 = n948 & n949;
  assign n951 = n946 & n950;
  assign n952 = n325 & n951;
  assign n953 = n944 & n952;
  assign n954 = n938 & n953;
  assign n955 = n923 & n954;
  assign n956 = ~n300 & n955;
  assign n957 = ~n255 & n956;
  assign n958 = ~n258 & n957;
  assign n959 = ~n553 & n958;
  assign n960 = ~n169 & ~n360;
  assign n961 = ~n447 & n960;
  assign n962 = ~n155 & n961;
  assign n963 = ~n350 & n962;
  assign n964 = ~n218 & n963;
  assign n965 = ~n234 & n964;
  assign n966 = ~n359 & n965;
  assign n967 = ~n357 & n966;
  assign n968 = ~n133 & ~n257;
  assign n969 = ~n368 & n968;
  assign n970 = ~n469 & ~n471;
  assign n971 = n969 & n970;
  assign n972 = ~n144 & n971;
  assign n973 = ~n327 & n972;
  assign n974 = ~n446 & n973;
  assign n975 = ~n315 & n974;
  assign n976 = ~n190 & ~n302;
  assign n977 = ~n174 & n976;
  assign n978 = ~n191 & n977;
  assign n979 = ~n168 & n978;
  assign n980 = ~n222 & ~n408;
  assign n981 = ~n394 & n980;
  assign n982 = ~n228 & n981;
  assign n983 = ~n417 & n982;
  assign n984 = ~n129 & ~n178;
  assign n985 = ~n196 & n984;
  assign n986 = ~n449 & n985;
  assign n987 = n256 & n986;
  assign n988 = n983 & n987;
  assign n989 = n926 & n988;
  assign n990 = ~n328 & n989;
  assign n991 = ~n176 & n990;
  assign n992 = ~n220 & n991;
  assign n993 = ~n172 & n992;
  assign n994 = n787 & n993;
  assign n995 = ~n223 & n994;
  assign n996 = ~n337 & n995;
  assign n997 = ~n175 & n996;
  assign n998 = ~n552 & n997;
  assign n999 = ~n351 & n998;
  assign n1000 = n979 & n999;
  assign n1001 = n141 & n1000;
  assign n1002 = n975 & n1001;
  assign n1003 = n967 & n1002;
  assign n1004 = n614 & n1003;
  assign n1005 = ~n299 & n1004;
  assign n1006 = ~n503 & n1005;
  assign n1007 = ~n367 & n1006;
  assign n1008 = ~n959 & ~n1007;
  assign n1009 = ~n786 & ~n1008;
  assign n1010 = ~\a[22]  & ~n56;
  assign n1011 = \a[7]  & ~n1010;
  assign n1012 = ~\a[7]  & n1010;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = ~n444 & ~n1013;
  assign n1015 = ~n1009 & n1014;
  assign n1016 = n1009 & ~n1014;
  assign n1017 = ~n1015 & ~n1016;
  assign n1018 = \a[8]  & \a[22] ;
  assign n1019 = \a[8]  & ~n57;
  assign n1020 = n829 & ~n1019;
  assign n1021 = ~n1018 & ~n1020;
  assign n1022 = n1017 & ~n1021;
  assign n1023 = ~n444 & n1022;
  assign n1024 = ~n1015 & ~n1023;
  assign n1025 = n905 & ~n1024;
  assign n1026 = n684 & ~n840;
  assign n1027 = n545 & n840;
  assign n1028 = n687 & n832;
  assign n1029 = n542 & ~n832;
  assign n1030 = ~n1028 & ~n1029;
  assign n1031 = ~n1027 & n1030;
  assign n1032 = ~n1026 & n1031;
  assign n1033 = ~n863 & ~n865;
  assign n1034 = ~n525 & n1033;
  assign n1035 = n525 & n868;
  assign n1036 = ~n828 & n863;
  assign n1037 = n529 & n1036;
  assign n1038 = ~n529 & n866;
  assign n1039 = ~n1037 & ~n1038;
  assign n1040 = ~n1035 & n1039;
  assign n1041 = ~n1034 & n1040;
  assign n1042 = ~n677 & n844;
  assign n1043 = n677 & n700;
  assign n1044 = n669 & n847;
  assign n1045 = ~n669 & n698;
  assign n1046 = ~n1044 & ~n1045;
  assign n1047 = ~n1043 & n1046;
  assign n1048 = ~n1042 & n1047;
  assign n1049 = n1041 & ~n1048;
  assign n1050 = ~n1041 & n1048;
  assign n1051 = ~n1049 & ~n1050;
  assign n1052 = n1032 & ~n1051;
  assign n1053 = n1041 & n1048;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = n905 & ~n1025;
  assign n1056 = ~n1024 & ~n1025;
  assign n1057 = ~n1055 & ~n1056;
  assign n1058 = ~n1054 & ~n1057;
  assign n1059 = ~n1025 & ~n1058;
  assign n1060 = ~n836 & ~n841;
  assign n1061 = ~n842 & ~n1060;
  assign n1062 = ~n1059 & n1061;
  assign n1063 = n1059 & ~n1061;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = n883 & ~n885;
  assign n1066 = ~n886 & ~n1065;
  assign n1067 = n1064 & n1066;
  assign n1068 = ~n1062 & ~n1067;
  assign n1069 = ~n891 & ~n894;
  assign n1070 = n893 & ~n894;
  assign n1071 = ~n1069 & ~n1070;
  assign n1072 = ~n1068 & n1071;
  assign n1073 = n1068 & ~n1071;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = ~n669 & n844;
  assign n1076 = n669 & n700;
  assign n1077 = n840 & n847;
  assign n1078 = n698 & ~n840;
  assign n1079 = ~n1077 & ~n1078;
  assign n1080 = ~n1076 & n1079;
  assign n1081 = ~n1075 & n1080;
  assign n1082 = n684 & ~n832;
  assign n1083 = n545 & n832;
  assign n1084 = n687 & n1021;
  assign n1085 = n542 & ~n1021;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = ~n1083 & n1086;
  assign n1088 = ~n1082 & n1087;
  assign n1089 = n1081 & n1088;
  assign n1090 = ~n348 & ~n495;
  assign n1091 = ~n335 & n1090;
  assign n1092 = ~n226 & ~n446;
  assign n1093 = ~n553 & n1092;
  assign n1094 = ~n175 & ~n343;
  assign n1095 = ~n503 & n1094;
  assign n1096 = ~n472 & n1095;
  assign n1097 = n1093 & n1096;
  assign n1098 = n1091 & n1097;
  assign n1099 = n983 & n1098;
  assign n1100 = n149 & n1099;
  assign n1101 = ~n196 & n1100;
  assign n1102 = ~n327 & n1101;
  assign n1103 = ~n212 & n1102;
  assign n1104 = ~n469 & n1103;
  assign n1105 = ~n118 & n395;
  assign n1106 = ~n235 & n1105;
  assign n1107 = n448 & n1106;
  assign n1108 = ~n224 & n1107;
  assign n1109 = n460 & ~n468;
  assign n1110 = ~n176 & n1109;
  assign n1111 = ~n214 & n1110;
  assign n1112 = ~n218 & n1111;
  assign n1113 = ~n504 & n1112;
  assign n1114 = ~n358 & n1113;
  assign n1115 = ~n345 & n1114;
  assign n1116 = ~n223 & ~n599;
  assign n1117 = ~n140 & ~n336;
  assign n1118 = n1116 & n1117;
  assign n1119 = n609 & n1118;
  assign n1120 = n558 & n1119;
  assign n1121 = n325 & n1120;
  assign n1122 = n1115 & n1121;
  assign n1123 = n1108 & n1122;
  assign n1124 = n311 & n1123;
  assign n1125 = n1104 & n1124;
  assign n1126 = ~n188 & n1125;
  assign n1127 = ~n133 & n1126;
  assign n1128 = ~n206 & n1127;
  assign n1129 = ~n166 & n1128;
  assign n1130 = ~n552 & n1129;
  assign n1131 = n459 & n1116;
  assign n1132 = n807 & n1131;
  assign n1133 = ~n220 & n1132;
  assign n1134 = ~n394 & n1133;
  assign n1135 = n646 & n948;
  assign n1136 = n314 & n1135;
  assign n1137 = n1108 & n1136;
  assign n1138 = n1134 & n1137;
  assign n1139 = ~n129 & n1138;
  assign n1140 = ~n196 & n1139;
  assign n1141 = ~n150 & n1140;
  assign n1142 = ~n213 & n1141;
  assign n1143 = ~n169 & n1142;
  assign n1144 = ~n315 & n1143;
  assign n1145 = ~n326 & n1144;
  assign n1146 = n637 & n911;
  assign n1147 = ~n194 & n1146;
  assign n1148 = ~n214 & n1147;
  assign n1149 = ~n348 & n1148;
  assign n1150 = ~n299 & n1149;
  assign n1151 = ~n552 & n1150;
  assign n1152 = ~n736 & n1151;
  assign n1153 = n560 & n969;
  assign n1154 = ~n324 & n1153;
  assign n1155 = n1152 & n1154;
  assign n1156 = n475 & n1155;
  assign n1157 = ~n167 & n1156;
  assign n1158 = ~n336 & n1157;
  assign n1159 = ~n258 & n1158;
  assign n1160 = ~n345 & n1159;
  assign n1161 = ~n154 & n1160;
  assign n1162 = ~n215 & n1161;
  assign n1163 = ~n208 & ~n408;
  assign n1164 = ~n142 & n1163;
  assign n1165 = ~n111 & n1164;
  assign n1166 = n760 & n1165;
  assign n1167 = n451 & n1166;
  assign n1168 = n505 & n1167;
  assign n1169 = n366 & n1168;
  assign n1170 = n141 & n1169;
  assign n1171 = n1162 & n1170;
  assign n1172 = n1145 & n1171;
  assign n1173 = ~n152 & n1172;
  assign n1174 = ~n219 & n1173;
  assign n1175 = ~n335 & n1174;
  assign n1176 = ~n1130 & ~n1175;
  assign n1177 = ~n959 & ~n1176;
  assign n1178 = n1130 & ~n1177;
  assign n1179 = ~n1130 & n1177;
  assign n1180 = \a[6]  & \a[22] ;
  assign n1181 = \a[6]  & ~n55;
  assign n1182 = n1010 & ~n1181;
  assign n1183 = ~n1180 & ~n1182;
  assign n1184 = ~n444 & ~n1183;
  assign n1185 = ~n1178 & n1184;
  assign n1186 = ~n1179 & n1185;
  assign n1187 = ~n1178 & ~n1186;
  assign n1188 = ~n1081 & ~n1088;
  assign n1189 = ~n1089 & ~n1188;
  assign n1190 = ~n1187 & n1189;
  assign n1191 = ~n1089 & ~n1190;
  assign n1192 = n959 & ~n1007;
  assign n1193 = ~n959 & n1007;
  assign n1194 = ~n1192 & ~n1193;
  assign n1195 = n959 & n1007;
  assign n1196 = n786 & ~n1195;
  assign n1197 = n1194 & ~n1196;
  assign n1198 = ~n525 & n1197;
  assign n1199 = ~n1009 & ~n1194;
  assign n1200 = n525 & ~n1009;
  assign n1201 = ~n1199 & ~n1200;
  assign n1202 = ~n1198 & n1201;
  assign n1203 = ~n1014 & n1202;
  assign n1204 = ~n529 & n1033;
  assign n1205 = n529 & n868;
  assign n1206 = n677 & n1036;
  assign n1207 = ~n677 & n866;
  assign n1208 = ~n1206 & ~n1207;
  assign n1209 = ~n1205 & n1208;
  assign n1210 = ~n1204 & n1209;
  assign n1211 = n1014 & ~n1202;
  assign n1212 = ~n1203 & ~n1211;
  assign n1213 = n1210 & n1212;
  assign n1214 = ~n1203 & ~n1213;
  assign n1215 = ~n1191 & ~n1214;
  assign n1216 = ~n1191 & ~n1215;
  assign n1217 = ~n1214 & ~n1215;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = ~n444 & ~n1023;
  assign n1220 = ~n1021 & n1219;
  assign n1221 = n1017 & ~n1023;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = ~n1218 & ~n1222;
  assign n1224 = ~n1215 & ~n1223;
  assign n1225 = ~n879 & ~n881;
  assign n1226 = ~n882 & ~n1225;
  assign n1227 = ~n1224 & n1226;
  assign n1228 = ~n1054 & ~n1058;
  assign n1229 = ~n1057 & ~n1058;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = n1224 & ~n1226;
  assign n1232 = ~n1227 & ~n1231;
  assign n1233 = ~n1230 & n1232;
  assign n1234 = ~n1227 & ~n1233;
  assign n1235 = ~n1064 & ~n1066;
  assign n1236 = ~n1067 & ~n1235;
  assign n1237 = ~n1234 & n1236;
  assign n1238 = n1232 & ~n1233;
  assign n1239 = ~n1230 & ~n1233;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = ~n1194 & ~n1196;
  assign n1242 = ~n525 & n1241;
  assign n1243 = n525 & n1199;
  assign n1244 = ~n1009 & n1194;
  assign n1245 = n529 & n1244;
  assign n1246 = ~n529 & n1197;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = ~n1243 & n1247;
  assign n1249 = ~n1242 & n1248;
  assign n1250 = ~n840 & n844;
  assign n1251 = n700 & n840;
  assign n1252 = n832 & n847;
  assign n1253 = n698 & ~n832;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = ~n1251 & n1254;
  assign n1256 = ~n1250 & n1255;
  assign n1257 = n684 & ~n1021;
  assign n1258 = n545 & n1021;
  assign n1259 = n687 & n1013;
  assign n1260 = n542 & ~n1013;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = ~n1258 & n1261;
  assign n1263 = ~n1257 & n1262;
  assign n1264 = n1256 & ~n1263;
  assign n1265 = ~n1256 & n1263;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = n1249 & ~n1266;
  assign n1268 = n1256 & n1263;
  assign n1269 = ~n1267 & ~n1268;
  assign n1270 = ~n1210 & ~n1212;
  assign n1271 = ~n1213 & ~n1270;
  assign n1272 = ~n1269 & n1271;
  assign n1273 = ~n1269 & ~n1272;
  assign n1274 = n1271 & ~n1272;
  assign n1275 = ~n1273 & ~n1274;
  assign n1276 = n1187 & ~n1189;
  assign n1277 = ~n1190 & ~n1276;
  assign n1278 = ~n1275 & n1277;
  assign n1279 = ~n1272 & ~n1278;
  assign n1280 = n1032 & ~n1052;
  assign n1281 = ~n1051 & ~n1052;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = ~n1279 & ~n1282;
  assign n1284 = ~n1279 & ~n1283;
  assign n1285 = ~n1282 & ~n1283;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = ~n1218 & ~n1223;
  assign n1288 = ~n1222 & ~n1223;
  assign n1289 = ~n1287 & ~n1288;
  assign n1290 = ~n1286 & ~n1289;
  assign n1291 = ~n1283 & ~n1290;
  assign n1292 = ~n1240 & ~n1291;
  assign n1293 = ~n1240 & ~n1292;
  assign n1294 = ~n1291 & ~n1292;
  assign n1295 = ~n1293 & ~n1294;
  assign n1296 = ~n677 & n1033;
  assign n1297 = n677 & n868;
  assign n1298 = n669 & n1036;
  assign n1299 = ~n669 & n866;
  assign n1300 = ~n1298 & ~n1299;
  assign n1301 = ~n1297 & n1300;
  assign n1302 = ~n1296 & n1301;
  assign n1303 = ~n1179 & n1187;
  assign n1304 = n1184 & ~n1186;
  assign n1305 = ~n1303 & ~n1304;
  assign n1306 = n1302 & ~n1305;
  assign n1307 = ~n275 & ~n444;
  assign n1308 = ~n1130 & n1307;
  assign n1309 = n1130 & ~n1307;
  assign n1310 = n1130 & ~n1175;
  assign n1311 = ~n1130 & n1175;
  assign n1312 = ~n1310 & ~n1311;
  assign n1313 = n1130 & n1175;
  assign n1314 = n959 & ~n1313;
  assign n1315 = n1312 & ~n1314;
  assign n1316 = ~n525 & n1315;
  assign n1317 = ~n1177 & ~n1312;
  assign n1318 = n525 & ~n1177;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = ~n1316 & n1319;
  assign n1321 = ~n1308 & n1320;
  assign n1322 = ~n1309 & n1321;
  assign n1323 = ~n1308 & ~n1322;
  assign n1324 = ~n1302 & n1305;
  assign n1325 = ~n1306 & ~n1324;
  assign n1326 = ~n1323 & n1325;
  assign n1327 = ~n1306 & ~n1326;
  assign n1328 = ~n529 & n1241;
  assign n1329 = n529 & n1199;
  assign n1330 = n677 & n1244;
  assign n1331 = ~n677 & n1197;
  assign n1332 = ~n1330 & ~n1331;
  assign n1333 = ~n1329 & n1332;
  assign n1334 = ~n1328 & n1333;
  assign n1335 = ~n669 & n1033;
  assign n1336 = n669 & n868;
  assign n1337 = n840 & n1036;
  assign n1338 = ~n840 & n866;
  assign n1339 = ~n1337 & ~n1338;
  assign n1340 = ~n1336 & n1339;
  assign n1341 = ~n1335 & n1340;
  assign n1342 = n1334 & n1341;
  assign n1343 = ~n832 & n844;
  assign n1344 = n700 & n832;
  assign n1345 = n847 & n1021;
  assign n1346 = n698 & ~n1021;
  assign n1347 = ~n1345 & ~n1346;
  assign n1348 = ~n1344 & n1347;
  assign n1349 = ~n1343 & n1348;
  assign n1350 = n1334 & ~n1341;
  assign n1351 = ~n1334 & n1341;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = n1349 & ~n1352;
  assign n1354 = ~n1342 & ~n1353;
  assign n1355 = ~n1249 & n1266;
  assign n1356 = ~n1267 & ~n1355;
  assign n1357 = ~n1354 & n1356;
  assign n1358 = n684 & ~n1013;
  assign n1359 = n545 & n1013;
  assign n1360 = n687 & n1183;
  assign n1361 = n542 & ~n1183;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = ~n1359 & n1362;
  assign n1364 = ~n1358 & n1363;
  assign n1365 = ~n279 & ~n444;
  assign n1366 = ~n1130 & n1365;
  assign n1367 = n1130 & ~n1365;
  assign n1368 = ~n1312 & ~n1314;
  assign n1369 = ~n525 & n1368;
  assign n1370 = n525 & n1317;
  assign n1371 = ~n1177 & n1312;
  assign n1372 = n529 & n1371;
  assign n1373 = ~n529 & n1315;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = ~n1370 & n1374;
  assign n1376 = ~n1369 & n1375;
  assign n1377 = ~n1366 & n1376;
  assign n1378 = ~n1367 & n1377;
  assign n1379 = ~n1366 & ~n1378;
  assign n1380 = n1364 & ~n1379;
  assign n1381 = ~n1364 & n1379;
  assign n1382 = ~n1380 & ~n1381;
  assign n1383 = ~n840 & n1033;
  assign n1384 = n840 & n868;
  assign n1385 = n832 & n1036;
  assign n1386 = ~n832 & n866;
  assign n1387 = ~n1385 & ~n1386;
  assign n1388 = ~n1384 & n1387;
  assign n1389 = ~n1383 & n1388;
  assign n1390 = ~n677 & n1241;
  assign n1391 = n677 & n1199;
  assign n1392 = n669 & n1244;
  assign n1393 = ~n669 & n1197;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = ~n1391 & n1394;
  assign n1396 = ~n1390 & n1395;
  assign n1397 = n1389 & n1396;
  assign n1398 = n844 & ~n1021;
  assign n1399 = n700 & n1021;
  assign n1400 = n847 & n1013;
  assign n1401 = n698 & ~n1013;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = ~n1399 & n1402;
  assign n1404 = ~n1398 & n1403;
  assign n1405 = ~n1389 & n1396;
  assign n1406 = n1389 & ~n1396;
  assign n1407 = ~n1405 & ~n1406;
  assign n1408 = n1404 & ~n1407;
  assign n1409 = ~n1397 & ~n1408;
  assign n1410 = n1382 & ~n1409;
  assign n1411 = ~n1380 & ~n1410;
  assign n1412 = n1354 & ~n1356;
  assign n1413 = ~n1357 & ~n1412;
  assign n1414 = ~n1411 & n1413;
  assign n1415 = ~n1357 & ~n1414;
  assign n1416 = ~n1327 & ~n1415;
  assign n1417 = ~n1327 & ~n1416;
  assign n1418 = ~n1415 & ~n1416;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = n1277 & ~n1278;
  assign n1421 = ~n1275 & ~n1278;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = ~n1419 & ~n1422;
  assign n1424 = ~n1416 & ~n1423;
  assign n1425 = ~n1286 & n1289;
  assign n1426 = n1286 & ~n1289;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = ~n1424 & ~n1427;
  assign n1429 = ~n1419 & ~n1423;
  assign n1430 = ~n1422 & ~n1423;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = ~n1309 & n1323;
  assign n1433 = n1320 & ~n1322;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = n1349 & ~n1353;
  assign n1436 = ~n1352 & ~n1353;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = ~n1434 & ~n1437;
  assign n1439 = ~n1434 & ~n1438;
  assign n1440 = ~n1437 & ~n1438;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = n684 & ~n1183;
  assign n1443 = n545 & n1183;
  assign n1444 = n275 & n687;
  assign n1445 = ~n275 & n542;
  assign n1446 = ~n1444 & ~n1445;
  assign n1447 = ~n1443 & n1446;
  assign n1448 = ~n1442 & n1447;
  assign n1449 = ~n286 & ~n444;
  assign n1450 = ~n221 & n809;
  assign n1451 = ~n174 & n1450;
  assign n1452 = ~n300 & n1451;
  assign n1453 = ~n123 & n1452;
  assign n1454 = ~n212 & n1453;
  assign n1455 = ~n347 & n1454;
  assign n1456 = ~n552 & n1455;
  assign n1457 = ~n553 & n1456;
  assign n1458 = ~n220 & ~n350;
  assign n1459 = ~n315 & n1458;
  assign n1460 = n432 & n584;
  assign n1461 = n1459 & n1460;
  assign n1462 = n968 & n1461;
  assign n1463 = n644 & n1462;
  assign n1464 = ~n337 & n1463;
  assign n1465 = ~n214 & n1464;
  assign n1466 = ~n417 & n1465;
  assign n1467 = ~n234 & n1466;
  assign n1468 = ~n367 & n1467;
  assign n1469 = ~n324 & ~n360;
  assign n1470 = ~n446 & n1469;
  assign n1471 = ~n172 & n1470;
  assign n1472 = ~n503 & n1471;
  assign n1473 = ~n356 & n1472;
  assign n1474 = ~n216 & n1473;
  assign n1475 = ~n342 & n1474;
  assign n1476 = ~n154 & n1475;
  assign n1477 = n373 & n1476;
  assign n1478 = n1468 & n1477;
  assign n1479 = n421 & n1478;
  assign n1480 = n1457 & n1479;
  assign n1481 = ~n178 & n1480;
  assign n1482 = ~n208 & n1481;
  assign n1483 = ~n118 & n1482;
  assign n1484 = ~n361 & n1483;
  assign n1485 = ~n258 & n1484;
  assign n1486 = ~n599 & n1485;
  assign n1487 = ~n211 & n1486;
  assign n1488 = ~n525 & n1487;
  assign n1489 = ~n1130 & ~n1488;
  assign n1490 = n1449 & n1489;
  assign n1491 = ~n529 & n1368;
  assign n1492 = n529 & n1317;
  assign n1493 = n677 & n1371;
  assign n1494 = ~n677 & n1315;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = ~n1492 & n1495;
  assign n1497 = ~n1491 & n1496;
  assign n1498 = ~n1449 & ~n1489;
  assign n1499 = ~n1490 & ~n1498;
  assign n1500 = n1497 & n1499;
  assign n1501 = ~n1490 & ~n1500;
  assign n1502 = n1448 & ~n1501;
  assign n1503 = ~n1448 & n1501;
  assign n1504 = ~n1502 & ~n1503;
  assign n1505 = ~n832 & n1033;
  assign n1506 = n832 & n868;
  assign n1507 = n1021 & n1036;
  assign n1508 = n866 & ~n1021;
  assign n1509 = ~n1507 & ~n1508;
  assign n1510 = ~n1506 & n1509;
  assign n1511 = ~n1505 & n1510;
  assign n1512 = ~n669 & n1241;
  assign n1513 = n669 & n1199;
  assign n1514 = n840 & n1244;
  assign n1515 = ~n840 & n1197;
  assign n1516 = ~n1514 & ~n1515;
  assign n1517 = ~n1513 & n1516;
  assign n1518 = ~n1512 & n1517;
  assign n1519 = n1511 & n1518;
  assign n1520 = n844 & ~n1013;
  assign n1521 = n700 & n1013;
  assign n1522 = n847 & n1183;
  assign n1523 = n698 & ~n1183;
  assign n1524 = ~n1522 & ~n1523;
  assign n1525 = ~n1521 & n1524;
  assign n1526 = ~n1520 & n1525;
  assign n1527 = ~n1511 & n1518;
  assign n1528 = n1511 & ~n1518;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = n1526 & ~n1529;
  assign n1531 = ~n1519 & ~n1530;
  assign n1532 = n1504 & ~n1531;
  assign n1533 = ~n1502 & ~n1532;
  assign n1534 = ~n1441 & ~n1533;
  assign n1535 = ~n1438 & ~n1534;
  assign n1536 = n1323 & ~n1325;
  assign n1537 = ~n1326 & ~n1536;
  assign n1538 = ~n1535 & n1537;
  assign n1539 = n1535 & ~n1537;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = n1411 & ~n1413;
  assign n1542 = ~n1414 & ~n1541;
  assign n1543 = n1540 & n1542;
  assign n1544 = ~n1538 & ~n1543;
  assign n1545 = ~n1431 & ~n1544;
  assign n1546 = n1431 & ~n1544;
  assign n1547 = ~n1431 & n1544;
  assign n1548 = ~n1546 & ~n1547;
  assign n1549 = n1130 & ~n1487;
  assign n1550 = ~n1487 & ~n1549;
  assign n1551 = ~n525 & n1550;
  assign n1552 = n525 & n1549;
  assign n1553 = n529 & ~n1130;
  assign n1554 = n1487 & ~n1553;
  assign n1555 = ~n1552 & ~n1554;
  assign n1556 = ~n1551 & n1555;
  assign n1557 = ~n286 & n684;
  assign n1558 = n286 & ~n544;
  assign n1559 = ~n687 & ~n1558;
  assign n1560 = ~n1557 & n1559;
  assign n1561 = n544 & n1560;
  assign n1562 = n1556 & n1561;
  assign n1563 = ~n275 & n684;
  assign n1564 = n275 & n545;
  assign n1565 = n279 & n687;
  assign n1566 = ~n279 & n542;
  assign n1567 = ~n1565 & ~n1566;
  assign n1568 = ~n1564 & n1567;
  assign n1569 = ~n1563 & n1568;
  assign n1570 = n1562 & n1569;
  assign n1571 = ~n840 & n1241;
  assign n1572 = n840 & n1199;
  assign n1573 = n832 & n1244;
  assign n1574 = ~n832 & n1197;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = ~n1572 & n1575;
  assign n1577 = ~n1571 & n1576;
  assign n1578 = ~n1021 & n1033;
  assign n1579 = n868 & n1021;
  assign n1580 = n1013 & n1036;
  assign n1581 = n866 & ~n1013;
  assign n1582 = ~n1580 & ~n1581;
  assign n1583 = ~n1579 & n1582;
  assign n1584 = ~n1578 & n1583;
  assign n1585 = n844 & ~n1183;
  assign n1586 = n700 & n1183;
  assign n1587 = n275 & n847;
  assign n1588 = ~n275 & n698;
  assign n1589 = ~n1587 & ~n1588;
  assign n1590 = ~n1586 & n1589;
  assign n1591 = ~n1585 & n1590;
  assign n1592 = n1584 & ~n1591;
  assign n1593 = ~n1584 & n1591;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = n1577 & ~n1594;
  assign n1596 = n1584 & n1591;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~n1562 & ~n1569;
  assign n1599 = ~n1570 & ~n1598;
  assign n1600 = ~n1597 & n1599;
  assign n1601 = ~n1570 & ~n1600;
  assign n1602 = ~n1367 & n1379;
  assign n1603 = n1376 & ~n1378;
  assign n1604 = ~n1602 & ~n1603;
  assign n1605 = n1601 & ~n1604;
  assign n1606 = ~n1601 & n1604;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = n1404 & ~n1408;
  assign n1609 = ~n1407 & ~n1408;
  assign n1610 = ~n1608 & ~n1609;
  assign n1611 = ~n1607 & ~n1610;
  assign n1612 = ~n1601 & ~n1604;
  assign n1613 = ~n1611 & ~n1612;
  assign n1614 = ~n1382 & n1409;
  assign n1615 = ~n1410 & ~n1614;
  assign n1616 = ~n1613 & n1615;
  assign n1617 = n1441 & ~n1533;
  assign n1618 = ~n1441 & n1533;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = n1613 & ~n1615;
  assign n1621 = ~n1616 & ~n1620;
  assign n1622 = ~n1619 & n1621;
  assign n1623 = ~n1616 & ~n1622;
  assign n1624 = ~n1540 & ~n1542;
  assign n1625 = ~n1543 & ~n1624;
  assign n1626 = ~n1623 & n1625;
  assign n1627 = ~n677 & n1368;
  assign n1628 = n677 & n1317;
  assign n1629 = n669 & n1371;
  assign n1630 = ~n669 & n1315;
  assign n1631 = ~n1629 & ~n1630;
  assign n1632 = ~n1628 & n1631;
  assign n1633 = ~n1627 & n1632;
  assign n1634 = ~n279 & n684;
  assign n1635 = n279 & n545;
  assign n1636 = n286 & n687;
  assign n1637 = ~n286 & n542;
  assign n1638 = ~n1636 & ~n1637;
  assign n1639 = ~n1635 & n1638;
  assign n1640 = ~n1634 & n1639;
  assign n1641 = n1633 & n1640;
  assign n1642 = ~n1556 & ~n1561;
  assign n1643 = ~n1562 & ~n1642;
  assign n1644 = ~n1633 & ~n1640;
  assign n1645 = ~n1641 & ~n1644;
  assign n1646 = n1643 & n1645;
  assign n1647 = ~n1641 & ~n1646;
  assign n1648 = ~n1497 & ~n1499;
  assign n1649 = ~n1500 & ~n1648;
  assign n1650 = ~n1647 & n1649;
  assign n1651 = n1647 & ~n1649;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = n1526 & ~n1530;
  assign n1654 = ~n1529 & ~n1530;
  assign n1655 = ~n1653 & ~n1654;
  assign n1656 = n1652 & ~n1655;
  assign n1657 = ~n1650 & ~n1656;
  assign n1658 = ~n1504 & n1531;
  assign n1659 = ~n1532 & ~n1658;
  assign n1660 = ~n1657 & n1659;
  assign n1661 = n1657 & ~n1659;
  assign n1662 = ~n1660 & ~n1661;
  assign n1663 = n1607 & n1610;
  assign n1664 = ~n1611 & ~n1663;
  assign n1665 = n1662 & n1664;
  assign n1666 = ~n1660 & ~n1665;
  assign n1667 = n1619 & ~n1621;
  assign n1668 = ~n1622 & ~n1667;
  assign n1669 = ~n1666 & n1668;
  assign n1670 = ~n677 & n1550;
  assign n1671 = n677 & n1549;
  assign n1672 = n669 & ~n1130;
  assign n1673 = n1487 & ~n1672;
  assign n1674 = ~n1671 & ~n1673;
  assign n1675 = ~n1670 & n1674;
  assign n1676 = ~n286 & n844;
  assign n1677 = n286 & ~n665;
  assign n1678 = ~n847 & ~n1677;
  assign n1679 = ~n1676 & n1678;
  assign n1680 = n665 & n1679;
  assign n1681 = n1675 & n1680;
  assign n1682 = ~n832 & n1241;
  assign n1683 = n832 & n1199;
  assign n1684 = n1021 & n1244;
  assign n1685 = ~n1021 & n1197;
  assign n1686 = ~n1684 & ~n1685;
  assign n1687 = ~n1683 & n1686;
  assign n1688 = ~n1682 & n1687;
  assign n1689 = ~n1013 & n1033;
  assign n1690 = n868 & n1013;
  assign n1691 = n1036 & n1183;
  assign n1692 = n866 & ~n1183;
  assign n1693 = ~n1691 & ~n1692;
  assign n1694 = ~n1690 & n1693;
  assign n1695 = ~n1689 & n1694;
  assign n1696 = n1688 & ~n1695;
  assign n1697 = ~n1688 & n1695;
  assign n1698 = ~n1696 & ~n1697;
  assign n1699 = n1681 & ~n1698;
  assign n1700 = n1688 & n1695;
  assign n1701 = ~n1699 & ~n1700;
  assign n1702 = ~n275 & n844;
  assign n1703 = n275 & n700;
  assign n1704 = n279 & n847;
  assign n1705 = ~n279 & n698;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = ~n1703 & n1706;
  assign n1708 = ~n1702 & n1707;
  assign n1709 = ~n529 & n1550;
  assign n1710 = n529 & n1549;
  assign n1711 = n677 & ~n1130;
  assign n1712 = n1487 & ~n1711;
  assign n1713 = ~n1710 & ~n1712;
  assign n1714 = ~n1709 & n1713;
  assign n1715 = ~n669 & n1368;
  assign n1716 = n669 & n1317;
  assign n1717 = n840 & n1371;
  assign n1718 = ~n840 & n1315;
  assign n1719 = ~n1717 & ~n1718;
  assign n1720 = ~n1716 & n1719;
  assign n1721 = ~n1715 & n1720;
  assign n1722 = n1714 & ~n1721;
  assign n1723 = ~n1714 & n1721;
  assign n1724 = ~n1722 & ~n1723;
  assign n1725 = n1708 & ~n1724;
  assign n1726 = n1714 & n1721;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = ~n1701 & ~n1727;
  assign n1729 = ~n1701 & ~n1728;
  assign n1730 = ~n1727 & ~n1728;
  assign n1731 = ~n1729 & ~n1730;
  assign n1732 = n1577 & ~n1595;
  assign n1733 = ~n1594 & ~n1595;
  assign n1734 = ~n1732 & ~n1733;
  assign n1735 = ~n1731 & ~n1734;
  assign n1736 = ~n1728 & ~n1735;
  assign n1737 = n1597 & ~n1599;
  assign n1738 = ~n1600 & ~n1737;
  assign n1739 = ~n1736 & n1738;
  assign n1740 = n1652 & ~n1656;
  assign n1741 = ~n1655 & ~n1656;
  assign n1742 = ~n1740 & ~n1741;
  assign n1743 = n1736 & ~n1738;
  assign n1744 = ~n1739 & ~n1743;
  assign n1745 = ~n1742 & n1744;
  assign n1746 = ~n1739 & ~n1745;
  assign n1747 = ~n1662 & ~n1664;
  assign n1748 = ~n1665 & ~n1747;
  assign n1749 = ~n1746 & n1748;
  assign n1750 = ~n544 & ~n1560;
  assign n1751 = ~n1021 & n1241;
  assign n1752 = n1021 & n1199;
  assign n1753 = n1013 & n1244;
  assign n1754 = ~n1013 & n1197;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = ~n1752 & n1755;
  assign n1757 = ~n1751 & n1756;
  assign n1758 = ~n840 & n1368;
  assign n1759 = n840 & n1317;
  assign n1760 = n832 & n1371;
  assign n1761 = ~n832 & n1315;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = ~n1759 & n1762;
  assign n1764 = ~n1758 & n1763;
  assign n1765 = n1033 & ~n1183;
  assign n1766 = n868 & n1183;
  assign n1767 = n275 & n1036;
  assign n1768 = ~n275 & n866;
  assign n1769 = ~n1767 & ~n1768;
  assign n1770 = ~n1766 & n1769;
  assign n1771 = ~n1765 & n1770;
  assign n1772 = n1764 & ~n1771;
  assign n1773 = ~n1764 & n1771;
  assign n1774 = ~n1772 & ~n1773;
  assign n1775 = n1757 & ~n1774;
  assign n1776 = n1764 & n1771;
  assign n1777 = ~n1775 & ~n1776;
  assign n1778 = ~n1561 & ~n1777;
  assign n1779 = ~n1750 & n1778;
  assign n1780 = ~n1561 & ~n1779;
  assign n1781 = ~n1750 & n1780;
  assign n1782 = ~n1777 & ~n1779;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = ~n1681 & n1698;
  assign n1785 = ~n1699 & ~n1784;
  assign n1786 = ~n1783 & n1785;
  assign n1787 = ~n1779 & ~n1786;
  assign n1788 = n1643 & ~n1646;
  assign n1789 = ~n1644 & n1647;
  assign n1790 = ~n1788 & ~n1789;
  assign n1791 = ~n1787 & n1790;
  assign n1792 = n1787 & ~n1790;
  assign n1793 = ~n1791 & ~n1792;
  assign n1794 = ~n1731 & ~n1735;
  assign n1795 = ~n1734 & ~n1735;
  assign n1796 = ~n1794 & ~n1795;
  assign n1797 = ~n1793 & ~n1796;
  assign n1798 = ~n1787 & ~n1790;
  assign n1799 = ~n1797 & ~n1798;
  assign n1800 = n1742 & ~n1744;
  assign n1801 = ~n1745 & ~n1800;
  assign n1802 = ~n1799 & n1801;
  assign n1803 = ~n669 & n1550;
  assign n1804 = n669 & n1549;
  assign n1805 = n840 & ~n1130;
  assign n1806 = n1487 & ~n1805;
  assign n1807 = ~n1804 & ~n1806;
  assign n1808 = ~n1803 & n1807;
  assign n1809 = ~n832 & n1368;
  assign n1810 = n832 & n1317;
  assign n1811 = n1021 & n1371;
  assign n1812 = ~n1021 & n1315;
  assign n1813 = ~n1811 & ~n1812;
  assign n1814 = ~n1810 & n1813;
  assign n1815 = ~n1809 & n1814;
  assign n1816 = n1808 & n1815;
  assign n1817 = ~n1013 & n1241;
  assign n1818 = n1013 & n1199;
  assign n1819 = n1183 & n1244;
  assign n1820 = ~n1183 & n1197;
  assign n1821 = ~n1819 & ~n1820;
  assign n1822 = ~n1818 & n1821;
  assign n1823 = ~n1817 & n1822;
  assign n1824 = n1808 & ~n1815;
  assign n1825 = ~n1808 & n1815;
  assign n1826 = ~n1824 & ~n1825;
  assign n1827 = n1823 & ~n1826;
  assign n1828 = ~n1816 & ~n1827;
  assign n1829 = ~n279 & n844;
  assign n1830 = n279 & n700;
  assign n1831 = n286 & n847;
  assign n1832 = ~n286 & n698;
  assign n1833 = ~n1831 & ~n1832;
  assign n1834 = ~n1830 & n1833;
  assign n1835 = ~n1829 & n1834;
  assign n1836 = ~n1675 & ~n1680;
  assign n1837 = ~n1681 & ~n1836;
  assign n1838 = n1835 & ~n1837;
  assign n1839 = ~n1835 & n1837;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = ~n1828 & ~n1840;
  assign n1842 = n1835 & n1837;
  assign n1843 = ~n1841 & ~n1842;
  assign n1844 = n1708 & ~n1725;
  assign n1845 = ~n1724 & ~n1725;
  assign n1846 = ~n1844 & ~n1845;
  assign n1847 = ~n1843 & ~n1846;
  assign n1848 = ~n1783 & ~n1786;
  assign n1849 = n1785 & ~n1786;
  assign n1850 = ~n1848 & ~n1849;
  assign n1851 = ~n1843 & ~n1847;
  assign n1852 = ~n1846 & ~n1847;
  assign n1853 = ~n1851 & ~n1852;
  assign n1854 = ~n1850 & ~n1853;
  assign n1855 = ~n1847 & ~n1854;
  assign n1856 = ~n275 & n1033;
  assign n1857 = n275 & n868;
  assign n1858 = n279 & n1036;
  assign n1859 = ~n279 & n866;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = ~n1857 & n1860;
  assign n1862 = ~n1856 & n1861;
  assign n1863 = ~n840 & n1550;
  assign n1864 = n840 & n1549;
  assign n1865 = n832 & ~n1130;
  assign n1866 = n1487 & ~n1865;
  assign n1867 = ~n1864 & ~n1866;
  assign n1868 = ~n1863 & n1867;
  assign n1869 = ~n286 & n1033;
  assign n1870 = n286 & ~n828;
  assign n1871 = ~n1036 & ~n1870;
  assign n1872 = ~n1869 & n1871;
  assign n1873 = n828 & n1872;
  assign n1874 = n1868 & n1873;
  assign n1875 = n1862 & n1874;
  assign n1876 = ~n1862 & n1874;
  assign n1877 = n1862 & ~n1874;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = ~n286 & ~n695;
  assign n1880 = ~n1878 & n1879;
  assign n1881 = ~n1875 & ~n1880;
  assign n1882 = ~n1757 & n1774;
  assign n1883 = ~n1775 & ~n1882;
  assign n1884 = ~n1881 & n1883;
  assign n1885 = n1881 & ~n1883;
  assign n1886 = ~n1884 & ~n1885;
  assign n1887 = n1828 & n1840;
  assign n1888 = ~n1841 & ~n1887;
  assign n1889 = ~n1886 & ~n1888;
  assign n1890 = n1886 & n1888;
  assign n1891 = ~n279 & n1033;
  assign n1892 = n279 & n868;
  assign n1893 = n286 & n1036;
  assign n1894 = ~n286 & n866;
  assign n1895 = ~n1893 & ~n1894;
  assign n1896 = ~n1892 & n1895;
  assign n1897 = ~n1891 & n1896;
  assign n1898 = ~n1021 & n1368;
  assign n1899 = n1021 & n1317;
  assign n1900 = n1013 & n1371;
  assign n1901 = ~n1013 & n1315;
  assign n1902 = ~n1900 & ~n1901;
  assign n1903 = ~n1899 & n1902;
  assign n1904 = ~n1898 & n1903;
  assign n1905 = ~n1183 & n1241;
  assign n1906 = n1183 & n1199;
  assign n1907 = n275 & n1244;
  assign n1908 = ~n275 & n1197;
  assign n1909 = ~n1907 & ~n1908;
  assign n1910 = ~n1906 & n1909;
  assign n1911 = ~n1905 & n1910;
  assign n1912 = n1904 & ~n1911;
  assign n1913 = ~n1904 & n1911;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = n1897 & ~n1914;
  assign n1916 = n1904 & n1911;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = ~n1823 & n1826;
  assign n1919 = ~n1827 & ~n1918;
  assign n1920 = ~n1917 & n1919;
  assign n1921 = n1878 & ~n1879;
  assign n1922 = ~n1880 & ~n1921;
  assign n1923 = ~n1917 & ~n1920;
  assign n1924 = n1919 & ~n1920;
  assign n1925 = ~n1923 & ~n1924;
  assign n1926 = n1922 & ~n1925;
  assign n1927 = ~n1920 & ~n1926;
  assign n1928 = ~n828 & ~n1872;
  assign n1929 = ~n1021 & n1550;
  assign n1930 = n1021 & n1549;
  assign n1931 = n1013 & ~n1130;
  assign n1932 = n1487 & ~n1931;
  assign n1933 = ~n1930 & ~n1932;
  assign n1934 = ~n1929 & n1933;
  assign n1935 = ~n286 & n1241;
  assign n1936 = n286 & ~n1009;
  assign n1937 = ~n1244 & ~n1936;
  assign n1938 = ~n1935 & n1937;
  assign n1939 = n1009 & n1938;
  assign n1940 = n1934 & n1939;
  assign n1941 = ~n1873 & n1940;
  assign n1942 = ~n1928 & n1941;
  assign n1943 = ~n1183 & n1368;
  assign n1944 = n1183 & n1317;
  assign n1945 = n275 & n1371;
  assign n1946 = ~n275 & n1315;
  assign n1947 = ~n1945 & ~n1946;
  assign n1948 = ~n1944 & n1947;
  assign n1949 = ~n1943 & n1948;
  assign n1950 = ~n279 & n1241;
  assign n1951 = n279 & n1199;
  assign n1952 = n286 & n1244;
  assign n1953 = ~n286 & n1197;
  assign n1954 = ~n1952 & ~n1953;
  assign n1955 = ~n1951 & n1954;
  assign n1956 = ~n1950 & n1955;
  assign n1957 = n1949 & n1956;
  assign n1958 = ~n1934 & ~n1939;
  assign n1959 = ~n1940 & ~n1958;
  assign n1960 = ~n1949 & ~n1956;
  assign n1961 = ~n1957 & ~n1960;
  assign n1962 = n1959 & n1961;
  assign n1963 = ~n1957 & ~n1962;
  assign n1964 = n1940 & ~n1942;
  assign n1965 = ~n1873 & ~n1942;
  assign n1966 = ~n1928 & n1965;
  assign n1967 = ~n1964 & ~n1966;
  assign n1968 = ~n1963 & ~n1967;
  assign n1969 = ~n1942 & ~n1968;
  assign n1970 = ~n275 & n1241;
  assign n1971 = n275 & n1199;
  assign n1972 = n279 & n1244;
  assign n1973 = ~n279 & n1197;
  assign n1974 = ~n1972 & ~n1973;
  assign n1975 = ~n1971 & n1974;
  assign n1976 = ~n1970 & n1975;
  assign n1977 = ~n1013 & n1368;
  assign n1978 = n1013 & n1317;
  assign n1979 = n1183 & n1371;
  assign n1980 = ~n1183 & n1315;
  assign n1981 = ~n1979 & ~n1980;
  assign n1982 = ~n1978 & n1981;
  assign n1983 = ~n1977 & n1982;
  assign n1984 = ~n832 & n1550;
  assign n1985 = n832 & n1549;
  assign n1986 = n1021 & ~n1130;
  assign n1987 = n1487 & ~n1986;
  assign n1988 = ~n1985 & ~n1987;
  assign n1989 = ~n1984 & n1988;
  assign n1990 = ~n1983 & n1989;
  assign n1991 = n1983 & ~n1989;
  assign n1992 = ~n1990 & ~n1991;
  assign n1993 = ~n1976 & n1992;
  assign n1994 = n1976 & ~n1992;
  assign n1995 = ~n1013 & n1550;
  assign n1996 = n1013 & n1549;
  assign n1997 = ~n1130 & n1183;
  assign n1998 = n1487 & ~n1997;
  assign n1999 = ~n1996 & ~n1998;
  assign n2000 = ~n1995 & n1999;
  assign n2001 = ~n275 & n1368;
  assign n2002 = n275 & n1317;
  assign n2003 = n279 & n1371;
  assign n2004 = ~n279 & n1315;
  assign n2005 = ~n2003 & ~n2004;
  assign n2006 = ~n2002 & n2005;
  assign n2007 = ~n2001 & n2006;
  assign n2008 = n2000 & ~n2007;
  assign n2009 = ~n2000 & n2007;
  assign n2010 = ~n2008 & ~n2009;
  assign n2011 = ~n1183 & n1550;
  assign n2012 = n1183 & n1549;
  assign n2013 = n275 & ~n1130;
  assign n2014 = n1487 & ~n2013;
  assign n2015 = ~n2012 & ~n2014;
  assign n2016 = ~n2011 & n2015;
  assign n2017 = ~n286 & n1368;
  assign n2018 = n286 & ~n1177;
  assign n2019 = ~n1371 & ~n2018;
  assign n2020 = ~n2017 & n2019;
  assign n2021 = n1177 & n2020;
  assign n2022 = n2016 & n2021;
  assign n2023 = n2010 & ~n2022;
  assign n2024 = ~n2010 & n2022;
  assign n2025 = ~n279 & n1368;
  assign n2026 = n279 & n1317;
  assign n2027 = ~n286 & n1315;
  assign n2028 = ~n1177 & ~n2020;
  assign n2029 = ~n275 & n1550;
  assign n2030 = n275 & n1549;
  assign n2031 = ~n279 & ~n1487;
  assign n2032 = n1130 & n1487;
  assign n2033 = n279 & ~n2032;
  assign n2034 = ~n2031 & ~n2033;
  assign n2035 = ~n2030 & ~n2034;
  assign n2036 = ~n2029 & n2035;
  assign n2037 = n286 & ~n1130;
  assign n2038 = ~n2031 & n2037;
  assign n2039 = ~n2036 & ~n2038;
  assign n2040 = ~n2021 & ~n2039;
  assign n2041 = ~n2028 & n2040;
  assign n2042 = n2036 & n2038;
  assign n2043 = ~n2041 & ~n2042;
  assign n2044 = ~n2016 & ~n2021;
  assign n2045 = ~n2022 & ~n2044;
  assign n2046 = n2043 & ~n2045;
  assign n2047 = n286 & n1371;
  assign n2048 = ~n2046 & ~n2047;
  assign n2049 = ~n2027 & n2048;
  assign n2050 = ~n2026 & n2049;
  assign n2051 = ~n2025 & n2050;
  assign n2052 = ~n2043 & n2045;
  assign n2053 = ~n2051 & ~n2052;
  assign n2054 = ~n286 & ~n1194;
  assign n2055 = n2053 & ~n2054;
  assign n2056 = ~n2024 & ~n2055;
  assign n2057 = ~n2023 & n2056;
  assign n2058 = ~n2053 & n2054;
  assign n2059 = ~n2057 & ~n2058;
  assign n2060 = n1959 & ~n1962;
  assign n2061 = ~n1960 & n1963;
  assign n2062 = ~n2060 & ~n2061;
  assign n2063 = n2059 & n2062;
  assign n2064 = n2000 & n2007;
  assign n2065 = ~n2024 & ~n2064;
  assign n2066 = ~n2063 & ~n2065;
  assign n2067 = ~n2059 & ~n2062;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = ~n1963 & ~n1968;
  assign n2070 = ~n1967 & ~n1968;
  assign n2071 = ~n2069 & ~n2070;
  assign n2072 = n2068 & n2071;
  assign n2073 = ~n1994 & ~n2072;
  assign n2074 = ~n1993 & n2073;
  assign n2075 = ~n2068 & ~n2071;
  assign n2076 = ~n2074 & ~n2075;
  assign n2077 = ~n1969 & ~n2076;
  assign n2078 = n1969 & n2076;
  assign n2079 = n1897 & ~n1915;
  assign n2080 = ~n1914 & ~n1915;
  assign n2081 = ~n2079 & ~n2080;
  assign n2082 = ~n1868 & ~n1873;
  assign n2083 = ~n1874 & ~n2082;
  assign n2084 = n1983 & n1989;
  assign n2085 = ~n1994 & ~n2084;
  assign n2086 = n2083 & ~n2085;
  assign n2087 = ~n2083 & n2085;
  assign n2088 = ~n2086 & ~n2087;
  assign n2089 = ~n2081 & n2088;
  assign n2090 = n2081 & ~n2088;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = ~n2078 & n2091;
  assign n2093 = ~n2077 & ~n2092;
  assign n2094 = ~n2086 & ~n2089;
  assign n2095 = ~n2093 & ~n2094;
  assign n2096 = n2093 & n2094;
  assign n2097 = ~n1922 & n1925;
  assign n2098 = ~n1926 & ~n2097;
  assign n2099 = ~n2096 & n2098;
  assign n2100 = ~n2095 & ~n2099;
  assign n2101 = n1927 & n2100;
  assign n2102 = ~n1890 & ~n2101;
  assign n2103 = ~n1889 & n2102;
  assign n2104 = ~n1927 & ~n2100;
  assign n2105 = ~n2103 & ~n2104;
  assign n2106 = ~n1884 & ~n1890;
  assign n2107 = ~n2105 & ~n2106;
  assign n2108 = n2105 & n2106;
  assign n2109 = n1850 & n1853;
  assign n2110 = ~n1854 & ~n2109;
  assign n2111 = ~n2108 & n2110;
  assign n2112 = ~n2107 & ~n2111;
  assign n2113 = n1855 & n2112;
  assign n2114 = n1793 & n1796;
  assign n2115 = ~n2113 & ~n2114;
  assign n2116 = ~n1797 & n2115;
  assign n2117 = ~n1855 & ~n2112;
  assign n2118 = ~n2116 & ~n2117;
  assign n2119 = n1799 & ~n1801;
  assign n2120 = ~n1802 & ~n2119;
  assign n2121 = ~n2118 & n2120;
  assign n2122 = ~n1802 & ~n2121;
  assign n2123 = n1746 & ~n1748;
  assign n2124 = ~n1749 & ~n2123;
  assign n2125 = ~n2122 & n2124;
  assign n2126 = ~n1749 & ~n2125;
  assign n2127 = n1666 & ~n1668;
  assign n2128 = ~n1669 & ~n2127;
  assign n2129 = ~n2126 & n2128;
  assign n2130 = ~n1669 & ~n2129;
  assign n2131 = n1623 & ~n1625;
  assign n2132 = ~n1626 & ~n2131;
  assign n2133 = ~n2130 & n2132;
  assign n2134 = ~n1626 & ~n2133;
  assign n2135 = ~n1548 & ~n2134;
  assign n2136 = ~n1545 & ~n2135;
  assign n2137 = n1424 & n1427;
  assign n2138 = ~n1428 & ~n2137;
  assign n2139 = ~n2136 & n2138;
  assign n2140 = ~n1428 & ~n2139;
  assign n2141 = ~n1295 & ~n2140;
  assign n2142 = ~n1292 & ~n2141;
  assign n2143 = n1234 & ~n1236;
  assign n2144 = ~n1237 & ~n2143;
  assign n2145 = ~n2142 & n2144;
  assign n2146 = ~n1237 & ~n2145;
  assign n2147 = ~n1074 & ~n2146;
  assign n2148 = ~n1068 & ~n1071;
  assign n2149 = ~n2147 & ~n2148;
  assign n2150 = n895 & ~n897;
  assign n2151 = ~n898 & ~n2150;
  assign n2152 = ~n2149 & n2151;
  assign n2153 = ~n898 & ~n2152;
  assign n2154 = ~n728 & ~n2153;
  assign n2155 = ~n722 & ~n725;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = n683 & ~n2156;
  assign n2158 = ~n683 & n2156;
  assign n2159 = ~n2157 & ~n2158;
  assign n2160 = n536 & n2159;
  assign n2161 = ~n536 & ~n2159;
  assign n2162 = ~n2160 & ~n2161;
  assign n2163 = ~n393 & ~n2162;
  assign n2164 = n393 & n2162;
  assign n2165 = ~n134 & ~n468;
  assign n2166 = ~n219 & n2165;
  assign n2167 = ~n254 & ~n329;
  assign n2168 = ~n358 & n2167;
  assign n2169 = ~n326 & n2168;
  assign n2170 = ~n342 & n2169;
  assign n2171 = n760 & n2170;
  assign n2172 = ~n226 & n2171;
  assign n2173 = ~n218 & n2172;
  assign n2174 = ~n167 & n2173;
  assign n2175 = ~n206 & n2174;
  assign n2176 = ~n190 & n2175;
  assign n2177 = ~n589 & n2176;
  assign n2178 = ~n736 & n2177;
  assign n2179 = ~n415 & n626;
  assign n2180 = ~n297 & n2179;
  assign n2181 = ~n356 & n2180;
  assign n2182 = ~n361 & n968;
  assign n2183 = ~n142 & n2182;
  assign n2184 = n555 & n2183;
  assign n2185 = n476 & n2184;
  assign n2186 = n1091 & n2185;
  assign n2187 = n2181 & n2186;
  assign n2188 = n986 & n2187;
  assign n2189 = n753 & n2188;
  assign n2190 = ~n154 & n2189;
  assign n2191 = ~n140 & n792;
  assign n2192 = ~n299 & n2191;
  assign n2193 = ~n458 & n2192;
  assign n2194 = ~n357 & n2193;
  assign n2195 = ~n148 & n2194;
  assign n2196 = ~n553 & n2195;
  assign n2197 = n153 & n808;
  assign n2198 = n397 & n2197;
  assign n2199 = n773 & n2198;
  assign n2200 = n2196 & n2199;
  assign n2201 = n2190 & n2200;
  assign n2202 = n2178 & n2201;
  assign n2203 = n2166 & n2202;
  assign n2204 = ~n328 & n2203;
  assign n2205 = ~n228 & n2204;
  assign n2206 = ~n177 & n2205;
  assign n2207 = ~n504 & n2206;
  assign n2208 = ~n367 & n2207;
  assign n2209 = ~n215 & n2208;
  assign n2210 = n728 & n2153;
  assign n2211 = ~n2154 & ~n2210;
  assign n2212 = ~n2209 & ~n2211;
  assign n2213 = n145 & n794;
  assign n2214 = n319 & n2213;
  assign n2215 = n474 & n2214;
  assign n2216 = n637 & n2215;
  assign n2217 = n739 & n2216;
  assign n2218 = n967 & n2217;
  assign n2219 = n606 & n2218;
  assign n2220 = n1104 & n2219;
  assign n2221 = ~n458 & n2220;
  assign n2222 = ~n297 & n2221;
  assign n2223 = ~n358 & n2222;
  assign n2224 = ~n168 & n2223;
  assign n2225 = ~n237 & n2224;
  assign n2226 = n2149 & ~n2151;
  assign n2227 = ~n2152 & ~n2226;
  assign n2228 = ~n2225 & ~n2227;
  assign n2229 = n2225 & n2227;
  assign n2230 = n331 & n2183;
  assign n2231 = n236 & n2230;
  assign n2232 = n301 & n2231;
  assign n2233 = n637 & n2232;
  assign n2234 = n2166 & n2233;
  assign n2235 = n355 & n2234;
  assign n2236 = ~n221 & n2235;
  assign n2237 = ~n394 & n2236;
  assign n2238 = ~n225 & n2237;
  assign n2239 = ~n206 & n2238;
  assign n2240 = ~n254 & n906;
  assign n2241 = ~n447 & n2240;
  assign n2242 = ~n148 & n2241;
  assign n2243 = ~n111 & n2242;
  assign n2244 = ~n238 & n2243;
  assign n2245 = n581 & n628;
  assign n2246 = n2244 & n2245;
  assign n2247 = ~n227 & n2246;
  assign n2248 = ~n417 & n2247;
  assign n2249 = ~n123 & n2248;
  assign n2250 = ~n736 & n2249;
  assign n2251 = ~n178 & ~n506;
  assign n2252 = ~n471 & n2251;
  assign n2253 = ~n302 & ~n313;
  assign n2254 = ~n445 & n2253;
  assign n2255 = n478 & n2254;
  assign n2256 = n2252 & n2255;
  assign n2257 = n156 & n2256;
  assign n2258 = n577 & n2257;
  assign n2259 = n644 & n2258;
  assign n2260 = n2250 & n2259;
  assign n2261 = n2239 & n2260;
  assign n2262 = ~n317 & n2261;
  assign n2263 = ~n336 & n2262;
  assign n2264 = ~n554 & n2263;
  assign n2265 = n1074 & n2146;
  assign n2266 = ~n2147 & ~n2265;
  assign n2267 = ~n2264 & ~n2266;
  assign n2268 = n396 & n2252;
  assign n2269 = n451 & n2268;
  assign n2270 = ~n139 & n2269;
  assign n2271 = ~n188 & n2270;
  assign n2272 = ~n129 & n2271;
  assign n2273 = ~n359 & n2272;
  assign n2274 = ~n335 & n2273;
  assign n2275 = ~n367 & n2274;
  assign n2276 = ~n599 & n2275;
  assign n2277 = ~n447 & ~n552;
  assign n2278 = ~n237 & n2277;
  assign n2279 = ~n152 & n2239;
  assign n2280 = ~n296 & n2279;
  assign n2281 = ~n215 & n2280;
  assign n2282 = n1459 & n2281;
  assign n2283 = n2278 & n2282;
  assign n2284 = n325 & n2283;
  assign n2285 = n2196 & n2284;
  assign n2286 = n2276 & n2285;
  assign n2287 = n980 & n2286;
  assign n2288 = ~n176 & n2287;
  assign n2289 = ~n343 & n2288;
  assign n2290 = ~n167 & n2289;
  assign n2291 = ~n360 & n2290;
  assign n2292 = ~n313 & n2291;
  assign n2293 = n2142 & ~n2144;
  assign n2294 = ~n2145 & ~n2293;
  assign n2295 = ~n2292 & ~n2294;
  assign n2296 = n2292 & n2294;
  assign n2297 = ~n138 & ~n227;
  assign n2298 = ~n123 & n2297;
  assign n2299 = ~n172 & n2298;
  assign n2300 = ~n234 & n2299;
  assign n2301 = ~n357 & n2300;
  assign n2302 = ~n216 & n2301;
  assign n2303 = ~n168 & n2302;
  assign n2304 = n141 & n1116;
  assign n2305 = n944 & n2304;
  assign n2306 = n644 & n2305;
  assign n2307 = n369 & n2306;
  assign n2308 = ~n337 & n2307;
  assign n2309 = ~n458 & n2308;
  assign n2310 = ~n447 & n2309;
  assign n2311 = ~n347 & n2310;
  assign n2312 = ~n106 & n923;
  assign n2313 = ~n326 & n2312;
  assign n2314 = ~n217 & ~n228;
  assign n2315 = ~n146 & n2314;
  assign n2316 = ~n211 & n2315;
  assign n2317 = ~n469 & n2316;
  assign n2318 = n2313 & n2317;
  assign n2319 = n2311 & n2318;
  assign n2320 = n2303 & n2319;
  assign n2321 = ~n328 & n2320;
  assign n2322 = ~n408 & n2321;
  assign n2323 = ~n194 & n2322;
  assign n2324 = ~n219 & n2323;
  assign n2325 = ~n298 & n2324;
  assign n2326 = n450 & n2325;
  assign n2327 = ~n445 & n2326;
  assign n2328 = n1295 & n2140;
  assign n2329 = ~n2141 & ~n2328;
  assign n2330 = ~n2327 & ~n2329;
  assign n2331 = ~n213 & n508;
  assign n2332 = ~n736 & n2331;
  assign n2333 = ~n345 & n2332;
  assign n2334 = n303 & n759;
  assign n2335 = n931 & n2334;
  assign n2336 = ~n169 & n2335;
  assign n2337 = ~n114 & n2336;
  assign n2338 = ~n326 & n2337;
  assign n2339 = ~n469 & n2338;
  assign n2340 = ~n138 & ~n146;
  assign n2341 = ~n106 & ~n348;
  assign n2342 = ~n238 & n2341;
  assign n2343 = n432 & n2342;
  assign n2344 = n2340 & n2343;
  assign n2345 = n1106 & n2344;
  assign n2346 = n344 & n2345;
  assign n2347 = n314 & n2346;
  assign n2348 = n2339 & n2347;
  assign n2349 = n995 & n2348;
  assign n2350 = n930 & n2349;
  assign n2351 = n2333 & n2350;
  assign n2352 = ~n152 & n2351;
  assign n2353 = ~n217 & n2352;
  assign n2354 = ~n495 & n2353;
  assign n2355 = n2136 & ~n2138;
  assign n2356 = ~n2139 & ~n2355;
  assign n2357 = ~n2354 & ~n2356;
  assign n2358 = n2354 & n2356;
  assign n2359 = n141 & ~n312;
  assign n2360 = ~n417 & n2359;
  assign n2361 = ~n313 & n2360;
  assign n2362 = ~n224 & n2361;
  assign n2363 = ~n553 & n2362;
  assign n2364 = ~n235 & n2363;
  assign n2365 = ~n255 & ~n449;
  assign n2366 = ~n554 & n2365;
  assign n2367 = ~n194 & ~n237;
  assign n2368 = n2366 & n2367;
  assign n2369 = n910 & n2368;
  assign n2370 = ~n188 & n2369;
  assign n2371 = ~n327 & n2370;
  assign n2372 = ~n348 & n2371;
  assign n2373 = ~n329 & n2372;
  assign n2374 = ~n191 & n2373;
  assign n2375 = ~n503 & n2374;
  assign n2376 = n382 & n448;
  assign n2377 = n2375 & n2376;
  assign n2378 = n753 & n2377;
  assign n2379 = n2364 & n2378;
  assign n2380 = ~n196 & n2379;
  assign n2381 = ~n221 & n2380;
  assign n2382 = ~n394 & n2381;
  assign n2383 = ~n167 & n2382;
  assign n2384 = ~n347 & n2383;
  assign n2385 = ~n472 & n2384;
  assign n2386 = n1548 & n2134;
  assign n2387 = ~n2135 & ~n2386;
  assign n2388 = ~n2385 & ~n2387;
  assign n2389 = n564 & n2254;
  assign n2390 = n906 & n2389;
  assign n2391 = n411 & n2390;
  assign n2392 = ~n360 & n2391;
  assign n2393 = ~n114 & n2392;
  assign n2394 = ~n326 & n2393;
  assign n2395 = ~n223 & n2394;
  assign n2396 = n416 & n473;
  assign n2397 = ~n298 & n2396;
  assign n2398 = ~n118 & n2397;
  assign n2399 = ~n224 & n2398;
  assign n2400 = ~n367 & n2399;
  assign n2401 = n590 & n2400;
  assign n2402 = n2395 & n2401;
  assign n2403 = n752 & n2402;
  assign n2404 = n986 & n2403;
  assign n2405 = n149 & n2404;
  assign n2406 = ~n228 & n2405;
  assign n2407 = ~n219 & n2406;
  assign n2408 = ~n226 & n2407;
  assign n2409 = ~n336 & n2408;
  assign n2410 = ~n234 & n2409;
  assign n2411 = ~n258 & n2410;
  assign n2412 = ~n554 & n2411;
  assign n2413 = ~n342 & n2412;
  assign n2414 = ~n296 & n2413;
  assign n2415 = n2130 & ~n2132;
  assign n2416 = ~n2133 & ~n2415;
  assign n2417 = ~n2414 & ~n2416;
  assign n2418 = ~n553 & ~n599;
  assign n2419 = ~n335 & n2418;
  assign n2420 = ~n111 & n2419;
  assign n2421 = ~n477 & n2420;
  assign n2422 = ~n296 & ~n449;
  assign n2423 = n970 & n2422;
  assign n2424 = n2421 & n2423;
  assign n2425 = n2278 & n2424;
  assign n2426 = n373 & n2425;
  assign n2427 = n2333 & n2426;
  assign n2428 = n926 & n2427;
  assign n2429 = ~n359 & n2428;
  assign n2430 = ~n358 & n2429;
  assign n2431 = ~n472 & n2430;
  assign n2432 = ~n223 & n2431;
  assign n2433 = ~n351 & ~n504;
  assign n2434 = n396 & n806;
  assign n2435 = n2433 & n2434;
  assign n2436 = n2400 & n2435;
  assign n2437 = n325 & n2436;
  assign n2438 = n323 & n2437;
  assign n2439 = n983 & n2438;
  assign n2440 = n2432 & n2439;
  assign n2441 = n165 & n2440;
  assign n2442 = ~n328 & n2441;
  assign n2443 = ~n214 & n2442;
  assign n2444 = ~n257 & n2443;
  assign n2445 = ~n360 & n2444;
  assign n2446 = ~n238 & n2445;
  assign n2447 = n2126 & ~n2128;
  assign n2448 = ~n2129 & ~n2447;
  assign n2449 = ~n2446 & ~n2448;
  assign n2450 = n2446 & n2448;
  assign n2451 = ~n152 & n1117;
  assign n2452 = ~n227 & n2451;
  assign n2453 = ~n347 & n2452;
  assign n2454 = ~n554 & n2453;
  assign n2455 = ~n176 & ~n312;
  assign n2456 = ~n370 & n2455;
  assign n2457 = ~n361 & n2456;
  assign n2458 = ~n132 & n2457;
  assign n2459 = n2454 & n2458;
  assign n2460 = ~n343 & n2459;
  assign n2461 = ~n458 & n2460;
  assign n2462 = ~n359 & n2461;
  assign n2463 = ~n552 & n2462;
  assign n2464 = ~n154 & n2463;
  assign n2465 = n256 & n2422;
  assign n2466 = n474 & n2465;
  assign n2467 = n2339 & n2466;
  assign n2468 = n2464 & n2467;
  assign n2469 = n789 & n2468;
  assign n2470 = ~n337 & n2469;
  assign n2471 = ~n208 & n2470;
  assign n2472 = ~n134 & n2471;
  assign n2473 = ~n192 & n2472;
  assign n2474 = ~n123 & n2473;
  assign n2475 = ~n224 & n2474;
  assign n2476 = ~n357 & n2475;
  assign n2477 = ~n445 & n2476;
  assign n2478 = n2122 & ~n2124;
  assign n2479 = ~n2125 & ~n2478;
  assign n2480 = ~n2477 & ~n2479;
  assign n2481 = n2477 & n2479;
  assign n2482 = ~n2118 & ~n2121;
  assign n2483 = n2120 & ~n2121;
  assign n2484 = ~n2482 & ~n2483;
  assign n2485 = n777 & n1096;
  assign n2486 = n914 & n2485;
  assign n2487 = n373 & n2486;
  assign n2488 = n2395 & n2487;
  assign n2489 = n739 & n2488;
  assign n2490 = n2190 & n2489;
  assign n2491 = ~n417 & n2490;
  assign n2492 = ~n192 & n2491;
  assign n2493 = ~n358 & n2492;
  assign n2494 = ~n190 & n2493;
  assign n2495 = ~n599 & n2494;
  assign n2496 = ~n2484 & n2495;
  assign n2497 = ~n2480 & ~n2496;
  assign n2498 = ~n2481 & n2497;
  assign n2499 = ~n2480 & ~n2498;
  assign n2500 = ~n2449 & ~n2499;
  assign n2501 = ~n2450 & n2500;
  assign n2502 = ~n2449 & ~n2501;
  assign n2503 = n2414 & n2416;
  assign n2504 = ~n2417 & ~n2503;
  assign n2505 = ~n2502 & n2504;
  assign n2506 = ~n2417 & ~n2505;
  assign n2507 = n2385 & n2387;
  assign n2508 = ~n2388 & ~n2507;
  assign n2509 = ~n2506 & n2508;
  assign n2510 = ~n2388 & ~n2509;
  assign n2511 = ~n2357 & ~n2510;
  assign n2512 = ~n2358 & n2511;
  assign n2513 = ~n2357 & ~n2512;
  assign n2514 = ~n2327 & ~n2330;
  assign n2515 = ~n2329 & ~n2330;
  assign n2516 = ~n2514 & ~n2515;
  assign n2517 = ~n2513 & ~n2516;
  assign n2518 = ~n2330 & ~n2517;
  assign n2519 = ~n2295 & ~n2518;
  assign n2520 = ~n2296 & n2519;
  assign n2521 = ~n2295 & ~n2520;
  assign n2522 = n2264 & n2266;
  assign n2523 = ~n2267 & ~n2522;
  assign n2524 = ~n2521 & n2523;
  assign n2525 = ~n2267 & ~n2524;
  assign n2526 = ~n2228 & ~n2525;
  assign n2527 = ~n2229 & n2526;
  assign n2528 = ~n2228 & ~n2527;
  assign n2529 = n2209 & n2211;
  assign n2530 = ~n2212 & ~n2529;
  assign n2531 = ~n2528 & n2530;
  assign n2532 = ~n2212 & ~n2531;
  assign n2533 = ~n2163 & ~n2532;
  assign n2534 = ~n2164 & n2533;
  assign n2535 = ~n2163 & ~n2534;
  assign n2536 = ~n408 & n796;
  assign n2537 = ~n188 & n2536;
  assign n2538 = ~n227 & n2537;
  assign n2539 = ~n174 & n2538;
  assign n2540 = ~n368 & n2539;
  assign n2541 = n478 & n1091;
  assign n2542 = n2339 & n2541;
  assign n2543 = n1468 & n2542;
  assign n2544 = n2540 & n2543;
  assign n2545 = n653 & n2544;
  assign n2546 = n149 & n2545;
  assign n2547 = ~n299 & n2546;
  assign n2548 = n945 & n2547;
  assign n2549 = ~n552 & n2548;
  assign n2550 = ~n554 & n2549;
  assign n2551 = ~n223 & n2550;
  assign n2552 = n2535 & n2551;
  assign n2553 = ~n2535 & ~n2551;
  assign n2554 = ~n2552 & ~n2553;
  assign n2555 = n295 & ~n2554;
  assign n2556 = ~n279 & n286;
  assign n2557 = n279 & ~n286;
  assign n2558 = ~n2556 & ~n2557;
  assign n2559 = ~n282 & n294;
  assign n2560 = n2558 & n2559;
  assign n2561 = n2528 & ~n2530;
  assign n2562 = ~n2531 & ~n2561;
  assign n2563 = n2560 & n2562;
  assign n2564 = ~n2532 & ~n2534;
  assign n2565 = ~n2164 & n2535;
  assign n2566 = ~n2564 & ~n2565;
  assign n2567 = n294 & ~n2558;
  assign n2568 = ~n2566 & n2567;
  assign n2569 = ~n2563 & ~n2568;
  assign n2570 = ~n2555 & n2569;
  assign n2571 = ~n282 & ~n294;
  assign n2572 = n2562 & ~n2566;
  assign n2573 = ~n2525 & ~n2527;
  assign n2574 = ~n2229 & n2528;
  assign n2575 = ~n2573 & ~n2574;
  assign n2576 = n2562 & ~n2575;
  assign n2577 = n2521 & ~n2523;
  assign n2578 = ~n2524 & ~n2577;
  assign n2579 = ~n2575 & n2578;
  assign n2580 = ~n2518 & ~n2520;
  assign n2581 = ~n2296 & n2521;
  assign n2582 = ~n2580 & ~n2581;
  assign n2583 = n2578 & ~n2582;
  assign n2584 = ~n2513 & ~n2517;
  assign n2585 = ~n2516 & ~n2517;
  assign n2586 = ~n2584 & ~n2585;
  assign n2587 = ~n2582 & ~n2586;
  assign n2588 = ~n2510 & ~n2512;
  assign n2589 = ~n2358 & n2513;
  assign n2590 = ~n2588 & ~n2589;
  assign n2591 = ~n2586 & ~n2590;
  assign n2592 = n2506 & ~n2508;
  assign n2593 = ~n2509 & ~n2592;
  assign n2594 = ~n2590 & n2593;
  assign n2595 = n2502 & ~n2504;
  assign n2596 = ~n2505 & ~n2595;
  assign n2597 = n2593 & n2596;
  assign n2598 = ~n2499 & ~n2501;
  assign n2599 = ~n2450 & n2502;
  assign n2600 = ~n2598 & ~n2599;
  assign n2601 = n2596 & ~n2600;
  assign n2602 = ~n2496 & ~n2498;
  assign n2603 = ~n2481 & n2499;
  assign n2604 = ~n2602 & ~n2603;
  assign n2605 = ~n2600 & ~n2604;
  assign n2606 = n2484 & ~n2495;
  assign n2607 = ~n2496 & ~n2606;
  assign n2608 = ~n2604 & ~n2607;
  assign n2609 = n2600 & n2608;
  assign n2610 = ~n2605 & ~n2609;
  assign n2611 = ~n2596 & n2600;
  assign n2612 = ~n2610 & ~n2611;
  assign n2613 = ~n2601 & n2612;
  assign n2614 = ~n2601 & ~n2613;
  assign n2615 = ~n2593 & ~n2596;
  assign n2616 = ~n2614 & ~n2615;
  assign n2617 = ~n2597 & n2616;
  assign n2618 = ~n2597 & ~n2617;
  assign n2619 = n2590 & ~n2593;
  assign n2620 = ~n2594 & ~n2619;
  assign n2621 = ~n2618 & n2620;
  assign n2622 = ~n2594 & ~n2621;
  assign n2623 = n2586 & n2590;
  assign n2624 = ~n2591 & ~n2623;
  assign n2625 = ~n2622 & n2624;
  assign n2626 = ~n2591 & ~n2625;
  assign n2627 = n2582 & n2586;
  assign n2628 = ~n2587 & ~n2627;
  assign n2629 = ~n2626 & n2628;
  assign n2630 = ~n2587 & ~n2629;
  assign n2631 = ~n2578 & n2582;
  assign n2632 = ~n2583 & ~n2631;
  assign n2633 = ~n2630 & n2632;
  assign n2634 = ~n2583 & ~n2633;
  assign n2635 = n2575 & ~n2578;
  assign n2636 = ~n2579 & ~n2635;
  assign n2637 = ~n2634 & n2636;
  assign n2638 = ~n2579 & ~n2637;
  assign n2639 = ~n2562 & n2575;
  assign n2640 = ~n2576 & ~n2639;
  assign n2641 = ~n2638 & n2640;
  assign n2642 = ~n2576 & ~n2641;
  assign n2643 = ~n2562 & n2566;
  assign n2644 = ~n2572 & ~n2643;
  assign n2645 = ~n2642 & n2644;
  assign n2646 = ~n2572 & ~n2645;
  assign n2647 = ~n2554 & ~n2566;
  assign n2648 = n2554 & n2566;
  assign n2649 = ~n2647 & ~n2648;
  assign n2650 = ~n2646 & n2649;
  assign n2651 = n2646 & ~n2649;
  assign n2652 = ~n2650 & ~n2651;
  assign n2653 = n2571 & n2652;
  assign n2654 = n2570 & ~n2653;
  assign n2655 = ~n275 & ~n2654;
  assign n2656 = n275 & n2654;
  assign n2657 = ~n2655 & ~n2656;
  assign n2658 = n669 & ~n677;
  assign n2659 = ~n669 & n677;
  assign n2660 = ~n2658 & ~n2659;
  assign n2661 = ~n2607 & ~n2660;
  assign n2662 = ~n525 & ~n2661;
  assign n2663 = n529 & ~n677;
  assign n2664 = ~n529 & n677;
  assign n2665 = ~n2663 & ~n2664;
  assign n2666 = n2660 & ~n2665;
  assign n2667 = ~n2607 & n2666;
  assign n2668 = n532 & ~n2660;
  assign n2669 = ~n2604 & n2668;
  assign n2670 = ~n2667 & ~n2669;
  assign n2671 = n2604 & ~n2607;
  assign n2672 = ~n2604 & n2607;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = ~n532 & ~n2660;
  assign n2675 = ~n2673 & n2674;
  assign n2676 = n2670 & ~n2675;
  assign n2677 = ~n525 & ~n2676;
  assign n2678 = ~n525 & ~n2677;
  assign n2679 = ~n2676 & ~n2677;
  assign n2680 = ~n2678 & ~n2679;
  assign n2681 = n2662 & ~n2680;
  assign n2682 = ~n2662 & n2680;
  assign n2683 = ~n2681 & ~n2682;
  assign n2684 = n832 & ~n1021;
  assign n2685 = ~n832 & n1021;
  assign n2686 = ~n2684 & ~n2685;
  assign n2687 = n669 & ~n840;
  assign n2688 = ~n669 & n840;
  assign n2689 = ~n2687 & ~n2688;
  assign n2690 = ~n2686 & ~n2689;
  assign n2691 = n832 & ~n840;
  assign n2692 = ~n832 & n840;
  assign n2693 = ~n2691 & ~n2692;
  assign n2694 = n2686 & ~n2689;
  assign n2695 = n2693 & n2694;
  assign n2696 = ~n2600 & n2695;
  assign n2697 = n2686 & ~n2693;
  assign n2698 = n2596 & n2697;
  assign n2699 = ~n2686 & n2689;
  assign n2700 = n2593 & n2699;
  assign n2701 = ~n2698 & ~n2700;
  assign n2702 = ~n2696 & n2701;
  assign n2703 = ~n2690 & n2702;
  assign n2704 = ~n2614 & ~n2617;
  assign n2705 = ~n2615 & n2618;
  assign n2706 = ~n2704 & ~n2705;
  assign n2707 = n2702 & n2706;
  assign n2708 = ~n2703 & ~n2707;
  assign n2709 = n669 & ~n2708;
  assign n2710 = ~n669 & n2708;
  assign n2711 = ~n2709 & ~n2710;
  assign n2712 = n2683 & n2711;
  assign n2713 = ~n2607 & ~n2686;
  assign n2714 = ~n669 & ~n2713;
  assign n2715 = ~n2607 & n2697;
  assign n2716 = ~n2604 & n2699;
  assign n2717 = ~n2715 & ~n2716;
  assign n2718 = ~n2673 & n2690;
  assign n2719 = n2717 & ~n2718;
  assign n2720 = ~n669 & ~n2719;
  assign n2721 = n669 & n2719;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = n2714 & n2722;
  assign n2724 = ~n2600 & n2699;
  assign n2725 = ~n2607 & n2695;
  assign n2726 = ~n2604 & n2697;
  assign n2727 = ~n2725 & ~n2726;
  assign n2728 = ~n2724 & n2727;
  assign n2729 = ~n2690 & n2728;
  assign n2730 = n2600 & ~n2672;
  assign n2731 = ~n2600 & n2672;
  assign n2732 = ~n2730 & ~n2731;
  assign n2733 = n2728 & ~n2732;
  assign n2734 = ~n2729 & ~n2733;
  assign n2735 = n669 & ~n2734;
  assign n2736 = ~n669 & n2734;
  assign n2737 = ~n2735 & ~n2736;
  assign n2738 = n2723 & n2737;
  assign n2739 = n2661 & n2738;
  assign n2740 = n2738 & ~n2739;
  assign n2741 = n2661 & ~n2739;
  assign n2742 = ~n2740 & ~n2741;
  assign n2743 = ~n2600 & n2697;
  assign n2744 = n2596 & n2699;
  assign n2745 = ~n2604 & n2695;
  assign n2746 = ~n2744 & ~n2745;
  assign n2747 = ~n2743 & n2746;
  assign n2748 = ~n2610 & ~n2613;
  assign n2749 = ~n2611 & n2614;
  assign n2750 = ~n2748 & ~n2749;
  assign n2751 = n2690 & ~n2750;
  assign n2752 = n2747 & ~n2751;
  assign n2753 = ~n669 & ~n2752;
  assign n2754 = n669 & n2752;
  assign n2755 = ~n2753 & ~n2754;
  assign n2756 = ~n2742 & n2755;
  assign n2757 = ~n2739 & ~n2756;
  assign n2758 = ~n2683 & ~n2711;
  assign n2759 = ~n2712 & ~n2758;
  assign n2760 = ~n2757 & n2759;
  assign n2761 = ~n2712 & ~n2760;
  assign n2762 = ~n2590 & n2699;
  assign n2763 = n2596 & n2695;
  assign n2764 = n2593 & n2697;
  assign n2765 = ~n2763 & ~n2764;
  assign n2766 = ~n2762 & n2765;
  assign n2767 = n2618 & ~n2620;
  assign n2768 = ~n2621 & ~n2767;
  assign n2769 = n2690 & n2768;
  assign n2770 = n2766 & ~n2769;
  assign n2771 = ~n669 & ~n2770;
  assign n2772 = n669 & n2770;
  assign n2773 = ~n2771 & ~n2772;
  assign n2774 = ~n2600 & n2668;
  assign n2775 = ~n532 & n2660;
  assign n2776 = n2665 & n2775;
  assign n2777 = ~n2607 & n2776;
  assign n2778 = ~n2604 & n2666;
  assign n2779 = ~n2777 & ~n2778;
  assign n2780 = ~n2774 & n2779;
  assign n2781 = ~n2674 & n2780;
  assign n2782 = ~n2732 & n2780;
  assign n2783 = ~n2781 & ~n2782;
  assign n2784 = n525 & ~n2783;
  assign n2785 = ~n525 & n2783;
  assign n2786 = ~n2784 & ~n2785;
  assign n2787 = n2681 & n2786;
  assign n2788 = ~n2681 & ~n2786;
  assign n2789 = ~n2787 & ~n2788;
  assign n2790 = n2773 & n2789;
  assign n2791 = ~n2773 & ~n2789;
  assign n2792 = ~n2790 & ~n2791;
  assign n2793 = n2761 & ~n2792;
  assign n2794 = ~n2761 & n2792;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = n1013 & ~n1021;
  assign n2797 = ~n1013 & n1021;
  assign n2798 = ~n2796 & ~n2797;
  assign n2799 = n275 & ~n1183;
  assign n2800 = ~n275 & n1183;
  assign n2801 = ~n2799 & ~n2800;
  assign n2802 = n2798 & ~n2801;
  assign n2803 = n2578 & n2802;
  assign n2804 = n1013 & ~n1183;
  assign n2805 = ~n1013 & n1183;
  assign n2806 = ~n2804 & ~n2805;
  assign n2807 = ~n2798 & n2801;
  assign n2808 = n2806 & n2807;
  assign n2809 = ~n2586 & n2808;
  assign n2810 = n2801 & ~n2806;
  assign n2811 = ~n2582 & n2810;
  assign n2812 = ~n2809 & ~n2811;
  assign n2813 = ~n2803 & n2812;
  assign n2814 = n2630 & ~n2632;
  assign n2815 = ~n2633 & ~n2814;
  assign n2816 = n2813 & ~n2815;
  assign n2817 = ~n2798 & ~n2801;
  assign n2818 = n2813 & ~n2817;
  assign n2819 = ~n2816 & ~n2818;
  assign n2820 = n1021 & ~n2819;
  assign n2821 = ~n1021 & n2819;
  assign n2822 = ~n2820 & ~n2821;
  assign n2823 = n2795 & n2822;
  assign n2824 = ~n2582 & n2802;
  assign n2825 = ~n2590 & n2808;
  assign n2826 = ~n2586 & n2810;
  assign n2827 = ~n2825 & ~n2826;
  assign n2828 = ~n2824 & n2827;
  assign n2829 = n2626 & ~n2628;
  assign n2830 = ~n2629 & ~n2829;
  assign n2831 = n2817 & n2830;
  assign n2832 = n2828 & ~n2831;
  assign n2833 = ~n1021 & ~n2832;
  assign n2834 = ~n2832 & ~n2833;
  assign n2835 = ~n1021 & ~n2833;
  assign n2836 = ~n2834 & ~n2835;
  assign n2837 = n2757 & ~n2759;
  assign n2838 = ~n2760 & ~n2837;
  assign n2839 = ~n2836 & n2838;
  assign n2840 = ~n2742 & ~n2756;
  assign n2841 = n2755 & ~n2756;
  assign n2842 = ~n2840 & ~n2841;
  assign n2843 = ~n2586 & n2802;
  assign n2844 = n2593 & n2808;
  assign n2845 = ~n2590 & n2810;
  assign n2846 = ~n2844 & ~n2845;
  assign n2847 = ~n2843 & n2846;
  assign n2848 = n2622 & ~n2624;
  assign n2849 = ~n2625 & ~n2848;
  assign n2850 = n2847 & ~n2849;
  assign n2851 = ~n2817 & n2847;
  assign n2852 = ~n2850 & ~n2851;
  assign n2853 = n1021 & ~n2852;
  assign n2854 = ~n1021 & n2852;
  assign n2855 = ~n2853 & ~n2854;
  assign n2856 = ~n2842 & n2855;
  assign n2857 = ~n2590 & n2802;
  assign n2858 = n2596 & n2808;
  assign n2859 = n2593 & n2810;
  assign n2860 = ~n2858 & ~n2859;
  assign n2861 = ~n2857 & n2860;
  assign n2862 = n2768 & n2817;
  assign n2863 = n2861 & ~n2862;
  assign n2864 = ~n1021 & ~n2863;
  assign n2865 = ~n2863 & ~n2864;
  assign n2866 = ~n1021 & ~n2864;
  assign n2867 = ~n2865 & ~n2866;
  assign n2868 = ~n2723 & ~n2737;
  assign n2869 = ~n2738 & ~n2868;
  assign n2870 = ~n2867 & n2869;
  assign n2871 = ~n2714 & ~n2722;
  assign n2872 = ~n2723 & ~n2871;
  assign n2873 = ~n2600 & n2808;
  assign n2874 = n2596 & n2810;
  assign n2875 = n2593 & n2802;
  assign n2876 = ~n2874 & ~n2875;
  assign n2877 = ~n2873 & n2876;
  assign n2878 = ~n2817 & n2877;
  assign n2879 = n2706 & n2877;
  assign n2880 = ~n2878 & ~n2879;
  assign n2881 = n1021 & ~n2880;
  assign n2882 = ~n1021 & n2880;
  assign n2883 = ~n2881 & ~n2882;
  assign n2884 = n2872 & n2883;
  assign n2885 = ~n2607 & n2810;
  assign n2886 = ~n2604 & n2802;
  assign n2887 = ~n2885 & ~n2886;
  assign n2888 = ~n2673 & n2817;
  assign n2889 = n2887 & ~n2888;
  assign n2890 = ~n1021 & ~n2889;
  assign n2891 = ~n1021 & ~n2890;
  assign n2892 = ~n2889 & ~n2890;
  assign n2893 = ~n2891 & ~n2892;
  assign n2894 = ~n2607 & ~n2801;
  assign n2895 = ~n1021 & ~n2894;
  assign n2896 = ~n2893 & n2895;
  assign n2897 = ~n2600 & n2802;
  assign n2898 = ~n2607 & n2808;
  assign n2899 = ~n2604 & n2810;
  assign n2900 = ~n2898 & ~n2899;
  assign n2901 = ~n2897 & n2900;
  assign n2902 = ~n2732 & n2901;
  assign n2903 = ~n2817 & n2901;
  assign n2904 = ~n2902 & ~n2903;
  assign n2905 = n1021 & ~n2904;
  assign n2906 = ~n1021 & n2904;
  assign n2907 = ~n2905 & ~n2906;
  assign n2908 = n2896 & n2907;
  assign n2909 = n2713 & n2908;
  assign n2910 = n2908 & ~n2909;
  assign n2911 = n2713 & ~n2909;
  assign n2912 = ~n2910 & ~n2911;
  assign n2913 = ~n2600 & n2810;
  assign n2914 = n2596 & n2802;
  assign n2915 = ~n2604 & n2808;
  assign n2916 = ~n2914 & ~n2915;
  assign n2917 = ~n2913 & n2916;
  assign n2918 = ~n2750 & n2817;
  assign n2919 = n2917 & ~n2918;
  assign n2920 = ~n1021 & ~n2919;
  assign n2921 = ~n1021 & ~n2920;
  assign n2922 = ~n2919 & ~n2920;
  assign n2923 = ~n2921 & ~n2922;
  assign n2924 = ~n2912 & ~n2923;
  assign n2925 = ~n2909 & ~n2924;
  assign n2926 = ~n2872 & ~n2883;
  assign n2927 = ~n2884 & ~n2926;
  assign n2928 = ~n2925 & n2927;
  assign n2929 = ~n2884 & ~n2928;
  assign n2930 = ~n2867 & ~n2870;
  assign n2931 = n2869 & ~n2870;
  assign n2932 = ~n2930 & ~n2931;
  assign n2933 = ~n2929 & ~n2932;
  assign n2934 = ~n2870 & ~n2933;
  assign n2935 = ~n2842 & ~n2856;
  assign n2936 = n2855 & ~n2856;
  assign n2937 = ~n2935 & ~n2936;
  assign n2938 = ~n2934 & ~n2937;
  assign n2939 = ~n2856 & ~n2938;
  assign n2940 = ~n2836 & ~n2839;
  assign n2941 = n2838 & ~n2839;
  assign n2942 = ~n2940 & ~n2941;
  assign n2943 = ~n2939 & ~n2942;
  assign n2944 = ~n2839 & ~n2943;
  assign n2945 = n2795 & ~n2823;
  assign n2946 = n2822 & ~n2823;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = ~n2944 & ~n2947;
  assign n2949 = ~n2823 & ~n2948;
  assign n2950 = ~n2586 & n2699;
  assign n2951 = n2593 & n2695;
  assign n2952 = ~n2590 & n2697;
  assign n2953 = ~n2951 & ~n2952;
  assign n2954 = ~n2950 & n2953;
  assign n2955 = n2690 & n2849;
  assign n2956 = n2954 & ~n2955;
  assign n2957 = ~n669 & ~n2956;
  assign n2958 = n669 & n2956;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = ~n2600 & n2666;
  assign n2961 = n2596 & n2668;
  assign n2962 = ~n2604 & n2776;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = ~n2960 & n2963;
  assign n2965 = n2674 & ~n2750;
  assign n2966 = n2964 & ~n2965;
  assign n2967 = ~n525 & ~n2966;
  assign n2968 = ~n2966 & ~n2967;
  assign n2969 = ~n525 & ~n2967;
  assign n2970 = ~n2968 & ~n2969;
  assign n2971 = ~n525 & ~n2607;
  assign n2972 = ~n2787 & ~n2971;
  assign n2973 = n2787 & n2971;
  assign n2974 = ~n2970 & ~n2973;
  assign n2975 = ~n2972 & n2974;
  assign n2976 = ~n2970 & ~n2975;
  assign n2977 = ~n2973 & ~n2975;
  assign n2978 = ~n2972 & n2977;
  assign n2979 = ~n2976 & ~n2978;
  assign n2980 = n2959 & ~n2979;
  assign n2981 = n2959 & ~n2980;
  assign n2982 = ~n2979 & ~n2980;
  assign n2983 = ~n2981 & ~n2982;
  assign n2984 = ~n2790 & ~n2794;
  assign n2985 = n2983 & n2984;
  assign n2986 = ~n2983 & ~n2984;
  assign n2987 = ~n2985 & ~n2986;
  assign n2988 = n2634 & ~n2636;
  assign n2989 = ~n2637 & ~n2988;
  assign n2990 = ~n2575 & n2802;
  assign n2991 = ~n2582 & n2808;
  assign n2992 = n2578 & n2810;
  assign n2993 = ~n2991 & ~n2992;
  assign n2994 = ~n2990 & n2993;
  assign n2995 = ~n2989 & n2994;
  assign n2996 = ~n2817 & n2994;
  assign n2997 = ~n2995 & ~n2996;
  assign n2998 = n1021 & ~n2997;
  assign n2999 = ~n1021 & n2997;
  assign n3000 = ~n2998 & ~n2999;
  assign n3001 = n2987 & n3000;
  assign n3002 = n2987 & ~n3001;
  assign n3003 = n3000 & ~n3001;
  assign n3004 = ~n3002 & ~n3003;
  assign n3005 = ~n2949 & ~n3004;
  assign n3006 = ~n2949 & ~n3005;
  assign n3007 = ~n3004 & ~n3005;
  assign n3008 = ~n3006 & ~n3007;
  assign n3009 = n2657 & ~n3008;
  assign n3010 = n2657 & ~n3009;
  assign n3011 = ~n3008 & ~n3009;
  assign n3012 = ~n3010 & ~n3011;
  assign n3013 = ~n2944 & ~n2948;
  assign n3014 = ~n2947 & ~n2948;
  assign n3015 = ~n3013 & ~n3014;
  assign n3016 = n295 & ~n2566;
  assign n3017 = n2560 & ~n2575;
  assign n3018 = n2562 & n2567;
  assign n3019 = ~n3017 & ~n3018;
  assign n3020 = ~n3016 & n3019;
  assign n3021 = n2642 & ~n2644;
  assign n3022 = ~n2645 & ~n3021;
  assign n3023 = n2571 & n3022;
  assign n3024 = n3020 & ~n3023;
  assign n3025 = ~n275 & ~n3024;
  assign n3026 = n275 & n3024;
  assign n3027 = ~n3025 & ~n3026;
  assign n3028 = ~n3015 & n3027;
  assign n3029 = n3027 & ~n3028;
  assign n3030 = ~n3015 & ~n3028;
  assign n3031 = ~n3029 & ~n3030;
  assign n3032 = ~n2939 & n2942;
  assign n3033 = n2939 & ~n2942;
  assign n3034 = ~n3032 & ~n3033;
  assign n3035 = n295 & n2562;
  assign n3036 = n2560 & n2578;
  assign n3037 = n2567 & ~n2575;
  assign n3038 = ~n3036 & ~n3037;
  assign n3039 = ~n3035 & n3038;
  assign n3040 = ~n2571 & n3039;
  assign n3041 = n2638 & ~n2640;
  assign n3042 = ~n2641 & ~n3041;
  assign n3043 = n3039 & ~n3042;
  assign n3044 = ~n3040 & ~n3043;
  assign n3045 = n275 & ~n3044;
  assign n3046 = ~n275 & n3044;
  assign n3047 = ~n3045 & ~n3046;
  assign n3048 = ~n3034 & n3047;
  assign n3049 = ~n2934 & ~n2938;
  assign n3050 = ~n2937 & ~n2938;
  assign n3051 = ~n3049 & ~n3050;
  assign n3052 = n295 & ~n2575;
  assign n3053 = n2560 & ~n2582;
  assign n3054 = n2567 & n2578;
  assign n3055 = ~n3053 & ~n3054;
  assign n3056 = ~n3052 & n3055;
  assign n3057 = ~n2571 & n3056;
  assign n3058 = ~n2989 & n3056;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = n275 & ~n3059;
  assign n3061 = ~n275 & n3059;
  assign n3062 = ~n3060 & ~n3061;
  assign n3063 = ~n3051 & n3062;
  assign n3064 = ~n2929 & n2932;
  assign n3065 = n2929 & ~n2932;
  assign n3066 = ~n3064 & ~n3065;
  assign n3067 = n295 & n2578;
  assign n3068 = n2560 & ~n2586;
  assign n3069 = n2567 & ~n2582;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = ~n3067 & n3070;
  assign n3072 = ~n2571 & n3071;
  assign n3073 = ~n2815 & n3071;
  assign n3074 = ~n3072 & ~n3073;
  assign n3075 = n275 & ~n3074;
  assign n3076 = ~n275 & n3074;
  assign n3077 = ~n3075 & ~n3076;
  assign n3078 = ~n3066 & n3077;
  assign n3079 = n295 & ~n2582;
  assign n3080 = n2560 & ~n2590;
  assign n3081 = n2567 & ~n2586;
  assign n3082 = ~n3080 & ~n3081;
  assign n3083 = ~n3079 & n3082;
  assign n3084 = n2571 & n2830;
  assign n3085 = n3083 & ~n3084;
  assign n3086 = ~n275 & ~n3085;
  assign n3087 = n275 & n3085;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = n2925 & ~n2927;
  assign n3090 = ~n2928 & ~n3089;
  assign n3091 = n3088 & n3090;
  assign n3092 = ~n2912 & ~n2924;
  assign n3093 = ~n2923 & ~n2924;
  assign n3094 = ~n3092 & ~n3093;
  assign n3095 = n295 & ~n2586;
  assign n3096 = n2560 & n2593;
  assign n3097 = n2567 & ~n2590;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = ~n3095 & n3098;
  assign n3100 = ~n2571 & n3099;
  assign n3101 = ~n2849 & n3099;
  assign n3102 = ~n3100 & ~n3101;
  assign n3103 = n275 & ~n3102;
  assign n3104 = ~n275 & n3102;
  assign n3105 = ~n3103 & ~n3104;
  assign n3106 = ~n3094 & n3105;
  assign n3107 = n295 & ~n2590;
  assign n3108 = n2560 & n2596;
  assign n3109 = n2567 & n2593;
  assign n3110 = ~n3108 & ~n3109;
  assign n3111 = ~n3107 & n3110;
  assign n3112 = n2571 & n2768;
  assign n3113 = n3111 & ~n3112;
  assign n3114 = ~n275 & ~n3113;
  assign n3115 = n275 & n3113;
  assign n3116 = ~n3114 & ~n3115;
  assign n3117 = ~n2896 & ~n2907;
  assign n3118 = ~n2908 & ~n3117;
  assign n3119 = n3116 & n3118;
  assign n3120 = n2893 & ~n2895;
  assign n3121 = ~n2896 & ~n3120;
  assign n3122 = n2560 & ~n2600;
  assign n3123 = n2567 & n2596;
  assign n3124 = n295 & n2593;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = ~n3122 & n3125;
  assign n3127 = ~n2571 & n3126;
  assign n3128 = n2706 & n3126;
  assign n3129 = ~n3127 & ~n3128;
  assign n3130 = n275 & ~n3129;
  assign n3131 = ~n275 & n3129;
  assign n3132 = ~n3130 & ~n3131;
  assign n3133 = n3121 & n3132;
  assign n3134 = ~n294 & ~n2607;
  assign n3135 = ~n275 & ~n3134;
  assign n3136 = n2567 & ~n2607;
  assign n3137 = n295 & ~n2604;
  assign n3138 = ~n3136 & ~n3137;
  assign n3139 = n2571 & ~n2673;
  assign n3140 = n3138 & ~n3139;
  assign n3141 = ~n275 & ~n3140;
  assign n3142 = n275 & n3140;
  assign n3143 = ~n3141 & ~n3142;
  assign n3144 = n3135 & n3143;
  assign n3145 = n295 & ~n2600;
  assign n3146 = n2560 & ~n2607;
  assign n3147 = n2567 & ~n2604;
  assign n3148 = ~n3146 & ~n3147;
  assign n3149 = ~n3145 & n3148;
  assign n3150 = ~n2571 & n3149;
  assign n3151 = ~n2732 & n3149;
  assign n3152 = ~n3150 & ~n3151;
  assign n3153 = n275 & ~n3152;
  assign n3154 = ~n275 & n3152;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = n3144 & n3155;
  assign n3157 = n2894 & n3156;
  assign n3158 = n3156 & ~n3157;
  assign n3159 = n2894 & ~n3157;
  assign n3160 = ~n3158 & ~n3159;
  assign n3161 = n2567 & ~n2600;
  assign n3162 = n295 & n2596;
  assign n3163 = n2560 & ~n2604;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = ~n3161 & n3164;
  assign n3166 = n2571 & ~n2750;
  assign n3167 = n3165 & ~n3166;
  assign n3168 = ~n275 & ~n3167;
  assign n3169 = n275 & n3167;
  assign n3170 = ~n3168 & ~n3169;
  assign n3171 = ~n3160 & n3170;
  assign n3172 = ~n3157 & ~n3171;
  assign n3173 = ~n3121 & ~n3132;
  assign n3174 = ~n3133 & ~n3173;
  assign n3175 = ~n3172 & n3174;
  assign n3176 = ~n3133 & ~n3175;
  assign n3177 = ~n3116 & ~n3118;
  assign n3178 = ~n3119 & ~n3177;
  assign n3179 = ~n3176 & n3178;
  assign n3180 = ~n3119 & ~n3179;
  assign n3181 = ~n3094 & ~n3106;
  assign n3182 = n3105 & ~n3106;
  assign n3183 = ~n3181 & ~n3182;
  assign n3184 = ~n3180 & ~n3183;
  assign n3185 = ~n3106 & ~n3184;
  assign n3186 = ~n3088 & ~n3090;
  assign n3187 = ~n3091 & ~n3186;
  assign n3188 = ~n3185 & n3187;
  assign n3189 = ~n3091 & ~n3188;
  assign n3190 = ~n3066 & ~n3078;
  assign n3191 = n3077 & ~n3078;
  assign n3192 = ~n3190 & ~n3191;
  assign n3193 = ~n3189 & ~n3192;
  assign n3194 = ~n3078 & ~n3193;
  assign n3195 = ~n3051 & ~n3063;
  assign n3196 = n3062 & ~n3063;
  assign n3197 = ~n3195 & ~n3196;
  assign n3198 = ~n3194 & ~n3197;
  assign n3199 = ~n3063 & ~n3198;
  assign n3200 = n3034 & ~n3047;
  assign n3201 = ~n3048 & ~n3200;
  assign n3202 = ~n3199 & n3201;
  assign n3203 = ~n3048 & ~n3202;
  assign n3204 = ~n3031 & ~n3203;
  assign n3205 = ~n3028 & ~n3204;
  assign n3206 = n3012 & n3205;
  assign n3207 = ~n3012 & ~n3205;
  assign n3208 = ~n3206 & ~n3207;
  assign n3209 = \a[0]  & ~\a[22] ;
  assign n3210 = \a[1]  & ~n3209;
  assign n3211 = ~\a[1]  & n3209;
  assign n3212 = ~n3210 & ~n3211;
  assign n3213 = ~n291 & n3212;
  assign n3214 = n291 & ~n3212;
  assign n3215 = ~n3213 & ~n3214;
  assign n3216 = \a[0]  & ~n3215;
  assign n3217 = \a[0]  & n3215;
  assign n3218 = ~n324 & n809;
  assign n3219 = n485 & n3218;
  assign n3220 = n431 & n3219;
  assign n3221 = n2244 & n3220;
  assign n3222 = n2333 & n3221;
  assign n3223 = n2418 & n3222;
  assign n3224 = n976 & n3223;
  assign n3225 = ~n504 & n3224;
  assign n3226 = ~n297 & n3225;
  assign n3227 = ~n212 & n3226;
  assign n3228 = ~n258 & n3227;
  assign n3229 = ~n237 & n3228;
  assign n3230 = ~n300 & n808;
  assign n3231 = ~n326 & n3230;
  assign n3232 = n200 & n3231;
  assign n3233 = n2166 & n3232;
  assign n3234 = ~n415 & n3233;
  assign n3235 = ~n226 & n3234;
  assign n3236 = ~n213 & n3235;
  assign n3237 = ~n370 & n3236;
  assign n3238 = ~n447 & n3237;
  assign n3239 = ~n335 & n3238;
  assign n3240 = ~n114 & n3239;
  assign n3241 = ~n358 & n3240;
  assign n3242 = ~n106 & n3241;
  assign n3243 = ~n342 & n3242;
  assign n3244 = n744 & n2366;
  assign n3245 = n156 & n3244;
  assign n3246 = n768 & n3245;
  assign n3247 = n3243 & n3246;
  assign n3248 = n210 & n3247;
  assign n3249 = ~n150 & n3248;
  assign n3250 = ~n176 & n3249;
  assign n3251 = ~n220 & n3250;
  assign n3252 = ~n227 & n3251;
  assign n3253 = ~n186 & n3252;
  assign n3254 = ~n446 & n3253;
  assign n3255 = ~n361 & n3254;
  assign n3256 = ~n477 & n3255;
  assign n3257 = n2552 & n3256;
  assign n3258 = n3229 & n3257;
  assign n3259 = ~n134 & ~n405;
  assign n3260 = n349 & n423;
  assign n3261 = n1165 & n3260;
  assign n3262 = n397 & n3261;
  assign n3263 = n437 & n3262;
  assign n3264 = n314 & n3263;
  assign n3265 = n485 & n3264;
  assign n3266 = n502 & n3265;
  assign n3267 = n453 & n3266;
  assign n3268 = n3259 & n3267;
  assign n3269 = ~n140 & n3268;
  assign n3270 = ~n3258 & n3269;
  assign n3271 = n3258 & ~n3269;
  assign n3272 = ~n3270 & ~n3271;
  assign n3273 = n3217 & n3272;
  assign n3274 = n288 & ~n3215;
  assign n3275 = ~n2552 & n3256;
  assign n3276 = n2552 & ~n3256;
  assign n3277 = ~n3275 & ~n3276;
  assign n3278 = n3274 & n3277;
  assign n3279 = ~n3229 & ~n3257;
  assign n3280 = ~n3258 & ~n3279;
  assign n3281 = ~\a[0]  & ~n3212;
  assign n3282 = ~n3280 & n3281;
  assign n3283 = ~n3278 & ~n3282;
  assign n3284 = ~n3273 & n3283;
  assign n3285 = ~n3216 & n3284;
  assign n3286 = n3277 & ~n3280;
  assign n3287 = ~n2554 & n3277;
  assign n3288 = ~n2647 & ~n2650;
  assign n3289 = n2554 & ~n3277;
  assign n3290 = ~n3287 & ~n3289;
  assign n3291 = ~n3288 & n3290;
  assign n3292 = ~n3287 & ~n3291;
  assign n3293 = ~n3277 & n3280;
  assign n3294 = ~n3286 & ~n3293;
  assign n3295 = ~n3292 & n3294;
  assign n3296 = ~n3286 & ~n3295;
  assign n3297 = ~n3272 & n3280;
  assign n3298 = n3272 & ~n3280;
  assign n3299 = ~n3297 & ~n3298;
  assign n3300 = ~n3296 & n3299;
  assign n3301 = n3296 & ~n3299;
  assign n3302 = ~n3300 & ~n3301;
  assign n3303 = n3284 & ~n3302;
  assign n3304 = ~n3285 & ~n3303;
  assign n3305 = n291 & ~n3304;
  assign n3306 = ~n291 & n3304;
  assign n3307 = ~n3305 & ~n3306;
  assign n3308 = n3208 & n3307;
  assign n3309 = n3031 & n3203;
  assign n3310 = ~n3204 & ~n3309;
  assign n3311 = n3217 & ~n3280;
  assign n3312 = ~n2554 & n3274;
  assign n3313 = n3277 & n3281;
  assign n3314 = ~n3312 & ~n3313;
  assign n3315 = ~n3311 & n3314;
  assign n3316 = ~n3216 & n3315;
  assign n3317 = n3292 & ~n3294;
  assign n3318 = ~n3295 & ~n3317;
  assign n3319 = n3315 & ~n3318;
  assign n3320 = ~n3316 & ~n3319;
  assign n3321 = n291 & ~n3320;
  assign n3322 = ~n291 & n3320;
  assign n3323 = ~n3321 & ~n3322;
  assign n3324 = n3310 & n3323;
  assign n3325 = n3199 & ~n3201;
  assign n3326 = n3217 & n3277;
  assign n3327 = ~n2566 & n3274;
  assign n3328 = ~n2554 & n3281;
  assign n3329 = ~n3327 & ~n3328;
  assign n3330 = ~n3326 & n3329;
  assign n3331 = n3288 & ~n3290;
  assign n3332 = ~n3291 & ~n3331;
  assign n3333 = n3216 & n3332;
  assign n3334 = n3330 & ~n3333;
  assign n3335 = ~n291 & ~n3334;
  assign n3336 = ~n3334 & ~n3335;
  assign n3337 = ~n291 & ~n3335;
  assign n3338 = ~n3336 & ~n3337;
  assign n3339 = n2562 & n3217;
  assign n3340 = n2578 & n3274;
  assign n3341 = ~n2575 & n3281;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = ~n3339 & n3342;
  assign n3344 = ~n291 & ~n3343;
  assign n3345 = n3042 & n3216;
  assign n3346 = n3343 & ~n3345;
  assign n3347 = n291 & n3346;
  assign n3348 = ~n291 & n3216;
  assign n3349 = n3042 & n3348;
  assign n3350 = ~n2575 & n3217;
  assign n3351 = ~n2582 & n3274;
  assign n3352 = n2578 & n3281;
  assign n3353 = ~n3351 & ~n3352;
  assign n3354 = ~n3350 & n3353;
  assign n3355 = ~n291 & ~n3354;
  assign n3356 = n2989 & n3216;
  assign n3357 = n3354 & ~n3356;
  assign n3358 = n291 & n3357;
  assign n3359 = n2989 & n3348;
  assign n3360 = n2578 & n3217;
  assign n3361 = ~n2586 & n3274;
  assign n3362 = ~n2582 & n3281;
  assign n3363 = ~n3361 & ~n3362;
  assign n3364 = ~n3360 & n3363;
  assign n3365 = ~n291 & ~n3364;
  assign n3366 = n2815 & n3216;
  assign n3367 = n3364 & ~n3366;
  assign n3368 = n291 & n3367;
  assign n3369 = n2815 & n3348;
  assign n3370 = n3172 & ~n3174;
  assign n3371 = ~n2586 & n3217;
  assign n3372 = n2593 & n3274;
  assign n3373 = ~n2590 & n3281;
  assign n3374 = ~n3372 & ~n3373;
  assign n3375 = ~n3371 & n3374;
  assign n3376 = ~n291 & ~n3375;
  assign n3377 = n2849 & n3216;
  assign n3378 = n3375 & ~n3377;
  assign n3379 = n291 & n3378;
  assign n3380 = n2849 & n3348;
  assign n3381 = ~n3144 & ~n3155;
  assign n3382 = ~n2600 & n3274;
  assign n3383 = n2596 & n3281;
  assign n3384 = n2593 & n3217;
  assign n3385 = ~n3383 & ~n3384;
  assign n3386 = ~n3382 & n3385;
  assign n3387 = ~n291 & ~n3386;
  assign n3388 = ~n2706 & n3216;
  assign n3389 = n3386 & ~n3388;
  assign n3390 = n291 & n3389;
  assign n3391 = ~n2706 & n3348;
  assign n3392 = \a[0]  & ~n2607;
  assign n3393 = n2732 & n3348;
  assign n3394 = ~n2600 & n3217;
  assign n3395 = ~n2607 & n3274;
  assign n3396 = ~n2604 & n3281;
  assign n3397 = ~n3395 & ~n3396;
  assign n3398 = ~n3394 & n3397;
  assign n3399 = ~n291 & ~n3398;
  assign n3400 = ~n2673 & n3348;
  assign n3401 = ~n2604 & n3217;
  assign n3402 = ~n2607 & n3281;
  assign n3403 = ~n291 & ~n3402;
  assign n3404 = ~n3401 & n3403;
  assign n3405 = ~n3400 & n3404;
  assign n3406 = ~n3399 & n3405;
  assign n3407 = ~n3393 & n3406;
  assign n3408 = ~n3392 & n3407;
  assign n3409 = ~n3134 & ~n3408;
  assign n3410 = ~n2600 & n3281;
  assign n3411 = n2596 & n3217;
  assign n3412 = ~n2604 & n3274;
  assign n3413 = ~n3411 & ~n3412;
  assign n3414 = ~n3410 & n3413;
  assign n3415 = ~n2750 & n3216;
  assign n3416 = n3414 & ~n3415;
  assign n3417 = ~n291 & ~n3416;
  assign n3418 = n291 & n3416;
  assign n3419 = ~n3417 & ~n3418;
  assign n3420 = ~n3409 & n3419;
  assign n3421 = n3134 & n3408;
  assign n3422 = ~n3420 & ~n3421;
  assign n3423 = ~n3135 & ~n3143;
  assign n3424 = ~n3144 & ~n3423;
  assign n3425 = n3422 & ~n3424;
  assign n3426 = ~n3391 & ~n3425;
  assign n3427 = ~n3390 & n3426;
  assign n3428 = ~n3387 & n3427;
  assign n3429 = ~n3422 & n3424;
  assign n3430 = ~n3428 & ~n3429;
  assign n3431 = ~n2590 & n3217;
  assign n3432 = n2596 & n3274;
  assign n3433 = n2593 & n3281;
  assign n3434 = ~n3432 & ~n3433;
  assign n3435 = ~n3431 & n3434;
  assign n3436 = n2768 & n3216;
  assign n3437 = n3435 & ~n3436;
  assign n3438 = ~n291 & ~n3437;
  assign n3439 = ~n3437 & ~n3438;
  assign n3440 = ~n291 & ~n3438;
  assign n3441 = ~n3439 & ~n3440;
  assign n3442 = n3430 & n3441;
  assign n3443 = ~n3156 & ~n3442;
  assign n3444 = ~n3381 & n3443;
  assign n3445 = ~n3430 & ~n3441;
  assign n3446 = ~n3444 & ~n3445;
  assign n3447 = ~n3160 & ~n3171;
  assign n3448 = n3170 & ~n3171;
  assign n3449 = ~n3447 & ~n3448;
  assign n3450 = n3446 & n3449;
  assign n3451 = ~n3380 & ~n3450;
  assign n3452 = ~n3379 & n3451;
  assign n3453 = ~n3376 & n3452;
  assign n3454 = ~n3446 & ~n3449;
  assign n3455 = ~n3453 & ~n3454;
  assign n3456 = ~n2582 & n3217;
  assign n3457 = ~n2590 & n3274;
  assign n3458 = ~n2586 & n3281;
  assign n3459 = ~n3457 & ~n3458;
  assign n3460 = ~n3456 & n3459;
  assign n3461 = n2830 & n3216;
  assign n3462 = n3460 & ~n3461;
  assign n3463 = ~n291 & ~n3462;
  assign n3464 = ~n3462 & ~n3463;
  assign n3465 = ~n291 & ~n3463;
  assign n3466 = ~n3464 & ~n3465;
  assign n3467 = n3455 & n3466;
  assign n3468 = ~n3175 & ~n3467;
  assign n3469 = ~n3370 & n3468;
  assign n3470 = ~n3455 & ~n3466;
  assign n3471 = ~n3469 & ~n3470;
  assign n3472 = n3176 & ~n3178;
  assign n3473 = ~n3179 & ~n3472;
  assign n3474 = n3471 & ~n3473;
  assign n3475 = ~n3369 & ~n3474;
  assign n3476 = ~n3368 & n3475;
  assign n3477 = ~n3365 & n3476;
  assign n3478 = ~n3471 & n3473;
  assign n3479 = ~n3477 & ~n3478;
  assign n3480 = ~n3180 & ~n3184;
  assign n3481 = ~n3183 & ~n3184;
  assign n3482 = ~n3480 & ~n3481;
  assign n3483 = n3479 & n3482;
  assign n3484 = ~n3359 & ~n3483;
  assign n3485 = ~n3358 & n3484;
  assign n3486 = ~n3355 & n3485;
  assign n3487 = ~n3479 & ~n3482;
  assign n3488 = ~n3486 & ~n3487;
  assign n3489 = n3185 & ~n3187;
  assign n3490 = ~n3188 & ~n3489;
  assign n3491 = n3488 & ~n3490;
  assign n3492 = ~n3349 & ~n3491;
  assign n3493 = ~n3347 & n3492;
  assign n3494 = ~n3344 & n3493;
  assign n3495 = ~n3488 & n3490;
  assign n3496 = ~n3494 & ~n3495;
  assign n3497 = n3189 & n3192;
  assign n3498 = ~n3193 & ~n3497;
  assign n3499 = ~n3496 & n3498;
  assign n3500 = ~n2566 & n3217;
  assign n3501 = ~n2575 & n3274;
  assign n3502 = n2562 & n3281;
  assign n3503 = ~n3501 & ~n3502;
  assign n3504 = ~n3500 & n3503;
  assign n3505 = n3022 & n3216;
  assign n3506 = n3504 & ~n3505;
  assign n3507 = n291 & ~n3506;
  assign n3508 = ~n291 & n3506;
  assign n3509 = ~n3507 & ~n3508;
  assign n3510 = ~n3499 & n3509;
  assign n3511 = n3496 & ~n3498;
  assign n3512 = ~n3510 & ~n3511;
  assign n3513 = n3194 & n3197;
  assign n3514 = ~n3198 & ~n3513;
  assign n3515 = ~n3512 & ~n3514;
  assign n3516 = ~n2554 & n3217;
  assign n3517 = n2562 & n3274;
  assign n3518 = ~n2566 & n3281;
  assign n3519 = ~n3517 & ~n3518;
  assign n3520 = ~n3516 & n3519;
  assign n3521 = n2652 & n3216;
  assign n3522 = n3520 & ~n3521;
  assign n3523 = ~n291 & ~n3522;
  assign n3524 = n291 & n3522;
  assign n3525 = ~n3523 & ~n3524;
  assign n3526 = ~n3515 & n3525;
  assign n3527 = n3512 & n3514;
  assign n3528 = ~n3526 & ~n3527;
  assign n3529 = n3338 & n3528;
  assign n3530 = ~n3202 & ~n3529;
  assign n3531 = ~n3325 & n3530;
  assign n3532 = ~n3338 & ~n3528;
  assign n3533 = ~n3531 & ~n3532;
  assign n3534 = n3310 & ~n3324;
  assign n3535 = n3323 & ~n3324;
  assign n3536 = ~n3534 & ~n3535;
  assign n3537 = ~n3533 & ~n3536;
  assign n3538 = ~n3324 & ~n3537;
  assign n3539 = n3208 & ~n3308;
  assign n3540 = n3307 & ~n3308;
  assign n3541 = ~n3539 & ~n3540;
  assign n3542 = ~n3538 & ~n3541;
  assign n3543 = ~n3308 & ~n3542;
  assign n3544 = ~n3009 & ~n3207;
  assign n3545 = n295 & n3277;
  assign n3546 = n2560 & ~n2566;
  assign n3547 = ~n2554 & n2567;
  assign n3548 = ~n3546 & ~n3547;
  assign n3549 = ~n3545 & n3548;
  assign n3550 = n2571 & n3332;
  assign n3551 = n3549 & ~n3550;
  assign n3552 = ~n275 & ~n3551;
  assign n3553 = n275 & n3551;
  assign n3554 = ~n3552 & ~n3553;
  assign n3555 = ~n3001 & ~n3005;
  assign n3556 = ~n2980 & ~n2986;
  assign n3557 = ~n2582 & n2699;
  assign n3558 = ~n2590 & n2695;
  assign n3559 = ~n2586 & n2697;
  assign n3560 = ~n3558 & ~n3559;
  assign n3561 = ~n3557 & n3560;
  assign n3562 = n2690 & n2830;
  assign n3563 = n3561 & ~n3562;
  assign n3564 = ~n669 & ~n3563;
  assign n3565 = n669 & n3563;
  assign n3566 = ~n3564 & ~n3565;
  assign n3567 = ~n525 & ~n2604;
  assign n3568 = ~n2600 & n2776;
  assign n3569 = n2596 & n2666;
  assign n3570 = n2593 & n2668;
  assign n3571 = ~n3569 & ~n3570;
  assign n3572 = ~n3568 & n3571;
  assign n3573 = n2674 & ~n2706;
  assign n3574 = n3572 & ~n3573;
  assign n3575 = ~n525 & ~n3574;
  assign n3576 = n3567 & ~n3575;
  assign n3577 = n3567 & ~n3576;
  assign n3578 = n525 & n3574;
  assign n3579 = ~n3575 & ~n3578;
  assign n3580 = ~n3576 & n3579;
  assign n3581 = ~n3577 & ~n3580;
  assign n3582 = ~n2977 & ~n3581;
  assign n3583 = ~n2977 & ~n3582;
  assign n3584 = ~n3581 & ~n3582;
  assign n3585 = ~n3583 & ~n3584;
  assign n3586 = n3566 & ~n3585;
  assign n3587 = n3566 & ~n3586;
  assign n3588 = ~n3585 & ~n3586;
  assign n3589 = ~n3587 & ~n3588;
  assign n3590 = ~n3556 & n3589;
  assign n3591 = n3556 & ~n3589;
  assign n3592 = ~n3590 & ~n3591;
  assign n3593 = n2562 & n2802;
  assign n3594 = n2578 & n2808;
  assign n3595 = ~n2575 & n2810;
  assign n3596 = ~n3594 & ~n3595;
  assign n3597 = ~n3593 & n3596;
  assign n3598 = ~n3042 & n3597;
  assign n3599 = ~n2817 & n3597;
  assign n3600 = ~n3598 & ~n3599;
  assign n3601 = n1021 & ~n3600;
  assign n3602 = ~n1021 & n3600;
  assign n3603 = ~n3601 & ~n3602;
  assign n3604 = ~n3592 & n3603;
  assign n3605 = n3592 & ~n3603;
  assign n3606 = ~n3604 & ~n3605;
  assign n3607 = ~n3555 & n3606;
  assign n3608 = n3555 & ~n3606;
  assign n3609 = ~n3607 & ~n3608;
  assign n3610 = n3554 & n3609;
  assign n3611 = ~n3554 & ~n3609;
  assign n3612 = ~n3610 & ~n3611;
  assign n3613 = ~n3544 & n3612;
  assign n3614 = n3544 & ~n3612;
  assign n3615 = ~n3613 & ~n3614;
  assign n3616 = ~n348 & n502;
  assign n3617 = ~n148 & n3616;
  assign n3618 = n514 & n3617;
  assign n3619 = n485 & n3618;
  assign n3620 = n414 & n3619;
  assign n3621 = n404 & n3620;
  assign n3622 = ~n188 & n3621;
  assign n3623 = ~n219 & n3622;
  assign n3624 = ~n224 & n3623;
  assign n3625 = n3258 & n3269;
  assign n3626 = ~n3624 & ~n3625;
  assign n3627 = n3624 & n3625;
  assign n3628 = ~n3626 & ~n3627;
  assign n3629 = n3217 & ~n3628;
  assign n3630 = n3274 & ~n3280;
  assign n3631 = n3272 & n3281;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = ~n3629 & n3632;
  assign n3634 = ~n3216 & n3633;
  assign n3635 = ~n3298 & ~n3300;
  assign n3636 = ~n3272 & n3628;
  assign n3637 = n3272 & ~n3628;
  assign n3638 = ~n3636 & ~n3637;
  assign n3639 = ~n3635 & n3638;
  assign n3640 = n3635 & ~n3638;
  assign n3641 = ~n3639 & ~n3640;
  assign n3642 = n3633 & ~n3641;
  assign n3643 = ~n3634 & ~n3642;
  assign n3644 = n291 & ~n3643;
  assign n3645 = ~n291 & n3643;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = n3615 & n3646;
  assign n3648 = ~n3615 & ~n3646;
  assign n3649 = ~n3647 & ~n3648;
  assign n3650 = ~n3543 & n3649;
  assign n3651 = n3543 & ~n3649;
  assign n3652 = ~n3650 & ~n3651;
  assign n3653 = ~n271 & n3652;
  assign n3654 = ~n114 & ~n506;
  assign n3655 = ~n736 & n3654;
  assign n3656 = ~n296 & n3655;
  assign n3657 = ~n154 & n3656;
  assign n3658 = n806 & n3657;
  assign n3659 = ~n139 & n3658;
  assign n3660 = ~n150 & n3659;
  assign n3661 = ~n186 & n3660;
  assign n3662 = ~n313 & n3661;
  assign n3663 = ~n133 & n3662;
  assign n3664 = ~n359 & n3663;
  assign n3665 = ~n142 & n3664;
  assign n3666 = ~n106 & n3665;
  assign n3667 = n372 & n505;
  assign n3668 = n1134 & n3667;
  assign n3669 = ~n217 & n3668;
  assign n3670 = ~n255 & n3669;
  assign n3671 = ~n495 & n3670;
  assign n3672 = ~n553 & n3671;
  assign n3673 = ~n445 & n3672;
  assign n3674 = ~n471 & n3673;
  assign n3675 = ~n215 & n3674;
  assign n3676 = n789 & n3675;
  assign n3677 = ~n417 & n3676;
  assign n3678 = ~n298 & n3677;
  assign n3679 = n2454 & n3678;
  assign n3680 = n3666 & n3679;
  assign n3681 = n980 & n3680;
  assign n3682 = ~n137 & n3681;
  assign n3683 = ~n254 & n3682;
  assign n3684 = ~n327 & n3683;
  assign n3685 = ~n446 & n3684;
  assign n3686 = ~n146 & n3685;
  assign n3687 = ~n297 & n3686;
  assign n3688 = ~n335 & n3687;
  assign n3689 = ~n470 & n3688;
  assign n3690 = ~n342 & n3689;
  assign n3691 = n3538 & ~n3540;
  assign n3692 = ~n3539 & n3691;
  assign n3693 = ~n3542 & ~n3692;
  assign n3694 = n397 & n2278;
  assign n3695 = n2303 & n3694;
  assign n3696 = ~n144 & n3695;
  assign n3697 = ~n503 & n3696;
  assign n3698 = ~n356 & n3697;
  assign n3699 = ~n477 & n3698;
  assign n3700 = n341 & n813;
  assign n3701 = ~n137 & n3700;
  assign n3702 = ~n155 & n3701;
  assign n3703 = n460 & n2422;
  assign n3704 = n2433 & n3703;
  assign n3705 = n344 & n3704;
  assign n3706 = n3702 & n3705;
  assign n3707 = n3699 & n3706;
  assign n3708 = n2364 & n3707;
  assign n3709 = ~n415 & n3708;
  assign n3710 = ~n150 & n3709;
  assign n3711 = ~n317 & n3710;
  assign n3712 = ~n219 & n3711;
  assign n3713 = ~n174 & n3712;
  assign n3714 = ~n218 & n3713;
  assign n3715 = ~n302 & n3714;
  assign n3716 = n3533 & n3536;
  assign n3717 = ~n3537 & ~n3716;
  assign n3718 = ~n3715 & n3717;
  assign n3719 = ~n3693 & ~n3718;
  assign n3720 = ~n3690 & ~n3719;
  assign n3721 = n3693 & n3718;
  assign n3722 = ~n3720 & ~n3721;
  assign n3723 = ~n271 & ~n3653;
  assign n3724 = n3652 & ~n3653;
  assign n3725 = ~n3723 & ~n3724;
  assign n3726 = ~n3722 & ~n3725;
  assign n3727 = ~n3653 & ~n3726;
  assign n3728 = n239 & n590;
  assign n3729 = ~n350 & n3728;
  assign n3730 = ~n123 & n3729;
  assign n3731 = ~n313 & n3730;
  assign n3732 = ~n207 & n3731;
  assign n3733 = ~n445 & n3732;
  assign n3734 = ~n469 & n3733;
  assign n3735 = n353 & ~n468;
  assign n3736 = n334 & n3735;
  assign n3737 = n1162 & n3736;
  assign n3738 = n3734 & n3737;
  assign n3739 = n2418 & n3738;
  assign n3740 = ~n222 & n3739;
  assign n3741 = ~n317 & n3740;
  assign n3742 = ~n177 & n3741;
  assign n3743 = ~n218 & n3742;
  assign n3744 = ~n554 & n3743;
  assign n3745 = ~n211 & n3744;
  assign n3746 = ~n132 & n3745;
  assign n3747 = ~n223 & n3746;
  assign n3748 = ~n3627 & n3747;
  assign n3749 = n3627 & ~n3747;
  assign n3750 = ~n3748 & ~n3749;
  assign n3751 = n3217 & n3750;
  assign n3752 = n3272 & n3274;
  assign n3753 = n3281 & ~n3628;
  assign n3754 = ~n3752 & ~n3753;
  assign n3755 = ~n3751 & n3754;
  assign n3756 = ~n3637 & ~n3639;
  assign n3757 = n3628 & ~n3750;
  assign n3758 = ~n3628 & n3750;
  assign n3759 = ~n3757 & ~n3758;
  assign n3760 = ~n3756 & n3759;
  assign n3761 = n3756 & ~n3759;
  assign n3762 = ~n3760 & ~n3761;
  assign n3763 = n3216 & n3762;
  assign n3764 = n3755 & ~n3763;
  assign n3765 = ~n291 & ~n3764;
  assign n3766 = ~n3764 & ~n3765;
  assign n3767 = ~n291 & ~n3765;
  assign n3768 = ~n3766 & ~n3767;
  assign n3769 = ~n3610 & ~n3613;
  assign n3770 = ~n2566 & n2802;
  assign n3771 = ~n2575 & n2808;
  assign n3772 = n2562 & n2810;
  assign n3773 = ~n3771 & ~n3772;
  assign n3774 = ~n3770 & n3773;
  assign n3775 = n2817 & n3022;
  assign n3776 = n3774 & ~n3775;
  assign n3777 = ~n1021 & ~n3776;
  assign n3778 = ~n3776 & ~n3777;
  assign n3779 = ~n1021 & ~n3777;
  assign n3780 = ~n3778 & ~n3779;
  assign n3781 = ~n3556 & ~n3589;
  assign n3782 = ~n3586 & ~n3781;
  assign n3783 = ~n3576 & ~n3582;
  assign n3784 = ~n2590 & n2668;
  assign n3785 = n2596 & n2776;
  assign n3786 = n2593 & n2666;
  assign n3787 = ~n3785 & ~n3786;
  assign n3788 = ~n3784 & n3787;
  assign n3789 = n2674 & n2768;
  assign n3790 = n3788 & ~n3789;
  assign n3791 = ~n525 & n2600;
  assign n3792 = ~n3790 & n3791;
  assign n3793 = n3790 & ~n3791;
  assign n3794 = ~n3792 & ~n3793;
  assign n3795 = ~n3783 & n3794;
  assign n3796 = n3783 & ~n3794;
  assign n3797 = ~n3795 & ~n3796;
  assign n3798 = n2578 & n2699;
  assign n3799 = ~n2586 & n2695;
  assign n3800 = ~n2582 & n2697;
  assign n3801 = ~n3799 & ~n3800;
  assign n3802 = ~n3798 & n3801;
  assign n3803 = ~n2690 & n3802;
  assign n3804 = ~n2815 & n3802;
  assign n3805 = ~n3803 & ~n3804;
  assign n3806 = n669 & ~n3805;
  assign n3807 = ~n669 & n3805;
  assign n3808 = ~n3806 & ~n3807;
  assign n3809 = n3797 & n3808;
  assign n3810 = n3797 & ~n3809;
  assign n3811 = n3808 & ~n3809;
  assign n3812 = ~n3810 & ~n3811;
  assign n3813 = ~n3782 & ~n3812;
  assign n3814 = ~n3782 & ~n3813;
  assign n3815 = ~n3812 & ~n3813;
  assign n3816 = ~n3814 & ~n3815;
  assign n3817 = ~n3780 & ~n3816;
  assign n3818 = ~n3780 & ~n3817;
  assign n3819 = ~n3816 & ~n3817;
  assign n3820 = ~n3818 & ~n3819;
  assign n3821 = ~n3604 & ~n3607;
  assign n3822 = n3820 & n3821;
  assign n3823 = ~n3820 & ~n3821;
  assign n3824 = ~n3822 & ~n3823;
  assign n3825 = n295 & ~n3280;
  assign n3826 = ~n2554 & n2560;
  assign n3827 = n2567 & n3277;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = ~n3825 & n3828;
  assign n3830 = ~n2571 & n3829;
  assign n3831 = ~n3318 & n3829;
  assign n3832 = ~n3830 & ~n3831;
  assign n3833 = n275 & ~n3832;
  assign n3834 = ~n275 & n3832;
  assign n3835 = ~n3833 & ~n3834;
  assign n3836 = n3824 & n3835;
  assign n3837 = n3824 & ~n3836;
  assign n3838 = n3835 & ~n3836;
  assign n3839 = ~n3837 & ~n3838;
  assign n3840 = ~n3769 & ~n3839;
  assign n3841 = ~n3769 & ~n3840;
  assign n3842 = ~n3839 & ~n3840;
  assign n3843 = ~n3841 & ~n3842;
  assign n3844 = ~n3768 & ~n3843;
  assign n3845 = ~n3768 & ~n3844;
  assign n3846 = ~n3843 & ~n3844;
  assign n3847 = ~n3845 & ~n3846;
  assign n3848 = ~n3647 & ~n3650;
  assign n3849 = n3847 & n3848;
  assign n3850 = ~n3847 & ~n3848;
  assign n3851 = ~n3849 & ~n3850;
  assign n3852 = n239 & n1093;
  assign n3853 = n806 & n3852;
  assign n3854 = n1459 & n3853;
  assign n3855 = n2311 & n3854;
  assign n3856 = n643 & n3855;
  assign n3857 = n623 & n3856;
  assign n3858 = n210 & n3857;
  assign n3859 = ~n255 & n3858;
  assign n3860 = ~n148 & n3859;
  assign n3861 = ~n345 & n3860;
  assign n3862 = ~n3851 & n3861;
  assign n3863 = n3851 & ~n3861;
  assign n3864 = ~n3862 & ~n3863;
  assign n3865 = ~n3727 & n3864;
  assign n3866 = n3727 & ~n3864;
  assign n3867 = ~n3865 & ~n3866;
  assign n3868 = ~n3722 & ~n3726;
  assign n3869 = ~n3725 & ~n3726;
  assign n3870 = ~n3868 & ~n3869;
  assign n3871 = n3867 & ~n3870;
  assign n3872 = n3867 & ~n3871;
  assign n3873 = ~n3870 & ~n3871;
  assign \sin[0]  = n3872 | n3873;
  assign n3875 = ~n3863 & ~n3865;
  assign n3876 = n3627 & n3747;
  assign n3877 = n236 & n2433;
  assign n3878 = n457 & n3877;
  assign n3879 = n753 & n3878;
  assign n3880 = ~n169 & n3879;
  assign n3881 = ~n118 & n3880;
  assign n3882 = ~n166 & n3881;
  assign n3883 = ~n168 & n3882;
  assign n3884 = n316 & n555;
  assign n3885 = n815 & n3884;
  assign n3886 = n1476 & n3885;
  assign n3887 = n3883 & n3886;
  assign n3888 = n2432 & n3887;
  assign n3889 = n976 & n3888;
  assign n3890 = ~n495 & n3889;
  assign n3891 = ~n470 & n3890;
  assign n3892 = ~n367 & n3891;
  assign n3893 = ~n326 & n3892;
  assign n3894 = ~n3876 & n3893;
  assign n3895 = n3876 & ~n3893;
  assign n3896 = ~n3894 & ~n3895;
  assign n3897 = n3217 & n3896;
  assign n3898 = n3274 & ~n3628;
  assign n3899 = n3281 & n3750;
  assign n3900 = ~n3898 & ~n3899;
  assign n3901 = ~n3897 & n3900;
  assign n3902 = ~n3758 & ~n3760;
  assign n3903 = ~n3750 & ~n3896;
  assign n3904 = n3750 & n3896;
  assign n3905 = ~n3903 & ~n3904;
  assign n3906 = ~n3902 & n3905;
  assign n3907 = n3902 & ~n3905;
  assign n3908 = ~n3906 & ~n3907;
  assign n3909 = n3216 & n3908;
  assign n3910 = n3901 & ~n3909;
  assign n3911 = ~n291 & ~n3910;
  assign n3912 = ~n3910 & ~n3911;
  assign n3913 = ~n291 & ~n3911;
  assign n3914 = ~n3912 & ~n3913;
  assign n3915 = ~n3836 & ~n3840;
  assign n3916 = ~n2554 & n2802;
  assign n3917 = n2562 & n2808;
  assign n3918 = ~n2566 & n2810;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = ~n3916 & n3919;
  assign n3921 = n2652 & n2817;
  assign n3922 = n3920 & ~n3921;
  assign n3923 = ~n1021 & ~n3922;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = ~n1021 & ~n3923;
  assign n3926 = ~n3924 & ~n3925;
  assign n3927 = ~n3809 & ~n3813;
  assign n3928 = ~n525 & ~n2600;
  assign n3929 = n3790 & n3928;
  assign n3930 = ~n3795 & ~n3929;
  assign n3931 = ~n2586 & n2668;
  assign n3932 = n2593 & n2776;
  assign n3933 = ~n2590 & n2666;
  assign n3934 = ~n3932 & ~n3933;
  assign n3935 = ~n3931 & n3934;
  assign n3936 = n2674 & n2849;
  assign n3937 = n3935 & ~n3936;
  assign n3938 = ~n525 & ~n2596;
  assign n3939 = ~n3937 & n3938;
  assign n3940 = n3937 & ~n3938;
  assign n3941 = ~n3939 & ~n3940;
  assign n3942 = ~n3930 & n3941;
  assign n3943 = ~n3930 & ~n3942;
  assign n3944 = n3941 & ~n3942;
  assign n3945 = ~n3943 & ~n3944;
  assign n3946 = ~n2575 & n2699;
  assign n3947 = ~n2582 & n2695;
  assign n3948 = n2578 & n2697;
  assign n3949 = ~n3947 & ~n3948;
  assign n3950 = ~n3946 & n3949;
  assign n3951 = ~n2690 & n3950;
  assign n3952 = ~n2989 & n3950;
  assign n3953 = ~n3951 & ~n3952;
  assign n3954 = n669 & ~n3953;
  assign n3955 = ~n669 & n3953;
  assign n3956 = ~n3954 & ~n3955;
  assign n3957 = ~n3945 & n3956;
  assign n3958 = ~n3945 & ~n3957;
  assign n3959 = n3956 & ~n3957;
  assign n3960 = ~n3958 & ~n3959;
  assign n3961 = ~n3927 & ~n3960;
  assign n3962 = ~n3927 & ~n3961;
  assign n3963 = ~n3960 & ~n3961;
  assign n3964 = ~n3962 & ~n3963;
  assign n3965 = ~n3926 & ~n3964;
  assign n3966 = ~n3926 & ~n3965;
  assign n3967 = ~n3964 & ~n3965;
  assign n3968 = ~n3966 & ~n3967;
  assign n3969 = ~n3817 & ~n3823;
  assign n3970 = n3968 & n3969;
  assign n3971 = ~n3968 & ~n3969;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = n295 & n3272;
  assign n3974 = n2560 & n3277;
  assign n3975 = n2567 & ~n3280;
  assign n3976 = ~n3974 & ~n3975;
  assign n3977 = ~n3973 & n3976;
  assign n3978 = ~n2571 & n3977;
  assign n3979 = ~n3302 & n3977;
  assign n3980 = ~n3978 & ~n3979;
  assign n3981 = n275 & ~n3980;
  assign n3982 = ~n275 & n3980;
  assign n3983 = ~n3981 & ~n3982;
  assign n3984 = n3972 & n3983;
  assign n3985 = n3972 & ~n3984;
  assign n3986 = n3983 & ~n3984;
  assign n3987 = ~n3985 & ~n3986;
  assign n3988 = ~n3915 & ~n3987;
  assign n3989 = ~n3915 & ~n3988;
  assign n3990 = ~n3987 & ~n3988;
  assign n3991 = ~n3989 & ~n3990;
  assign n3992 = ~n3914 & ~n3991;
  assign n3993 = ~n3914 & ~n3992;
  assign n3994 = ~n3991 & ~n3992;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = ~n3844 & ~n3850;
  assign n3997 = n3995 & n3996;
  assign n3998 = ~n3995 & ~n3996;
  assign n3999 = ~n3997 & ~n3998;
  assign n4000 = ~n140 & ~n405;
  assign n4001 = ~n361 & n4000;
  assign n4002 = ~n258 & n4001;
  assign n4003 = n637 & n2340;
  assign n4004 = n2276 & n4003;
  assign n4005 = n249 & n4004;
  assign n4006 = n753 & n4005;
  assign n4007 = n4002 & n4006;
  assign n4008 = n210 & n4007;
  assign n4009 = n3231 & n4008;
  assign n4010 = ~n175 & n4009;
  assign n4011 = ~n155 & n4010;
  assign n4012 = ~n327 & n4011;
  assign n4013 = ~n191 & n4012;
  assign n4014 = ~n118 & n4013;
  assign n4015 = ~n445 & n4014;
  assign n4016 = ~n3999 & n4015;
  assign n4017 = n3999 & ~n4015;
  assign n4018 = ~n4016 & ~n4017;
  assign n4019 = ~n3875 & n4018;
  assign n4020 = n3875 & ~n4018;
  assign n4021 = ~n4019 & ~n4020;
  assign n4022 = n3871 & n4021;
  assign n4023 = ~n3871 & ~n4021;
  assign n4024 = ~n4022 & ~n4023;
  assign n4025 = \a[22]  & ~\a[23] ;
  assign n4026 = ~\a[22]  & \a[23] ;
  assign n4027 = ~n4025 & ~n4026;
  assign n4028 = \sin[0]  & ~n4027;
  assign n4029 = ~n4024 & n4028;
  assign n4030 = n4024 & ~n4028;
  assign \sin[1]  = n4029 | n4030;
  assign n4032 = ~n4017 & ~n4019;
  assign n4033 = n346 & ~n408;
  assign n4034 = ~n129 & n4033;
  assign n4035 = ~n228 & n4034;
  assign n4036 = ~n142 & n4035;
  assign n4037 = ~n132 & n4036;
  assign n4038 = n416 & n608;
  assign n4039 = n805 & n4038;
  assign n4040 = n4037 & n4039;
  assign n4041 = n3699 & n4040;
  assign n4042 = ~n313 & n4041;
  assign n4043 = ~n458 & n4042;
  assign n4044 = ~n504 & n4043;
  assign n4045 = ~n298 & n4044;
  assign n4046 = ~n146 & n4045;
  assign n4047 = ~n506 & n4046;
  assign n4048 = ~n326 & n4047;
  assign n4049 = ~n3992 & ~n3998;
  assign n4050 = n3274 & n3750;
  assign n4051 = n3281 & n3896;
  assign n4052 = ~n4050 & ~n4051;
  assign n4053 = ~n3750 & ~n3906;
  assign n4054 = n3896 & ~n4053;
  assign n4055 = ~n3896 & ~n3906;
  assign n4056 = ~n4054 & ~n4055;
  assign n4057 = n3216 & n4056;
  assign n4058 = n4052 & ~n4057;
  assign n4059 = ~n291 & ~n4058;
  assign n4060 = ~n4058 & ~n4059;
  assign n4061 = ~n291 & ~n4059;
  assign n4062 = ~n4060 & ~n4061;
  assign n4063 = ~n3984 & ~n3988;
  assign n4064 = n2802 & n3277;
  assign n4065 = ~n2566 & n2808;
  assign n4066 = ~n2554 & n2810;
  assign n4067 = ~n4065 & ~n4066;
  assign n4068 = ~n4064 & n4067;
  assign n4069 = n2817 & n3332;
  assign n4070 = n4068 & ~n4069;
  assign n4071 = ~n1021 & ~n4070;
  assign n4072 = ~n4070 & ~n4071;
  assign n4073 = ~n1021 & ~n4071;
  assign n4074 = ~n4072 & ~n4073;
  assign n4075 = ~n3957 & ~n3961;
  assign n4076 = ~n525 & n3937;
  assign n4077 = n2596 & n4076;
  assign n4078 = ~n3942 & ~n4077;
  assign n4079 = ~n2582 & n2668;
  assign n4080 = ~n2590 & n2776;
  assign n4081 = ~n2586 & n2666;
  assign n4082 = ~n4080 & ~n4081;
  assign n4083 = ~n4079 & n4082;
  assign n4084 = n2674 & n2830;
  assign n4085 = n4083 & ~n4084;
  assign n4086 = ~n525 & ~n2593;
  assign n4087 = ~n4085 & n4086;
  assign n4088 = n4085 & ~n4086;
  assign n4089 = ~n4087 & ~n4088;
  assign n4090 = ~n4078 & n4089;
  assign n4091 = ~n4078 & ~n4090;
  assign n4092 = n4089 & ~n4090;
  assign n4093 = ~n4091 & ~n4092;
  assign n4094 = n2562 & n2699;
  assign n4095 = n2578 & n2695;
  assign n4096 = ~n2575 & n2697;
  assign n4097 = ~n4095 & ~n4096;
  assign n4098 = ~n4094 & n4097;
  assign n4099 = ~n2690 & n4098;
  assign n4100 = ~n3042 & n4098;
  assign n4101 = ~n4099 & ~n4100;
  assign n4102 = n669 & ~n4101;
  assign n4103 = ~n669 & n4101;
  assign n4104 = ~n4102 & ~n4103;
  assign n4105 = ~n4093 & n4104;
  assign n4106 = ~n4093 & ~n4105;
  assign n4107 = n4104 & ~n4105;
  assign n4108 = ~n4106 & ~n4107;
  assign n4109 = ~n4075 & ~n4108;
  assign n4110 = ~n4075 & ~n4109;
  assign n4111 = ~n4108 & ~n4109;
  assign n4112 = ~n4110 & ~n4111;
  assign n4113 = ~n4074 & ~n4112;
  assign n4114 = ~n4074 & ~n4113;
  assign n4115 = ~n4112 & ~n4113;
  assign n4116 = ~n4114 & ~n4115;
  assign n4117 = ~n3965 & ~n3971;
  assign n4118 = n4116 & n4117;
  assign n4119 = ~n4116 & ~n4117;
  assign n4120 = ~n4118 & ~n4119;
  assign n4121 = n295 & ~n3628;
  assign n4122 = n2560 & ~n3280;
  assign n4123 = n2567 & n3272;
  assign n4124 = ~n4122 & ~n4123;
  assign n4125 = ~n4121 & n4124;
  assign n4126 = ~n2571 & n4125;
  assign n4127 = ~n3641 & n4125;
  assign n4128 = ~n4126 & ~n4127;
  assign n4129 = n275 & ~n4128;
  assign n4130 = ~n275 & n4128;
  assign n4131 = ~n4129 & ~n4130;
  assign n4132 = n4120 & n4131;
  assign n4133 = n4120 & ~n4132;
  assign n4134 = n4131 & ~n4132;
  assign n4135 = ~n4133 & ~n4134;
  assign n4136 = ~n4063 & ~n4135;
  assign n4137 = ~n4063 & ~n4136;
  assign n4138 = ~n4135 & ~n4136;
  assign n4139 = ~n4137 & ~n4138;
  assign n4140 = ~n4062 & ~n4139;
  assign n4141 = ~n4062 & ~n4140;
  assign n4142 = ~n4139 & ~n4140;
  assign n4143 = ~n4141 & ~n4142;
  assign n4144 = ~n4049 & n4143;
  assign n4145 = n4049 & ~n4143;
  assign n4146 = ~n4144 & ~n4145;
  assign n4147 = ~n4048 & ~n4146;
  assign n4148 = n4048 & n4146;
  assign n4149 = ~n4032 & ~n4148;
  assign n4150 = ~n4147 & n4149;
  assign n4151 = ~n4032 & ~n4150;
  assign n4152 = ~n4147 & ~n4150;
  assign n4153 = ~n4148 & n4152;
  assign n4154 = ~n4151 & ~n4153;
  assign n4155 = ~n4022 & n4154;
  assign n4156 = n4022 & ~n4154;
  assign n4157 = ~n4155 & ~n4156;
  assign n4158 = ~\sin[0]  & ~n4024;
  assign n4159 = ~n4027 & ~n4158;
  assign n4160 = ~n4157 & n4159;
  assign n4161 = n4157 & ~n4159;
  assign \sin[2]  = n4160 | n4161;
  assign n4163 = n2340 & n3657;
  assign n4164 = n397 & n4163;
  assign n4165 = n946 & n4164;
  assign n4166 = n2196 & n4165;
  assign n4167 = n1468 & n4166;
  assign n4168 = n735 & n4167;
  assign n4169 = n355 & n4168;
  assign n4170 = ~n317 & n4169;
  assign n4171 = ~n175 & n4170;
  assign n4172 = ~n370 & n4171;
  assign n4173 = ~n111 & n4172;
  assign n4174 = ~n258 & n4173;
  assign n4175 = ~n238 & n4174;
  assign n4176 = ~n4049 & ~n4143;
  assign n4177 = ~n4140 & ~n4176;
  assign n4178 = ~n4132 & ~n4136;
  assign n4179 = n3274 & n3896;
  assign n4180 = n3216 & n4054;
  assign n4181 = ~n4179 & ~n4180;
  assign n4182 = ~n291 & ~n4181;
  assign n4183 = ~n4181 & ~n4182;
  assign n4184 = ~n291 & ~n4182;
  assign n4185 = ~n4183 & ~n4184;
  assign n4186 = n2802 & ~n3280;
  assign n4187 = ~n2554 & n2808;
  assign n4188 = n2810 & n3277;
  assign n4189 = ~n4187 & ~n4188;
  assign n4190 = ~n4186 & n4189;
  assign n4191 = n2817 & n3318;
  assign n4192 = n4190 & ~n4191;
  assign n4193 = ~n1021 & ~n4192;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = ~n1021 & ~n4193;
  assign n4196 = ~n4194 & ~n4195;
  assign n4197 = ~n4105 & ~n4109;
  assign n4198 = ~n525 & n4085;
  assign n4199 = n2593 & n4198;
  assign n4200 = ~n4090 & ~n4199;
  assign n4201 = n2578 & n2668;
  assign n4202 = ~n2586 & n2776;
  assign n4203 = ~n2582 & n2666;
  assign n4204 = ~n4202 & ~n4203;
  assign n4205 = ~n4201 & n4204;
  assign n4206 = n2674 & n2815;
  assign n4207 = n4205 & ~n4206;
  assign n4208 = ~n525 & n2590;
  assign n4209 = ~n4207 & n4208;
  assign n4210 = n4207 & ~n4208;
  assign n4211 = ~n4209 & ~n4210;
  assign n4212 = ~n4200 & n4211;
  assign n4213 = ~n4200 & ~n4212;
  assign n4214 = n4211 & ~n4212;
  assign n4215 = ~n4213 & ~n4214;
  assign n4216 = ~n2566 & n2699;
  assign n4217 = ~n2575 & n2695;
  assign n4218 = n2562 & n2697;
  assign n4219 = ~n4217 & ~n4218;
  assign n4220 = ~n4216 & n4219;
  assign n4221 = ~n2690 & n4220;
  assign n4222 = ~n3022 & n4220;
  assign n4223 = ~n4221 & ~n4222;
  assign n4224 = n669 & ~n4223;
  assign n4225 = ~n669 & n4223;
  assign n4226 = ~n4224 & ~n4225;
  assign n4227 = ~n4215 & n4226;
  assign n4228 = n4215 & ~n4226;
  assign n4229 = ~n4227 & ~n4228;
  assign n4230 = ~n4197 & n4229;
  assign n4231 = n4197 & ~n4229;
  assign n4232 = ~n4230 & ~n4231;
  assign n4233 = ~n4196 & n4232;
  assign n4234 = ~n4196 & ~n4233;
  assign n4235 = n4232 & ~n4233;
  assign n4236 = ~n4234 & ~n4235;
  assign n4237 = ~n4113 & ~n4119;
  assign n4238 = n4236 & n4237;
  assign n4239 = ~n4236 & ~n4237;
  assign n4240 = ~n4238 & ~n4239;
  assign n4241 = n295 & n3750;
  assign n4242 = n2560 & n3272;
  assign n4243 = n2567 & ~n3628;
  assign n4244 = ~n4242 & ~n4243;
  assign n4245 = ~n4241 & n4244;
  assign n4246 = ~n2571 & n4245;
  assign n4247 = ~n3762 & n4245;
  assign n4248 = ~n4246 & ~n4247;
  assign n4249 = n275 & ~n4248;
  assign n4250 = ~n275 & n4248;
  assign n4251 = ~n4249 & ~n4250;
  assign n4252 = n4240 & n4251;
  assign n4253 = ~n4240 & ~n4251;
  assign n4254 = ~n4252 & ~n4253;
  assign n4255 = ~n4185 & n4254;
  assign n4256 = n4185 & ~n4254;
  assign n4257 = ~n4255 & ~n4256;
  assign n4258 = ~n4178 & n4257;
  assign n4259 = n4178 & ~n4257;
  assign n4260 = ~n4258 & ~n4259;
  assign n4261 = ~n4177 & n4260;
  assign n4262 = n4177 & ~n4260;
  assign n4263 = ~n4261 & ~n4262;
  assign n4264 = ~n4175 & n4263;
  assign n4265 = ~n4175 & ~n4264;
  assign n4266 = n4263 & ~n4264;
  assign n4267 = ~n4265 & ~n4266;
  assign n4268 = ~n4152 & ~n4267;
  assign n4269 = n4152 & ~n4266;
  assign n4270 = ~n4265 & n4269;
  assign n4271 = ~n4268 & ~n4270;
  assign n4272 = n4156 & n4271;
  assign n4273 = n4271 & ~n4272;
  assign n4274 = n4156 & ~n4272;
  assign n4275 = ~n4273 & ~n4274;
  assign n4276 = ~n4157 & n4158;
  assign n4277 = ~n4027 & ~n4276;
  assign n4278 = ~n4275 & n4277;
  assign n4279 = n4275 & ~n4277;
  assign \sin[3]  = ~n4278 & ~n4279;
  assign n4281 = ~n4264 & ~n4268;
  assign n4282 = n346 & n496;
  assign n4283 = n301 & n4282;
  assign n4284 = n2464 & n4283;
  assign n4285 = n975 & n4284;
  assign n4286 = n752 & n4285;
  assign n4287 = n644 & n4286;
  assign n4288 = n2418 & n4287;
  assign n4289 = ~n178 & n4288;
  assign n4290 = ~n194 & n4289;
  assign n4291 = ~n589 & n4290;
  assign n4292 = ~n4258 & ~n4261;
  assign n4293 = ~n4252 & ~n4255;
  assign n4294 = ~n4233 & ~n4239;
  assign n4295 = ~n4227 & ~n4230;
  assign n4296 = ~n2575 & n2668;
  assign n4297 = ~n2582 & n2776;
  assign n4298 = n2578 & n2666;
  assign n4299 = ~n4297 & ~n4298;
  assign n4300 = ~n4296 & n4299;
  assign n4301 = n2674 & n2989;
  assign n4302 = n4300 & ~n4301;
  assign n4303 = ~n525 & ~n4302;
  assign n4304 = ~n4302 & ~n4303;
  assign n4305 = ~n525 & ~n4303;
  assign n4306 = ~n4304 & ~n4305;
  assign n4307 = ~n291 & ~n525;
  assign n4308 = ~n2586 & n4307;
  assign n4309 = ~n291 & ~n4308;
  assign n4310 = ~n2586 & ~n4308;
  assign n4311 = ~n525 & n4310;
  assign n4312 = ~n4309 & ~n4311;
  assign n4313 = ~n4306 & ~n4312;
  assign n4314 = ~n4306 & ~n4313;
  assign n4315 = ~n4312 & ~n4313;
  assign n4316 = ~n4314 & ~n4315;
  assign n4317 = ~n525 & ~n2590;
  assign n4318 = n4207 & n4317;
  assign n4319 = ~n4212 & ~n4318;
  assign n4320 = n4316 & ~n4319;
  assign n4321 = ~n4316 & n4319;
  assign n4322 = ~n4320 & ~n4321;
  assign n4323 = ~n2554 & n2699;
  assign n4324 = n2562 & n2695;
  assign n4325 = ~n2566 & n2697;
  assign n4326 = ~n4324 & ~n4325;
  assign n4327 = ~n4323 & n4326;
  assign n4328 = n2652 & n2690;
  assign n4329 = n4327 & ~n4328;
  assign n4330 = ~n669 & ~n4329;
  assign n4331 = n669 & n4329;
  assign n4332 = ~n4330 & ~n4331;
  assign n4333 = ~n4322 & n4332;
  assign n4334 = ~n4322 & ~n4333;
  assign n4335 = n4332 & ~n4333;
  assign n4336 = ~n4334 & ~n4335;
  assign n4337 = ~n4295 & n4336;
  assign n4338 = n4295 & ~n4336;
  assign n4339 = ~n4337 & ~n4338;
  assign n4340 = n2802 & n3272;
  assign n4341 = n2808 & n3277;
  assign n4342 = n2810 & ~n3280;
  assign n4343 = ~n4341 & ~n4342;
  assign n4344 = ~n4340 & n4343;
  assign n4345 = n2817 & n3302;
  assign n4346 = n4344 & ~n4345;
  assign n4347 = ~n1021 & ~n4346;
  assign n4348 = ~n1021 & ~n4347;
  assign n4349 = ~n4346 & ~n4347;
  assign n4350 = ~n4348 & ~n4349;
  assign n4351 = ~n4339 & ~n4350;
  assign n4352 = n4339 & n4350;
  assign n4353 = ~n4351 & ~n4352;
  assign n4354 = ~n4294 & n4353;
  assign n4355 = n4294 & ~n4353;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = n295 & n3896;
  assign n4358 = n2560 & ~n3628;
  assign n4359 = n2567 & n3750;
  assign n4360 = ~n4358 & ~n4359;
  assign n4361 = ~n4357 & n4360;
  assign n4362 = n2571 & n3908;
  assign n4363 = n4361 & ~n4362;
  assign n4364 = ~n275 & ~n4363;
  assign n4365 = n275 & n4363;
  assign n4366 = ~n4364 & ~n4365;
  assign n4367 = n4356 & n4366;
  assign n4368 = ~n4356 & ~n4366;
  assign n4369 = ~n4367 & ~n4368;
  assign n4370 = ~n4293 & n4369;
  assign n4371 = n4293 & ~n4369;
  assign n4372 = ~n4370 & ~n4371;
  assign n4373 = n4292 & ~n4372;
  assign n4374 = ~n4292 & n4372;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = n4291 & ~n4375;
  assign n4377 = ~n4291 & n4375;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = ~n4281 & n4378;
  assign n4380 = n4281 & ~n4378;
  assign n4381 = ~n4379 & ~n4380;
  assign n4382 = ~n4272 & ~n4381;
  assign n4383 = n4272 & n4381;
  assign n4384 = ~n4382 & ~n4383;
  assign n4385 = n4275 & n4276;
  assign n4386 = ~n4027 & ~n4385;
  assign n4387 = ~n4384 & n4386;
  assign n4388 = n4384 & ~n4386;
  assign \sin[4]  = n4387 | n4388;
  assign n4390 = ~n4377 & ~n4379;
  assign n4391 = ~n317 & ~n359;
  assign n4392 = ~n472 & n4391;
  assign n4393 = n189 & n807;
  assign n4394 = n4392 & n4393;
  assign n4395 = n2317 & n4394;
  assign n4396 = n314 & n4395;
  assign n4397 = n3883 & n4396;
  assign n4398 = n3243 & n4397;
  assign n4399 = n4002 & n4398;
  assign n4400 = n369 & n4399;
  assign n4401 = ~n178 & n4400;
  assign n4402 = ~n417 & n4401;
  assign n4403 = ~n299 & n4402;
  assign n4404 = ~n237 & n4403;
  assign n4405 = ~n4370 & ~n4374;
  assign n4406 = ~n4354 & ~n4367;
  assign n4407 = ~n4295 & ~n4336;
  assign n4408 = ~n4351 & ~n4407;
  assign n4409 = n2802 & ~n3628;
  assign n4410 = n2808 & ~n3280;
  assign n4411 = n2810 & n3272;
  assign n4412 = ~n4410 & ~n4411;
  assign n4413 = ~n4409 & n4412;
  assign n4414 = n2817 & n3641;
  assign n4415 = n4413 & ~n4414;
  assign n4416 = ~n1021 & ~n4415;
  assign n4417 = ~n4415 & ~n4416;
  assign n4418 = ~n1021 & ~n4416;
  assign n4419 = ~n4417 & ~n4418;
  assign n4420 = ~n4316 & ~n4319;
  assign n4421 = ~n4333 & ~n4420;
  assign n4422 = ~n4308 & ~n4313;
  assign n4423 = ~n2582 & n4307;
  assign n4424 = ~n291 & ~n4423;
  assign n4425 = ~n2582 & ~n4423;
  assign n4426 = ~n525 & n4425;
  assign n4427 = ~n4424 & ~n4426;
  assign n4428 = ~n4422 & ~n4427;
  assign n4429 = ~n4422 & ~n4428;
  assign n4430 = ~n4427 & ~n4428;
  assign n4431 = ~n4429 & ~n4430;
  assign n4432 = n2562 & n2668;
  assign n4433 = n2578 & n2776;
  assign n4434 = ~n2575 & n2666;
  assign n4435 = ~n4433 & ~n4434;
  assign n4436 = ~n4432 & n4435;
  assign n4437 = ~n2674 & n4436;
  assign n4438 = ~n3042 & n4436;
  assign n4439 = ~n4437 & ~n4438;
  assign n4440 = n525 & ~n4439;
  assign n4441 = ~n525 & n4439;
  assign n4442 = ~n4440 & ~n4441;
  assign n4443 = ~n4431 & n4442;
  assign n4444 = ~n4431 & ~n4443;
  assign n4445 = n4442 & ~n4443;
  assign n4446 = ~n4444 & ~n4445;
  assign n4447 = n2699 & n3277;
  assign n4448 = ~n2566 & n2695;
  assign n4449 = ~n2554 & n2697;
  assign n4450 = ~n4448 & ~n4449;
  assign n4451 = ~n4447 & n4450;
  assign n4452 = n2690 & n3332;
  assign n4453 = n4451 & ~n4452;
  assign n4454 = ~n669 & ~n4453;
  assign n4455 = n669 & n4453;
  assign n4456 = ~n4454 & ~n4455;
  assign n4457 = ~n4446 & n4456;
  assign n4458 = ~n4445 & ~n4456;
  assign n4459 = ~n4444 & n4458;
  assign n4460 = ~n4457 & ~n4459;
  assign n4461 = ~n4421 & n4460;
  assign n4462 = ~n4421 & ~n4461;
  assign n4463 = n4460 & ~n4461;
  assign n4464 = ~n4462 & ~n4463;
  assign n4465 = ~n4419 & ~n4464;
  assign n4466 = n4419 & ~n4463;
  assign n4467 = ~n4462 & n4466;
  assign n4468 = ~n4465 & ~n4467;
  assign n4469 = ~n4408 & n4468;
  assign n4470 = ~n4408 & ~n4469;
  assign n4471 = n4468 & ~n4469;
  assign n4472 = ~n4470 & ~n4471;
  assign n4473 = n2560 & n3750;
  assign n4474 = n2567 & n3896;
  assign n4475 = ~n4473 & ~n4474;
  assign n4476 = n2571 & n4056;
  assign n4477 = n4475 & ~n4476;
  assign n4478 = ~n275 & ~n4477;
  assign n4479 = n275 & n4477;
  assign n4480 = ~n4478 & ~n4479;
  assign n4481 = ~n4472 & n4480;
  assign n4482 = ~n4471 & ~n4480;
  assign n4483 = ~n4470 & n4482;
  assign n4484 = ~n4481 & ~n4483;
  assign n4485 = ~n4406 & n4484;
  assign n4486 = n4406 & ~n4484;
  assign n4487 = ~n4485 & ~n4486;
  assign n4488 = ~n4405 & n4487;
  assign n4489 = n4405 & ~n4487;
  assign n4490 = ~n4488 & ~n4489;
  assign n4491 = n4404 & ~n4490;
  assign n4492 = ~n4404 & n4490;
  assign n4493 = ~n4491 & ~n4492;
  assign n4494 = ~n4390 & n4493;
  assign n4495 = n4390 & ~n4493;
  assign n4496 = ~n4494 & ~n4495;
  assign n4497 = ~n4383 & ~n4496;
  assign n4498 = n4383 & n4496;
  assign n4499 = ~n4497 & ~n4498;
  assign n4500 = ~n4384 & n4385;
  assign n4501 = ~n4027 & ~n4500;
  assign n4502 = ~n4499 & n4501;
  assign n4503 = n4499 & ~n4501;
  assign \sin[5]  = n4502 | n4503;
  assign n4505 = ~n4492 & ~n4494;
  assign n4506 = n316 & n1117;
  assign n4507 = n586 & n4506;
  assign n4508 = n2421 & n4507;
  assign n4509 = n2340 & n4508;
  assign n4510 = n156 & n4509;
  assign n4511 = n369 & n4510;
  assign n4512 = n976 & n4511;
  assign n4513 = ~n357 & n4512;
  assign n4514 = n253 & n970;
  assign n4515 = n2458 & n4514;
  assign n4516 = n3259 & n4515;
  assign n4517 = n4513 & n4516;
  assign n4518 = ~n337 & n4517;
  assign n4519 = ~n150 & n4518;
  assign n4520 = ~n172 & n4519;
  assign n4521 = ~n169 & n4520;
  assign n4522 = ~n447 & n4521;
  assign n4523 = ~n148 & n4522;
  assign n4524 = ~n4485 & ~n4488;
  assign n4525 = ~n4469 & ~n4481;
  assign n4526 = ~n4461 & ~n4465;
  assign n4527 = n2560 & n3896;
  assign n4528 = n2571 & n4054;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = n275 & ~n4529;
  assign n4531 = ~n275 & n4529;
  assign n4532 = ~n4530 & ~n4531;
  assign n4533 = ~n4526 & ~n4532;
  assign n4534 = n4526 & n4532;
  assign n4535 = ~n4533 & ~n4534;
  assign n4536 = n2802 & n3750;
  assign n4537 = n2808 & n3272;
  assign n4538 = n2810 & ~n3628;
  assign n4539 = ~n4537 & ~n4538;
  assign n4540 = ~n4536 & n4539;
  assign n4541 = n2817 & n3762;
  assign n4542 = n4540 & ~n4541;
  assign n4543 = ~n1021 & ~n4542;
  assign n4544 = ~n4542 & ~n4543;
  assign n4545 = ~n1021 & ~n4543;
  assign n4546 = ~n4544 & ~n4545;
  assign n4547 = ~n4443 & ~n4457;
  assign n4548 = ~n4423 & ~n4428;
  assign n4549 = n2578 & n4307;
  assign n4550 = ~n291 & ~n4549;
  assign n4551 = n2578 & ~n4549;
  assign n4552 = ~n525 & n4551;
  assign n4553 = ~n4550 & ~n4552;
  assign n4554 = ~n4548 & ~n4553;
  assign n4555 = ~n4548 & ~n4554;
  assign n4556 = ~n4553 & ~n4554;
  assign n4557 = ~n4555 & ~n4556;
  assign n4558 = ~n2566 & n2668;
  assign n4559 = ~n2575 & n2776;
  assign n4560 = n2562 & n2666;
  assign n4561 = ~n4559 & ~n4560;
  assign n4562 = ~n4558 & n4561;
  assign n4563 = ~n2674 & n4562;
  assign n4564 = ~n3022 & n4562;
  assign n4565 = ~n4563 & ~n4564;
  assign n4566 = n525 & ~n4565;
  assign n4567 = ~n525 & n4565;
  assign n4568 = ~n4566 & ~n4567;
  assign n4569 = ~n4557 & n4568;
  assign n4570 = ~n4557 & ~n4569;
  assign n4571 = n4568 & ~n4569;
  assign n4572 = ~n4570 & ~n4571;
  assign n4573 = n2699 & ~n3280;
  assign n4574 = ~n2554 & n2695;
  assign n4575 = n2697 & n3277;
  assign n4576 = ~n4574 & ~n4575;
  assign n4577 = ~n4573 & n4576;
  assign n4578 = n2690 & n3318;
  assign n4579 = n4577 & ~n4578;
  assign n4580 = ~n669 & ~n4579;
  assign n4581 = n669 & n4579;
  assign n4582 = ~n4580 & ~n4581;
  assign n4583 = ~n4572 & n4582;
  assign n4584 = ~n4571 & ~n4582;
  assign n4585 = ~n4570 & n4584;
  assign n4586 = ~n4583 & ~n4585;
  assign n4587 = ~n4547 & n4586;
  assign n4588 = ~n4547 & ~n4587;
  assign n4589 = n4586 & ~n4587;
  assign n4590 = ~n4588 & ~n4589;
  assign n4591 = ~n4546 & ~n4590;
  assign n4592 = n4546 & ~n4589;
  assign n4593 = ~n4588 & n4592;
  assign n4594 = ~n4591 & ~n4593;
  assign n4595 = n4535 & n4594;
  assign n4596 = ~n4535 & ~n4594;
  assign n4597 = ~n4595 & ~n4596;
  assign n4598 = ~n4525 & n4597;
  assign n4599 = n4525 & ~n4597;
  assign n4600 = ~n4598 & ~n4599;
  assign n4601 = ~n4524 & n4600;
  assign n4602 = n4524 & ~n4600;
  assign n4603 = ~n4601 & ~n4602;
  assign n4604 = n4523 & ~n4603;
  assign n4605 = ~n4523 & n4603;
  assign n4606 = ~n4604 & ~n4605;
  assign n4607 = ~n4505 & n4606;
  assign n4608 = n4505 & ~n4606;
  assign n4609 = ~n4607 & ~n4608;
  assign n4610 = ~n4498 & ~n4609;
  assign n4611 = n4498 & n4609;
  assign n4612 = ~n4610 & ~n4611;
  assign n4613 = ~n4499 & n4500;
  assign n4614 = ~n4027 & ~n4613;
  assign n4615 = ~n4612 & n4614;
  assign n4616 = n4612 & ~n4614;
  assign \sin[6]  = n4615 | n4616;
  assign n4618 = ~n4605 & ~n4607;
  assign n4619 = ~n4533 & ~n4595;
  assign n4620 = ~n4587 & ~n4591;
  assign n4621 = n2802 & n3896;
  assign n4622 = n2808 & ~n3628;
  assign n4623 = n2810 & n3750;
  assign n4624 = ~n4622 & ~n4623;
  assign n4625 = ~n4621 & n4624;
  assign n4626 = ~n3908 & n4625;
  assign n4627 = ~n2817 & n4625;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = n1021 & ~n4628;
  assign n4630 = ~n1021 & n4628;
  assign n4631 = ~n4629 & ~n4630;
  assign n4632 = ~n4620 & n4631;
  assign n4633 = n4620 & ~n4631;
  assign n4634 = ~n4632 & ~n4633;
  assign n4635 = ~n4569 & ~n4583;
  assign n4636 = ~n4549 & ~n4554;
  assign n4637 = ~n2554 & n2668;
  assign n4638 = n2562 & n2776;
  assign n4639 = ~n2566 & n2666;
  assign n4640 = ~n4638 & ~n4639;
  assign n4641 = ~n4637 & n4640;
  assign n4642 = n2652 & n2674;
  assign n4643 = n4641 & ~n4642;
  assign n4644 = ~n525 & ~n4643;
  assign n4645 = ~n4643 & ~n4644;
  assign n4646 = ~n525 & ~n4644;
  assign n4647 = ~n4645 & ~n4646;
  assign n4648 = ~n525 & ~n2575;
  assign n4649 = n275 & n291;
  assign n4650 = ~n275 & ~n291;
  assign n4651 = ~n4649 & ~n4650;
  assign n4652 = n4648 & n4651;
  assign n4653 = ~n4648 & ~n4651;
  assign n4654 = ~n4652 & ~n4653;
  assign n4655 = ~n4647 & n4654;
  assign n4656 = ~n4647 & ~n4655;
  assign n4657 = n4654 & ~n4655;
  assign n4658 = ~n4656 & ~n4657;
  assign n4659 = ~n4636 & n4658;
  assign n4660 = n4636 & ~n4658;
  assign n4661 = ~n4659 & ~n4660;
  assign n4662 = n2699 & n3272;
  assign n4663 = n2695 & n3277;
  assign n4664 = n2697 & ~n3280;
  assign n4665 = ~n4663 & ~n4664;
  assign n4666 = ~n4662 & n4665;
  assign n4667 = ~n2690 & n4666;
  assign n4668 = ~n3302 & n4666;
  assign n4669 = ~n4667 & ~n4668;
  assign n4670 = n669 & ~n4669;
  assign n4671 = ~n669 & n4669;
  assign n4672 = ~n4670 & ~n4671;
  assign n4673 = ~n4661 & n4672;
  assign n4674 = ~n4661 & ~n4673;
  assign n4675 = n4672 & ~n4673;
  assign n4676 = ~n4674 & ~n4675;
  assign n4677 = ~n4635 & ~n4676;
  assign n4678 = ~n4635 & ~n4677;
  assign n4679 = ~n4676 & ~n4677;
  assign n4680 = ~n4678 & ~n4679;
  assign n4681 = n4634 & ~n4680;
  assign n4682 = n4634 & ~n4681;
  assign n4683 = ~n4680 & ~n4681;
  assign n4684 = ~n4682 & ~n4683;
  assign n4685 = ~n4619 & n4684;
  assign n4686 = n4619 & ~n4684;
  assign n4687 = ~n4685 & ~n4686;
  assign n4688 = ~n4598 & ~n4601;
  assign n4689 = n4687 & n4688;
  assign n4690 = ~n4687 & ~n4688;
  assign n4691 = ~n4689 & ~n4690;
  assign n4692 = n931 & n2281;
  assign n4693 = n4392 & n4692;
  assign n4694 = n809 & n4693;
  assign n4695 = n4513 & n4694;
  assign n4696 = ~n129 & n4695;
  assign n4697 = ~n194 & n4696;
  assign n4698 = ~n137 & n4697;
  assign n4699 = ~n218 & n4698;
  assign n4700 = n1090 & n4699;
  assign n4701 = ~n168 & n4700;
  assign n4702 = ~n445 & n4701;
  assign n4703 = n4691 & ~n4702;
  assign n4704 = ~n4691 & n4702;
  assign n4705 = ~n4703 & ~n4704;
  assign n4706 = ~n4618 & n4705;
  assign n4707 = n4618 & ~n4705;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = n4611 & n4708;
  assign n4710 = ~n4611 & ~n4708;
  assign n4711 = ~n4709 & ~n4710;
  assign n4712 = ~n4612 & n4613;
  assign n4713 = ~n4027 & ~n4712;
  assign n4714 = ~n4711 & n4713;
  assign n4715 = n4711 & ~n4713;
  assign \sin[7]  = n4714 | n4715;
  assign n4717 = ~n4703 & ~n4706;
  assign n4718 = n609 & n2181;
  assign n4719 = n165 & n4718;
  assign n4720 = ~n221 & n4719;
  assign n4721 = ~n219 & n4720;
  assign n4722 = ~n167 & n4721;
  assign n4723 = ~n225 & n4722;
  assign n4724 = ~n446 & n4723;
  assign n4725 = ~n111 & n4724;
  assign n4726 = ~n211 & n4725;
  assign n4727 = n961 & n2342;
  assign n4728 = n979 & n4727;
  assign n4729 = n3678 & n4728;
  assign n4730 = n4726 & n4729;
  assign n4731 = ~n408 & n4730;
  assign n4732 = ~n257 & n4731;
  assign n4733 = ~n207 & n4732;
  assign n4734 = ~n361 & n4733;
  assign n4735 = ~n224 & n4734;
  assign n4736 = ~n326 & n4735;
  assign n4737 = ~n469 & n4736;
  assign n4738 = ~n4619 & ~n4684;
  assign n4739 = ~n4690 & ~n4738;
  assign n4740 = ~n4632 & ~n4681;
  assign n4741 = n2808 & n3750;
  assign n4742 = n2810 & n3896;
  assign n4743 = ~n4741 & ~n4742;
  assign n4744 = n2817 & n4056;
  assign n4745 = n4743 & ~n4744;
  assign n4746 = ~n1021 & ~n4745;
  assign n4747 = ~n4745 & ~n4746;
  assign n4748 = ~n1021 & ~n4746;
  assign n4749 = ~n4747 & ~n4748;
  assign n4750 = ~n4673 & ~n4677;
  assign n4751 = ~n4636 & ~n4658;
  assign n4752 = ~n4655 & ~n4751;
  assign n4753 = ~n525 & n2562;
  assign n4754 = ~n4649 & ~n4652;
  assign n4755 = ~n4753 & ~n4754;
  assign n4756 = ~n4753 & ~n4755;
  assign n4757 = ~n4754 & ~n4755;
  assign n4758 = ~n4756 & ~n4757;
  assign n4759 = n2668 & n3277;
  assign n4760 = ~n2566 & n2776;
  assign n4761 = ~n2554 & n2666;
  assign n4762 = ~n4760 & ~n4761;
  assign n4763 = ~n4759 & n4762;
  assign n4764 = ~n2674 & n4763;
  assign n4765 = ~n3332 & n4763;
  assign n4766 = ~n4764 & ~n4765;
  assign n4767 = n525 & ~n4766;
  assign n4768 = ~n525 & n4766;
  assign n4769 = ~n4767 & ~n4768;
  assign n4770 = ~n4758 & n4769;
  assign n4771 = n4758 & ~n4769;
  assign n4772 = ~n4770 & ~n4771;
  assign n4773 = ~n4752 & n4772;
  assign n4774 = ~n4752 & ~n4773;
  assign n4775 = n4772 & ~n4773;
  assign n4776 = ~n4774 & ~n4775;
  assign n4777 = n2699 & ~n3628;
  assign n4778 = n2695 & ~n3280;
  assign n4779 = n2697 & n3272;
  assign n4780 = ~n4778 & ~n4779;
  assign n4781 = ~n4777 & n4780;
  assign n4782 = n2690 & n3641;
  assign n4783 = n4781 & ~n4782;
  assign n4784 = ~n669 & ~n4783;
  assign n4785 = n669 & n4783;
  assign n4786 = ~n4784 & ~n4785;
  assign n4787 = ~n4776 & n4786;
  assign n4788 = ~n4775 & ~n4786;
  assign n4789 = ~n4774 & n4788;
  assign n4790 = ~n4787 & ~n4789;
  assign n4791 = ~n4750 & n4790;
  assign n4792 = n4750 & ~n4790;
  assign n4793 = ~n4791 & ~n4792;
  assign n4794 = ~n4749 & n4793;
  assign n4795 = n4749 & ~n4793;
  assign n4796 = ~n4794 & ~n4795;
  assign n4797 = ~n4740 & n4796;
  assign n4798 = n4740 & ~n4796;
  assign n4799 = ~n4797 & ~n4798;
  assign n4800 = ~n4739 & n4799;
  assign n4801 = n4739 & ~n4799;
  assign n4802 = ~n4800 & ~n4801;
  assign n4803 = n4737 & ~n4802;
  assign n4804 = ~n4737 & n4802;
  assign n4805 = ~n4803 & ~n4804;
  assign n4806 = ~n4717 & n4805;
  assign n4807 = n4717 & ~n4805;
  assign n4808 = ~n4806 & ~n4807;
  assign n4809 = ~n4709 & ~n4808;
  assign n4810 = n4709 & n4808;
  assign n4811 = ~n4809 & ~n4810;
  assign n4812 = ~n4711 & n4712;
  assign n4813 = ~n4027 & ~n4812;
  assign n4814 = ~n4811 & n4813;
  assign n4815 = n4811 & ~n4813;
  assign \sin[8]  = n4814 | n4815;
  assign n4817 = ~n4804 & ~n4806;
  assign n4818 = n757 & n809;
  assign n4819 = n204 & n4818;
  assign n4820 = n3231 & n4819;
  assign n4821 = n2432 & n4820;
  assign n4822 = n3259 & n4821;
  assign n4823 = ~n337 & n4822;
  assign n4824 = ~n327 & n4823;
  assign n4825 = ~n225 & n4824;
  assign n4826 = ~n133 & n4825;
  assign n4827 = ~n234 & n4826;
  assign n4828 = ~n356 & n4827;
  assign n4829 = ~n216 & n4828;
  assign n4830 = ~n4791 & ~n4794;
  assign n4831 = ~n4755 & ~n4770;
  assign n4832 = n2668 & ~n3280;
  assign n4833 = ~n2554 & n2776;
  assign n4834 = n2666 & n3277;
  assign n4835 = ~n4833 & ~n4834;
  assign n4836 = ~n4832 & n4835;
  assign n4837 = n2674 & n3318;
  assign n4838 = n4836 & ~n4837;
  assign n4839 = ~n525 & ~n4838;
  assign n4840 = ~n4838 & ~n4839;
  assign n4841 = ~n525 & ~n4839;
  assign n4842 = ~n4840 & ~n4841;
  assign n4843 = ~n525 & n2644;
  assign n4844 = ~n4842 & ~n4843;
  assign n4845 = ~n4842 & ~n4844;
  assign n4846 = ~n4843 & ~n4844;
  assign n4847 = ~n4845 & ~n4846;
  assign n4848 = ~n4831 & n4847;
  assign n4849 = n4831 & ~n4847;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = n2699 & n3750;
  assign n4852 = n2695 & n3272;
  assign n4853 = n2697 & ~n3628;
  assign n4854 = ~n4852 & ~n4853;
  assign n4855 = ~n4851 & n4854;
  assign n4856 = n2690 & n3762;
  assign n4857 = n4855 & ~n4856;
  assign n4858 = ~n669 & ~n4857;
  assign n4859 = n669 & n4857;
  assign n4860 = ~n4858 & ~n4859;
  assign n4861 = ~n4850 & n4860;
  assign n4862 = ~n4850 & ~n4861;
  assign n4863 = n4860 & ~n4861;
  assign n4864 = ~n4862 & ~n4863;
  assign n4865 = ~n4773 & ~n4787;
  assign n4866 = n2808 & n3896;
  assign n4867 = n2817 & n4054;
  assign n4868 = ~n4866 & ~n4867;
  assign n4869 = ~n1021 & n4868;
  assign n4870 = n1021 & ~n4868;
  assign n4871 = ~n4869 & ~n4870;
  assign n4872 = ~n4865 & ~n4871;
  assign n4873 = n4865 & n4871;
  assign n4874 = ~n4872 & ~n4873;
  assign n4875 = ~n4864 & n4874;
  assign n4876 = ~n4864 & ~n4875;
  assign n4877 = n4874 & ~n4875;
  assign n4878 = ~n4876 & ~n4877;
  assign n4879 = ~n4830 & n4878;
  assign n4880 = n4830 & ~n4878;
  assign n4881 = ~n4879 & ~n4880;
  assign n4882 = ~n4797 & ~n4800;
  assign n4883 = n4881 & n4882;
  assign n4884 = ~n4881 & ~n4882;
  assign n4885 = ~n4883 & ~n4884;
  assign n4886 = n4829 & ~n4885;
  assign n4887 = ~n4829 & n4885;
  assign n4888 = ~n4886 & ~n4887;
  assign n4889 = ~n4817 & n4888;
  assign n4890 = n4817 & ~n4888;
  assign n4891 = ~n4889 & ~n4890;
  assign n4892 = ~n4810 & ~n4891;
  assign n4893 = n4810 & n4891;
  assign n4894 = ~n4892 & ~n4893;
  assign n4895 = ~n4811 & n4812;
  assign n4896 = ~n4027 & ~n4895;
  assign n4897 = ~n4894 & n4896;
  assign n4898 = n4894 & ~n4896;
  assign \sin[9]  = n4897 | n4898;
  assign n4900 = ~n4887 & ~n4889;
  assign n4901 = n259 & n655;
  assign n4902 = n476 & n4901;
  assign n4903 = n505 & n4902;
  assign n4904 = n210 & n4903;
  assign n4905 = n3666 & n4904;
  assign n4906 = n1104 & n4905;
  assign n4907 = n3259 & n4906;
  assign n4908 = n977 & n4907;
  assign n4909 = ~n312 & n4908;
  assign n4910 = ~n192 & n4909;
  assign n4911 = ~n315 & n4910;
  assign n4912 = ~n4830 & ~n4878;
  assign n4913 = ~n4884 & ~n4912;
  assign n4914 = ~n4872 & ~n4875;
  assign n4915 = ~n2566 & ~n4753;
  assign n4916 = ~n525 & n4915;
  assign n4917 = ~n4844 & ~n4916;
  assign n4918 = ~n525 & ~n2554;
  assign n4919 = ~n1021 & ~n4918;
  assign n4920 = n1021 & n4918;
  assign n4921 = n4753 & ~n4920;
  assign n4922 = ~n4919 & n4921;
  assign n4923 = n4753 & ~n4922;
  assign n4924 = ~n4920 & ~n4922;
  assign n4925 = ~n4919 & n4924;
  assign n4926 = ~n4923 & ~n4925;
  assign n4927 = ~n4917 & ~n4926;
  assign n4928 = ~n4917 & ~n4927;
  assign n4929 = ~n4926 & ~n4927;
  assign n4930 = ~n4928 & ~n4929;
  assign n4931 = n2668 & n3272;
  assign n4932 = n2776 & n3277;
  assign n4933 = n2666 & ~n3280;
  assign n4934 = ~n4932 & ~n4933;
  assign n4935 = ~n4931 & n4934;
  assign n4936 = n2674 & n3302;
  assign n4937 = n4935 & ~n4936;
  assign n4938 = ~n525 & ~n4937;
  assign n4939 = ~n525 & ~n4938;
  assign n4940 = ~n4937 & ~n4938;
  assign n4941 = ~n4939 & ~n4940;
  assign n4942 = ~n4930 & ~n4941;
  assign n4943 = ~n4930 & ~n4942;
  assign n4944 = ~n4941 & ~n4942;
  assign n4945 = ~n4943 & ~n4944;
  assign n4946 = ~n4831 & ~n4847;
  assign n4947 = ~n4861 & ~n4946;
  assign n4948 = n2699 & n3896;
  assign n4949 = n2695 & ~n3628;
  assign n4950 = n2697 & n3750;
  assign n4951 = ~n4949 & ~n4950;
  assign n4952 = ~n4948 & n4951;
  assign n4953 = ~n2690 & n4952;
  assign n4954 = ~n3908 & n4952;
  assign n4955 = ~n4953 & ~n4954;
  assign n4956 = n669 & ~n4955;
  assign n4957 = ~n669 & n4955;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = ~n4947 & n4958;
  assign n4960 = ~n4947 & ~n4959;
  assign n4961 = n4958 & ~n4959;
  assign n4962 = ~n4960 & ~n4961;
  assign n4963 = ~n4945 & ~n4962;
  assign n4964 = n4945 & ~n4961;
  assign n4965 = ~n4960 & n4964;
  assign n4966 = ~n4963 & ~n4965;
  assign n4967 = ~n4914 & n4966;
  assign n4968 = n4914 & ~n4966;
  assign n4969 = ~n4967 & ~n4968;
  assign n4970 = ~n4913 & n4969;
  assign n4971 = n4913 & ~n4969;
  assign n4972 = ~n4970 & ~n4971;
  assign n4973 = n4911 & ~n4972;
  assign n4974 = ~n4911 & n4972;
  assign n4975 = ~n4973 & ~n4974;
  assign n4976 = ~n4900 & n4975;
  assign n4977 = n4900 & ~n4975;
  assign n4978 = ~n4976 & ~n4977;
  assign n4979 = ~n4893 & ~n4978;
  assign n4980 = n4893 & n4978;
  assign n4981 = ~n4979 & ~n4980;
  assign n4982 = ~n4894 & n4895;
  assign n4983 = ~n4027 & ~n4982;
  assign n4984 = ~n4981 & n4983;
  assign n4985 = n4981 & ~n4983;
  assign \sin[10]  = n4984 | n4985;
  assign n4987 = ~n4974 & ~n4976;
  assign n4988 = n911 & n969;
  assign n4989 = n499 & n4988;
  assign n4990 = n3734 & n4989;
  assign n4991 = n636 & n4990;
  assign n4992 = n453 & n4991;
  assign n4993 = ~n336 & n4992;
  assign n4994 = ~n4967 & ~n4970;
  assign n4995 = ~n4959 & ~n4963;
  assign n4996 = ~n4927 & ~n4942;
  assign n4997 = ~n525 & n3277;
  assign n4998 = ~n4924 & n4997;
  assign n4999 = n4924 & ~n4997;
  assign n5000 = ~n4998 & ~n4999;
  assign n5001 = n2668 & ~n3628;
  assign n5002 = n2776 & ~n3280;
  assign n5003 = n2666 & n3272;
  assign n5004 = ~n5002 & ~n5003;
  assign n5005 = ~n5001 & n5004;
  assign n5006 = ~n2674 & n5005;
  assign n5007 = ~n3641 & n5005;
  assign n5008 = ~n5006 & ~n5007;
  assign n5009 = n525 & ~n5008;
  assign n5010 = ~n525 & n5008;
  assign n5011 = ~n5009 & ~n5010;
  assign n5012 = ~n5000 & n5011;
  assign n5013 = n5000 & ~n5011;
  assign n5014 = ~n5012 & ~n5013;
  assign n5015 = ~n4996 & n5014;
  assign n5016 = ~n4996 & ~n5015;
  assign n5017 = n5014 & ~n5015;
  assign n5018 = ~n5016 & ~n5017;
  assign n5019 = n2695 & n3750;
  assign n5020 = n2697 & n3896;
  assign n5021 = ~n5019 & ~n5020;
  assign n5022 = n2690 & n4056;
  assign n5023 = n5021 & ~n5022;
  assign n5024 = ~n669 & ~n5023;
  assign n5025 = n669 & n5023;
  assign n5026 = ~n5024 & ~n5025;
  assign n5027 = ~n5018 & n5026;
  assign n5028 = ~n5017 & ~n5026;
  assign n5029 = ~n5016 & n5028;
  assign n5030 = ~n5027 & ~n5029;
  assign n5031 = ~n4995 & n5030;
  assign n5032 = n4995 & ~n5030;
  assign n5033 = ~n5031 & ~n5032;
  assign n5034 = ~n4994 & n5033;
  assign n5035 = n4994 & ~n5033;
  assign n5036 = ~n5034 & ~n5035;
  assign n5037 = n4993 & ~n5036;
  assign n5038 = ~n4993 & n5036;
  assign n5039 = ~n5037 & ~n5038;
  assign n5040 = ~n4987 & n5039;
  assign n5041 = n4987 & ~n5039;
  assign n5042 = ~n5040 & ~n5041;
  assign n5043 = ~n4980 & ~n5042;
  assign n5044 = n4980 & n5042;
  assign n5045 = ~n5043 & ~n5044;
  assign n5046 = ~n4981 & n4982;
  assign n5047 = ~n4027 & ~n5046;
  assign n5048 = ~n5045 & n5047;
  assign n5049 = n5045 & ~n5047;
  assign \sin[11]  = n5048 | n5049;
  assign n5051 = ~n5038 & ~n5040;
  assign n5052 = ~n177 & ~n186;
  assign n5053 = ~n207 & n5052;
  assign n5054 = ~n234 & n5053;
  assign n5055 = ~n335 & n5054;
  assign n5056 = n2367 & n5055;
  assign n5057 = n946 & n5056;
  assign n5058 = n4037 & n5057;
  assign n5059 = n2250 & n5058;
  assign n5060 = n380 & n5059;
  assign n5061 = ~n139 & n5060;
  assign n5062 = ~n134 & n5061;
  assign n5063 = ~n211 & n5062;
  assign n5064 = ~n5031 & ~n5034;
  assign n5065 = ~n5015 & ~n5027;
  assign n5066 = n2695 & n3896;
  assign n5067 = n2690 & n4054;
  assign n5068 = ~n5066 & ~n5067;
  assign n5069 = ~n669 & ~n5068;
  assign n5070 = n669 & n5068;
  assign n5071 = ~n5069 & ~n5070;
  assign n5072 = n2668 & n3750;
  assign n5073 = n2776 & n3272;
  assign n5074 = n2666 & ~n3628;
  assign n5075 = ~n5073 & ~n5074;
  assign n5076 = ~n5072 & n5075;
  assign n5077 = n2674 & n3762;
  assign n5078 = n5076 & ~n5077;
  assign n5079 = ~n525 & ~n5078;
  assign n5080 = ~n525 & ~n5079;
  assign n5081 = ~n5078 & ~n5079;
  assign n5082 = ~n5080 & ~n5081;
  assign n5083 = n5071 & ~n5082;
  assign n5084 = n5071 & ~n5083;
  assign n5085 = ~n5082 & ~n5083;
  assign n5086 = ~n5084 & ~n5085;
  assign n5087 = ~n4924 & ~n4997;
  assign n5088 = ~n5012 & ~n5087;
  assign n5089 = ~n525 & ~n3280;
  assign n5090 = ~n4997 & n5089;
  assign n5091 = n4997 & ~n5089;
  assign n5092 = ~n5088 & ~n5091;
  assign n5093 = ~n5090 & n5092;
  assign n5094 = ~n5088 & ~n5093;
  assign n5095 = ~n5091 & ~n5093;
  assign n5096 = ~n5090 & n5095;
  assign n5097 = ~n5094 & ~n5096;
  assign n5098 = ~n5086 & n5097;
  assign n5099 = n5086 & ~n5097;
  assign n5100 = ~n5098 & ~n5099;
  assign n5101 = ~n5065 & ~n5100;
  assign n5102 = n5065 & n5100;
  assign n5103 = ~n5101 & ~n5102;
  assign n5104 = ~n5064 & n5103;
  assign n5105 = n5064 & ~n5103;
  assign n5106 = ~n5104 & ~n5105;
  assign n5107 = n5063 & ~n5106;
  assign n5108 = ~n5063 & n5106;
  assign n5109 = ~n5107 & ~n5108;
  assign n5110 = ~n5051 & n5109;
  assign n5111 = n5051 & ~n5109;
  assign n5112 = ~n5110 & ~n5111;
  assign n5113 = ~n5044 & ~n5112;
  assign n5114 = n5044 & n5112;
  assign n5115 = ~n5113 & ~n5114;
  assign n5116 = ~n5045 & n5046;
  assign n5117 = ~n4027 & ~n5116;
  assign n5118 = ~n5115 & n5117;
  assign n5119 = n5115 & ~n5117;
  assign \sin[12]  = n5118 | n5119;
  assign n5121 = ~n5108 & ~n5110;
  assign n5122 = ~n194 & ~n394;
  assign n5123 = ~n255 & n5122;
  assign n5124 = ~n360 & n5123;
  assign n5125 = ~n118 & n5124;
  assign n5126 = n156 & n5125;
  assign n5127 = n4002 & n5126;
  assign n5128 = n311 & n5127;
  assign n5129 = n2178 & n5128;
  assign n5130 = n980 & n5129;
  assign n5131 = n3699 & n5130;
  assign n5132 = ~n196 & n5131;
  assign n5133 = ~n343 & n5132;
  assign n5134 = ~n257 & n5133;
  assign n5135 = ~n169 & n5134;
  assign n5136 = ~n142 & n5135;
  assign n5137 = ~n470 & n5136;
  assign n5138 = ~n351 & n5137;
  assign n5139 = ~n5101 & ~n5104;
  assign n5140 = n2668 & n3896;
  assign n5141 = n2776 & ~n3628;
  assign n5142 = n2666 & n3750;
  assign n5143 = ~n5141 & ~n5142;
  assign n5144 = ~n5140 & n5143;
  assign n5145 = n2674 & n3908;
  assign n5146 = n5144 & ~n5145;
  assign n5147 = ~n525 & ~n5146;
  assign n5148 = ~n5146 & ~n5147;
  assign n5149 = ~n525 & ~n5147;
  assign n5150 = ~n5148 & ~n5149;
  assign n5151 = n669 & n5089;
  assign n5152 = ~n669 & ~n5089;
  assign n5153 = ~n5151 & ~n5152;
  assign n5154 = ~n525 & n3272;
  assign n5155 = n5153 & n5154;
  assign n5156 = ~n5153 & ~n5154;
  assign n5157 = ~n5155 & ~n5156;
  assign n5158 = ~n5150 & n5157;
  assign n5159 = ~n5150 & ~n5158;
  assign n5160 = n5157 & ~n5158;
  assign n5161 = ~n5159 & ~n5160;
  assign n5162 = ~n5095 & n5161;
  assign n5163 = n5095 & ~n5161;
  assign n5164 = ~n5162 & ~n5163;
  assign n5165 = ~n5086 & ~n5097;
  assign n5166 = ~n5083 & ~n5165;
  assign n5167 = ~n5164 & ~n5166;
  assign n5168 = n5164 & n5166;
  assign n5169 = ~n5167 & ~n5168;
  assign n5170 = ~n5139 & n5169;
  assign n5171 = n5139 & ~n5169;
  assign n5172 = ~n5170 & ~n5171;
  assign n5173 = ~n5138 & n5172;
  assign n5174 = n5138 & ~n5172;
  assign n5175 = ~n5121 & ~n5174;
  assign n5176 = ~n5173 & n5175;
  assign n5177 = ~n5121 & ~n5176;
  assign n5178 = ~n5173 & ~n5176;
  assign n5179 = ~n5174 & n5178;
  assign n5180 = ~n5177 & ~n5179;
  assign n5181 = ~n5114 & n5180;
  assign n5182 = n5114 & ~n5180;
  assign n5183 = ~n5181 & ~n5182;
  assign n5184 = ~n5115 & n5116;
  assign n5185 = ~n4027 & ~n5184;
  assign n5186 = ~n5183 & n5185;
  assign n5187 = n5183 & ~n5185;
  assign \sin[13]  = n5186 | n5187;
  assign n5189 = n2367 & n2433;
  assign n5190 = n473 & n5189;
  assign n5191 = n967 & n5190;
  assign n5192 = n2190 & n5191;
  assign n5193 = n1457 & n5192;
  assign n5194 = n983 & n5193;
  assign n5195 = n3259 & n5194;
  assign n5196 = ~n138 & n5195;
  assign n5197 = ~n176 & n5196;
  assign n5198 = ~n127 & n5197;
  assign n5199 = ~n343 & n5198;
  assign n5200 = ~n370 & n5199;
  assign n5201 = ~n336 & n5200;
  assign n5202 = ~n506 & n5201;
  assign n5203 = ~n5167 & ~n5170;
  assign n5204 = ~n5095 & ~n5161;
  assign n5205 = ~n5158 & ~n5204;
  assign n5206 = ~n525 & ~n3628;
  assign n5207 = ~n5151 & ~n5155;
  assign n5208 = ~n5206 & ~n5207;
  assign n5209 = ~n5206 & ~n5208;
  assign n5210 = ~n5207 & ~n5208;
  assign n5211 = ~n5209 & ~n5210;
  assign n5212 = n2776 & n3750;
  assign n5213 = n2666 & n3896;
  assign n5214 = ~n5212 & ~n5213;
  assign n5215 = ~n2674 & n5214;
  assign n5216 = ~n4056 & n5214;
  assign n5217 = ~n5215 & ~n5216;
  assign n5218 = n525 & ~n5217;
  assign n5219 = ~n525 & n5217;
  assign n5220 = ~n5218 & ~n5219;
  assign n5221 = ~n5211 & n5220;
  assign n5222 = n5211 & ~n5220;
  assign n5223 = ~n5221 & ~n5222;
  assign n5224 = ~n5205 & n5223;
  assign n5225 = n5205 & ~n5223;
  assign n5226 = ~n5224 & ~n5225;
  assign n5227 = ~n5203 & n5226;
  assign n5228 = n5203 & ~n5226;
  assign n5229 = ~n5227 & ~n5228;
  assign n5230 = n5202 & ~n5229;
  assign n5231 = ~n5202 & n5229;
  assign n5232 = ~n5230 & ~n5231;
  assign n5233 = ~n5178 & n5232;
  assign n5234 = n5178 & ~n5232;
  assign n5235 = ~n5233 & ~n5234;
  assign n5236 = ~n5182 & ~n5235;
  assign n5237 = n5182 & n5235;
  assign n5238 = ~n5236 & ~n5237;
  assign n5239 = ~n5183 & n5184;
  assign n5240 = ~n4027 & ~n5239;
  assign n5241 = ~n5238 & n5240;
  assign n5242 = n5238 & ~n5240;
  assign \sin[14]  = n5241 | n5242;
  assign n5244 = ~n5231 & ~n5233;
  assign n5245 = ~n337 & n1145;
  assign n5246 = ~n328 & n5245;
  assign n5247 = ~n254 & n5246;
  assign n5248 = n970 & n5247;
  assign n5249 = n344 & n5248;
  assign n5250 = n5055 & n5249;
  assign n5251 = n2375 & n5250;
  assign n5252 = n1115 & n5251;
  assign n5253 = ~n127 & n5252;
  assign n5254 = ~n226 & n5253;
  assign n5255 = ~n217 & n5254;
  assign n5256 = ~n356 & n5255;
  assign n5257 = ~n506 & n5256;
  assign n5258 = ~n736 & n5257;
  assign n5259 = n2776 & n3896;
  assign n5260 = n2674 & n4054;
  assign n5261 = ~n5259 & ~n5260;
  assign n5262 = ~n525 & ~n5261;
  assign n5263 = ~n5261 & ~n5262;
  assign n5264 = ~n525 & ~n5262;
  assign n5265 = ~n5263 & ~n5264;
  assign n5266 = ~n525 & n3759;
  assign n5267 = ~n5265 & ~n5266;
  assign n5268 = ~n5265 & ~n5267;
  assign n5269 = ~n5266 & ~n5267;
  assign n5270 = ~n5268 & ~n5269;
  assign n5271 = ~n5208 & ~n5221;
  assign n5272 = n5270 & n5271;
  assign n5273 = ~n5270 & ~n5271;
  assign n5274 = ~n5272 & ~n5273;
  assign n5275 = ~n5224 & ~n5227;
  assign n5276 = ~n5274 & n5275;
  assign n5277 = n5274 & ~n5275;
  assign n5278 = ~n5276 & ~n5277;
  assign n5279 = ~n5258 & n5278;
  assign n5280 = n5258 & ~n5278;
  assign n5281 = ~n5244 & ~n5280;
  assign n5282 = ~n5279 & n5281;
  assign n5283 = ~n5244 & ~n5282;
  assign n5284 = ~n5279 & ~n5282;
  assign n5285 = ~n5280 & n5284;
  assign n5286 = ~n5283 & ~n5285;
  assign n5287 = ~n5237 & n5286;
  assign n5288 = n5237 & ~n5286;
  assign n5289 = ~n5287 & ~n5288;
  assign n5290 = ~n5238 & n5239;
  assign n5291 = ~n4027 & ~n5290;
  assign n5292 = ~n5289 & n5291;
  assign n5293 = n5289 & ~n5291;
  assign \sin[15]  = n5292 | n5293;
  assign n5295 = n638 & n2313;
  assign n5296 = n2252 & n5295;
  assign n5297 = n5125 & n5296;
  assign n5298 = n233 & n5297;
  assign n5299 = n475 & n5298;
  assign n5300 = n3702 & n5299;
  assign n5301 = ~n208 & n5300;
  assign n5302 = ~n447 & n5301;
  assign n5303 = ~n477 & n5302;
  assign n5304 = ~n5273 & ~n5277;
  assign n5305 = n3750 & ~n5206;
  assign n5306 = ~n525 & n5305;
  assign n5307 = ~n5267 & ~n5306;
  assign n5308 = ~n5304 & n5307;
  assign n5309 = n5304 & ~n5307;
  assign n5310 = ~n5308 & ~n5309;
  assign n5311 = n3896 & ~n5206;
  assign n5312 = ~n3896 & n5206;
  assign n5313 = ~n5311 & ~n5312;
  assign n5314 = ~n525 & n5313;
  assign n5315 = n5310 & ~n5314;
  assign n5316 = ~n5310 & n5314;
  assign n5317 = ~n5315 & ~n5316;
  assign n5318 = ~n5303 & ~n5317;
  assign n5319 = n5303 & n5317;
  assign n5320 = ~n5284 & ~n5319;
  assign n5321 = ~n5318 & n5320;
  assign n5322 = ~n5284 & ~n5321;
  assign n5323 = ~n5318 & ~n5321;
  assign n5324 = ~n5319 & n5323;
  assign n5325 = ~n5322 & ~n5324;
  assign n5326 = ~n5288 & n5325;
  assign n5327 = n5288 & ~n5325;
  assign n5328 = ~n5326 & ~n5327;
  assign n5329 = ~n5289 & n5290;
  assign n5330 = ~n4027 & ~n5329;
  assign n5331 = ~n5328 & n5330;
  assign n5332 = n5328 & ~n5330;
  assign \sin[16]  = n5331 | n5332;
  assign n5334 = n158 & n775;
  assign n5335 = n906 & n5334;
  assign n5336 = n259 & n5335;
  assign n5337 = n3243 & n5336;
  assign n5338 = n571 & n5337;
  assign n5339 = n980 & n5338;
  assign n5340 = ~n139 & n5339;
  assign n5341 = ~n207 & n5340;
  assign n5342 = ~n297 & n5341;
  assign n5343 = ~n368 & n5342;
  assign n5344 = ~n215 & n5343;
  assign n5345 = ~n5323 & ~n5344;
  assign n5346 = n5323 & n5344;
  assign n5347 = ~n5345 & ~n5346;
  assign n5348 = ~n5327 & n5347;
  assign n5349 = n5327 & ~n5347;
  assign n5350 = ~n5348 & ~n5349;
  assign n5351 = ~n5328 & n5329;
  assign n5352 = ~n4027 & ~n5351;
  assign n5353 = ~n5350 & n5352;
  assign n5354 = n5350 & ~n5352;
  assign \sin[17]  = ~n5353 & ~n5354;
  assign n5356 = n5327 & n5347;
  assign n5357 = n588 & n2170;
  assign n5358 = n608 & n5357;
  assign n5359 = n1152 & n5358;
  assign n5360 = n1108 & n5359;
  assign n5361 = n986 & n5360;
  assign n5362 = n3675 & n5361;
  assign n5363 = ~n176 & n5362;
  assign n5364 = ~n227 & n5363;
  assign n5365 = ~n207 & n5364;
  assign n5366 = ~n357 & n5365;
  assign n5367 = ~n238 & n5366;
  assign n5368 = n5345 & ~n5367;
  assign n5369 = ~n5345 & n5367;
  assign n5370 = ~n5368 & ~n5369;
  assign n5371 = ~n5356 & ~n5370;
  assign n5372 = n5356 & ~n5369;
  assign n5373 = ~n5371 & ~n5372;
  assign n5374 = n5350 & n5351;
  assign n5375 = ~n4027 & ~n5374;
  assign n5376 = ~n5373 & n5375;
  assign n5377 = n5373 & ~n5375;
  assign \sin[18]  = n5376 | n5377;
  assign n5379 = n4392 & n5247;
  assign n5380 = n373 & n5379;
  assign n5381 = n2540 & n5380;
  assign n5382 = n938 & n5381;
  assign n5383 = ~n144 & n5382;
  assign n5384 = ~n152 & n5383;
  assign n5385 = ~n208 & n5384;
  assign n5386 = ~n140 & n5385;
  assign n5387 = ~n446 & n5386;
  assign n5388 = ~n298 & n5387;
  assign n5389 = ~n206 & n5388;
  assign n5390 = ~n5368 & n5389;
  assign n5391 = n5368 & ~n5389;
  assign n5392 = ~n5390 & ~n5391;
  assign n5393 = ~n5372 & ~n5392;
  assign n5394 = n5372 & n5392;
  assign n5395 = ~n5393 & ~n5394;
  assign n5396 = ~n5373 & n5374;
  assign n5397 = ~n4027 & ~n5396;
  assign n5398 = ~n5395 & n5397;
  assign n5399 = n5395 & ~n5397;
  assign \sin[19]  = n5398 | n5399;
  assign n5401 = n189 & n459;
  assign n5402 = n999 & n5401;
  assign n5403 = n502 & n5402;
  assign n5404 = n4726 & n5403;
  assign n5405 = n369 & n5404;
  assign n5406 = ~n194 & n5405;
  assign n5407 = ~n227 & n5406;
  assign n5408 = ~n312 & n5407;
  assign n5409 = ~n218 & n5408;
  assign n5410 = ~n213 & n5409;
  assign n5411 = ~n212 & n5410;
  assign n5412 = ~n554 & n5411;
  assign n5413 = n5391 & ~n5412;
  assign n5414 = ~n5391 & n5412;
  assign n5415 = ~n5413 & ~n5414;
  assign n5416 = ~n5394 & ~n5415;
  assign n5417 = n5394 & ~n5414;
  assign n5418 = ~n5416 & ~n5417;
  assign n5419 = ~n5395 & n5396;
  assign n5420 = ~n4027 & ~n5419;
  assign n5421 = ~n5418 & n5420;
  assign n5422 = n5418 & ~n5420;
  assign \sin[20]  = n5421 | n5422;
  assign n5424 = n489 & n3617;
  assign n5425 = n444 & n5424;
  assign n5426 = ~n343 & n5425;
  assign n5427 = ~n360 & n5426;
  assign n5428 = ~n5413 & n5427;
  assign n5429 = n5413 & ~n5427;
  assign n5430 = ~n5428 & ~n5429;
  assign n5431 = ~n5417 & ~n5430;
  assign n5432 = n5417 & n5430;
  assign n5433 = ~n5431 & ~n5432;
  assign n5434 = ~n5418 & n5419;
  assign n5435 = ~n4027 & ~n5434;
  assign n5436 = ~n5433 & n5435;
  assign n5437 = n5433 & ~n5435;
  assign \sin[21]  = n5436 | n5437;
  assign n5439 = n444 & n517;
  assign n5440 = n5429 & ~n5439;
  assign n5441 = ~n5429 & n5439;
  assign n5442 = ~n5440 & ~n5441;
  assign n5443 = ~n5432 & ~n5442;
  assign n5444 = n5432 & ~n5441;
  assign n5445 = ~n5443 & ~n5444;
  assign n5446 = ~n5433 & n5434;
  assign n5447 = ~n4027 & ~n5446;
  assign n5448 = ~n5445 & n5447;
  assign n5449 = n5445 & ~n5447;
  assign \sin[22]  = n5448 | n5449;
  assign n5451 = ~\a[22]  & n71;
  assign n5452 = ~n5440 & ~n5444;
  assign n5453 = n5440 & n5444;
  assign n5454 = ~n5452 & ~n5453;
  assign n5455 = ~n5445 & n5446;
  assign n5456 = ~n4027 & ~n5455;
  assign n5457 = n5454 & ~n5456;
  assign n5458 = ~n5454 & n5456;
  assign n5459 = ~n5457 & ~n5458;
  assign \sin[23]  = n5451 | ~n5459;
  assign n5461 = ~n5452 & n5455;
  assign n5462 = ~n5453 & ~n5455;
  assign n5463 = ~n5461 & ~n5462;
  assign n5464 = ~n5451 & n5463;
  assign \sin[24]  = ~n4027 & ~n5464;
endmodule

