extern function void send(input_tx t);                                    

int save_pnt = 5;
logic [15:0] tx_save [0:5];
int init_flag = 1;