--
--
--
--
library ieee;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity ram0 is
 port (Clock: in std_logic;
       AddressBus: in std_logic_vector(11 downto 0);
       DataOut: out std_logic_vector(11 downto 0);
       DataIn: in std_logic_vector(11 downto 0);
       MemoryRead: in std_logic);
end ram0;

architecture syn of ram0 is

type memory_type is array (0 to 4127) of std_logic_vector(11 downto 0);
constant Bz : std_logic_vector(11 downto 0) := O"0000";

signal memory : memory_type :=
(


O"0000",O"5001",O"0002",O"0003",O"4500",O"2331",O"2324",O"0000",O"4005",O"2222",O"0000",O"1004",O"7773",O"1723",O"1021",O"0000",O"7777",O"3777",O"5777",O"6777",O"7377",O"7577",O"7677",O"7737",O"0000",O"7757",O"7767",O"7773",O"7775",O"7776",O"0000",O"1777",
O"0777",O"0377",O"0177",O"0077",O"0037",O"0017",O"0007",O"0003",O"0000",O"0001",O"4400",O"4577",O"2525",O"6666",O"4444",O"7070",O"0707",O"5252",O"1111",O"5252",O"0004",O"0244",O"0100",O"0336",O"0407",O"5472",O"3600",O"0212",O"0400",O"5476",O"3550",O"7700",
O"0330",O"0306",O"0564",O"1754",O"0527",O"0300",O"1676",O"7404",O"0000",O"7402",O"7401",O"7403",O"1610",O"7400",O"0526",O"0200",O"0430",O"5522",O"3530",O"7762",O"0450",O"5526",O"3510",O"7756",O"0510",O"5532",O"3470",O"1000",O"7744",O"1113",O"0370",O"1001",
O"0645",O"1532",O"2326",O"0651",O"1645",O"7410",O"0766",O"1600",O"0637",O"1655",O"0701",O"1163",O"7740",O"0012",O"1327",O"0363",O"0777",O"1166",O"7607",O"0256",O"0004",O"0077",O"7772",O"7746",O"7477",O"7766",O"0176",O"0172",O"0173",O"0174",O"0175",O"1234",
O"0000",O"7200",O"1052",O"3377",O"7440",O"7402",O"1052",O"7410",O"0000",O"7041",O"1377",O"7440",O"7402",O"7200",O"1053",O"3200",O"7440",O"7402",O"1053",O"7041",O"1200",O"7440",O"7402",O"7200",O"1020",O"3200",O"7440",O"7402",O"1200",O"7040",O"7440",O"7402",
O"7200",O"1036",O"3200",O"7440",O"7402",O"1200",O"7440",O"7402",O"7200",O"1054",O"3200",O"7440",O"7402",O"1054",O"7041",O"1200",O"7440",O"7402",O"7200",O"1055",O"3200",O"7440",O"7402",O"1055",O"7041",O"1200",O"7440",O"7402",O"7200",O"1056",O"3377",O"7440",
O"7402",O"1056",O"7041",O"1377",O"7440",O"7402",O"7200",O"1057",O"3377",O"7440",O"7402",O"1057",O"7041",O"1377",O"7440",O"7402",O"7200",O"1060",O"3000",O"7440",O"7402",O"1060",O"7041",O"1000",O"7440",O"7402",O"7200",O"1061",O"3000",O"7440",O"7402",O"1061",
O"7041",O"1000",O"7440",O"7402",O"7200",O"1062",O"3000",O"7440",O"7402",O"1062",O"7041",O"1000",O"7440",O"7402",O"7200",O"1063",O"3000",O"7440",O"7402",O"1063",O"7041",O"1000",O"7440",O"7402",O"5374",O"0610",O"5773",O"3450",O"7000",O"7000",O"7410",O"0000",
O"7200",O"1442",O"7041",O"1177",O"7440",O"7402",O"7200",O"7410",O"0000",O"1020",O"0442",O"7041",O"1177",O"7440",O"7402",O"7200",O"1020",O"3000",O"2436",O"7402",O"1000",O"7440",O"7402",O"7200",O"1572",O"7041",O"1176",O"7440",O"7402",O"7200",O"1020",O"0572",
O"7041",O"1176",O"7440",O"7402",O"7200",O"1172",O"3000",O"2436",O"7410",O"7402",O"1000",O"7041",O"1172",O"7040",O"7440",O"7402",O"7200",O"1573",O"7041",O"1172",O"7440",O"7402",O"7200",O"1020",O"0573",O"7041",O"1172",O"7440",O"7402",O"7200",O"1173",O"3000",
O"2436",O"7410",O"7402",O"1000",O"7041",O"1173",O"7040",O"7440",O"7402",O"7200",O"1574",O"7041",O"1173",O"7440",O"7402",O"7200",O"1020",O"0574",O"7041",O"1173",O"7440",O"7402",O"7200",O"1174",O"3000",O"2436",O"7410",O"7402",O"1000",O"7041",O"1174",O"7040",
O"7440",O"7402",O"7200",O"1575",O"7041",O"1174",O"7440",O"7402",O"7200",O"1020",O"0575",O"7041",O"1174",O"7440",O"7402",O"7200",O"1175",O"3000",O"2436",O"7410",O"7402",O"1000",O"7041",O"1175",O"7040",O"7440",O"7402",O"5377",O"0610",O"5776",O"3430",O"7000",
O"7200",O"1576",O"7041",O"1175",O"7440",O"7402",O"7200",O"1036",O"3010",O"0410",O"1010",O"1035",O"7040",O"7440",O"7402",O"7200",O"1035",O"3010",O"0410",O"1010",O"1036",O"7040",O"7440",O"7402",O"7200",O"1034",O"3010",O"3410",O"1010",O"1051",O"7040",O"7440",
O"7402",O"7200",O"1033",O"3010",O"1410",O"7200",O"1010",O"1047",O"7040",O"7440",O"7402",O"7200",O"1032",O"3010",O"0410",O"1010",O"1046",O"7040",O"7440",O"7402",O"7200",O"1031",O"3010",O"0410",O"1010",O"1045",O"7040",O"7440",O"7402",O"7200",O"1027",O"3010",
O"0410",O"1010",O"1044",O"7040",O"7440",O"7402",O"7200",O"1026",O"3010",O"0410",O"1010",O"1043",O"7040",O"7440",O"7402",O"7200",O"1025",O"3010",O"0410",O"1010",O"1042",O"7040",O"7440",O"7402",O"7200",O"1024",O"3010",O"0410",O"1010",O"1041",O"7040",O"7440",
O"7402",O"7200",O"1023",O"3010",O"0410",O"1010",O"1040",O"7040",O"7440",O"7402",O"7200",O"1022",O"3010",O"2410",O"7000",O"1010",O"1037",O"7040",O"7440",O"7402",O"7200",O"1021",O"3010",O"0410",O"1010",O"1021",O"7040",O"7440",O"7402",O"7000",O"7000",O"7000",
O"7200",O"1020",O"3010",O"0410",O"1010",O"1020",O"7040",O"7410",O"0000",O"7440",O"7402",O"7200",O"1036",O"3011",O"0411",O"1011",O"1035",O"7040",O"7440",O"7402",O"7200",O"1035",O"3011",O"0411",O"1011",O"1036",O"7040",O"7440",O"7402",O"7200",O"1034",O"3011",
O"3411",O"1011",O"1051",O"7040",O"7440",O"7402",O"7200",O"1033",O"3011",O"1411",O"7200",O"1011",O"1047",O"7040",O"7440",O"7402",O"7200",O"1032",O"3011",O"0411",O"1011",O"1046",O"7040",O"7440",O"7402",O"7200",O"1031",O"3011",O"0411",O"1011",O"1045",O"7040",
O"7440",O"7402",O"7200",O"1027",O"3011",O"0411",O"1011",O"1044",O"7040",O"7440",O"7402",O"7200",O"1026",O"3011",O"0411",O"1011",O"1043",O"7040",O"7440",O"7402",O"7200",O"1025",O"3011",O"0411",O"1011",O"1042",O"7040",O"7440",O"7402",O"7200",O"1024",O"3011",
O"0411",O"1011",O"1041",O"7040",O"7440",O"7402",O"7200",O"1023",O"3011",O"0411",O"1011",O"1040",O"7040",O"7440",O"7402",O"7200",O"1022",O"3011",O"2411",O"7000",O"1011",O"1037",O"7040",O"7440",O"7402",O"7000",O"5376",O"0610",O"5775",O"3410",O"7000",O"7000",
O"7200",O"1021",O"3011",O"0411",O"1011",O"1021",O"7040",O"7440",O"7402",O"7200",O"1020",O"3011",O"0411",O"1011",O"1020",O"7040",O"7440",O"7402",O"7200",O"1036",O"3012",O"0412",O"1012",O"1035",O"7040",O"7440",O"7402",O"7200",O"1035",O"3012",O"0412",O"1012",
O"1036",O"7040",O"7440",O"7402",O"7200",O"1034",O"3012",O"3412",O"1012",O"1051",O"7040",O"7440",O"7402",O"7200",O"1033",O"3012",O"1412",O"7200",O"1012",O"1047",O"7040",O"7440",O"7402",O"7200",O"1032",O"3012",O"0412",O"1012",O"1046",O"7040",O"7440",O"7402",
O"7200",O"1031",O"3012",O"0412",O"1012",O"1045",O"7040",O"7440",O"7402",O"7200",O"1027",O"3012",O"0412",O"1012",O"1044",O"7040",O"7440",O"7402",O"7200",O"1026",O"3012",O"0412",O"1012",O"1043",O"7040",O"7440",O"7402",O"7200",O"1025",O"3012",O"0412",O"1012",
O"1042",O"7040",O"7440",O"7402",O"7200",O"1024",O"3012",O"0412",O"1012",O"1041",O"7040",O"7440",O"7402",O"7200",O"1023",O"3012",O"0412",O"1012",O"1040",O"7040",O"7440",O"7402",O"7200",O"1022",O"3012",O"2412",O"7000",O"1012",O"1037",O"7040",O"7440",O"7402",
O"7200",O"1021",O"3012",O"0412",O"1012",O"1021",O"7040",O"7440",O"7402",O"7200",O"1020",O"3012",O"0412",O"1012",O"1020",O"7040",O"7440",O"7402",O"7200",O"1036",O"3013",O"0413",O"1013",O"1035",O"7040",O"7440",O"7402",O"7200",O"1035",O"3013",O"0413",O"1013",
O"1036",O"7040",O"7440",O"7402",O"7200",O"1034",O"3013",O"3413",O"1013",O"1051",O"7040",O"7440",O"7402",O"7200",O"1033",O"3013",O"1413",O"7200",O"1013",O"1047",O"7040",O"7440",O"7402",O"7200",O"1032",O"3013",O"0413",O"1013",O"1046",O"7040",O"7440",O"7402",
O"7200",O"1031",O"3013",O"0413",O"1013",O"1045",O"7040",O"7440",O"7402",O"7200",O"1027",O"3013",O"0413",O"1013",O"1044",O"7040",O"7440",O"7402",O"7200",O"1026",O"3013",O"0413",O"1013",O"1043",O"7040",O"7440",O"7402",O"7200",O"1025",O"3013",O"0413",O"1013",
O"1042",O"7040",O"7440",O"7402",O"7200",O"1024",O"3013",O"0413",O"1013",O"1041",O"7040",O"7440",O"7402",O"7200",O"1023",O"3013",O"0413",O"1013",O"1040",O"7040",O"7440",O"7402",O"7200",O"1022",O"3013",O"2413",O"7000",O"1013",O"1037",O"7040",O"7440",O"7402",
O"7200",O"1021",O"3013",O"0413",O"1013",O"1021",O"7040",O"7440",O"7402",O"7200",O"1020",O"3013",O"0413",O"1013",O"1020",O"7040",O"7440",O"7402",O"7200",O"1036",O"3014",O"0414",O"1014",O"1035",O"7040",O"7440",O"7402",O"7200",O"1035",O"3014",O"0414",O"1014",
O"1036",O"7040",O"7440",O"7402",O"7200",O"1034",O"3014",O"3414",O"1014",O"1051",O"7040",O"7440",O"7402",O"7200",O"1033",O"3014",O"1414",O"7200",O"1014",O"1047",O"7040",O"7440",O"7402",O"7200",O"1032",O"3014",O"0414",O"1014",O"1046",O"7040",O"7440",O"7402",
O"7200",O"1031",O"3014",O"0414",O"1014",O"1045",O"7040",O"7440",O"7402",O"7200",O"1027",O"3014",O"0414",O"1014",O"1044",O"7040",O"7440",O"7402",O"7200",O"1026",O"3014",O"0414",O"1014",O"1043",O"7040",O"7440",O"7402",O"7200",O"1025",O"3014",O"0414",O"1014",
O"1042",O"7040",O"7440",O"7402",O"7200",O"1024",O"3014",O"0414",O"1014",O"1041",O"7040",O"7440",O"7402",O"7200",O"1023",O"3014",O"0414",O"1014",O"1040",O"7040",O"7440",O"7402",O"7200",O"1022",O"3014",O"2414",O"7000",O"1014",O"1037",O"7040",O"7440",O"7402",
O"7200",O"1021",O"3014",O"0414",O"1014",O"1021",O"7040",O"7410",O"0000",O"7440",O"7402",O"7200",O"1020",O"3014",O"0414",O"1014",O"1020",O"7040",O"7440",O"7402",O"7200",O"1036",O"3015",O"0415",O"1015",O"1035",O"7040",O"7440",O"7402",O"7200",O"1035",O"3015",
O"0415",O"1015",O"1036",O"7040",O"7440",O"7402",O"7200",O"1034",O"3015",O"3415",O"1015",O"1051",O"7040",O"7440",O"7402",O"7200",O"1033",O"3015",O"1415",O"7200",O"1015",O"1047",O"7040",O"7440",O"7402",O"7200",O"1032",O"3015",O"0415",O"1015",O"1046",O"7040",
O"7440",O"7402",O"7200",O"1031",O"3015",O"0415",O"1015",O"1045",O"7040",O"7440",O"7402",O"7200",O"1027",O"3015",O"0415",O"1015",O"1044",O"7040",O"7440",O"7402",O"7200",O"1026",O"3015",O"0415",O"1015",O"1043",O"7040",O"7440",O"7402",O"7200",O"1025",O"3015",
O"0415",O"1015",O"1042",O"7040",O"7440",O"7402",O"7200",O"1024",O"3015",O"0415",O"1015",O"1041",O"7040",O"7440",O"7402",O"7200",O"1023",O"3015",O"0415",O"1015",O"1040",O"7040",O"7440",O"7402",O"7000",O"7000",O"5376",O"0610",O"5775",O"3370",O"7000",O"7000",
O"7200",O"1022",O"3015",O"2415",O"7000",O"1015",O"1037",O"7040",O"7440",O"7402",O"7200",O"1021",O"3015",O"0415",O"1015",O"1021",O"7040",O"7440",O"7402",O"7200",O"1020",O"3015",O"0415",O"1015",O"1020",O"7040",O"7440",O"7402",O"7200",O"1036",O"3016",O"0416",
O"1016",O"1035",O"7040",O"7440",O"7402",O"7200",O"1035",O"3016",O"0416",O"1016",O"1036",O"7040",O"7440",O"7402",O"7200",O"1034",O"3016",O"3416",O"1016",O"1051",O"7040",O"7440",O"7402",O"7200",O"1033",O"3016",O"1416",O"7200",O"1016",O"1047",O"7040",O"7440",
O"7402",O"7200",O"1032",O"3016",O"0416",O"1016",O"1046",O"7040",O"7440",O"7402",O"7200",O"1031",O"3016",O"0416",O"1016",O"1045",O"7040",O"7440",O"7402",O"7200",O"1027",O"3016",O"0416",O"1016",O"1044",O"7040",O"7440",O"7402",O"7200",O"1026",O"3016",O"0416",
O"1016",O"1043",O"7040",O"7440",O"7402",O"7200",O"1025",O"3016",O"0416",O"1016",O"1042",O"7040",O"7440",O"7402",O"7200",O"1024",O"3016",O"0416",O"1016",O"1041",O"7040",O"7440",O"7402",O"7200",O"1023",O"3016",O"0416",O"1016",O"1040",O"7040",O"7440",O"7402",
O"7200",O"1022",O"3016",O"2416",O"7000",O"1016",O"1037",O"7040",O"7440",O"7402",O"7200",O"1021",O"3016",O"0416",O"1016",O"1021",O"7040",O"7440",O"7402",O"7200",O"1020",O"3016",O"0416",O"1016",O"1020",O"7040",O"7440",O"7402",O"7200",O"1036",O"3017",O"0417",
O"1017",O"1035",O"7040",O"7440",O"7402",O"7200",O"1035",O"3017",O"0417",O"1017",O"1036",O"7040",O"7440",O"7402",O"7200",O"1034",O"3017",O"3417",O"1017",O"1051",O"7040",O"7440",O"7402",O"7200",O"1033",O"3017",O"1417",O"7200",O"1017",O"1047",O"7040",O"7440",
O"7402",O"7200",O"1032",O"3017",O"0417",O"1017",O"1046",O"7040",O"7440",O"7402",O"7200",O"1031",O"3017",O"0417",O"1017",O"1045",O"7040",O"7440",O"7402",O"7200",O"1027",O"3017",O"0417",O"1017",O"1044",O"7040",O"7440",O"7402",O"7200",O"1026",O"3017",O"0417",
O"1017",O"1043",O"7040",O"7440",O"7402",O"7200",O"1025",O"3017",O"0417",O"1017",O"1042",O"7040",O"7440",O"7402",O"7200",O"1024",O"3017",O"0417",O"1017",O"1041",O"7040",O"7440",O"7402",O"7200",O"1023",O"3017",O"0417",O"1017",O"1040",O"7040",O"7440",O"7402",
O"7200",O"1022",O"3017",O"2417",O"7000",O"1017",O"1037",O"7040",O"7440",O"7402",O"7200",O"1021",O"3017",O"0417",O"1017",O"1021",O"7040",O"7440",O"7402",O"7200",O"1020",O"3017",O"0417",O"1017",O"1020",O"7040",O"7440",O"7402",O"5236",O"7402",O"7410",O"2644",
O"1237",O"3010",O"5410",O"7402",O"7402",O"4247",O"7402",O"7402",O"1247",O"7410",O"2646",O"7041",O"1252",O"7440",O"7402",O"7410",O"2664",O"1260",O"3010",O"4410",O"7402",O"7402",O"1265",O"7410",O"2664",O"7041",O"1270",O"7440",O"7402",O"4676",O"4011",O"6041",
O"6046",O"6041",O"5301",O"7200",O"1312",O"3002",O"6001",O"7000",O"7402",O"2710",O"2713",O"7440",O"7402",O"1000",O"7041",O"1311",O"7640",O"7402",O"1041",O"6041",O"6046",O"6041",O"5325",O"7200",O"1336",O"3002",O"6001",O"1020",O"7402",O"2734",O"2737",O"7040",
O"7440",O"7402",O"1000",O"7041",O"1335",O"7640",O"7402",O"1041",O"6041",O"6046",O"6041",O"5352",O"7200",O"1364",O"3002",O"1020",O"6001",O"0020",O"7402",O"2762",O"2765",O"7040",O"7440",O"7402",O"1000",O"7041",O"1363",O"7640",O"7402",O"7000",O"7000",O"7000",
O"1041",O"6041",O"6046",O"6041",O"5203",O"7200",O"1215",O"3002",O"1020",O"6001",O"3003",O"7402",O"3013",O"3016",O"7440",O"7402",O"1003",O"7040",O"7440",O"7402",O"3003",O"1000",O"7041",O"1214",O"7640",O"7402",O"1041",O"6041",O"6046",O"6041",O"5235",O"7200",
O"1250",O"3002",O"1035",O"3003",O"6001",O"2003",O"7402",O"3046",O"3051",O"7440",O"7402",O"1003",O"7040",O"7440",O"7402",O"3003",O"1000",O"7041",O"1247",O"7640",O"7402",O"1041",O"6041",O"6046",O"6041",O"5270",O"7200",O"1304",O"3002",O"1020",O"3003",O"6001",
O"2003",O"7402",O"7402",O"3102",O"3105",O"7440",O"7402",O"1003",O"7440",O"7402",O"3003",O"1000",O"7041",O"1303",O"7640",O"7402",O"1041",O"6041",O"6046",O"6041",O"5323",O"7200",O"1334",O"3002",O"6001",O"5331",O"7402",O"3131",O"3135",O"7440",O"7402",O"1000",
O"7041",O"1333",O"7640",O"7402",O"1041",O"6041",O"6046",O"6041",O"5347",O"7200",O"1360",O"3002",O"6001",O"4003",O"7402",O"3156",O"3161",O"7440",O"7402",O"1003",O"7041",O"1357",O"7440",O"7402",O"1000",O"7041",O"1064",O"7640",O"7402",O"7000",O"7000",O"7000",
O"1041",O"6041",O"6046",O"6041",O"5203",O"7200",O"1215",O"3002",O"1020",O"6001",O"7200",O"7402",O"3213",O"3216",O"7440",O"7402",O"1000",O"7041",O"1214",O"7640",O"7402",O"1041",O"6041",O"6046",O"6041",O"5230",O"7200",O"1242",O"3002",O"6001",O"6041",O"7402",
O"7402",O"3240",O"3243",O"7440",O"7402",O"1000",O"7041",O"1241",O"7640",O"7402",O"1041",O"6041",O"6046",O"6041",O"5255",O"7200",O"1317",O"3002",O"6001",O"6002",O"6001",O"6002",O"6001",O"6002",O"6001",O"6002",O"6001",O"6002",O"6001",O"6002",O"6001",O"6002",
O"6001",O"6002",O"6001",O"6002",O"6001",O"6002",O"6001",O"6002",O"6001",O"6002",O"6001",O"6002",O"6041",O"7402",O"7410",O"3321",O"7410",O"7402",O"6042",O"7200",O"1334",O"3002",O"6001",O"7000",O"7000",O"7000",O"7000",O"7410",O"3336",O"7410",O"7402",O"6002",
O"7200",O"5742",O"4000",O"4010",O"7777",O"7777",O"7777",O"7777",O"1743",O"7440",O"7402",O"7200",O"3743",O"7200",O"5757",O"2173",O"2010",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"1760",O"7440",O"7402",O"5774",O"3400",O"7777",O"7777",O"7777",
O"7200",O"5602",O"1173",O"1010",O"7777",O"7777",O"7777",O"7777",O"1603",O"7440",O"7402",O"7200",O"3603",O"7200",O"5617",O"0574",O"0410",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"1620",O"7440",O"7402",O"7200",O"3620",O"7200",O"5637",O"0371",
O"0210",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"1640",O"7440",O"7402",O"7200",O"3640",O"7200",O"5657",O"0130",O"0110",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"1660",O"7440",O"7402",O"7200",O"3110",O"7200",O"5677",O"0124",
O"0050",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"1700",O"7440",O"7402",O"7200",O"3050",O"7200",O"5717",O"0120",O"0030",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"1720",O"7440",O"7402",O"7200",O"3030",O"7200",O"3000",O"5740",
O"0074",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"1436",O"7440",O"7402",O"7200",O"3000",O"7200",O"5757",O"0070",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"1446",O"7440",O"7402",O"7200",O"3007",O"1223",O"7001",O"3223",O"1223",O"1224",O"7640",O"5622",O"3223",O"1225",O"6046",O"6041",O"5217",O"5622",O"0201",O"0000",O"7730",O"0207",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"0610",O"5602",O"3350",O"0000",O"2405",O"2324",O"5606",O"2400",O"0000",O"0000",O"1221",O"3001",O"3002",O"3003",O"1041",O"2211",O"5611",O"5402",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",
O"1234",O"0000",O"0000",O"0000",O"0411",O"2320",O"5620",O"0100",O"1101",O"1456",O"2001",O"0000",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",
O"1234",O"0000",O"2754",O"0000",O"3024",O"6256",O"0216",O"5707",O"7562",O"6065",O"0000",O"0000",O"0000",O"0700",O"7005",O"5620",O"0100",O"0556",O"2001",O"0000",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",
O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",O"7136",O"2745",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",
O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777",O"7777"
);
begin

-- DataOut <= memory(conv_integer(unsigned(AddressBus))) when (MemoryRequest = '1' and MemoryRead = '1') else (others => 'Z');

process (Clock)
begin
   if(Clock'event and Clock = '0' and MemoryRead = '0') then 
      memory(conv_integer(unsigned(AddressBus))) <= DataIn;
   end if;
   if(Clock'event and Clock = '0' and MemoryRead = '1') then 
      DataOut <= memory(conv_integer(unsigned(AddressBus)));
   end if;
end process;

end syn;
