// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: rca_driver.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2016-04-18-EP on Tue Mar 19 21:50:30 2019
//=============================================================================
// Description: Driver for rca
//=============================================================================

`ifndef RCA_DRIVER_SV
`define RCA_DRIVER_SV

// You can insert code here by setting driver_inc_before_class in file rca.tpl

class rca_driver extends uvm_driver #(trans);

  `uvm_component_utils(rca_driver)

  virtual rca_if vif;

  extern function new(string name, uvm_component parent);

  // Methods run_phase and do_drive generated by setting driver_inc in file rca.tpl
  extern task run_phase(uvm_phase phase);
  extern task do_drive();

  // You can insert code here by setting driver_inc_inside_class in file rca.tpl

endclass : rca_driver 


function rca_driver::new(string name, uvm_component parent);
  super.new(name, parent);
endfunction : new


task rca_driver::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)

  forever
  begin
    seq_item_port.get_next_item(req);
      `uvm_info(get_type_name(), {"req item\n",req.sprint}, UVM_HIGH)
    do_drive();
    seq_item_port.item_done();
  end
endtask : run_phase


// Start of inlined include file generated_tb/tb/include/rca_driver_inc.sv
task rca_driver::do_drive();
  vif.a <= req.input1;
  vif.b <= req.input2;
  vif.ci <= req.carryinput;
  @(posedge vif.clk);
endtask// End of inlined include file

// You can insert code here by setting driver_inc_after_class in file rca.tpl

`endif // RCA_DRIVER_SV

