// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: top_pkg.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2016-04-18-EP on Sat Apr 27 13:59:59 2019
//=============================================================================
// Description: Package for top
//=============================================================================

package top_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  import data_input_pkg::*;
  import data_output_pkg::*;

  `include "top_config.sv"
  `include "top_seq_lib.sv"
  `include "port_converter.sv"
  `include "reference.sv"
  `include "top_env.sv"

endpackage : top_pkg

