module design7_20_35_top #(parameter WIDTH=32,CHANNEL=20) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	reg [WIDTH-1:0] d_in10;
	reg [WIDTH-1:0] d_in11;
	reg [WIDTH-1:0] d_in12;
	reg [WIDTH-1:0] d_in13;
	reg [WIDTH-1:0] d_in14;
	reg [WIDTH-1:0] d_in15;
	reg [WIDTH-1:0] d_in16;
	reg [WIDTH-1:0] d_in17;
	reg [WIDTH-1:0] d_in18;
	reg [WIDTH-1:0] d_in19;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;
	wire [WIDTH-1:0] d_out10;
	wire [WIDTH-1:0] d_out11;
	wire [WIDTH-1:0] d_out12;
	wire [WIDTH-1:0] d_out13;
	wire [WIDTH-1:0] d_out14;
	wire [WIDTH-1:0] d_out15;
	wire [WIDTH-1:0] d_out16;
	wire [WIDTH-1:0] d_out17;
	wire [WIDTH-1:0] d_out18;
	wire [WIDTH-1:0] d_out19;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH+1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 = tmp[WIDTH-1:0];
		d_in1 = tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 = tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 = tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 = tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 = tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 = tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 = tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 = tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 = tmp[(WIDTH*10)-1:WIDTH*9];
		d_in10 = tmp[(WIDTH*11)-1:WIDTH*10];
		d_in11 = tmp[(WIDTH*12)-1:WIDTH*11];
		d_in12 = tmp[(WIDTH*13)-1:WIDTH*12];
		d_in13 = tmp[(WIDTH*14)-1:WIDTH*13];
		d_in14 = tmp[(WIDTH*15)-1:WIDTH*14];
		d_in15 = tmp[(WIDTH*16)-1:WIDTH*15];
		d_in16 = tmp[(WIDTH*17)-1:WIDTH*16];
		d_in17 = tmp[(WIDTH*18)-1:WIDTH*17];
		d_in18 = tmp[(WIDTH*19)-1:WIDTH*18];
		d_in19 = tmp[(WIDTH*20)-1:WIDTH*19];
	end

	design7_20_35 #(.WIDTH(WIDTH)) design7_20_35_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_in10(d_in10),.d_in11(d_in11),.d_in12(d_in12),.d_in13(d_in13),.d_in14(d_in14),.d_in15(d_in15),.d_in16(d_in16),.d_in17(d_in17),.d_in18(d_in18),.d_in19(d_in19),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.d_out10(d_out10),.d_out11(d_out11),.d_out12(d_out12),.d_out13(d_out13),.d_out14(d_out14),.d_out15(d_out15),.d_out16(d_out16),.d_out17(d_out17),.d_out18(d_out18),.d_out19(d_out19),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9^d_out10^d_out11^d_out12^d_out13^d_out14^d_out15^d_out16^d_out17^d_out18^d_out19;

endmodule

module design7_20_35 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_in10, d_in11, d_in12, d_in13, d_in14, d_in15, d_in16, d_in17, d_in18, d_in19, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, d_out10, d_out11, d_out12, d_out13, d_out14, d_out15, d_out16, d_out17, d_out18, d_out19, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	input [WIDTH-1:0] d_in10; 
	input [WIDTH-1:0] d_in11; 
	input [WIDTH-1:0] d_in12; 
	input [WIDTH-1:0] d_in13; 
	input [WIDTH-1:0] d_in14; 
	input [WIDTH-1:0] d_in15; 
	input [WIDTH-1:0] d_in16; 
	input [WIDTH-1:0] d_in17; 
	input [WIDTH-1:0] d_in18; 
	input [WIDTH-1:0] d_in19; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 
	output [WIDTH-1:0] d_out10; 
	output [WIDTH-1:0] d_out11; 
	output [WIDTH-1:0] d_out12; 
	output [WIDTH-1:0] d_out13; 
	output [WIDTH-1:0] d_out14; 
	output [WIDTH-1:0] d_out15; 
	output [WIDTH-1:0] d_out16; 
	output [WIDTH-1:0] d_out17; 
	output [WIDTH-1:0] d_out18; 
	output [WIDTH-1:0] d_out19; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d0_29;
	wire [WIDTH-1:0] wire_d0_30;
	wire [WIDTH-1:0] wire_d0_31;
	wire [WIDTH-1:0] wire_d0_32;
	wire [WIDTH-1:0] wire_d0_33;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d1_29;
	wire [WIDTH-1:0] wire_d1_30;
	wire [WIDTH-1:0] wire_d1_31;
	wire [WIDTH-1:0] wire_d1_32;
	wire [WIDTH-1:0] wire_d1_33;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d2_29;
	wire [WIDTH-1:0] wire_d2_30;
	wire [WIDTH-1:0] wire_d2_31;
	wire [WIDTH-1:0] wire_d2_32;
	wire [WIDTH-1:0] wire_d2_33;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d3_29;
	wire [WIDTH-1:0] wire_d3_30;
	wire [WIDTH-1:0] wire_d3_31;
	wire [WIDTH-1:0] wire_d3_32;
	wire [WIDTH-1:0] wire_d3_33;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d4_29;
	wire [WIDTH-1:0] wire_d4_30;
	wire [WIDTH-1:0] wire_d4_31;
	wire [WIDTH-1:0] wire_d4_32;
	wire [WIDTH-1:0] wire_d4_33;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d5_29;
	wire [WIDTH-1:0] wire_d5_30;
	wire [WIDTH-1:0] wire_d5_31;
	wire [WIDTH-1:0] wire_d5_32;
	wire [WIDTH-1:0] wire_d5_33;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d6_29;
	wire [WIDTH-1:0] wire_d6_30;
	wire [WIDTH-1:0] wire_d6_31;
	wire [WIDTH-1:0] wire_d6_32;
	wire [WIDTH-1:0] wire_d6_33;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d7_29;
	wire [WIDTH-1:0] wire_d7_30;
	wire [WIDTH-1:0] wire_d7_31;
	wire [WIDTH-1:0] wire_d7_32;
	wire [WIDTH-1:0] wire_d7_33;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d8_29;
	wire [WIDTH-1:0] wire_d8_30;
	wire [WIDTH-1:0] wire_d8_31;
	wire [WIDTH-1:0] wire_d8_32;
	wire [WIDTH-1:0] wire_d8_33;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d9_29;
	wire [WIDTH-1:0] wire_d9_30;
	wire [WIDTH-1:0] wire_d9_31;
	wire [WIDTH-1:0] wire_d9_32;
	wire [WIDTH-1:0] wire_d9_33;
	wire [WIDTH-1:0] wire_d10_0;
	wire [WIDTH-1:0] wire_d10_1;
	wire [WIDTH-1:0] wire_d10_2;
	wire [WIDTH-1:0] wire_d10_3;
	wire [WIDTH-1:0] wire_d10_4;
	wire [WIDTH-1:0] wire_d10_5;
	wire [WIDTH-1:0] wire_d10_6;
	wire [WIDTH-1:0] wire_d10_7;
	wire [WIDTH-1:0] wire_d10_8;
	wire [WIDTH-1:0] wire_d10_9;
	wire [WIDTH-1:0] wire_d10_10;
	wire [WIDTH-1:0] wire_d10_11;
	wire [WIDTH-1:0] wire_d10_12;
	wire [WIDTH-1:0] wire_d10_13;
	wire [WIDTH-1:0] wire_d10_14;
	wire [WIDTH-1:0] wire_d10_15;
	wire [WIDTH-1:0] wire_d10_16;
	wire [WIDTH-1:0] wire_d10_17;
	wire [WIDTH-1:0] wire_d10_18;
	wire [WIDTH-1:0] wire_d10_19;
	wire [WIDTH-1:0] wire_d10_20;
	wire [WIDTH-1:0] wire_d10_21;
	wire [WIDTH-1:0] wire_d10_22;
	wire [WIDTH-1:0] wire_d10_23;
	wire [WIDTH-1:0] wire_d10_24;
	wire [WIDTH-1:0] wire_d10_25;
	wire [WIDTH-1:0] wire_d10_26;
	wire [WIDTH-1:0] wire_d10_27;
	wire [WIDTH-1:0] wire_d10_28;
	wire [WIDTH-1:0] wire_d10_29;
	wire [WIDTH-1:0] wire_d10_30;
	wire [WIDTH-1:0] wire_d10_31;
	wire [WIDTH-1:0] wire_d10_32;
	wire [WIDTH-1:0] wire_d10_33;
	wire [WIDTH-1:0] wire_d11_0;
	wire [WIDTH-1:0] wire_d11_1;
	wire [WIDTH-1:0] wire_d11_2;
	wire [WIDTH-1:0] wire_d11_3;
	wire [WIDTH-1:0] wire_d11_4;
	wire [WIDTH-1:0] wire_d11_5;
	wire [WIDTH-1:0] wire_d11_6;
	wire [WIDTH-1:0] wire_d11_7;
	wire [WIDTH-1:0] wire_d11_8;
	wire [WIDTH-1:0] wire_d11_9;
	wire [WIDTH-1:0] wire_d11_10;
	wire [WIDTH-1:0] wire_d11_11;
	wire [WIDTH-1:0] wire_d11_12;
	wire [WIDTH-1:0] wire_d11_13;
	wire [WIDTH-1:0] wire_d11_14;
	wire [WIDTH-1:0] wire_d11_15;
	wire [WIDTH-1:0] wire_d11_16;
	wire [WIDTH-1:0] wire_d11_17;
	wire [WIDTH-1:0] wire_d11_18;
	wire [WIDTH-1:0] wire_d11_19;
	wire [WIDTH-1:0] wire_d11_20;
	wire [WIDTH-1:0] wire_d11_21;
	wire [WIDTH-1:0] wire_d11_22;
	wire [WIDTH-1:0] wire_d11_23;
	wire [WIDTH-1:0] wire_d11_24;
	wire [WIDTH-1:0] wire_d11_25;
	wire [WIDTH-1:0] wire_d11_26;
	wire [WIDTH-1:0] wire_d11_27;
	wire [WIDTH-1:0] wire_d11_28;
	wire [WIDTH-1:0] wire_d11_29;
	wire [WIDTH-1:0] wire_d11_30;
	wire [WIDTH-1:0] wire_d11_31;
	wire [WIDTH-1:0] wire_d11_32;
	wire [WIDTH-1:0] wire_d11_33;
	wire [WIDTH-1:0] wire_d12_0;
	wire [WIDTH-1:0] wire_d12_1;
	wire [WIDTH-1:0] wire_d12_2;
	wire [WIDTH-1:0] wire_d12_3;
	wire [WIDTH-1:0] wire_d12_4;
	wire [WIDTH-1:0] wire_d12_5;
	wire [WIDTH-1:0] wire_d12_6;
	wire [WIDTH-1:0] wire_d12_7;
	wire [WIDTH-1:0] wire_d12_8;
	wire [WIDTH-1:0] wire_d12_9;
	wire [WIDTH-1:0] wire_d12_10;
	wire [WIDTH-1:0] wire_d12_11;
	wire [WIDTH-1:0] wire_d12_12;
	wire [WIDTH-1:0] wire_d12_13;
	wire [WIDTH-1:0] wire_d12_14;
	wire [WIDTH-1:0] wire_d12_15;
	wire [WIDTH-1:0] wire_d12_16;
	wire [WIDTH-1:0] wire_d12_17;
	wire [WIDTH-1:0] wire_d12_18;
	wire [WIDTH-1:0] wire_d12_19;
	wire [WIDTH-1:0] wire_d12_20;
	wire [WIDTH-1:0] wire_d12_21;
	wire [WIDTH-1:0] wire_d12_22;
	wire [WIDTH-1:0] wire_d12_23;
	wire [WIDTH-1:0] wire_d12_24;
	wire [WIDTH-1:0] wire_d12_25;
	wire [WIDTH-1:0] wire_d12_26;
	wire [WIDTH-1:0] wire_d12_27;
	wire [WIDTH-1:0] wire_d12_28;
	wire [WIDTH-1:0] wire_d12_29;
	wire [WIDTH-1:0] wire_d12_30;
	wire [WIDTH-1:0] wire_d12_31;
	wire [WIDTH-1:0] wire_d12_32;
	wire [WIDTH-1:0] wire_d12_33;
	wire [WIDTH-1:0] wire_d13_0;
	wire [WIDTH-1:0] wire_d13_1;
	wire [WIDTH-1:0] wire_d13_2;
	wire [WIDTH-1:0] wire_d13_3;
	wire [WIDTH-1:0] wire_d13_4;
	wire [WIDTH-1:0] wire_d13_5;
	wire [WIDTH-1:0] wire_d13_6;
	wire [WIDTH-1:0] wire_d13_7;
	wire [WIDTH-1:0] wire_d13_8;
	wire [WIDTH-1:0] wire_d13_9;
	wire [WIDTH-1:0] wire_d13_10;
	wire [WIDTH-1:0] wire_d13_11;
	wire [WIDTH-1:0] wire_d13_12;
	wire [WIDTH-1:0] wire_d13_13;
	wire [WIDTH-1:0] wire_d13_14;
	wire [WIDTH-1:0] wire_d13_15;
	wire [WIDTH-1:0] wire_d13_16;
	wire [WIDTH-1:0] wire_d13_17;
	wire [WIDTH-1:0] wire_d13_18;
	wire [WIDTH-1:0] wire_d13_19;
	wire [WIDTH-1:0] wire_d13_20;
	wire [WIDTH-1:0] wire_d13_21;
	wire [WIDTH-1:0] wire_d13_22;
	wire [WIDTH-1:0] wire_d13_23;
	wire [WIDTH-1:0] wire_d13_24;
	wire [WIDTH-1:0] wire_d13_25;
	wire [WIDTH-1:0] wire_d13_26;
	wire [WIDTH-1:0] wire_d13_27;
	wire [WIDTH-1:0] wire_d13_28;
	wire [WIDTH-1:0] wire_d13_29;
	wire [WIDTH-1:0] wire_d13_30;
	wire [WIDTH-1:0] wire_d13_31;
	wire [WIDTH-1:0] wire_d13_32;
	wire [WIDTH-1:0] wire_d13_33;
	wire [WIDTH-1:0] wire_d14_0;
	wire [WIDTH-1:0] wire_d14_1;
	wire [WIDTH-1:0] wire_d14_2;
	wire [WIDTH-1:0] wire_d14_3;
	wire [WIDTH-1:0] wire_d14_4;
	wire [WIDTH-1:0] wire_d14_5;
	wire [WIDTH-1:0] wire_d14_6;
	wire [WIDTH-1:0] wire_d14_7;
	wire [WIDTH-1:0] wire_d14_8;
	wire [WIDTH-1:0] wire_d14_9;
	wire [WIDTH-1:0] wire_d14_10;
	wire [WIDTH-1:0] wire_d14_11;
	wire [WIDTH-1:0] wire_d14_12;
	wire [WIDTH-1:0] wire_d14_13;
	wire [WIDTH-1:0] wire_d14_14;
	wire [WIDTH-1:0] wire_d14_15;
	wire [WIDTH-1:0] wire_d14_16;
	wire [WIDTH-1:0] wire_d14_17;
	wire [WIDTH-1:0] wire_d14_18;
	wire [WIDTH-1:0] wire_d14_19;
	wire [WIDTH-1:0] wire_d14_20;
	wire [WIDTH-1:0] wire_d14_21;
	wire [WIDTH-1:0] wire_d14_22;
	wire [WIDTH-1:0] wire_d14_23;
	wire [WIDTH-1:0] wire_d14_24;
	wire [WIDTH-1:0] wire_d14_25;
	wire [WIDTH-1:0] wire_d14_26;
	wire [WIDTH-1:0] wire_d14_27;
	wire [WIDTH-1:0] wire_d14_28;
	wire [WIDTH-1:0] wire_d14_29;
	wire [WIDTH-1:0] wire_d14_30;
	wire [WIDTH-1:0] wire_d14_31;
	wire [WIDTH-1:0] wire_d14_32;
	wire [WIDTH-1:0] wire_d14_33;
	wire [WIDTH-1:0] wire_d15_0;
	wire [WIDTH-1:0] wire_d15_1;
	wire [WIDTH-1:0] wire_d15_2;
	wire [WIDTH-1:0] wire_d15_3;
	wire [WIDTH-1:0] wire_d15_4;
	wire [WIDTH-1:0] wire_d15_5;
	wire [WIDTH-1:0] wire_d15_6;
	wire [WIDTH-1:0] wire_d15_7;
	wire [WIDTH-1:0] wire_d15_8;
	wire [WIDTH-1:0] wire_d15_9;
	wire [WIDTH-1:0] wire_d15_10;
	wire [WIDTH-1:0] wire_d15_11;
	wire [WIDTH-1:0] wire_d15_12;
	wire [WIDTH-1:0] wire_d15_13;
	wire [WIDTH-1:0] wire_d15_14;
	wire [WIDTH-1:0] wire_d15_15;
	wire [WIDTH-1:0] wire_d15_16;
	wire [WIDTH-1:0] wire_d15_17;
	wire [WIDTH-1:0] wire_d15_18;
	wire [WIDTH-1:0] wire_d15_19;
	wire [WIDTH-1:0] wire_d15_20;
	wire [WIDTH-1:0] wire_d15_21;
	wire [WIDTH-1:0] wire_d15_22;
	wire [WIDTH-1:0] wire_d15_23;
	wire [WIDTH-1:0] wire_d15_24;
	wire [WIDTH-1:0] wire_d15_25;
	wire [WIDTH-1:0] wire_d15_26;
	wire [WIDTH-1:0] wire_d15_27;
	wire [WIDTH-1:0] wire_d15_28;
	wire [WIDTH-1:0] wire_d15_29;
	wire [WIDTH-1:0] wire_d15_30;
	wire [WIDTH-1:0] wire_d15_31;
	wire [WIDTH-1:0] wire_d15_32;
	wire [WIDTH-1:0] wire_d15_33;
	wire [WIDTH-1:0] wire_d16_0;
	wire [WIDTH-1:0] wire_d16_1;
	wire [WIDTH-1:0] wire_d16_2;
	wire [WIDTH-1:0] wire_d16_3;
	wire [WIDTH-1:0] wire_d16_4;
	wire [WIDTH-1:0] wire_d16_5;
	wire [WIDTH-1:0] wire_d16_6;
	wire [WIDTH-1:0] wire_d16_7;
	wire [WIDTH-1:0] wire_d16_8;
	wire [WIDTH-1:0] wire_d16_9;
	wire [WIDTH-1:0] wire_d16_10;
	wire [WIDTH-1:0] wire_d16_11;
	wire [WIDTH-1:0] wire_d16_12;
	wire [WIDTH-1:0] wire_d16_13;
	wire [WIDTH-1:0] wire_d16_14;
	wire [WIDTH-1:0] wire_d16_15;
	wire [WIDTH-1:0] wire_d16_16;
	wire [WIDTH-1:0] wire_d16_17;
	wire [WIDTH-1:0] wire_d16_18;
	wire [WIDTH-1:0] wire_d16_19;
	wire [WIDTH-1:0] wire_d16_20;
	wire [WIDTH-1:0] wire_d16_21;
	wire [WIDTH-1:0] wire_d16_22;
	wire [WIDTH-1:0] wire_d16_23;
	wire [WIDTH-1:0] wire_d16_24;
	wire [WIDTH-1:0] wire_d16_25;
	wire [WIDTH-1:0] wire_d16_26;
	wire [WIDTH-1:0] wire_d16_27;
	wire [WIDTH-1:0] wire_d16_28;
	wire [WIDTH-1:0] wire_d16_29;
	wire [WIDTH-1:0] wire_d16_30;
	wire [WIDTH-1:0] wire_d16_31;
	wire [WIDTH-1:0] wire_d16_32;
	wire [WIDTH-1:0] wire_d16_33;
	wire [WIDTH-1:0] wire_d17_0;
	wire [WIDTH-1:0] wire_d17_1;
	wire [WIDTH-1:0] wire_d17_2;
	wire [WIDTH-1:0] wire_d17_3;
	wire [WIDTH-1:0] wire_d17_4;
	wire [WIDTH-1:0] wire_d17_5;
	wire [WIDTH-1:0] wire_d17_6;
	wire [WIDTH-1:0] wire_d17_7;
	wire [WIDTH-1:0] wire_d17_8;
	wire [WIDTH-1:0] wire_d17_9;
	wire [WIDTH-1:0] wire_d17_10;
	wire [WIDTH-1:0] wire_d17_11;
	wire [WIDTH-1:0] wire_d17_12;
	wire [WIDTH-1:0] wire_d17_13;
	wire [WIDTH-1:0] wire_d17_14;
	wire [WIDTH-1:0] wire_d17_15;
	wire [WIDTH-1:0] wire_d17_16;
	wire [WIDTH-1:0] wire_d17_17;
	wire [WIDTH-1:0] wire_d17_18;
	wire [WIDTH-1:0] wire_d17_19;
	wire [WIDTH-1:0] wire_d17_20;
	wire [WIDTH-1:0] wire_d17_21;
	wire [WIDTH-1:0] wire_d17_22;
	wire [WIDTH-1:0] wire_d17_23;
	wire [WIDTH-1:0] wire_d17_24;
	wire [WIDTH-1:0] wire_d17_25;
	wire [WIDTH-1:0] wire_d17_26;
	wire [WIDTH-1:0] wire_d17_27;
	wire [WIDTH-1:0] wire_d17_28;
	wire [WIDTH-1:0] wire_d17_29;
	wire [WIDTH-1:0] wire_d17_30;
	wire [WIDTH-1:0] wire_d17_31;
	wire [WIDTH-1:0] wire_d17_32;
	wire [WIDTH-1:0] wire_d17_33;
	wire [WIDTH-1:0] wire_d18_0;
	wire [WIDTH-1:0] wire_d18_1;
	wire [WIDTH-1:0] wire_d18_2;
	wire [WIDTH-1:0] wire_d18_3;
	wire [WIDTH-1:0] wire_d18_4;
	wire [WIDTH-1:0] wire_d18_5;
	wire [WIDTH-1:0] wire_d18_6;
	wire [WIDTH-1:0] wire_d18_7;
	wire [WIDTH-1:0] wire_d18_8;
	wire [WIDTH-1:0] wire_d18_9;
	wire [WIDTH-1:0] wire_d18_10;
	wire [WIDTH-1:0] wire_d18_11;
	wire [WIDTH-1:0] wire_d18_12;
	wire [WIDTH-1:0] wire_d18_13;
	wire [WIDTH-1:0] wire_d18_14;
	wire [WIDTH-1:0] wire_d18_15;
	wire [WIDTH-1:0] wire_d18_16;
	wire [WIDTH-1:0] wire_d18_17;
	wire [WIDTH-1:0] wire_d18_18;
	wire [WIDTH-1:0] wire_d18_19;
	wire [WIDTH-1:0] wire_d18_20;
	wire [WIDTH-1:0] wire_d18_21;
	wire [WIDTH-1:0] wire_d18_22;
	wire [WIDTH-1:0] wire_d18_23;
	wire [WIDTH-1:0] wire_d18_24;
	wire [WIDTH-1:0] wire_d18_25;
	wire [WIDTH-1:0] wire_d18_26;
	wire [WIDTH-1:0] wire_d18_27;
	wire [WIDTH-1:0] wire_d18_28;
	wire [WIDTH-1:0] wire_d18_29;
	wire [WIDTH-1:0] wire_d18_30;
	wire [WIDTH-1:0] wire_d18_31;
	wire [WIDTH-1:0] wire_d18_32;
	wire [WIDTH-1:0] wire_d18_33;
	wire [WIDTH-1:0] wire_d19_0;
	wire [WIDTH-1:0] wire_d19_1;
	wire [WIDTH-1:0] wire_d19_2;
	wire [WIDTH-1:0] wire_d19_3;
	wire [WIDTH-1:0] wire_d19_4;
	wire [WIDTH-1:0] wire_d19_5;
	wire [WIDTH-1:0] wire_d19_6;
	wire [WIDTH-1:0] wire_d19_7;
	wire [WIDTH-1:0] wire_d19_8;
	wire [WIDTH-1:0] wire_d19_9;
	wire [WIDTH-1:0] wire_d19_10;
	wire [WIDTH-1:0] wire_d19_11;
	wire [WIDTH-1:0] wire_d19_12;
	wire [WIDTH-1:0] wire_d19_13;
	wire [WIDTH-1:0] wire_d19_14;
	wire [WIDTH-1:0] wire_d19_15;
	wire [WIDTH-1:0] wire_d19_16;
	wire [WIDTH-1:0] wire_d19_17;
	wire [WIDTH-1:0] wire_d19_18;
	wire [WIDTH-1:0] wire_d19_19;
	wire [WIDTH-1:0] wire_d19_20;
	wire [WIDTH-1:0] wire_d19_21;
	wire [WIDTH-1:0] wire_d19_22;
	wire [WIDTH-1:0] wire_d19_23;
	wire [WIDTH-1:0] wire_d19_24;
	wire [WIDTH-1:0] wire_d19_25;
	wire [WIDTH-1:0] wire_d19_26;
	wire [WIDTH-1:0] wire_d19_27;
	wire [WIDTH-1:0] wire_d19_28;
	wire [WIDTH-1:0] wire_d19_29;
	wire [WIDTH-1:0] wire_d19_30;
	wire [WIDTH-1:0] wire_d19_31;
	wire [WIDTH-1:0] wire_d19_32;
	wire [WIDTH-1:0] wire_d19_33;

	invertion #(.WIDTH(WIDTH)) invertion_instance00(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	encoder #(.WIDTH(WIDTH)) encoder_instance01(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance02(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance03(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance04(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance05(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance06(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance07(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance08(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance09(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance029(.data_in(wire_d0_28),.data_out(wire_d0_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance030(.data_in(wire_d0_29),.data_out(wire_d0_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance031(.data_in(wire_d0_30),.data_out(wire_d0_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance032(.data_in(wire_d0_31),.data_out(wire_d0_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance033(.data_in(wire_d0_32),.data_out(wire_d0_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance034(.data_in(wire_d0_33),.data_out(d_out0),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance10(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	encoder #(.WIDTH(WIDTH)) encoder_instance11(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance12(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance13(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance14(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance15(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance17(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance19(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance129(.data_in(wire_d1_28),.data_out(wire_d1_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance130(.data_in(wire_d1_29),.data_out(wire_d1_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131(.data_in(wire_d1_30),.data_out(wire_d1_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance132(.data_in(wire_d1_31),.data_out(wire_d1_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance133(.data_in(wire_d1_32),.data_out(wire_d1_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance134(.data_in(wire_d1_33),.data_out(d_out1),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance20(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	invertion #(.WIDTH(WIDTH)) invertion_instance21(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance22(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance23(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance24(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance25(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance26(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance27(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance28(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance29(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance229(.data_in(wire_d2_28),.data_out(wire_d2_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance230(.data_in(wire_d2_29),.data_out(wire_d2_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance231(.data_in(wire_d2_30),.data_out(wire_d2_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232(.data_in(wire_d2_31),.data_out(wire_d2_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance233(.data_in(wire_d2_32),.data_out(wire_d2_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance234(.data_in(wire_d2_33),.data_out(d_out2),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance30(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	invertion #(.WIDTH(WIDTH)) invertion_instance31(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance32(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance33(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance34(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance35(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance36(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance37(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance38(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance39(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance329(.data_in(wire_d3_28),.data_out(wire_d3_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance330(.data_in(wire_d3_29),.data_out(wire_d3_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance331(.data_in(wire_d3_30),.data_out(wire_d3_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance332(.data_in(wire_d3_31),.data_out(wire_d3_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333(.data_in(wire_d3_32),.data_out(wire_d3_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance334(.data_in(wire_d3_33),.data_out(d_out3),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance40(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	encoder #(.WIDTH(WIDTH)) encoder_instance41(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance42(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance43(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance44(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance45(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance46(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance47(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance48(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance49(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance429(.data_in(wire_d4_28),.data_out(wire_d4_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance430(.data_in(wire_d4_29),.data_out(wire_d4_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance431(.data_in(wire_d4_30),.data_out(wire_d4_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance432(.data_in(wire_d4_31),.data_out(wire_d4_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance433(.data_in(wire_d4_32),.data_out(wire_d4_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434(.data_in(wire_d4_33),.data_out(d_out4),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance50(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	register #(.WIDTH(WIDTH)) register_instance51(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance52(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance53(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance55(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance56(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance57(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance58(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance59(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance529(.data_in(wire_d5_28),.data_out(wire_d5_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance530(.data_in(wire_d5_29),.data_out(wire_d5_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance531(.data_in(wire_d5_30),.data_out(wire_d5_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance532(.data_in(wire_d5_31),.data_out(wire_d5_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance533(.data_in(wire_d5_32),.data_out(wire_d5_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance534(.data_in(wire_d5_33),.data_out(d_out5),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance60(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance61(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance62(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance63(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance64(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance65(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance66(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance67(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance68(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance69(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance629(.data_in(wire_d6_28),.data_out(wire_d6_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance630(.data_in(wire_d6_29),.data_out(wire_d6_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance631(.data_in(wire_d6_30),.data_out(wire_d6_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance632(.data_in(wire_d6_31),.data_out(wire_d6_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance633(.data_in(wire_d6_32),.data_out(wire_d6_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance634(.data_in(wire_d6_33),.data_out(d_out6),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance70(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	large_mux #(.WIDTH(WIDTH)) large_mux_instance71(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance72(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance73(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance74(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance75(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance76(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance77(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance78(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance79(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance729(.data_in(wire_d7_28),.data_out(wire_d7_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance730(.data_in(wire_d7_29),.data_out(wire_d7_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance731(.data_in(wire_d7_30),.data_out(wire_d7_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance732(.data_in(wire_d7_31),.data_out(wire_d7_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance733(.data_in(wire_d7_32),.data_out(wire_d7_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance734(.data_in(wire_d7_33),.data_out(d_out7),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance80(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance81(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance82(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance83(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance84(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance85(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance86(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance88(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance89(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance829(.data_in(wire_d8_28),.data_out(wire_d8_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance830(.data_in(wire_d8_29),.data_out(wire_d8_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance831(.data_in(wire_d8_30),.data_out(wire_d8_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance832(.data_in(wire_d8_31),.data_out(wire_d8_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance833(.data_in(wire_d8_32),.data_out(wire_d8_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance834(.data_in(wire_d8_33),.data_out(d_out8),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance90(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance91(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance92(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance93(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance94(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance95(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance96(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance97(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance98(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance99(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance929(.data_in(wire_d9_28),.data_out(wire_d9_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance930(.data_in(wire_d9_29),.data_out(wire_d9_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance931(.data_in(wire_d9_30),.data_out(wire_d9_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance932(.data_in(wire_d9_31),.data_out(wire_d9_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance933(.data_in(wire_d9_32),.data_out(wire_d9_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance934(.data_in(wire_d9_33),.data_out(d_out9),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100(.data_in(d_in10),.data_out(wire_d10_0),.clk(clk),.rst(rst));            //channel 11
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance101(.data_in(wire_d10_0),.data_out(wire_d10_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance102(.data_in(wire_d10_1),.data_out(wire_d10_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance103(.data_in(wire_d10_2),.data_out(wire_d10_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance104(.data_in(wire_d10_3),.data_out(wire_d10_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance105(.data_in(wire_d10_4),.data_out(wire_d10_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance106(.data_in(wire_d10_5),.data_out(wire_d10_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance107(.data_in(wire_d10_6),.data_out(wire_d10_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance108(.data_in(wire_d10_7),.data_out(wire_d10_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance109(.data_in(wire_d10_8),.data_out(wire_d10_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1010(.data_in(wire_d10_9),.data_out(wire_d10_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1011(.data_in(wire_d10_10),.data_out(wire_d10_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1012(.data_in(wire_d10_11),.data_out(wire_d10_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1013(.data_in(wire_d10_12),.data_out(wire_d10_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1014(.data_in(wire_d10_13),.data_out(wire_d10_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1015(.data_in(wire_d10_14),.data_out(wire_d10_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1016(.data_in(wire_d10_15),.data_out(wire_d10_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1017(.data_in(wire_d10_16),.data_out(wire_d10_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1018(.data_in(wire_d10_17),.data_out(wire_d10_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1019(.data_in(wire_d10_18),.data_out(wire_d10_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1020(.data_in(wire_d10_19),.data_out(wire_d10_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1021(.data_in(wire_d10_20),.data_out(wire_d10_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1022(.data_in(wire_d10_21),.data_out(wire_d10_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1023(.data_in(wire_d10_22),.data_out(wire_d10_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1024(.data_in(wire_d10_23),.data_out(wire_d10_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1025(.data_in(wire_d10_24),.data_out(wire_d10_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1026(.data_in(wire_d10_25),.data_out(wire_d10_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1027(.data_in(wire_d10_26),.data_out(wire_d10_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1028(.data_in(wire_d10_27),.data_out(wire_d10_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1029(.data_in(wire_d10_28),.data_out(wire_d10_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1030(.data_in(wire_d10_29),.data_out(wire_d10_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1031(.data_in(wire_d10_30),.data_out(wire_d10_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1032(.data_in(wire_d10_31),.data_out(wire_d10_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1033(.data_in(wire_d10_32),.data_out(wire_d10_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1034(.data_in(wire_d10_33),.data_out(d_out10),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance110(.data_in(d_in11),.data_out(wire_d11_0),.clk(clk),.rst(rst));            //channel 12
	encoder #(.WIDTH(WIDTH)) encoder_instance111(.data_in(wire_d11_0),.data_out(wire_d11_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance112(.data_in(wire_d11_1),.data_out(wire_d11_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance113(.data_in(wire_d11_2),.data_out(wire_d11_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance114(.data_in(wire_d11_3),.data_out(wire_d11_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance115(.data_in(wire_d11_4),.data_out(wire_d11_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance116(.data_in(wire_d11_5),.data_out(wire_d11_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance117(.data_in(wire_d11_6),.data_out(wire_d11_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance118(.data_in(wire_d11_7),.data_out(wire_d11_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance119(.data_in(wire_d11_8),.data_out(wire_d11_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1110(.data_in(wire_d11_9),.data_out(wire_d11_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1111(.data_in(wire_d11_10),.data_out(wire_d11_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1112(.data_in(wire_d11_11),.data_out(wire_d11_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1113(.data_in(wire_d11_12),.data_out(wire_d11_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1114(.data_in(wire_d11_13),.data_out(wire_d11_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1115(.data_in(wire_d11_14),.data_out(wire_d11_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1116(.data_in(wire_d11_15),.data_out(wire_d11_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1117(.data_in(wire_d11_16),.data_out(wire_d11_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1118(.data_in(wire_d11_17),.data_out(wire_d11_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1119(.data_in(wire_d11_18),.data_out(wire_d11_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1120(.data_in(wire_d11_19),.data_out(wire_d11_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1121(.data_in(wire_d11_20),.data_out(wire_d11_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1122(.data_in(wire_d11_21),.data_out(wire_d11_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1123(.data_in(wire_d11_22),.data_out(wire_d11_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1124(.data_in(wire_d11_23),.data_out(wire_d11_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1125(.data_in(wire_d11_24),.data_out(wire_d11_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1126(.data_in(wire_d11_25),.data_out(wire_d11_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1127(.data_in(wire_d11_26),.data_out(wire_d11_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1128(.data_in(wire_d11_27),.data_out(wire_d11_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1129(.data_in(wire_d11_28),.data_out(wire_d11_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1130(.data_in(wire_d11_29),.data_out(wire_d11_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1131(.data_in(wire_d11_30),.data_out(wire_d11_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1132(.data_in(wire_d11_31),.data_out(wire_d11_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1133(.data_in(wire_d11_32),.data_out(wire_d11_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1134(.data_in(wire_d11_33),.data_out(d_out11),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance120(.data_in(d_in12),.data_out(wire_d12_0),.clk(clk),.rst(rst));            //channel 13
	invertion #(.WIDTH(WIDTH)) invertion_instance121(.data_in(wire_d12_0),.data_out(wire_d12_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance122(.data_in(wire_d12_1),.data_out(wire_d12_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance123(.data_in(wire_d12_2),.data_out(wire_d12_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance124(.data_in(wire_d12_3),.data_out(wire_d12_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance125(.data_in(wire_d12_4),.data_out(wire_d12_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance126(.data_in(wire_d12_5),.data_out(wire_d12_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance127(.data_in(wire_d12_6),.data_out(wire_d12_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance128(.data_in(wire_d12_7),.data_out(wire_d12_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance129(.data_in(wire_d12_8),.data_out(wire_d12_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1210(.data_in(wire_d12_9),.data_out(wire_d12_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1211(.data_in(wire_d12_10),.data_out(wire_d12_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1212(.data_in(wire_d12_11),.data_out(wire_d12_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1213(.data_in(wire_d12_12),.data_out(wire_d12_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1214(.data_in(wire_d12_13),.data_out(wire_d12_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1215(.data_in(wire_d12_14),.data_out(wire_d12_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1216(.data_in(wire_d12_15),.data_out(wire_d12_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1217(.data_in(wire_d12_16),.data_out(wire_d12_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1218(.data_in(wire_d12_17),.data_out(wire_d12_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1219(.data_in(wire_d12_18),.data_out(wire_d12_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1220(.data_in(wire_d12_19),.data_out(wire_d12_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1221(.data_in(wire_d12_20),.data_out(wire_d12_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1222(.data_in(wire_d12_21),.data_out(wire_d12_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1223(.data_in(wire_d12_22),.data_out(wire_d12_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1224(.data_in(wire_d12_23),.data_out(wire_d12_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1225(.data_in(wire_d12_24),.data_out(wire_d12_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1226(.data_in(wire_d12_25),.data_out(wire_d12_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1227(.data_in(wire_d12_26),.data_out(wire_d12_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1228(.data_in(wire_d12_27),.data_out(wire_d12_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1229(.data_in(wire_d12_28),.data_out(wire_d12_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1230(.data_in(wire_d12_29),.data_out(wire_d12_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1231(.data_in(wire_d12_30),.data_out(wire_d12_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1232(.data_in(wire_d12_31),.data_out(wire_d12_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1233(.data_in(wire_d12_32),.data_out(wire_d12_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1234(.data_in(wire_d12_33),.data_out(d_out12),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance130(.data_in(d_in13),.data_out(wire_d13_0),.clk(clk),.rst(rst));            //channel 14
	encoder #(.WIDTH(WIDTH)) encoder_instance131(.data_in(wire_d13_0),.data_out(wire_d13_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance132(.data_in(wire_d13_1),.data_out(wire_d13_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance133(.data_in(wire_d13_2),.data_out(wire_d13_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance134(.data_in(wire_d13_3),.data_out(wire_d13_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance135(.data_in(wire_d13_4),.data_out(wire_d13_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance136(.data_in(wire_d13_5),.data_out(wire_d13_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance137(.data_in(wire_d13_6),.data_out(wire_d13_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance138(.data_in(wire_d13_7),.data_out(wire_d13_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance139(.data_in(wire_d13_8),.data_out(wire_d13_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1310(.data_in(wire_d13_9),.data_out(wire_d13_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1311(.data_in(wire_d13_10),.data_out(wire_d13_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1312(.data_in(wire_d13_11),.data_out(wire_d13_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1313(.data_in(wire_d13_12),.data_out(wire_d13_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1314(.data_in(wire_d13_13),.data_out(wire_d13_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1315(.data_in(wire_d13_14),.data_out(wire_d13_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1316(.data_in(wire_d13_15),.data_out(wire_d13_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1317(.data_in(wire_d13_16),.data_out(wire_d13_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1318(.data_in(wire_d13_17),.data_out(wire_d13_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1319(.data_in(wire_d13_18),.data_out(wire_d13_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1320(.data_in(wire_d13_19),.data_out(wire_d13_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1321(.data_in(wire_d13_20),.data_out(wire_d13_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1322(.data_in(wire_d13_21),.data_out(wire_d13_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1323(.data_in(wire_d13_22),.data_out(wire_d13_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1324(.data_in(wire_d13_23),.data_out(wire_d13_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1325(.data_in(wire_d13_24),.data_out(wire_d13_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1326(.data_in(wire_d13_25),.data_out(wire_d13_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1327(.data_in(wire_d13_26),.data_out(wire_d13_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1328(.data_in(wire_d13_27),.data_out(wire_d13_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1329(.data_in(wire_d13_28),.data_out(wire_d13_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1330(.data_in(wire_d13_29),.data_out(wire_d13_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1331(.data_in(wire_d13_30),.data_out(wire_d13_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1332(.data_in(wire_d13_31),.data_out(wire_d13_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1333(.data_in(wire_d13_32),.data_out(wire_d13_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1334(.data_in(wire_d13_33),.data_out(d_out13),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance140(.data_in(d_in14),.data_out(wire_d14_0),.clk(clk),.rst(rst));            //channel 15
	encoder #(.WIDTH(WIDTH)) encoder_instance141(.data_in(wire_d14_0),.data_out(wire_d14_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance142(.data_in(wire_d14_1),.data_out(wire_d14_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance143(.data_in(wire_d14_2),.data_out(wire_d14_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance144(.data_in(wire_d14_3),.data_out(wire_d14_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance145(.data_in(wire_d14_4),.data_out(wire_d14_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance146(.data_in(wire_d14_5),.data_out(wire_d14_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance147(.data_in(wire_d14_6),.data_out(wire_d14_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance148(.data_in(wire_d14_7),.data_out(wire_d14_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance149(.data_in(wire_d14_8),.data_out(wire_d14_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1410(.data_in(wire_d14_9),.data_out(wire_d14_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1411(.data_in(wire_d14_10),.data_out(wire_d14_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1412(.data_in(wire_d14_11),.data_out(wire_d14_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1413(.data_in(wire_d14_12),.data_out(wire_d14_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1414(.data_in(wire_d14_13),.data_out(wire_d14_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1415(.data_in(wire_d14_14),.data_out(wire_d14_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1416(.data_in(wire_d14_15),.data_out(wire_d14_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1417(.data_in(wire_d14_16),.data_out(wire_d14_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1418(.data_in(wire_d14_17),.data_out(wire_d14_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1419(.data_in(wire_d14_18),.data_out(wire_d14_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1420(.data_in(wire_d14_19),.data_out(wire_d14_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1421(.data_in(wire_d14_20),.data_out(wire_d14_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1422(.data_in(wire_d14_21),.data_out(wire_d14_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1423(.data_in(wire_d14_22),.data_out(wire_d14_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1424(.data_in(wire_d14_23),.data_out(wire_d14_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1425(.data_in(wire_d14_24),.data_out(wire_d14_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1426(.data_in(wire_d14_25),.data_out(wire_d14_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1427(.data_in(wire_d14_26),.data_out(wire_d14_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1428(.data_in(wire_d14_27),.data_out(wire_d14_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1429(.data_in(wire_d14_28),.data_out(wire_d14_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1430(.data_in(wire_d14_29),.data_out(wire_d14_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1431(.data_in(wire_d14_30),.data_out(wire_d14_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1432(.data_in(wire_d14_31),.data_out(wire_d14_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1433(.data_in(wire_d14_32),.data_out(wire_d14_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1434(.data_in(wire_d14_33),.data_out(d_out14),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance150(.data_in(d_in15),.data_out(wire_d15_0),.clk(clk),.rst(rst));            //channel 16
	invertion #(.WIDTH(WIDTH)) invertion_instance151(.data_in(wire_d15_0),.data_out(wire_d15_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance152(.data_in(wire_d15_1),.data_out(wire_d15_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance153(.data_in(wire_d15_2),.data_out(wire_d15_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance154(.data_in(wire_d15_3),.data_out(wire_d15_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance155(.data_in(wire_d15_4),.data_out(wire_d15_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance156(.data_in(wire_d15_5),.data_out(wire_d15_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance157(.data_in(wire_d15_6),.data_out(wire_d15_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance158(.data_in(wire_d15_7),.data_out(wire_d15_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance159(.data_in(wire_d15_8),.data_out(wire_d15_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1510(.data_in(wire_d15_9),.data_out(wire_d15_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1511(.data_in(wire_d15_10),.data_out(wire_d15_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1512(.data_in(wire_d15_11),.data_out(wire_d15_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1513(.data_in(wire_d15_12),.data_out(wire_d15_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1514(.data_in(wire_d15_13),.data_out(wire_d15_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1515(.data_in(wire_d15_14),.data_out(wire_d15_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1516(.data_in(wire_d15_15),.data_out(wire_d15_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1517(.data_in(wire_d15_16),.data_out(wire_d15_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1518(.data_in(wire_d15_17),.data_out(wire_d15_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1519(.data_in(wire_d15_18),.data_out(wire_d15_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1520(.data_in(wire_d15_19),.data_out(wire_d15_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1521(.data_in(wire_d15_20),.data_out(wire_d15_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1522(.data_in(wire_d15_21),.data_out(wire_d15_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1523(.data_in(wire_d15_22),.data_out(wire_d15_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1524(.data_in(wire_d15_23),.data_out(wire_d15_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1525(.data_in(wire_d15_24),.data_out(wire_d15_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1526(.data_in(wire_d15_25),.data_out(wire_d15_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1527(.data_in(wire_d15_26),.data_out(wire_d15_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1528(.data_in(wire_d15_27),.data_out(wire_d15_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1529(.data_in(wire_d15_28),.data_out(wire_d15_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1530(.data_in(wire_d15_29),.data_out(wire_d15_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1531(.data_in(wire_d15_30),.data_out(wire_d15_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1532(.data_in(wire_d15_31),.data_out(wire_d15_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1533(.data_in(wire_d15_32),.data_out(wire_d15_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1534(.data_in(wire_d15_33),.data_out(d_out15),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance160(.data_in(d_in16),.data_out(wire_d16_0),.clk(clk),.rst(rst));            //channel 17
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161(.data_in(wire_d16_0),.data_out(wire_d16_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance162(.data_in(wire_d16_1),.data_out(wire_d16_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance163(.data_in(wire_d16_2),.data_out(wire_d16_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance164(.data_in(wire_d16_3),.data_out(wire_d16_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance165(.data_in(wire_d16_4),.data_out(wire_d16_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance166(.data_in(wire_d16_5),.data_out(wire_d16_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance167(.data_in(wire_d16_6),.data_out(wire_d16_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance168(.data_in(wire_d16_7),.data_out(wire_d16_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance169(.data_in(wire_d16_8),.data_out(wire_d16_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1610(.data_in(wire_d16_9),.data_out(wire_d16_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1611(.data_in(wire_d16_10),.data_out(wire_d16_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1612(.data_in(wire_d16_11),.data_out(wire_d16_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1613(.data_in(wire_d16_12),.data_out(wire_d16_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1614(.data_in(wire_d16_13),.data_out(wire_d16_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1615(.data_in(wire_d16_14),.data_out(wire_d16_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1616(.data_in(wire_d16_15),.data_out(wire_d16_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1617(.data_in(wire_d16_16),.data_out(wire_d16_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1618(.data_in(wire_d16_17),.data_out(wire_d16_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1619(.data_in(wire_d16_18),.data_out(wire_d16_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1620(.data_in(wire_d16_19),.data_out(wire_d16_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1621(.data_in(wire_d16_20),.data_out(wire_d16_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1622(.data_in(wire_d16_21),.data_out(wire_d16_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1623(.data_in(wire_d16_22),.data_out(wire_d16_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1624(.data_in(wire_d16_23),.data_out(wire_d16_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1625(.data_in(wire_d16_24),.data_out(wire_d16_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1626(.data_in(wire_d16_25),.data_out(wire_d16_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1627(.data_in(wire_d16_26),.data_out(wire_d16_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1628(.data_in(wire_d16_27),.data_out(wire_d16_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1629(.data_in(wire_d16_28),.data_out(wire_d16_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1630(.data_in(wire_d16_29),.data_out(wire_d16_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1631(.data_in(wire_d16_30),.data_out(wire_d16_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1632(.data_in(wire_d16_31),.data_out(wire_d16_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1633(.data_in(wire_d16_32),.data_out(wire_d16_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1634(.data_in(wire_d16_33),.data_out(d_out16),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance170(.data_in(d_in17),.data_out(wire_d17_0),.clk(clk),.rst(rst));            //channel 18
	encoder #(.WIDTH(WIDTH)) encoder_instance171(.data_in(wire_d17_0),.data_out(wire_d17_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance172(.data_in(wire_d17_1),.data_out(wire_d17_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance173(.data_in(wire_d17_2),.data_out(wire_d17_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance174(.data_in(wire_d17_3),.data_out(wire_d17_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance175(.data_in(wire_d17_4),.data_out(wire_d17_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance176(.data_in(wire_d17_5),.data_out(wire_d17_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance177(.data_in(wire_d17_6),.data_out(wire_d17_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance178(.data_in(wire_d17_7),.data_out(wire_d17_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance179(.data_in(wire_d17_8),.data_out(wire_d17_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1710(.data_in(wire_d17_9),.data_out(wire_d17_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1711(.data_in(wire_d17_10),.data_out(wire_d17_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1712(.data_in(wire_d17_11),.data_out(wire_d17_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1713(.data_in(wire_d17_12),.data_out(wire_d17_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1714(.data_in(wire_d17_13),.data_out(wire_d17_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1715(.data_in(wire_d17_14),.data_out(wire_d17_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1716(.data_in(wire_d17_15),.data_out(wire_d17_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1717(.data_in(wire_d17_16),.data_out(wire_d17_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1718(.data_in(wire_d17_17),.data_out(wire_d17_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1719(.data_in(wire_d17_18),.data_out(wire_d17_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1720(.data_in(wire_d17_19),.data_out(wire_d17_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1721(.data_in(wire_d17_20),.data_out(wire_d17_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1722(.data_in(wire_d17_21),.data_out(wire_d17_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1723(.data_in(wire_d17_22),.data_out(wire_d17_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1724(.data_in(wire_d17_23),.data_out(wire_d17_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1725(.data_in(wire_d17_24),.data_out(wire_d17_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1726(.data_in(wire_d17_25),.data_out(wire_d17_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1727(.data_in(wire_d17_26),.data_out(wire_d17_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1728(.data_in(wire_d17_27),.data_out(wire_d17_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1729(.data_in(wire_d17_28),.data_out(wire_d17_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1730(.data_in(wire_d17_29),.data_out(wire_d17_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1731(.data_in(wire_d17_30),.data_out(wire_d17_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1732(.data_in(wire_d17_31),.data_out(wire_d17_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1733(.data_in(wire_d17_32),.data_out(wire_d17_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1734(.data_in(wire_d17_33),.data_out(d_out17),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance180(.data_in(d_in18),.data_out(wire_d18_0),.clk(clk),.rst(rst));            //channel 19
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181(.data_in(wire_d18_0),.data_out(wire_d18_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance182(.data_in(wire_d18_1),.data_out(wire_d18_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance183(.data_in(wire_d18_2),.data_out(wire_d18_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance184(.data_in(wire_d18_3),.data_out(wire_d18_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance185(.data_in(wire_d18_4),.data_out(wire_d18_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance186(.data_in(wire_d18_5),.data_out(wire_d18_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance187(.data_in(wire_d18_6),.data_out(wire_d18_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance188(.data_in(wire_d18_7),.data_out(wire_d18_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance189(.data_in(wire_d18_8),.data_out(wire_d18_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1810(.data_in(wire_d18_9),.data_out(wire_d18_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1811(.data_in(wire_d18_10),.data_out(wire_d18_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1812(.data_in(wire_d18_11),.data_out(wire_d18_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1813(.data_in(wire_d18_12),.data_out(wire_d18_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1814(.data_in(wire_d18_13),.data_out(wire_d18_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1815(.data_in(wire_d18_14),.data_out(wire_d18_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1816(.data_in(wire_d18_15),.data_out(wire_d18_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1817(.data_in(wire_d18_16),.data_out(wire_d18_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1818(.data_in(wire_d18_17),.data_out(wire_d18_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1819(.data_in(wire_d18_18),.data_out(wire_d18_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1820(.data_in(wire_d18_19),.data_out(wire_d18_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1821(.data_in(wire_d18_20),.data_out(wire_d18_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1822(.data_in(wire_d18_21),.data_out(wire_d18_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1823(.data_in(wire_d18_22),.data_out(wire_d18_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1824(.data_in(wire_d18_23),.data_out(wire_d18_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1825(.data_in(wire_d18_24),.data_out(wire_d18_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1826(.data_in(wire_d18_25),.data_out(wire_d18_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1827(.data_in(wire_d18_26),.data_out(wire_d18_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1828(.data_in(wire_d18_27),.data_out(wire_d18_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1829(.data_in(wire_d18_28),.data_out(wire_d18_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1830(.data_in(wire_d18_29),.data_out(wire_d18_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1831(.data_in(wire_d18_30),.data_out(wire_d18_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1832(.data_in(wire_d18_31),.data_out(wire_d18_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1833(.data_in(wire_d18_32),.data_out(wire_d18_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1834(.data_in(wire_d18_33),.data_out(d_out18),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance190(.data_in(d_in19),.data_out(wire_d19_0),.clk(clk),.rst(rst));            //channel 20
	invertion #(.WIDTH(WIDTH)) invertion_instance191(.data_in(wire_d19_0),.data_out(wire_d19_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance192(.data_in(wire_d19_1),.data_out(wire_d19_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance193(.data_in(wire_d19_2),.data_out(wire_d19_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance194(.data_in(wire_d19_3),.data_out(wire_d19_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance195(.data_in(wire_d19_4),.data_out(wire_d19_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance196(.data_in(wire_d19_5),.data_out(wire_d19_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance197(.data_in(wire_d19_6),.data_out(wire_d19_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance198(.data_in(wire_d19_7),.data_out(wire_d19_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance199(.data_in(wire_d19_8),.data_out(wire_d19_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1910(.data_in(wire_d19_9),.data_out(wire_d19_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1911(.data_in(wire_d19_10),.data_out(wire_d19_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1912(.data_in(wire_d19_11),.data_out(wire_d19_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1913(.data_in(wire_d19_12),.data_out(wire_d19_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1914(.data_in(wire_d19_13),.data_out(wire_d19_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1915(.data_in(wire_d19_14),.data_out(wire_d19_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1916(.data_in(wire_d19_15),.data_out(wire_d19_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1917(.data_in(wire_d19_16),.data_out(wire_d19_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1918(.data_in(wire_d19_17),.data_out(wire_d19_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1919(.data_in(wire_d19_18),.data_out(wire_d19_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1920(.data_in(wire_d19_19),.data_out(wire_d19_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1921(.data_in(wire_d19_20),.data_out(wire_d19_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1922(.data_in(wire_d19_21),.data_out(wire_d19_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1923(.data_in(wire_d19_22),.data_out(wire_d19_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1924(.data_in(wire_d19_23),.data_out(wire_d19_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1925(.data_in(wire_d19_24),.data_out(wire_d19_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1926(.data_in(wire_d19_25),.data_out(wire_d19_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1927(.data_in(wire_d19_26),.data_out(wire_d19_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1928(.data_in(wire_d19_27),.data_out(wire_d19_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1929(.data_in(wire_d19_28),.data_out(wire_d19_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1930(.data_in(wire_d19_29),.data_out(wire_d19_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1931(.data_in(wire_d19_30),.data_out(wire_d19_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1932(.data_in(wire_d19_31),.data_out(wire_d19_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1933(.data_in(wire_d19_32),.data_out(wire_d19_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1934(.data_in(wire_d19_33),.data_out(d_out19),.clk(clk),.rst(rst));


endmodule