// SPDX-License-Identifier: Apache-2.0
// Copyright 2019-2020 Western Digital Corporation or its affiliates.
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
// http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

//********************************************************************************
// $Id$
//
// Function: SweRVolf tech-agnostic toplevel
// Comments:
//
//********************************************************************************

`default_nettype none
module swervolf_core
  #(parameter bootrom_file  = "",
    parameter clk_freq_hz = 0)
   (input wire 	clk,
    input wire 	       rstn,
    input wire 	       dmi_reg_en,
    input wire [6:0]   dmi_reg_addr,
    input wire 	       dmi_reg_wr_en,
    input wire [31:0]  dmi_reg_wdata,
    output wire [31:0] dmi_reg_rdata,
    input wire 	       dmi_hard_reset,
    output wire        o_flash_sclk,
    output wire        o_flash_cs_n,
    output wire        o_flash_mosi,
    input wire 	       i_flash_miso,
    input wire 	       i_uart_rx,
    output wire        o_uart_tx,
    output wire [5:0]  o_ram_awid,
    output wire [31:0] o_ram_awaddr,
    output wire [7:0]  o_ram_awlen,
    output wire [2:0]  o_ram_awsize,
    output wire [1:0]  o_ram_awburst,
    output wire        o_ram_awlock,
    output wire [3:0]  o_ram_awcache,
    output wire [2:0]  o_ram_awprot,
    output wire [3:0]  o_ram_awregion,
    output wire [3:0]  o_ram_awqos,
    output wire        o_ram_awvalid,
    input wire 	       i_ram_awready,
    output wire [5:0]  o_ram_arid,
    output wire [31:0] o_ram_araddr,
    output wire [7:0]  o_ram_arlen,
    output wire [2:0]  o_ram_arsize,
    output wire [1:0]  o_ram_arburst,
    output wire        o_ram_arlock,
    output wire [3:0]  o_ram_arcache,
    output wire [2:0]  o_ram_arprot,
    output wire [3:0]  o_ram_arregion,
    output wire [3:0]  o_ram_arqos,
    output wire        o_ram_arvalid,
    input wire 	       i_ram_arready,
    output wire [63:0] o_ram_wdata,
    output wire [7:0]  o_ram_wstrb,
    output wire        o_ram_wlast,
    output wire        o_ram_wvalid,
    input wire 	       i_ram_wready,
    input wire [5:0]   i_ram_bid,
    input wire [1:0]   i_ram_bresp,
    input wire 	       i_ram_bvalid,
    output wire        o_ram_bready,
    input wire [5:0]   i_ram_rid,
    input wire [63:0]  i_ram_rdata,
    input wire [1:0]   i_ram_rresp,
    input wire 	       i_ram_rlast,
    input wire 	       i_ram_rvalid,
    output wire        o_ram_rready,
    input wire 	       i_ram_init_done,
    input wire 	       i_ram_init_error,
    input wire [63:0]  i_gpio,
    output wire [63:0] o_gpio);

   localparam BOOTROM_SIZE = 32'h1000;

   wire        rst_n = rstn;
   wire        timer_irq;
   wire        uart_irq;
   wire        spi0_irq;
   wire        sw_irq4;
   wire        sw_irq3;
   wire        nmi_int;
   
    wire [5:0]  ram_awid;
     wire [31:0] ram_awaddr;
     wire [7:0]  ram_awlen;
     wire [2:0]  ram_awsize;
     wire [1:0]  ram_awburst;
     wire        ram_awlock;
     wire [3:0]  ram_awcache;
     wire [2:0]  ram_awprot;
     wire [3:0]  ram_awregion;
     wire [3:0]  ram_awqos;
     wire        ram_awvalid;
     wire        ram_awready;
     wire [5:0]  ram_arid;
     wire [31:0] ram_araddr;
     wire [7:0]  ram_arlen;
     wire [2:0]  ram_arsize;
     wire [1:0]  ram_arburst;
     wire        ram_arlock;
     wire [3:0]  ram_arcache;
     wire [2:0]  ram_arprot;
     wire [3:0]  ram_arregion;
     wire [3:0]  ram_arqos;
     wire        ram_arvalid;
     wire        ram_arready;
     wire [63:0] ram_wdata;
     wire [7:0]  ram_wstrb;
     wire        ram_wlast;
     wire        ram_wvalid;
     wire        ram_wready;
     wire [5:0]  ram_bid;
     wire [1:0]  ram_bresp;
     wire        ram_bvalid;
     wire        ram_bready;
     wire [5:0]  ram_rid;
     wire [63:0] ram_rdata;
     wire [1:0]  ram_rresp;
     wire        ram_rlast;
     wire        ram_rvalid;
     wire        ram_rready;
  
 //    wire        dmi_reg_en;
 //    wire [6:0]  dmi_reg_addr;
 //    wire        dmi_reg_wr_en;
 //    wire [31:0] dmi_reg_wdata;
 //    wire [31:0] dmi_reg_rdata;
  //   wire        dmi_hard_reset;
   
   
   wire [31:0] nmi_vec;

//`include "axi_intercon.vh"

   assign o_ram_awid     = ram_awid;
   assign o_ram_awaddr   = ram_awaddr;
   assign o_ram_awlen    = ram_awlen;
   assign o_ram_awsize   = ram_awsize;
   assign o_ram_awburst  = ram_awburst;
   assign o_ram_awlock   = ram_awlock;
   assign o_ram_awcache  = ram_awcache;
   assign o_ram_awprot   = ram_awprot;
   assign o_ram_awregion = ram_awregion;
   assign o_ram_awqos    = ram_awqos;
   assign o_ram_awvalid  = ram_awvalid;
   assign ram_awready    = i_ram_awready;
   assign o_ram_arid     = ram_arid;
   assign o_ram_araddr   = ram_araddr;
   assign o_ram_arlen    = ram_arlen;
   assign o_ram_arsize   = ram_arsize;
   assign o_ram_arburst  = ram_arburst;
   assign o_ram_arlock   = ram_arlock;
   assign o_ram_arcache  = ram_arcache;
   assign o_ram_arprot   = ram_arprot;
   assign o_ram_arregion = ram_arregion;
   assign o_ram_arqos    = ram_arqos;
   assign o_ram_arvalid  = ram_arvalid;
   assign ram_arready    = i_ram_arready;
   assign o_ram_wdata    = ram_wdata;
   assign o_ram_wstrb    = ram_wstrb;
   assign o_ram_wlast    = ram_wlast;
   assign o_ram_wvalid   = ram_wvalid;
   assign ram_wready     = i_ram_wready;
   assign ram_bid        = i_ram_bid;
   assign ram_bresp      = i_ram_bresp;
   assign ram_bvalid     = i_ram_bvalid;
   assign o_ram_bready   = ram_bready;
   assign ram_rid        = i_ram_rid;
   assign ram_rdata      = i_ram_rdata;
   assign ram_rresp      = i_ram_rresp;
   assign ram_rlast      = i_ram_rlast;
   assign ram_rvalid     = i_ram_rvalid;
   assign o_ram_rready   = ram_rready;

   wire 		      wb_clk = clk;
   wire 		      wb_rst = ~rst_n;

//`include "wb_intercon.vh"

   wire [15:2] 		       wb_adr;
   wire wb_m2s_io_adr;
   wire wb_m2s_io_cti;
   wire wb_m2s_io_bte;
   
   
   assign wb_m2s_io_adr = {16'd0,wb_adr,2'b00};
   assign wb_m2s_io_cti = 3'b000;
   assign wb_m2s_io_bte = 2'b00;

wire wb_m2s_io_dat;
wire wb_m2s_io_sel;
wire wb_m2s_io_we;
wire wb_m2s_io_cyc;
wire wb_m2s_io_stb;
wire wb_s2m_io_dat;
wire wb_s2m_io_ack;
wire wb_s2m_io_err;

wire wb_s2m_io;


wire  io_awaddr;
wire io_awid;
wire io_awvalid;
wire io_awready;

wire [15:0] io_araddr;
wire io_arid;
wire io_arvalid;
wire io_arready;

wire io_wdata;
wire io_wstrb;
wire io_wvalid;
wire io_wready;

wire io_bid;
wire io_bresp;
wire io_bvalid;
wire io_bready;

wire io_rdata;
wire io_rid;
wire io_rresp;
wire io_rlast;
wire io_rvalid;
wire io_rready;

wire    wb_mem_wrapper;


   axi2wb
     #(.AW (16),
       .IW (4+3))
   axi2wb
     (
      .i_clk       (clk),
      .i_rst       (~rst_n),
      .o_wb_adr    (wb_adr),
      .o_wb_dat    (wb_m2s_io_dat),
      .o_wb_sel    (wb_m2s_io_sel),
      .o_wb_we     (wb_m2s_io_we),
      .o_wb_cyc    (wb_m2s_io_cyc),
      .o_wb_stb    (wb_m2s_io_stb),
      .i_wb_rdt    (wb_s2m_io_dat),
      .i_wb_ack    (wb_s2m_io_ack),
      .i_wb_err    (wb_s2m_io_err),

      .i_awaddr    (io_awaddr),
      .i_awid      (io_awid),
      .i_awvalid   (io_awvalid),
      .o_awready   (io_awready),

      .i_araddr    (io_araddr[15:0]),
      .i_arid      (io_arid),
      .i_arvalid   (io_arvalid),
      .o_arready   (io_arready),

      .i_wdata     (io_wdata),
      .i_wstrb     (io_wstrb),
      .i_wvalid    (io_wvalid),
      .o_wready    (io_wready),

      .o_bid       (io_bid),
      .o_bresp     (io_bresp),
      .o_bvalid    (io_bvalid),
      .i_bready    (io_bready),

      .o_rdata     (io_rdata),
      .o_rid       (io_rid),
      .o_rresp     (io_rresp),
      .o_rlast     (io_rlast),
      .o_rvalid    (io_rvalid),
      .i_rready    (io_rready));

wire wb_m2s_rom_adr;
wire wb_m2s_rom_dat;
wire wb_m2s_rom_sel;
wire wb_m2s_rom_we;
wire wb_m2s_rom_cyc;
wire wb_m2s_rom_stb;
wire wb_s2m_rom_dat;
wire wb_s2m_rom_ack;


   wb_mem_wrapper
     #(.MEM_SIZE  (BOOTROM_SIZE),
       .INIT_FILE (bootrom_file))
   bootrom
     (.i_clk    (wb_clk),
      .i_rst    (wb_rst),
   //   .i_wb_adr (wb_m2s_rom_adr[$clog2(BOOTROM_SIZE)-1:2]),
      .i_wb_dat (wb_m2s_rom_dat),
      .i_wb_sel (wb_m2s_rom_sel),
      .i_wb_we  (wb_m2s_rom_we),
      .i_wb_cyc (wb_m2s_rom_cyc),
      .i_wb_stb (wb_m2s_rom_stb),
      .o_wb_rdt (wb_s2m_rom_dat),
      .o_wb_ack (wb_s2m_rom_ack));

wire wb_s2m_rom_err;
wire wb_s2m_rom_rty;

wire wb_m2s_sys_adr;
wire wb_m2s_sys_dat;
wire wb_m2s_sys_sel;
wire wb_m2s_sys_we;
wire wb_m2s_sys_cyc;
wire wb_m2s_sys_stb;
wire wb_s2m_sys_dat;
wire wb_s2m_sys_ack;
   assign wb_s2m_rom_err = 1'b0;
   assign wb_s2m_rom_rty = 1'b0;

   swervolf_syscon
     #(.clk_freq_hz (clk_freq_hz))
   syscon
     (.i_clk            (clk),
      .i_rst            (wb_rst),

      .i_gpio           (i_gpio),
      .o_gpio           (o_gpio),
      .o_timer_irq      (timer_irq),
      .o_sw_irq3        (sw_irq3),
      .o_sw_irq4        (sw_irq4),
      .i_ram_init_done  (i_ram_init_done),
      .i_ram_init_error (i_ram_init_error),
      .o_nmi_vec        (nmi_vec),
      .o_nmi_int        (nmi_int),

//      .i_wb_adr         (wb_m2s_sys_adr[5:0]),
      .i_wb_dat         (wb_m2s_sys_dat),
      .i_wb_sel         (wb_m2s_sys_sel),
      .i_wb_we          (wb_m2s_sys_we),
      .i_wb_cyc         (wb_m2s_sys_cyc),
      .i_wb_stb         (wb_m2s_sys_stb),
      .o_wb_rdt         (wb_s2m_sys_dat),
      .o_wb_ack         (wb_s2m_sys_ack));


wire wb_s2m_sys_err;
wire wb_s2m_sys_rty;
wire wb_s2m_spi_flash_dat;


wire wb_m2s_spi_flash_we;
wire wb_m2s_spi_flash_cyc;
wire wb_m2s_spi_flash_stb;

wire wb_s2m_spi_flash_ack;


   assign wb_s2m_sys_err = 1'b0;
   assign wb_s2m_sys_rty = 1'b0;

   wire [7:0] 		       spi_rdt;
   assign wb_s2m_spi_flash_dat = {24'd0,spi_rdt};

   simple_spi spi
     (// Wishbone slave interface
      .clk_i  (clk),
      .rst_i  (wb_rst),
      /* Note! Below is a horrible hack that needs some explanation

       The AXI bus is 64-bit and there is no support for telling the slave
       that it just wants to read a part of a 64-bit word.

       On the slave side, the SPI controller has an 8-bit databus.
       So in order to ensure that only one register gets accessed by the 64-bit
       master, the registers are placed 64 bits apart from each other, at
       addresses 0x0, 0x8, 0x10, 0x18 and 0x20 instead of the original 0x0, 0x1,
       0x2, 0x3 and 0x4. This works easy enough by just cutting of the three
       least significant bits of the address before passing it to the slave.

       Now, to complicate things, there is an wb2axi bridge that converts 64-bit
       datapath into 32 bits between the master and slave. Since the master
       can't indicate what part of the 64-bit word it actually wants to read,
       every 64-bit read gets turned into two consecutive 32-bit reads on the
       wishbone side.

       E.g. a read from address 0x8 on the 64-bit AXI side gets turned into two
       read operations from 0x8 and 0xc on the 32-bit Wishbone side.

       Usually this is not a real problem. Just a bit inefficient. But in this
       case we have the SPDR register that holds the incoming data. When we
       read a byte from that register, it is removed from the SPI FIFO and
       can't be read again. Now, if we read from this register two times, every
       time we just want to read a byte, this means that we throw away half of
       our received data and things break down.

       Writes are no problem since, there is a byte mask that tells which
       bytes to really write

       In order to work around this issue, we look at bit 2. Why? Because a
       64-bit read to any of the mapped registers (which are 64-bit aligned)
       will get turned into two read operations. First, one against the actual
       register, and then an additional read from address+4, i.e. address, but
       with bit 2 set as well. We still need to respond to the second read but
       it doesn't matter what data it contains since no one should look at it.

       So, when we see a read with bit 2 set, we redirect this access to
       register zero. Doesn't really matter which register as long as we pick
       a non-volatile one.

       TODO: Make something sensible here instead
       */
 //     .adr_i  (wb_m2s_spi_flash_adr[2] ? 3'd0 : wb_m2s_spi_flash_adr[5:3]),
 //     .dat_i  (wb_m2s_spi_flash_dat[7:0]),
      .we_i   (wb_m2s_spi_flash_we),
      .cyc_i  (wb_m2s_spi_flash_cyc),
      .stb_i  (wb_m2s_spi_flash_stb),
      .dat_o  (spi_rdt),
      .ack_o  (wb_s2m_spi_flash_ack),
      .inta_o (spi0_irq),
      // SPI interface
      .sck_o  (o_flash_sclk),
     // .ss_o   (o_flash_cs_n),
      .mosi_o (o_flash_mosi),
      .miso_i (i_flash_miso));
wire wb_s2m_spi_flash_err;
wire wb_s2m_spi_flash_rty;
   assign wb_s2m_spi_flash_err = 1'b0;
   assign wb_s2m_spi_flash_rty = 1'b0;

   wire [7:0] 		       uart_rdt;
   
   wire wb_s2m_uart_dat;
   wire wb_s2m_uart_err;
   wire wb_s2m_uart_rty;
   
   
   assign wb_s2m_uart_dat = {24'd0, uart_rdt};
   assign wb_s2m_uart_err = 1'b0;
   assign wb_s2m_uart_rty = 1'b0;

   uart_top uart16550_0
     (// Wishbone slave interface
      .wb_clk_i	(clk),
      .wb_rst_i	(~rst_n),
  //    .wb_adr_i	(wb_m2s_uart_adr[4:2]),
 //     .wb_dat_i	(wb_m2s_uart_dat[7:0]),
 // //    .wb_we_i	(wb_m2s_uart_we),
 //     .wb_cyc_i	(wb_m2s_uart_cyc),
 //     .wb_stb_i	(wb_m2s_uart_stb),
      .wb_sel_i	(4'b0), // Not used in 8-bit mode
      .wb_dat_o	(uart_rdt),
 //     .wb_ack_o	(wb_s2m_uart_ack),

      // Outputs
      .int_o     (uart_irq),
      .stx_pad_o (o_uart_tx),
      .rts_pad_o (),
      .dtr_pad_o (),

      // Inputs
      .srx_pad_i (i_uart_rx),
      .cts_pad_i (1'b0),
      .dsr_pad_i (1'b0),
      .ri_pad_i  (1'b0),
      .dcd_pad_i (1'b0));

  //  swerv_wrapper_dmi rvtop
  //    (
  //     .clk     (clk),
  //     .rst_l   (rstn),
  //     .dbg_rst_l   (rstn),
  //     .rst_vec (31'h40000000),
  //     .nmi_int (nmi_int),
  //     .nmi_vec (nmi_vec[31:1]),
// 
  //     .trace_rv_i_insn_ip      (),
  //     .trace_rv_i_address_ip   (),
  //     .trace_rv_i_valid_ip     (),
  //     .trace_rv_i_exception_ip (),
  //     .trace_rv_i_ecause_ip    (),
  //     .trace_rv_i_interrupt_ip (),
  //     .trace_rv_i_tval_ip      (),

      // Bus signals
      //-------------------------- LSU AXI signals--------------------------
  //    .lsu_axi_awvalid  (lsu_awvalid),
  //    .lsu_axi_awready  (lsu_awready),
   //   .lsu_axi_awid     (lsu_awid   ),
   //   .lsu_axi_awaddr   (lsu_awaddr ),
  //    .lsu_axi_awregion (lsu_awregion),
  //    .lsu_axi_awlen    (lsu_awlen  ),
  //    .lsu_axi_awsize   (lsu_awsize ),
 //     .lsu_axi_awburst  (lsu_awburst),
 //     .lsu_axi_awlock   (lsu_awlock ),
  //    .lsu_axi_awcache  (lsu_awcache),
  //    .lsu_axi_awprot   (lsu_awprot ),
  //    .lsu_axi_awqos    (lsu_awqos  ),

  //    .lsu_axi_wvalid   (lsu_wvalid),
   //   .lsu_axi_wready   (lsu_wready),
   //   .lsu_axi_wdata    (lsu_wdata),
   //   .lsu_axi_wstrb    (lsu_wstrb),
   //   .lsu_axi_wlast    (lsu_wlast),

  //    .lsu_axi_bvalid   (lsu_bvalid),
  //    .lsu_axi_bready   (lsu_bready),
  //    .lsu_axi_bresp    (lsu_bresp ),
   //   .lsu_axi_bid      (lsu_bid   ),

 //     .lsu_axi_arvalid  (lsu_arvalid ),
 //     .lsu_axi_arready  (lsu_arready ),
 //     .lsu_axi_arid     (lsu_arid    ),
  //    .lsu_axi_araddr   (lsu_araddr  ),
  //    .lsu_axi_arregion (lsu_arregion),
  //    .lsu_axi_arlen    (lsu_arlen   ),
  //    .lsu_axi_arsize   (lsu_arsize  ),
  //    .lsu_axi_arburst  (lsu_arburst ),
  //    .lsu_axi_arlock   (lsu_arlock  ),
 //     .lsu_axi_arcache  (lsu_arcache ),
  //    .lsu_axi_arprot   (lsu_arprot  ),
//      .lsu_axi_arqos    (lsu_arqos   ),

 //     .lsu_axi_rvalid   (lsu_rvalid),
 //     .lsu_axi_rready   (lsu_rready),
 //     .lsu_axi_rid      (lsu_rid   ),
 //     .lsu_axi_rdata    (lsu_rdata ),
 //     .lsu_axi_rresp    (lsu_rresp ),
 //     .lsu_axi_rlast    (lsu_rlast ),

//       //-------------------------- IFU AXI signals--------------------------
//       .ifu_axi_awvalid  (),
//       .ifu_axi_awready  (1'b0),
//       .ifu_axi_awid     (),
//       .ifu_axi_awaddr   (),
//       .ifu_axi_awregion (),
//       .ifu_axi_awlen    (),
//       .ifu_axi_awsize   (),
//       .ifu_axi_awburst  (),
//       .ifu_axi_awlock   (),
//       .ifu_axi_awcache  (),
//       .ifu_axi_awprot   (),
//       .ifu_axi_awqos    (),
// 
//       .ifu_axi_wvalid   (),
//       .ifu_axi_wready   (1'b0),
//       .ifu_axi_wdata    (),
//       .ifu_axi_wstrb    (),
//       .ifu_axi_wlast    (),
// 
//       .ifu_axi_bvalid   (1'b0),
//       .ifu_axi_bready   (),
//       .ifu_axi_bresp    (2'b00),
//       .ifu_axi_bid      (3'd0),
// 
//   //    .ifu_axi_arvalid  (ifu_arvalid ),
//   //    .ifu_axi_arready  (ifu_arready ),
//   //    .ifu_axi_arid     (ifu_arid    ),
//   //    .ifu_axi_araddr   (ifu_araddr  ),
//   //    .ifu_axi_arregion (ifu_arregion),
//   //    .ifu_axi_arlen    (ifu_arlen   ),
//   //    .ifu_axi_arsize   (ifu_arsize  ),
//   //    .ifu_axi_arburst  (ifu_arburst ),
//   //    .ifu_axi_arlock   (ifu_arlock  ),
//   //    .ifu_axi_arcache  (ifu_arcache ),
//   //    .ifu_axi_arprot   (ifu_arprot  ),
//    //   .ifu_axi_arqos    (ifu_arqos   ),
// 
// //      .ifu_axi_rvalid   (ifu_rvalid),
// //      .ifu_axi_rready   (ifu_rready),
// //ifu_axi_rid      (ifu_rid   ),
// //      .ifu_axi_rdata    (ifu_rdata ),
//  //     .ifu_axi_rresp    (ifu_rresp ),
//   //    .ifu_axi_rlast    (ifu_rlast ),
// 
//       //-------------------------- SB AXI signals-------------------------
//  //     .sb_axi_awvalid  (sb_awvalid ),
//  //     .sb_axi_awready  (sb_awready ),
//  //     .sb_axi_awid     (sb_awid    ),
// //      .sb_axi_awaddr   (sb_awaddr  ),
//  //     .sb_axi_awregion (sb_awregion),
//  //     .sb_axi_awlen    (sb_awlen   ),
//  //     .sb_axi_awsize   (sb_awsize  ),
//  //     .sb_axi_awburst  (sb_awburst ),
//  //     .sb_axi_awlock   (sb_awlock  ),
//  //     .sb_axi_awcache  (sb_awcache ),
//   //    .sb_axi_awprot   (sb_awprot  ),
//  //     .sb_axi_awqos    (sb_awqos   ),
//   //    .sb_axi_wvalid   (sb_wvalid  ),
// //      .sb_axi_wready   (sb_wready  ),
// //      .sb_axi_wdata    (sb_wdata   ),
// //      .sb_axi_wstrb    (sb_wstrb   ),
// //      .sb_axi_wlast    (sb_wlast   ),
// //      .sb_axi_bvalid   (sb_bvalid  ),
// //      .sb_axi_bready   (sb_bready  ),
//  //     .sb_axi_bresp    (sb_bresp   ),
// //      .sb_axi_bid      (sb_bid     ),
// //      .sb_axi_arvalid  (sb_arvalid ),
//  //     .sb_axi_arready  (sb_arready ),
//     //  .sb_axi_arid     (sb_arid    ),
//   //    .sb_axi_araddr   (sb_araddr  ),
//   //    .sb_axi_arregion (sb_arregion),
//   //    .sb_axi_arlen    (sb_arlen   ),
//   //    .sb_axi_arsize   (sb_arsize  ),
//   //    .sb_axi_arburst  (sb_arburst ),
//   //    .sb_axi_arlock   (sb_arlock  ),
//   //    .sb_axi_arcache  (sb_arcache ),
//   //    .sb_axi_arprot   (sb_arprot  ),
//   //    .sb_axi_arqos    (sb_arqos   ),
// //.sb_axi_rvalid   (sb_rvalid  ),
// //      .sb_axi_rready   (sb_rready  ),
// //.sb_axi_rid      (sb_rid     ),
//  //     .sb_axi_rdata    (sb_rdata   ),
//  //     .sb_axi_rresp    (sb_rresp   ),
//  //     .sb_axi_rlast    (sb_rlast   ),
// 
//       //-------------------------- DMA AXI signals--------------------------
//       .dma_axi_awvalid  (1'b0),
//       .dma_axi_awready  (),
//       .dma_axi_awid     (1'd0),
//       .dma_axi_awaddr   (32'd0),
//       .dma_axi_awsize   (3'd0),
//       .dma_axi_awprot   (3'd0),
//       .dma_axi_awlen    (8'd0),
//       .dma_axi_awburst  (2'd0),
// 
//       .dma_axi_wvalid   (1'b0),
//       .dma_axi_wready   (),
//       .dma_axi_wdata    (64'd0),
//       .dma_axi_wstrb    (8'd0),
//       .dma_axi_wlast    (1'b0),
// 
//       .dma_axi_bvalid   (),
//       .dma_axi_bready   (1'b0),
//       .dma_axi_bresp    (),
//       .dma_axi_bid      (),
// 
//       .dma_axi_arvalid  (1'b0),
//       .dma_axi_arready  (),
//       .dma_axi_arid     (1'd0),
//       .dma_axi_araddr   (32'd0),
//       .dma_axi_arsize   (3'd0),
//       .dma_axi_arprot   (3'd0),
//       .dma_axi_arlen    (8'd0),
//       .dma_axi_arburst  (2'd0),
// 
//       .dma_axi_rvalid   (),
//       .dma_axi_rready   (1'b0),
//       .dma_axi_rid      (),
//       .dma_axi_rdata    (),
//       .dma_axi_rresp    (),
//       .dma_axi_rlast    (),
// 
//       // clk ratio signals
//       .lsu_bus_clk_en (1'b1),
//       .ifu_bus_clk_en (1'b1),
//       .dbg_bus_clk_en (1'b1),
//       .dma_bus_clk_en (1'b1),
// 
//       .timer_int (timer_irq),
//       .extintsrc_req ({4'd0, sw_irq4, sw_irq3, spi0_irq, uart_irq}),
// 
//       .dec_tlu_perfcnt0 (),
//       .dec_tlu_perfcnt1 (),
//       .dec_tlu_perfcnt2 (),
//       .dec_tlu_perfcnt3 (),
// 
//       .dmi_reg_rdata    (dmi_reg_rdata),
//       .dmi_reg_wdata    (dmi_reg_wdata),
//       .dmi_reg_addr     (dmi_reg_addr),
//       .dmi_reg_en       (dmi_reg_en),
//       .dmi_reg_wr_en    (dmi_reg_wr_en),
//       .dmi_hard_reset   (dmi_hard_reset),
// 
//       .mpc_debug_halt_req (1'b0),
//       .mpc_debug_run_req  (1'b0),
//       .mpc_reset_run_req  (1'b1),
//       .mpc_debug_halt_ack (),
//       .mpc_debug_run_ack  (),
//       .debug_brkpt_status (),
// 
//       .i_cpu_halt_req      (1'b0),
//       .o_cpu_halt_ack      (),
//       .o_cpu_halt_status   (),
//       .o_debug_mode_status (),
//       .i_cpu_run_req       (1'b0),
//       .o_cpu_run_ack       (),
// 
//       .scan_mode  (1'b0),
//       .mbist_mode (1'b0));
// 
 endmodule
