`define CLB_X 66
`define CLB_Y 78
`define A2F_BWID  20 * 2 *`CLB_X + 20 * 2 * `CLB_Y
`define DEF_BWID  40 * 2 *`CLB_X + 40 * 2 * `CLB_Y
`define PLL_NUM 4
`define SCAN_NUM 9
//*************************
`define FAB_IO_NUM 380  
`define FAB_GBOX_NUM `FAB_IO_NUM 
//*************************
`define GBOX_DWID 10
`define FAB_GBOX_DWID `FAB_GBOX_NUM * `GBOX_DWID
//*************************

