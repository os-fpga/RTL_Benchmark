-------------------------------------------------------------------------------
--
-- GCpad controller core
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- $Id: gcpad_sampler-c.vhd,v 1.1 2004-10-08 21:19:17 arniml Exp $
--
-------------------------------------------------------------------------------

configuration gcpad_sampler_rtl_c0 of gcpad_sampler is

  for rtl
  end for;

end gcpad_sampler_rtl_c0;
