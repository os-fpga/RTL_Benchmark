//------------------------------------------------------------------------
// Filename     : atcbusdec200_config.vh
// Description  : specify AHB-Lite slave configurations
//------------------------------------------------------------------------
`ifdef ATCBUSDEC200_CONFIG_VH
`else
`define ATCBUSDEC200_CONFIG_VH

// Specify AHB slaves according to the SoC configuration
`include "ae350_config.vh"
`include "ae350_const.vh"


`define	ATCBUSDEC200_ADDR_DECODE_WIDTH 29
//`define ATCBUSDEC200_DATA_WIDTH_64
//`define ATCBUSDEC200_DATA_WIDTH_128

`define ATCBUSDEC200_SLV0_SUPPORT
`define ATCBUSDEC200_SLV1_SUPPORT
`ifdef AE350_SMC_SUPPORT
	`define ATCBUSDEC200_SLV2_SUPPORT
`endif
`ifdef AE350_LCDC_SUPPORT
	`define ATCBUSDEC200_SLV3_SUPPORT
`endif
`ifdef AE350_MAC_SUPPORT
	`define ATCBUSDEC200_SLV4_SUPPORT
`endif

//`define ATCBUSDEC200_SLV5_SUPPORT
//`define ATCBUSDEC200_SLV6_SUPPORT
//`define ATCBUSDEC200_SLV7_SUPPORT
//`define ATCBUSDEC200_SLV8_SUPPORT
//`define ATCBUSDEC200_SLV9_SUPPORT


//-------------------------------------------------
// AHB Slave Base Address
//-------------------------------------------------
`define ATCBUSDEC200_SLV0_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0000_0000 //1MB
`define ATCBUSDEC200_SLV1_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h10000000
`define ATCBUSDEC200_SLV2_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0040_0000 //1MB	SMC
`define ATCBUSDEC200_SLV3_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0020_0000 //1MB	LCDC
`define ATCBUSDEC200_SLV4_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0010_0000 //1MB	MAC
//`define ATCBUSDEC200_SLV5_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0050_0000 //1MB	L2C Control Slave Port
//`define ATCBUSDEC200_SLV6_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0400_0000 //32MB 	PLIC
//`define ATCBUSDEC200_SLV7_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0600_0000 //1MB	PLMT
//`define ATCBUSDEC200_SLV8_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0680_0000 //1MB	PLDM
//`define ATCBUSDEC200_SLV9_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0640_0000 //4MB	PLIC_SW
 // 64
//`define ATCBUSDEC200_SLV9_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0400_0000  //16MB
//`define ATCBUSDEC200_SLV10_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0500_0000 //16MB
//`define ATCBUSDEC200_SLV11_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0040_0000 //1MB
//`define ATCBUSDEC200_SLV12_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0700_0000 //4MB
//`define ATCBUSDEC200_SLV13_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0740_0000 //4MB
//`define ATCBUSDEC200_SLV14_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0780_0000 //4MB 
//`define ATCBUSDEC200_SLV15_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h07c0_0000 //4MB
//// 128
//`define ATCBUSDEC200_SLV16_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0800_0000 //8MB
//`define ATCBUSDEC200_SLV17_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0880_0000 //8MB
//`define ATCBUSDEC200_SLV18_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0900_0000 //8MB
//`define ATCBUSDEC200_SLV19_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0980_0000 //8MB
//`define ATCBUSDEC200_SLV20_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0a00_0000 //8MB
//`define ATCBUSDEC200_SLV21_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0a80_0000 //8MB
//`define ATCBUSDEC200_SLV22_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0b00_0000 //8MB
//`define ATCBUSDEC200_SLV23_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0b80_0000 //8MB
//`define ATCBUSDEC200_SLV24_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0c00_0000 //8MB 
//`define ATCBUSDEC200_SLV25_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0c80_0000 //8MB
//`define ATCBUSDEC200_SLV26_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0d00_0000 //8MB
//`define ATCBUSDEC200_SLV27_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0d80_0000 //8MB
//`define ATCBUSDEC200_SLV28_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0e00_0000 //8MB
//`define ATCBUSDEC200_SLV29_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0e80_0000 //8MB
//`define ATCBUSDEC200_SLV30_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0f00_0000 //8MB
//`define ATCBUSDEC200_SLV31_OFFSET `ATCBUSDEC200_ADDR_DECODE_WIDTH'h0f80_0000 //8MB
`define  ATCBUSDEC200_SLV1_SIZE 9
`define  ATCBUSDEC200_SLV2_SIZE 1
`define  ATCBUSDEC200_SLV3_SIZE 1
`define  ATCBUSDEC200_SLV4_SIZE 1
`define  ATCBUSDEC200_SLV5_SIZE 1
//`define  ATCBUSDEC200_SLV6_SIZE 6
//`define  ATCBUSDEC200_SLV7_SIZE 1
//`define  ATCBUSDEC200_SLV8_SIZE 1
//`define  ATCBUSDEC200_SLV9_SIZE 3
//`define  ATCBUSDEC200_SLV9_SIZE 5
//`define ATCBUSDEC200_SLV10_SIZE 5
//`define ATCBUSDEC200_SLV11_SIZE 5
//`define ATCBUSDEC200_SLV12_SIZE 5
//`define ATCBUSDEC200_SLV13_SIZE 5
//`define ATCBUSDEC200_SLV14_SIZE 3
//`define ATCBUSDEC200_SLV15_SIZE 3
//`define ATCBUSDEC200_SLV16_SIZE 3
//`define ATCBUSDEC200_SLV17_SIZE 3
//`define ATCBUSDEC200_SLV18_SIZE 4
//`define ATCBUSDEC200_SLV19_SIZE 4
//`define ATCBUSDEC200_SLV20_SIZE 4
//`define ATCBUSDEC200_SLV21_SIZE 4
//`define ATCBUSDEC200_SLV22_SIZE 4
//`define ATCBUSDEC200_SLV23_SIZE 4
//`define ATCBUSDEC200_SLV24_SIZE 4
//`define ATCBUSDEC200_SLV25_SIZE 4
//`define ATCBUSDEC200_SLV26_SIZE 4
//`define ATCBUSDEC200_SLV27_SIZE 4
//`define ATCBUSDEC200_SLV28_SIZE 4
//`define ATCBUSDEC200_SLV29_SIZE 4
//`define ATCBUSDEC200_SLV30_SIZE 4
//`define ATCBUSDEC200_SLV31_SIZE 4
`endif //ATCBUSDEC200_CONFIG_VH
