parameter imwidth=512;
parameter imheight=512;
