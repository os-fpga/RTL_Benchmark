--
--  Copyright (c) 2003 Launchbird Design Systems, Inc.
--  All rights reserved.
--  
--  Redistribution and use in source and binary forms, with or without modification, are permitted provided that the following conditions are met:
--    Redistributions of source code must retain the above copyright notice, this list of conditions and the following disclaimer.
--    Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the following disclaimer in the documentation and/or other materials provided with the distribution.
--  
--  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES,
--  INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.
--  IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY,
--  OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
--  OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
--  (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--  
--  Overview:
--  
--    Reconfigurable Computing Array (RCA) is a fine-grained array of programmable tiles.
--    Similar to FPGA CLBs, a tile can implement a wide variety of logic functions.
--    But unlike most FPGAs, RCA can be partially reconfigured dynamically.
--  
--    Also, RCA has no routing fabric.  Instead, the square tiles communicate directly
--    with their nearest neighbor (N, S, W, E), providing fast, deterministic timing and 
--    far greater logic density compared with FPGAs.
--  
--    Each tile implements a programmable 4-bit input to 4-bit output function.
--  
--  Interface:
--  
--    Each side of the array comprises 2 N-bit data buses for a total of 8 buses:
--    north_i, north_o, south_i, south_o, west_i, west_o, east_i, and east_o.
--    The 0 bit in each bus corresponds to northern most or western most tile.
--    All tile registers are synchronized on clock_main_c.
--  
--    Device programming is controlled via the configuration bus.  Each directional datapath
--    of each tile is addressable for configuration.  The configuration addressing format follows:
--  
--      ConfigAddr = {RowSelect, ColSelect, DirSelect} where
--      DirSelect  : 00=north, 01=south, 10=west, 11=east.
--  
--    The configuration data format follows:
--  
--      ConfigData[17]    : Output Select (0=direct, 1=registered)
--      ConfigData[16:14] : Input Select 2  (000=north_in, 001=south_in, 010=west_in, 011=east_in, 100=north_state, 101=south_state, 110=west_state, 111=east_state
--      ConfigData[13:11] : Input Select 1
--      ConfigData[10:8]  : Input Select 0
--      ConfigData[7:0]   : LUT data  {f(7), f(6), f(5), f(4), f(3), f(2), f(1), f(0)}
--  
--  
--  Generated by Confluence 0.6.3  --  Launchbird Design Systems, Inc.  --  www.launchbird.com
--  
--  Build Date : Thu Aug 21 15:06:59 CDT 2003
--  
--  Interface
--  
--    Build Name    : cf_rca_16
--    Clock Domains : clock_config_c  clock_main_c  
--    Vector Input  : config_write_i(1)
--    Vector Input  : config_addr_i(10)
--    Vector Input  : config_data_i(18)
--    Vector Input  : north_i(16)
--    Vector Input  : south_i(16)
--    Vector Input  : west_i(16)
--    Vector Input  : east_i(16)
--    Vector Output : north_o(16)
--    Vector Output : south_o(16)
--    Vector Output : west_o(16)
--    Vector Output : east_o(16)
--  
--  
--  

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end entity cf_rca_16_38;
architecture rtl of cf_rca_16_38 is
signal n1 : unsigned(15 downto 0);
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(15 downto 0);
signal n5 : unsigned(15 downto 0);
signal n6 : unsigned(15 downto 0);
signal n7 : unsigned(15 downto 0);
signal n8 : unsigned(15 downto 0);
signal n9 : unsigned(15 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(15 downto 0);
signal n16 : unsigned(15 downto 0);
begin
n1 <= "1000000000000000";
n2 <= "0100000000000000";
n3 <= "0010000000000000";
n4 <= "0001000000000000";
n5 <= "0000100000000000";
n6 <= "0000010000000000";
n7 <= "0000001000000000";
n8 <= "0000000100000000";
n9 <= "0000000010000000";
n10 <= "0000000001000000";
n11 <= "0000000000100000";
n12 <= "0000000000010000";
n13 <= "0000000000001000";
n14 <= "0000000000000100";
n15 <= "0000000000000010";
n16 <= "0000000000000001";
o16 <= n16;
o15 <= n15;
o14 <= n14;
o13 <= n13;
o12 <= n12;
o11 <= n11;
o10 <= n10;
o9 <= n9;
o8 <= n8;
o7 <= n7;
o6 <= n6;
o5 <= n5;
o4 <= n4;
o3 <= n3;
o2 <= n2;
o1 <= n1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_37 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end entity cf_rca_16_37;
architecture rtl of cf_rca_16_37 is
signal n1 : unsigned(4 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(4 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(4 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(4 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(4 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(15 downto 0);
signal n16 : unsigned(15 downto 0);
signal n17 : unsigned(15 downto 0);
signal n18 : unsigned(15 downto 0);
begin
n1 <= "11001";
n2 <= "1" when i1 = n1 else "0";
n3 <= "11010";
n4 <= "1" when i1 = n3 else "0";
n5 <= "11011";
n6 <= "1" when i1 = n5 else "0";
n7 <= "11100";
n8 <= "1" when i1 = n7 else "0";
n9 <= "11101";
n10 <= "1" when i1 = n9 else "0";
n11 <= "11110";
n12 <= "1" when i1 = n11 else "0";
n13 <= i3 when n12 = "1" else i2;
n14 <= i4 when n10 = "1" else n13;
n15 <= i5 when n8 = "1" else n14;
n16 <= i6 when n6 = "1" else n15;
n17 <= i7 when n4 = "1" else n16;
n18 <= i8 when n2 = "1" else n17;
o1 <= n18;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_36 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end entity cf_rca_16_36;
architecture rtl of cf_rca_16_36 is
signal n1 : unsigned(4 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(4 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(4 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(4 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(15 downto 0);
signal s16_1 : unsigned(15 downto 0);
component cf_rca_16_37 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_37;
begin
n1 <= "10100";
n2 <= "1" when i1 = n1 else "0";
n3 <= "10101";
n4 <= "1" when i1 = n3 else "0";
n5 <= "10110";
n6 <= "1" when i1 = n5 else "0";
n7 <= "10111";
n8 <= "1" when i1 = n7 else "0";
n9 <= "11000";
n10 <= "1" when i1 = n9 else "0";
n11 <= i9 when n10 = "1" else s16_1;
n12 <= i10 when n8 = "1" else n11;
n13 <= i11 when n6 = "1" else n12;
n14 <= i12 when n4 = "1" else n13;
n15 <= i13 when n2 = "1" else n14;
s16 : cf_rca_16_37 port map (i1, i2, i3, i4, i5, i6, i7, i8, s16_1);
o1 <= n15;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_35 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end entity cf_rca_16_35;
architecture rtl of cf_rca_16_35 is
signal n1 : unsigned(4 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(4 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(4 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(4 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(15 downto 0);
signal s16_1 : unsigned(15 downto 0);
component cf_rca_16_36 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_36;
begin
n1 <= "01111";
n2 <= "1" when i1 = n1 else "0";
n3 <= "10000";
n4 <= "1" when i1 = n3 else "0";
n5 <= "10001";
n6 <= "1" when i1 = n5 else "0";
n7 <= "10010";
n8 <= "1" when i1 = n7 else "0";
n9 <= "10011";
n10 <= "1" when i1 = n9 else "0";
n11 <= i14 when n10 = "1" else s16_1;
n12 <= i15 when n8 = "1" else n11;
n13 <= i16 when n6 = "1" else n12;
n14 <= i17 when n4 = "1" else n13;
n15 <= i18 when n2 = "1" else n14;
s16 : cf_rca_16_36 port map (i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, s16_1);
o1 <= n15;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_34 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end entity cf_rca_16_34;
architecture rtl of cf_rca_16_34 is
signal n1 : unsigned(4 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(4 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(4 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(4 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(15 downto 0);
signal s16_1 : unsigned(15 downto 0);
component cf_rca_16_35 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_35;
begin
n1 <= "01010";
n2 <= "1" when i1 = n1 else "0";
n3 <= "01011";
n4 <= "1" when i1 = n3 else "0";
n5 <= "01100";
n6 <= "1" when i1 = n5 else "0";
n7 <= "01101";
n8 <= "1" when i1 = n7 else "0";
n9 <= "01110";
n10 <= "1" when i1 = n9 else "0";
n11 <= i18 when n10 = "1" else s16_1;
n12 <= i18 when n8 = "1" else n11;
n13 <= i18 when n6 = "1" else n12;
n14 <= i18 when n4 = "1" else n13;
n15 <= i18 when n2 = "1" else n14;
s16 : cf_rca_16_35 port map (i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, s16_1);
o1 <= n15;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_33 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end entity cf_rca_16_33;
architecture rtl of cf_rca_16_33 is
signal n1 : unsigned(4 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(4 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(4 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(4 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(15 downto 0);
signal s16_1 : unsigned(15 downto 0);
component cf_rca_16_34 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_34;
begin
n1 <= "00101";
n2 <= "1" when i1 = n1 else "0";
n3 <= "00110";
n4 <= "1" when i1 = n3 else "0";
n5 <= "00111";
n6 <= "1" when i1 = n5 else "0";
n7 <= "01000";
n8 <= "1" when i1 = n7 else "0";
n9 <= "01001";
n10 <= "1" when i1 = n9 else "0";
n11 <= i18 when n10 = "1" else s16_1;
n12 <= i18 when n8 = "1" else n11;
n13 <= i18 when n6 = "1" else n12;
n14 <= i18 when n4 = "1" else n13;
n15 <= i18 when n2 = "1" else n14;
s16 : cf_rca_16_34 port map (i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, s16_1);
o1 <= n15;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end entity cf_rca_16_32;
architecture rtl of cf_rca_16_32 is
signal n1 : unsigned(4 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(4 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(4 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(4 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(15 downto 0);
signal n13 : unsigned(15 downto 0);
signal n14 : unsigned(15 downto 0);
signal n15 : unsigned(15 downto 0);
signal s16_1 : unsigned(15 downto 0);
component cf_rca_16_33 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_33;
begin
n1 <= "00000";
n2 <= "1" when i1 = n1 else "0";
n3 <= "00001";
n4 <= "1" when i1 = n3 else "0";
n5 <= "00010";
n6 <= "1" when i1 = n5 else "0";
n7 <= "00011";
n8 <= "1" when i1 = n7 else "0";
n9 <= "00100";
n10 <= "1" when i1 = n9 else "0";
n11 <= i18 when n10 = "1" else s16_1;
n12 <= i18 when n8 = "1" else n11;
n13 <= i18 when n6 = "1" else n12;
n14 <= i18 when n4 = "1" else n13;
n15 <= i18 when n2 = "1" else n14;
s16 : cf_rca_16_33 port map (i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, s16_1);
o1 <= n15;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_31 is
port (
i1 : in  unsigned(2 downto 0);
i2 : in  unsigned(3 downto 0);
i3 : in  unsigned(3 downto 0);
i4 : in  unsigned(3 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(3 downto 0);
o1 : out unsigned(3 downto 0));
end entity cf_rca_16_31;
architecture rtl of cf_rca_16_31 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(2 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(2 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(2 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(3 downto 0);
signal n14 : unsigned(3 downto 0);
signal n15 : unsigned(3 downto 0);
signal n16 : unsigned(3 downto 0);
signal n17 : unsigned(3 downto 0);
signal n18 : unsigned(3 downto 0);
begin
n1 <= "001";
n2 <= "1" when i1 = n1 else "0";
n3 <= "010";
n4 <= "1" when i1 = n3 else "0";
n5 <= "011";
n6 <= "1" when i1 = n5 else "0";
n7 <= "100";
n8 <= "1" when i1 = n7 else "0";
n9 <= "101";
n10 <= "1" when i1 = n9 else "0";
n11 <= "110";
n12 <= "1" when i1 = n11 else "0";
n13 <= i3 when n12 = "1" else i2;
n14 <= i4 when n10 = "1" else n13;
n15 <= i5 when n8 = "1" else n14;
n16 <= i6 when n6 = "1" else n15;
n17 <= i6 when n4 = "1" else n16;
n18 <= i6 when n2 = "1" else n17;
o1 <= n18;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_30 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end entity cf_rca_16_30;
architecture rtl of cf_rca_16_30 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(3 downto 0);
signal n3 : unsigned(3 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(3 downto 0);
signal n6 : unsigned(3 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(3 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(17 downto 0) := "000000000000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(2 downto 0);
signal n14 : unsigned(2 downto 0);
signal n15 : unsigned(2 downto 0);
signal n16 : unsigned(7 downto 0);
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(17 downto 0) := "000000000000000000";
signal n19 : unsigned(0 downto 0);
signal n20 : unsigned(2 downto 0);
signal n21 : unsigned(2 downto 0);
signal n22 : unsigned(2 downto 0);
signal n23 : unsigned(7 downto 0);
signal n24 : unsigned(0 downto 0);
signal n25 : unsigned(17 downto 0) := "000000000000000000";
signal n26 : unsigned(0 downto 0);
signal n27 : unsigned(2 downto 0);
signal n28 : unsigned(2 downto 0);
signal n29 : unsigned(2 downto 0);
signal n30 : unsigned(7 downto 0);
signal n31 : unsigned(0 downto 0);
signal n32 : unsigned(17 downto 0) := "000000000000000000";
signal n33 : unsigned(0 downto 0);
signal n34 : unsigned(2 downto 0);
signal n35 : unsigned(2 downto 0);
signal n36 : unsigned(2 downto 0);
signal n37 : unsigned(7 downto 0);
signal n38 : unsigned(0 downto 0) := "0";
signal n39 : unsigned(0 downto 0) := "0";
signal n40 : unsigned(0 downto 0);
signal n41 : unsigned(6 downto 0);
signal n42 : unsigned(0 downto 0);
signal n43 : unsigned(5 downto 0);
signal n44 : unsigned(0 downto 0);
signal n45 : unsigned(4 downto 0);
signal n46 : unsigned(0 downto 0);
signal n47 : unsigned(3 downto 0);
signal n48 : unsigned(0 downto 0);
signal n49 : unsigned(2 downto 0);
signal n50 : unsigned(0 downto 0);
signal n51 : unsigned(1 downto 0);
signal n52 : unsigned(0 downto 0);
signal n53 : unsigned(0 downto 0);
signal n54 : unsigned(0 downto 0);
signal n55 : unsigned(0 downto 0);
signal n56 : unsigned(6 downto 0);
signal n57 : unsigned(0 downto 0);
signal n58 : unsigned(5 downto 0);
signal n59 : unsigned(0 downto 0);
signal n60 : unsigned(4 downto 0);
signal n61 : unsigned(0 downto 0);
signal n62 : unsigned(3 downto 0);
signal n63 : unsigned(0 downto 0);
signal n64 : unsigned(2 downto 0);
signal n65 : unsigned(0 downto 0);
signal n66 : unsigned(1 downto 0);
signal n67 : unsigned(0 downto 0);
signal n68 : unsigned(0 downto 0);
signal n69 : unsigned(0 downto 0);
signal n70 : unsigned(0 downto 0);
signal n71 : unsigned(6 downto 0);
signal n72 : unsigned(0 downto 0);
signal n73 : unsigned(5 downto 0);
signal n74 : unsigned(0 downto 0);
signal n75 : unsigned(4 downto 0);
signal n76 : unsigned(0 downto 0);
signal n77 : unsigned(3 downto 0);
signal n78 : unsigned(0 downto 0);
signal n79 : unsigned(2 downto 0);
signal n80 : unsigned(0 downto 0);
signal n81 : unsigned(1 downto 0);
signal n82 : unsigned(0 downto 0);
signal n83 : unsigned(0 downto 0);
signal n84 : unsigned(0 downto 0);
signal n85 : unsigned(0 downto 0);
signal n86 : unsigned(6 downto 0);
signal n87 : unsigned(0 downto 0);
signal n88 : unsigned(5 downto 0);
signal n89 : unsigned(0 downto 0);
signal n90 : unsigned(4 downto 0);
signal n91 : unsigned(0 downto 0);
signal n92 : unsigned(3 downto 0);
signal n93 : unsigned(0 downto 0);
signal n94 : unsigned(2 downto 0);
signal n95 : unsigned(0 downto 0);
signal n96 : unsigned(1 downto 0);
signal n97 : unsigned(0 downto 0);
signal n98 : unsigned(0 downto 0);
signal n99 : unsigned(0 downto 0);
signal n100 : unsigned(1 downto 0);
signal n101 : unsigned(0 downto 0);
signal n102 : unsigned(0 downto 0);
signal n103 : unsigned(0 downto 0);
signal n104 : unsigned(0 downto 0);
signal n105 : unsigned(0 downto 0);
signal n106 : unsigned(0 downto 0);
signal n107 : unsigned(0 downto 0);
signal n108 : unsigned(0 downto 0);
signal n109 : unsigned(0 downto 0);
signal n110 : unsigned(0 downto 0);
signal n111 : unsigned(0 downto 0);
signal n112 : unsigned(1 downto 0);
signal n113 : unsigned(0 downto 0);
signal n114 : unsigned(0 downto 0);
signal n115 : unsigned(0 downto 0);
signal n116 : unsigned(0 downto 0);
signal n117 : unsigned(0 downto 0);
signal n118 : unsigned(0 downto 0);
signal n119 : unsigned(0 downto 0);
signal n120 : unsigned(0 downto 0);
signal n121 : unsigned(0 downto 0);
signal n122 : unsigned(0 downto 0);
signal n123 : unsigned(0 downto 0);
signal n124 : unsigned(1 downto 0);
signal n125 : unsigned(0 downto 0);
signal n126 : unsigned(0 downto 0);
signal n127 : unsigned(0 downto 0);
signal n128 : unsigned(0 downto 0);
signal n129 : unsigned(0 downto 0);
signal n130 : unsigned(0 downto 0);
signal n131 : unsigned(0 downto 0);
signal n132 : unsigned(0 downto 0);
signal n133 : unsigned(0 downto 0);
signal n134 : unsigned(0 downto 0);
signal n135 : unsigned(0 downto 0);
signal n136 : unsigned(1 downto 0);
signal n137 : unsigned(2 downto 0);
signal n138 : unsigned(1 downto 0);
signal n139 : unsigned(0 downto 0);
signal n140 : unsigned(0 downto 0);
signal n141 : unsigned(0 downto 0);
signal n142 : unsigned(0 downto 0);
signal n143 : unsigned(0 downto 0);
signal n144 : unsigned(0 downto 0);
signal n145 : unsigned(0 downto 0);
signal n146 : unsigned(0 downto 0);
signal n147 : unsigned(0 downto 0);
signal n148 : unsigned(0 downto 0);
signal n149 : unsigned(0 downto 0);
signal n150 : unsigned(0 downto 0) := "0";
signal n151 : unsigned(1 downto 0);
signal n152 : unsigned(0 downto 0);
signal n153 : unsigned(0 downto 0);
signal n154 : unsigned(0 downto 0);
signal n155 : unsigned(0 downto 0);
signal n156 : unsigned(0 downto 0);
signal n157 : unsigned(0 downto 0);
signal n158 : unsigned(0 downto 0);
signal n159 : unsigned(0 downto 0);
signal n160 : unsigned(0 downto 0);
signal n161 : unsigned(0 downto 0);
signal n162 : unsigned(0 downto 0);
signal n163 : unsigned(1 downto 0);
signal n164 : unsigned(0 downto 0);
signal n165 : unsigned(0 downto 0);
signal n166 : unsigned(0 downto 0);
signal n167 : unsigned(0 downto 0);
signal n168 : unsigned(0 downto 0);
signal n169 : unsigned(0 downto 0);
signal n170 : unsigned(0 downto 0);
signal n171 : unsigned(0 downto 0);
signal n172 : unsigned(0 downto 0);
signal n173 : unsigned(0 downto 0);
signal n174 : unsigned(0 downto 0);
signal n175 : unsigned(1 downto 0);
signal n176 : unsigned(0 downto 0);
signal n177 : unsigned(0 downto 0);
signal n178 : unsigned(0 downto 0);
signal n179 : unsigned(0 downto 0);
signal n180 : unsigned(0 downto 0);
signal n181 : unsigned(0 downto 0);
signal n182 : unsigned(0 downto 0);
signal n183 : unsigned(0 downto 0);
signal n184 : unsigned(0 downto 0);
signal n185 : unsigned(0 downto 0);
signal n186 : unsigned(0 downto 0);
signal n187 : unsigned(1 downto 0);
signal n188 : unsigned(2 downto 0);
signal n189 : unsigned(1 downto 0);
signal n190 : unsigned(0 downto 0);
signal n191 : unsigned(0 downto 0);
signal n192 : unsigned(0 downto 0);
signal n193 : unsigned(0 downto 0);
signal n194 : unsigned(0 downto 0);
signal n195 : unsigned(0 downto 0);
signal n196 : unsigned(0 downto 0);
signal n197 : unsigned(0 downto 0);
signal n198 : unsigned(0 downto 0);
signal n199 : unsigned(0 downto 0);
signal n200 : unsigned(0 downto 0);
signal n201 : unsigned(0 downto 0) := "0";
signal n202 : unsigned(1 downto 0);
signal n203 : unsigned(0 downto 0);
signal n204 : unsigned(0 downto 0);
signal n205 : unsigned(0 downto 0);
signal n206 : unsigned(0 downto 0);
signal n207 : unsigned(0 downto 0);
signal n208 : unsigned(0 downto 0);
signal n209 : unsigned(0 downto 0);
signal n210 : unsigned(0 downto 0);
signal n211 : unsigned(0 downto 0);
signal n212 : unsigned(0 downto 0);
signal n213 : unsigned(0 downto 0);
signal n214 : unsigned(1 downto 0);
signal n215 : unsigned(0 downto 0);
signal n216 : unsigned(0 downto 0);
signal n217 : unsigned(0 downto 0);
signal n218 : unsigned(0 downto 0);
signal n219 : unsigned(0 downto 0);
signal n220 : unsigned(0 downto 0);
signal n221 : unsigned(0 downto 0);
signal n222 : unsigned(0 downto 0);
signal n223 : unsigned(0 downto 0);
signal n224 : unsigned(0 downto 0);
signal n225 : unsigned(0 downto 0);
signal n226 : unsigned(1 downto 0);
signal n227 : unsigned(0 downto 0);
signal n228 : unsigned(0 downto 0);
signal n229 : unsigned(0 downto 0);
signal n230 : unsigned(0 downto 0);
signal n231 : unsigned(0 downto 0);
signal n232 : unsigned(0 downto 0);
signal n233 : unsigned(0 downto 0);
signal n234 : unsigned(0 downto 0);
signal n235 : unsigned(0 downto 0);
signal n236 : unsigned(0 downto 0);
signal n237 : unsigned(0 downto 0);
signal n238 : unsigned(1 downto 0);
signal n239 : unsigned(2 downto 0);
signal n240 : unsigned(1 downto 0);
signal n241 : unsigned(0 downto 0);
signal n242 : unsigned(0 downto 0);
signal n243 : unsigned(0 downto 0);
signal n244 : unsigned(0 downto 0);
signal n245 : unsigned(0 downto 0);
signal n246 : unsigned(0 downto 0);
signal n247 : unsigned(0 downto 0);
signal n248 : unsigned(0 downto 0);
signal n249 : unsigned(0 downto 0);
signal n250 : unsigned(0 downto 0);
signal n251 : unsigned(0 downto 0);
signal n252 : unsigned(0 downto 0) := "0";
signal n253 : unsigned(1 downto 0);
signal n254 : unsigned(0 downto 0);
signal n255 : unsigned(0 downto 0);
signal n256 : unsigned(0 downto 0);
signal n257 : unsigned(0 downto 0);
signal n258 : unsigned(0 downto 0);
signal n259 : unsigned(0 downto 0);
signal n260 : unsigned(0 downto 0);
signal n261 : unsigned(0 downto 0);
signal n262 : unsigned(0 downto 0);
signal n263 : unsigned(0 downto 0);
signal n264 : unsigned(0 downto 0);
signal n265 : unsigned(1 downto 0);
signal n266 : unsigned(0 downto 0);
signal n267 : unsigned(0 downto 0);
signal n268 : unsigned(0 downto 0);
signal n269 : unsigned(0 downto 0);
signal n270 : unsigned(0 downto 0);
signal n271 : unsigned(0 downto 0);
signal n272 : unsigned(0 downto 0);
signal n273 : unsigned(0 downto 0);
signal n274 : unsigned(0 downto 0);
signal n275 : unsigned(0 downto 0);
signal n276 : unsigned(0 downto 0);
signal n277 : unsigned(1 downto 0);
signal n278 : unsigned(0 downto 0);
signal n279 : unsigned(0 downto 0);
signal n280 : unsigned(0 downto 0);
signal n281 : unsigned(0 downto 0);
signal n282 : unsigned(0 downto 0);
signal n283 : unsigned(0 downto 0);
signal n284 : unsigned(0 downto 0);
signal n285 : unsigned(0 downto 0);
signal n286 : unsigned(0 downto 0);
signal n287 : unsigned(0 downto 0);
signal n288 : unsigned(0 downto 0);
signal n289 : unsigned(1 downto 0);
signal n290 : unsigned(2 downto 0);
signal n291 : unsigned(1 downto 0);
signal n292 : unsigned(0 downto 0);
signal n293 : unsigned(0 downto 0);
signal n294 : unsigned(0 downto 0);
signal n295 : unsigned(0 downto 0);
signal n296 : unsigned(0 downto 0);
signal n297 : unsigned(0 downto 0);
signal n298 : unsigned(0 downto 0);
signal n299 : unsigned(0 downto 0);
signal n300 : unsigned(0 downto 0);
signal n301 : unsigned(0 downto 0);
signal n302 : unsigned(0 downto 0);
signal n303 : unsigned(0 downto 0) := "0";
signal n304 : unsigned(0 downto 0);
signal n305 : unsigned(0 downto 0);
signal n306 : unsigned(0 downto 0);
signal n307 : unsigned(0 downto 0);
signal n308 : unsigned(0 downto 0) := "0";
signal n309 : unsigned(0 downto 0) := "0";
signal s310_1 : unsigned(3 downto 0);
component cf_rca_16_31 is
port (
i1 : in  unsigned(2 downto 0);
i2 : in  unsigned(3 downto 0);
i3 : in  unsigned(3 downto 0);
i4 : in  unsigned(3 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(3 downto 0);
o1 : out unsigned(3 downto 0));
end component cf_rca_16_31;
begin
n1 <= i7 & i4;
n2 <= "1000";
n3 <= "0100";
n4 <= "0010";
n5 <= "0001";
n6 <= "0000";
n7 <= "000";
n8 <= "1" when n1 = n7 else "0";
n9 <= n6 when n8 = "1" else s310_1;
n10 <= n9(0 downto 0);
process (clock_config_c) begin
  if rising_edge(clock_config_c) then
    if i2 = "1" then
      n11 <= "000000000000000000";
    elsif n10 = "1" then
      n11 <= i3;
    end if;
  end if;
end process;
n12 <= n11(17 downto 17);
n13 <= n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14);
n14 <= n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11);
n15 <= n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8);
n16 <= n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n17 <= n9(1 downto 1);
process (clock_config_c) begin
  if rising_edge(clock_config_c) then
    if i2 = "1" then
      n18 <= "000000000000000000";
    elsif n17 = "1" then
      n18 <= i3;
    end if;
  end if;
end process;
n19 <= n18(17 downto 17);
n20 <= n18(16 downto 16) &
  n18(15 downto 15) &
  n18(14 downto 14);
n21 <= n18(13 downto 13) &
  n18(12 downto 12) &
  n18(11 downto 11);
n22 <= n18(10 downto 10) &
  n18(9 downto 9) &
  n18(8 downto 8);
n23 <= n18(7 downto 7) &
  n18(6 downto 6) &
  n18(5 downto 5) &
  n18(4 downto 4) &
  n18(3 downto 3) &
  n18(2 downto 2) &
  n18(1 downto 1) &
  n18(0 downto 0);
n24 <= n9(2 downto 2);
process (clock_config_c) begin
  if rising_edge(clock_config_c) then
    if i2 = "1" then
      n25 <= "000000000000000000";
    elsif n24 = "1" then
      n25 <= i3;
    end if;
  end if;
end process;
n26 <= n25(17 downto 17);
n27 <= n25(16 downto 16) &
  n25(15 downto 15) &
  n25(14 downto 14);
n28 <= n25(13 downto 13) &
  n25(12 downto 12) &
  n25(11 downto 11);
n29 <= n25(10 downto 10) &
  n25(9 downto 9) &
  n25(8 downto 8);
n30 <= n25(7 downto 7) &
  n25(6 downto 6) &
  n25(5 downto 5) &
  n25(4 downto 4) &
  n25(3 downto 3) &
  n25(2 downto 2) &
  n25(1 downto 1) &
  n25(0 downto 0);
n31 <= n9(3 downto 3);
process (clock_config_c) begin
  if rising_edge(clock_config_c) then
    if i2 = "1" then
      n32 <= "000000000000000000";
    elsif n31 = "1" then
      n32 <= i3;
    end if;
  end if;
end process;
n33 <= n32(17 downto 17);
n34 <= n32(16 downto 16) &
  n32(15 downto 15) &
  n32(14 downto 14);
n35 <= n32(13 downto 13) &
  n32(12 downto 12) &
  n32(11 downto 11);
n36 <= n32(10 downto 10) &
  n32(9 downto 9) &
  n32(8 downto 8);
n37 <= n32(7 downto 7) &
  n32(6 downto 6) &
  n32(5 downto 5) &
  n32(4 downto 4) &
  n32(3 downto 3) &
  n32(2 downto 2) &
  n32(1 downto 1) &
  n32(0 downto 0);
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n38 <= "0";
    elsif i1 = "1" then
      n38 <= i8;
    end if;
  end if;
end process;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n39 <= "0";
    elsif i1 = "1" then
      n39 <= i6;
    end if;
  end if;
end process;
n40 <= n16(7 downto 7);
n41 <= n16(6 downto 6) &
  n16(5 downto 5) &
  n16(4 downto 4) &
  n16(3 downto 3) &
  n16(2 downto 2) &
  n16(1 downto 1) &
  n16(0 downto 0);
n42 <= n41(6 downto 6);
n43 <= n41(5 downto 5) &
  n41(4 downto 4) &
  n41(3 downto 3) &
  n41(2 downto 2) &
  n41(1 downto 1) &
  n41(0 downto 0);
n44 <= n43(5 downto 5);
n45 <= n43(4 downto 4) &
  n43(3 downto 3) &
  n43(2 downto 2) &
  n43(1 downto 1) &
  n43(0 downto 0);
n46 <= n45(4 downto 4);
n47 <= n45(3 downto 3) &
  n45(2 downto 2) &
  n45(1 downto 1) &
  n45(0 downto 0);
n48 <= n47(3 downto 3);
n49 <= n47(2 downto 2) &
  n47(1 downto 1) &
  n47(0 downto 0);
n50 <= n49(2 downto 2);
n51 <= n49(1 downto 1) &
  n49(0 downto 0);
n52 <= n51(1 downto 1);
n53 <= n51(0 downto 0);
n54 <= n53(0 downto 0);
n55 <= n23(7 downto 7);
n56 <= n23(6 downto 6) &
  n23(5 downto 5) &
  n23(4 downto 4) &
  n23(3 downto 3) &
  n23(2 downto 2) &
  n23(1 downto 1) &
  n23(0 downto 0);
n57 <= n56(6 downto 6);
n58 <= n56(5 downto 5) &
  n56(4 downto 4) &
  n56(3 downto 3) &
  n56(2 downto 2) &
  n56(1 downto 1) &
  n56(0 downto 0);
n59 <= n58(5 downto 5);
n60 <= n58(4 downto 4) &
  n58(3 downto 3) &
  n58(2 downto 2) &
  n58(1 downto 1) &
  n58(0 downto 0);
n61 <= n60(4 downto 4);
n62 <= n60(3 downto 3) &
  n60(2 downto 2) &
  n60(1 downto 1) &
  n60(0 downto 0);
n63 <= n62(3 downto 3);
n64 <= n62(2 downto 2) &
  n62(1 downto 1) &
  n62(0 downto 0);
n65 <= n64(2 downto 2);
n66 <= n64(1 downto 1) &
  n64(0 downto 0);
n67 <= n66(1 downto 1);
n68 <= n66(0 downto 0);
n69 <= n68(0 downto 0);
n70 <= n30(7 downto 7);
n71 <= n30(6 downto 6) &
  n30(5 downto 5) &
  n30(4 downto 4) &
  n30(3 downto 3) &
  n30(2 downto 2) &
  n30(1 downto 1) &
  n30(0 downto 0);
n72 <= n71(6 downto 6);
n73 <= n71(5 downto 5) &
  n71(4 downto 4) &
  n71(3 downto 3) &
  n71(2 downto 2) &
  n71(1 downto 1) &
  n71(0 downto 0);
n74 <= n73(5 downto 5);
n75 <= n73(4 downto 4) &
  n73(3 downto 3) &
  n73(2 downto 2) &
  n73(1 downto 1) &
  n73(0 downto 0);
n76 <= n75(4 downto 4);
n77 <= n75(3 downto 3) &
  n75(2 downto 2) &
  n75(1 downto 1) &
  n75(0 downto 0);
n78 <= n77(3 downto 3);
n79 <= n77(2 downto 2) &
  n77(1 downto 1) &
  n77(0 downto 0);
n80 <= n79(2 downto 2);
n81 <= n79(1 downto 1) &
  n79(0 downto 0);
n82 <= n81(1 downto 1);
n83 <= n81(0 downto 0);
n84 <= n83(0 downto 0);
n85 <= n37(7 downto 7);
n86 <= n37(6 downto 6) &
  n37(5 downto 5) &
  n37(4 downto 4) &
  n37(3 downto 3) &
  n37(2 downto 2) &
  n37(1 downto 1) &
  n37(0 downto 0);
n87 <= n86(6 downto 6);
n88 <= n86(5 downto 5) &
  n86(4 downto 4) &
  n86(3 downto 3) &
  n86(2 downto 2) &
  n86(1 downto 1) &
  n86(0 downto 0);
n89 <= n88(5 downto 5);
n90 <= n88(4 downto 4) &
  n88(3 downto 3) &
  n88(2 downto 2) &
  n88(1 downto 1) &
  n88(0 downto 0);
n91 <= n90(4 downto 4);
n92 <= n90(3 downto 3) &
  n90(2 downto 2) &
  n90(1 downto 1) &
  n90(0 downto 0);
n93 <= n92(3 downto 3);
n94 <= n92(2 downto 2) &
  n92(1 downto 1) &
  n92(0 downto 0);
n95 <= n94(2 downto 2);
n96 <= n94(1 downto 1) &
  n94(0 downto 0);
n97 <= n96(1 downto 1);
n98 <= n96(0 downto 0);
n99 <= n98(0 downto 0);
n100 <= n13(2 downto 2) &
  n13(1 downto 1);
n101 <= n13(0 downto 0);
n102 <= n309 when n101 = "1" else n38;
n103 <= n308 when n101 = "1" else n39;
n104 <= n201 when n101 = "1" else n150;
n105 <= n303 when n101 = "1" else n252;
n106 <= n100(1 downto 1);
n107 <= n100(0 downto 0);
n108 <= n103 when n107 = "1" else n102;
n109 <= n105 when n107 = "1" else n104;
n110 <= n106(0 downto 0);
n111 <= n109 when n110 = "1" else n108;
n112 <= n14(2 downto 2) &
  n14(1 downto 1);
n113 <= n14(0 downto 0);
n114 <= n309 when n113 = "1" else n38;
n115 <= n308 when n113 = "1" else n39;
n116 <= n201 when n113 = "1" else n150;
n117 <= n303 when n113 = "1" else n252;
n118 <= n112(1 downto 1);
n119 <= n112(0 downto 0);
n120 <= n115 when n119 = "1" else n114;
n121 <= n117 when n119 = "1" else n116;
n122 <= n118(0 downto 0);
n123 <= n121 when n122 = "1" else n120;
n124 <= n15(2 downto 2) &
  n15(1 downto 1);
n125 <= n15(0 downto 0);
n126 <= n309 when n125 = "1" else n38;
n127 <= n308 when n125 = "1" else n39;
n128 <= n201 when n125 = "1" else n150;
n129 <= n303 when n125 = "1" else n252;
n130 <= n124(1 downto 1);
n131 <= n124(0 downto 0);
n132 <= n127 when n131 = "1" else n126;
n133 <= n129 when n131 = "1" else n128;
n134 <= n130(0 downto 0);
n135 <= n133 when n134 = "1" else n132;
n136 <= n123 & n135;
n137 <= n111 & n136;
n138 <= n137(2 downto 2) &
  n137(1 downto 1);
n139 <= n137(0 downto 0);
n140 <= n52 when n139 = "1" else n54;
n141 <= n48 when n139 = "1" else n50;
n142 <= n44 when n139 = "1" else n46;
n143 <= n40 when n139 = "1" else n42;
n144 <= n138(1 downto 1);
n145 <= n138(0 downto 0);
n146 <= n141 when n145 = "1" else n140;
n147 <= n143 when n145 = "1" else n142;
n148 <= n144(0 downto 0);
n149 <= n147 when n148 = "1" else n146;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n150 <= "0";
    elsif i1 = "1" then
      n150 <= n149;
    end if;
  end if;
end process;
n151 <= n20(2 downto 2) &
  n20(1 downto 1);
n152 <= n20(0 downto 0);
n153 <= n309 when n152 = "1" else n38;
n154 <= n308 when n152 = "1" else n39;
n155 <= n201 when n152 = "1" else n150;
n156 <= n303 when n152 = "1" else n252;
n157 <= n151(1 downto 1);
n158 <= n151(0 downto 0);
n159 <= n154 when n158 = "1" else n153;
n160 <= n156 when n158 = "1" else n155;
n161 <= n157(0 downto 0);
n162 <= n160 when n161 = "1" else n159;
n163 <= n21(2 downto 2) &
  n21(1 downto 1);
n164 <= n21(0 downto 0);
n165 <= n309 when n164 = "1" else n38;
n166 <= n308 when n164 = "1" else n39;
n167 <= n201 when n164 = "1" else n150;
n168 <= n303 when n164 = "1" else n252;
n169 <= n163(1 downto 1);
n170 <= n163(0 downto 0);
n171 <= n166 when n170 = "1" else n165;
n172 <= n168 when n170 = "1" else n167;
n173 <= n169(0 downto 0);
n174 <= n172 when n173 = "1" else n171;
n175 <= n22(2 downto 2) &
  n22(1 downto 1);
n176 <= n22(0 downto 0);
n177 <= n309 when n176 = "1" else n38;
n178 <= n308 when n176 = "1" else n39;
n179 <= n201 when n176 = "1" else n150;
n180 <= n303 when n176 = "1" else n252;
n181 <= n175(1 downto 1);
n182 <= n175(0 downto 0);
n183 <= n178 when n182 = "1" else n177;
n184 <= n180 when n182 = "1" else n179;
n185 <= n181(0 downto 0);
n186 <= n184 when n185 = "1" else n183;
n187 <= n174 & n186;
n188 <= n162 & n187;
n189 <= n188(2 downto 2) &
  n188(1 downto 1);
n190 <= n188(0 downto 0);
n191 <= n67 when n190 = "1" else n69;
n192 <= n63 when n190 = "1" else n65;
n193 <= n59 when n190 = "1" else n61;
n194 <= n55 when n190 = "1" else n57;
n195 <= n189(1 downto 1);
n196 <= n189(0 downto 0);
n197 <= n192 when n196 = "1" else n191;
n198 <= n194 when n196 = "1" else n193;
n199 <= n195(0 downto 0);
n200 <= n198 when n199 = "1" else n197;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n201 <= "0";
    elsif i1 = "1" then
      n201 <= n200;
    end if;
  end if;
end process;
n202 <= n27(2 downto 2) &
  n27(1 downto 1);
n203 <= n27(0 downto 0);
n204 <= n309 when n203 = "1" else n38;
n205 <= n308 when n203 = "1" else n39;
n206 <= n201 when n203 = "1" else n150;
n207 <= n303 when n203 = "1" else n252;
n208 <= n202(1 downto 1);
n209 <= n202(0 downto 0);
n210 <= n205 when n209 = "1" else n204;
n211 <= n207 when n209 = "1" else n206;
n212 <= n208(0 downto 0);
n213 <= n211 when n212 = "1" else n210;
n214 <= n28(2 downto 2) &
  n28(1 downto 1);
n215 <= n28(0 downto 0);
n216 <= n309 when n215 = "1" else n38;
n217 <= n308 when n215 = "1" else n39;
n218 <= n201 when n215 = "1" else n150;
n219 <= n303 when n215 = "1" else n252;
n220 <= n214(1 downto 1);
n221 <= n214(0 downto 0);
n222 <= n217 when n221 = "1" else n216;
n223 <= n219 when n221 = "1" else n218;
n224 <= n220(0 downto 0);
n225 <= n223 when n224 = "1" else n222;
n226 <= n29(2 downto 2) &
  n29(1 downto 1);
n227 <= n29(0 downto 0);
n228 <= n309 when n227 = "1" else n38;
n229 <= n308 when n227 = "1" else n39;
n230 <= n201 when n227 = "1" else n150;
n231 <= n303 when n227 = "1" else n252;
n232 <= n226(1 downto 1);
n233 <= n226(0 downto 0);
n234 <= n229 when n233 = "1" else n228;
n235 <= n231 when n233 = "1" else n230;
n236 <= n232(0 downto 0);
n237 <= n235 when n236 = "1" else n234;
n238 <= n225 & n237;
n239 <= n213 & n238;
n240 <= n239(2 downto 2) &
  n239(1 downto 1);
n241 <= n239(0 downto 0);
n242 <= n82 when n241 = "1" else n84;
n243 <= n78 when n241 = "1" else n80;
n244 <= n74 when n241 = "1" else n76;
n245 <= n70 when n241 = "1" else n72;
n246 <= n240(1 downto 1);
n247 <= n240(0 downto 0);
n248 <= n243 when n247 = "1" else n242;
n249 <= n245 when n247 = "1" else n244;
n250 <= n246(0 downto 0);
n251 <= n249 when n250 = "1" else n248;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n252 <= "0";
    elsif i1 = "1" then
      n252 <= n251;
    end if;
  end if;
end process;
n253 <= n34(2 downto 2) &
  n34(1 downto 1);
n254 <= n34(0 downto 0);
n255 <= n309 when n254 = "1" else n38;
n256 <= n308 when n254 = "1" else n39;
n257 <= n201 when n254 = "1" else n150;
n258 <= n303 when n254 = "1" else n252;
n259 <= n253(1 downto 1);
n260 <= n253(0 downto 0);
n261 <= n256 when n260 = "1" else n255;
n262 <= n258 when n260 = "1" else n257;
n263 <= n259(0 downto 0);
n264 <= n262 when n263 = "1" else n261;
n265 <= n35(2 downto 2) &
  n35(1 downto 1);
n266 <= n35(0 downto 0);
n267 <= n309 when n266 = "1" else n38;
n268 <= n308 when n266 = "1" else n39;
n269 <= n201 when n266 = "1" else n150;
n270 <= n303 when n266 = "1" else n252;
n271 <= n265(1 downto 1);
n272 <= n265(0 downto 0);
n273 <= n268 when n272 = "1" else n267;
n274 <= n270 when n272 = "1" else n269;
n275 <= n271(0 downto 0);
n276 <= n274 when n275 = "1" else n273;
n277 <= n36(2 downto 2) &
  n36(1 downto 1);
n278 <= n36(0 downto 0);
n279 <= n309 when n278 = "1" else n38;
n280 <= n308 when n278 = "1" else n39;
n281 <= n201 when n278 = "1" else n150;
n282 <= n303 when n278 = "1" else n252;
n283 <= n277(1 downto 1);
n284 <= n277(0 downto 0);
n285 <= n280 when n284 = "1" else n279;
n286 <= n282 when n284 = "1" else n281;
n287 <= n283(0 downto 0);
n288 <= n286 when n287 = "1" else n285;
n289 <= n276 & n288;
n290 <= n264 & n289;
n291 <= n290(2 downto 2) &
  n290(1 downto 1);
n292 <= n290(0 downto 0);
n293 <= n97 when n292 = "1" else n99;
n294 <= n93 when n292 = "1" else n95;
n295 <= n89 when n292 = "1" else n91;
n296 <= n85 when n292 = "1" else n87;
n297 <= n291(1 downto 1);
n298 <= n291(0 downto 0);
n299 <= n294 when n298 = "1" else n293;
n300 <= n296 when n298 = "1" else n295;
n301 <= n297(0 downto 0);
n302 <= n300 when n301 = "1" else n299;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n303 <= "0";
    elsif i1 = "1" then
      n303 <= n302;
    end if;
  end if;
end process;
n304 <= n150 when n12 = "1" else n149;
n305 <= n201 when n19 = "1" else n200;
n306 <= n252 when n26 = "1" else n251;
n307 <= n303 when n33 = "1" else n302;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n308 <= "0";
    elsif i1 = "1" then
      n308 <= i5;
    end if;
  end if;
end process;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n309 <= "0";
    elsif i1 = "1" then
      n309 <= i9;
    end if;
  end if;
end process;
s310 : cf_rca_16_31 port map (n1, n2, n3, n4, n5, n6, s310_1);
o4 <= n307;
o3 <= n306;
o2 <= n305;
o1 <= n304;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end entity cf_rca_16_29;
architecture rtl of cf_rca_16_29 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(3 downto 0);
signal n3 : unsigned(3 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(3 downto 0);
signal n6 : unsigned(3 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(3 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(17 downto 0) := "000000000000000000";
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(2 downto 0);
signal n14 : unsigned(2 downto 0);
signal n15 : unsigned(2 downto 0);
signal n16 : unsigned(7 downto 0);
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(17 downto 0) := "000000000000000000";
signal n19 : unsigned(0 downto 0);
signal n20 : unsigned(2 downto 0);
signal n21 : unsigned(2 downto 0);
signal n22 : unsigned(2 downto 0);
signal n23 : unsigned(7 downto 0);
signal n24 : unsigned(0 downto 0);
signal n25 : unsigned(17 downto 0) := "000000000000000000";
signal n26 : unsigned(0 downto 0);
signal n27 : unsigned(2 downto 0);
signal n28 : unsigned(2 downto 0);
signal n29 : unsigned(2 downto 0);
signal n30 : unsigned(7 downto 0);
signal n31 : unsigned(0 downto 0);
signal n32 : unsigned(17 downto 0) := "000000000000000000";
signal n33 : unsigned(0 downto 0);
signal n34 : unsigned(2 downto 0);
signal n35 : unsigned(2 downto 0);
signal n36 : unsigned(2 downto 0);
signal n37 : unsigned(7 downto 0);
signal n38 : unsigned(0 downto 0) := "0";
signal n39 : unsigned(0 downto 0) := "0";
signal n40 : unsigned(0 downto 0);
signal n41 : unsigned(6 downto 0);
signal n42 : unsigned(0 downto 0);
signal n43 : unsigned(5 downto 0);
signal n44 : unsigned(0 downto 0);
signal n45 : unsigned(4 downto 0);
signal n46 : unsigned(0 downto 0);
signal n47 : unsigned(3 downto 0);
signal n48 : unsigned(0 downto 0);
signal n49 : unsigned(2 downto 0);
signal n50 : unsigned(0 downto 0);
signal n51 : unsigned(1 downto 0);
signal n52 : unsigned(0 downto 0);
signal n53 : unsigned(0 downto 0);
signal n54 : unsigned(0 downto 0);
signal n55 : unsigned(0 downto 0);
signal n56 : unsigned(6 downto 0);
signal n57 : unsigned(0 downto 0);
signal n58 : unsigned(5 downto 0);
signal n59 : unsigned(0 downto 0);
signal n60 : unsigned(4 downto 0);
signal n61 : unsigned(0 downto 0);
signal n62 : unsigned(3 downto 0);
signal n63 : unsigned(0 downto 0);
signal n64 : unsigned(2 downto 0);
signal n65 : unsigned(0 downto 0);
signal n66 : unsigned(1 downto 0);
signal n67 : unsigned(0 downto 0);
signal n68 : unsigned(0 downto 0);
signal n69 : unsigned(0 downto 0);
signal n70 : unsigned(0 downto 0);
signal n71 : unsigned(6 downto 0);
signal n72 : unsigned(0 downto 0);
signal n73 : unsigned(5 downto 0);
signal n74 : unsigned(0 downto 0);
signal n75 : unsigned(4 downto 0);
signal n76 : unsigned(0 downto 0);
signal n77 : unsigned(3 downto 0);
signal n78 : unsigned(0 downto 0);
signal n79 : unsigned(2 downto 0);
signal n80 : unsigned(0 downto 0);
signal n81 : unsigned(1 downto 0);
signal n82 : unsigned(0 downto 0);
signal n83 : unsigned(0 downto 0);
signal n84 : unsigned(0 downto 0);
signal n85 : unsigned(0 downto 0);
signal n86 : unsigned(6 downto 0);
signal n87 : unsigned(0 downto 0);
signal n88 : unsigned(5 downto 0);
signal n89 : unsigned(0 downto 0);
signal n90 : unsigned(4 downto 0);
signal n91 : unsigned(0 downto 0);
signal n92 : unsigned(3 downto 0);
signal n93 : unsigned(0 downto 0);
signal n94 : unsigned(2 downto 0);
signal n95 : unsigned(0 downto 0);
signal n96 : unsigned(1 downto 0);
signal n97 : unsigned(0 downto 0);
signal n98 : unsigned(0 downto 0);
signal n99 : unsigned(0 downto 0);
signal n100 : unsigned(1 downto 0);
signal n101 : unsigned(0 downto 0);
signal n102 : unsigned(0 downto 0);
signal n103 : unsigned(0 downto 0);
signal n104 : unsigned(0 downto 0);
signal n105 : unsigned(0 downto 0);
signal n106 : unsigned(0 downto 0);
signal n107 : unsigned(0 downto 0);
signal n108 : unsigned(0 downto 0);
signal n109 : unsigned(0 downto 0);
signal n110 : unsigned(0 downto 0);
signal n111 : unsigned(0 downto 0);
signal n112 : unsigned(1 downto 0);
signal n113 : unsigned(0 downto 0);
signal n114 : unsigned(0 downto 0);
signal n115 : unsigned(0 downto 0);
signal n116 : unsigned(0 downto 0);
signal n117 : unsigned(0 downto 0);
signal n118 : unsigned(0 downto 0);
signal n119 : unsigned(0 downto 0);
signal n120 : unsigned(0 downto 0);
signal n121 : unsigned(0 downto 0);
signal n122 : unsigned(0 downto 0);
signal n123 : unsigned(0 downto 0);
signal n124 : unsigned(1 downto 0);
signal n125 : unsigned(0 downto 0);
signal n126 : unsigned(0 downto 0);
signal n127 : unsigned(0 downto 0);
signal n128 : unsigned(0 downto 0);
signal n129 : unsigned(0 downto 0);
signal n130 : unsigned(0 downto 0);
signal n131 : unsigned(0 downto 0);
signal n132 : unsigned(0 downto 0);
signal n133 : unsigned(0 downto 0);
signal n134 : unsigned(0 downto 0);
signal n135 : unsigned(0 downto 0);
signal n136 : unsigned(1 downto 0);
signal n137 : unsigned(2 downto 0);
signal n138 : unsigned(1 downto 0);
signal n139 : unsigned(0 downto 0);
signal n140 : unsigned(0 downto 0);
signal n141 : unsigned(0 downto 0);
signal n142 : unsigned(0 downto 0);
signal n143 : unsigned(0 downto 0);
signal n144 : unsigned(0 downto 0);
signal n145 : unsigned(0 downto 0);
signal n146 : unsigned(0 downto 0);
signal n147 : unsigned(0 downto 0);
signal n148 : unsigned(0 downto 0);
signal n149 : unsigned(0 downto 0);
signal n150 : unsigned(0 downto 0) := "0";
signal n151 : unsigned(1 downto 0);
signal n152 : unsigned(0 downto 0);
signal n153 : unsigned(0 downto 0);
signal n154 : unsigned(0 downto 0);
signal n155 : unsigned(0 downto 0);
signal n156 : unsigned(0 downto 0);
signal n157 : unsigned(0 downto 0);
signal n158 : unsigned(0 downto 0);
signal n159 : unsigned(0 downto 0);
signal n160 : unsigned(0 downto 0);
signal n161 : unsigned(0 downto 0);
signal n162 : unsigned(0 downto 0);
signal n163 : unsigned(1 downto 0);
signal n164 : unsigned(0 downto 0);
signal n165 : unsigned(0 downto 0);
signal n166 : unsigned(0 downto 0);
signal n167 : unsigned(0 downto 0);
signal n168 : unsigned(0 downto 0);
signal n169 : unsigned(0 downto 0);
signal n170 : unsigned(0 downto 0);
signal n171 : unsigned(0 downto 0);
signal n172 : unsigned(0 downto 0);
signal n173 : unsigned(0 downto 0);
signal n174 : unsigned(0 downto 0);
signal n175 : unsigned(1 downto 0);
signal n176 : unsigned(0 downto 0);
signal n177 : unsigned(0 downto 0);
signal n178 : unsigned(0 downto 0);
signal n179 : unsigned(0 downto 0);
signal n180 : unsigned(0 downto 0);
signal n181 : unsigned(0 downto 0);
signal n182 : unsigned(0 downto 0);
signal n183 : unsigned(0 downto 0);
signal n184 : unsigned(0 downto 0);
signal n185 : unsigned(0 downto 0);
signal n186 : unsigned(0 downto 0);
signal n187 : unsigned(1 downto 0);
signal n188 : unsigned(2 downto 0);
signal n189 : unsigned(1 downto 0);
signal n190 : unsigned(0 downto 0);
signal n191 : unsigned(0 downto 0);
signal n192 : unsigned(0 downto 0);
signal n193 : unsigned(0 downto 0);
signal n194 : unsigned(0 downto 0);
signal n195 : unsigned(0 downto 0);
signal n196 : unsigned(0 downto 0);
signal n197 : unsigned(0 downto 0);
signal n198 : unsigned(0 downto 0);
signal n199 : unsigned(0 downto 0);
signal n200 : unsigned(0 downto 0);
signal n201 : unsigned(0 downto 0) := "0";
signal n202 : unsigned(1 downto 0);
signal n203 : unsigned(0 downto 0);
signal n204 : unsigned(0 downto 0);
signal n205 : unsigned(0 downto 0);
signal n206 : unsigned(0 downto 0);
signal n207 : unsigned(0 downto 0);
signal n208 : unsigned(0 downto 0);
signal n209 : unsigned(0 downto 0);
signal n210 : unsigned(0 downto 0);
signal n211 : unsigned(0 downto 0);
signal n212 : unsigned(0 downto 0);
signal n213 : unsigned(0 downto 0);
signal n214 : unsigned(1 downto 0);
signal n215 : unsigned(0 downto 0);
signal n216 : unsigned(0 downto 0);
signal n217 : unsigned(0 downto 0);
signal n218 : unsigned(0 downto 0);
signal n219 : unsigned(0 downto 0);
signal n220 : unsigned(0 downto 0);
signal n221 : unsigned(0 downto 0);
signal n222 : unsigned(0 downto 0);
signal n223 : unsigned(0 downto 0);
signal n224 : unsigned(0 downto 0);
signal n225 : unsigned(0 downto 0);
signal n226 : unsigned(1 downto 0);
signal n227 : unsigned(0 downto 0);
signal n228 : unsigned(0 downto 0);
signal n229 : unsigned(0 downto 0);
signal n230 : unsigned(0 downto 0);
signal n231 : unsigned(0 downto 0);
signal n232 : unsigned(0 downto 0);
signal n233 : unsigned(0 downto 0);
signal n234 : unsigned(0 downto 0);
signal n235 : unsigned(0 downto 0);
signal n236 : unsigned(0 downto 0);
signal n237 : unsigned(0 downto 0);
signal n238 : unsigned(1 downto 0);
signal n239 : unsigned(2 downto 0);
signal n240 : unsigned(1 downto 0);
signal n241 : unsigned(0 downto 0);
signal n242 : unsigned(0 downto 0);
signal n243 : unsigned(0 downto 0);
signal n244 : unsigned(0 downto 0);
signal n245 : unsigned(0 downto 0);
signal n246 : unsigned(0 downto 0);
signal n247 : unsigned(0 downto 0);
signal n248 : unsigned(0 downto 0);
signal n249 : unsigned(0 downto 0);
signal n250 : unsigned(0 downto 0);
signal n251 : unsigned(0 downto 0);
signal n252 : unsigned(0 downto 0) := "0";
signal n253 : unsigned(1 downto 0);
signal n254 : unsigned(0 downto 0);
signal n255 : unsigned(0 downto 0);
signal n256 : unsigned(0 downto 0);
signal n257 : unsigned(0 downto 0);
signal n258 : unsigned(0 downto 0);
signal n259 : unsigned(0 downto 0);
signal n260 : unsigned(0 downto 0);
signal n261 : unsigned(0 downto 0);
signal n262 : unsigned(0 downto 0);
signal n263 : unsigned(0 downto 0);
signal n264 : unsigned(0 downto 0);
signal n265 : unsigned(1 downto 0);
signal n266 : unsigned(0 downto 0);
signal n267 : unsigned(0 downto 0);
signal n268 : unsigned(0 downto 0);
signal n269 : unsigned(0 downto 0);
signal n270 : unsigned(0 downto 0);
signal n271 : unsigned(0 downto 0);
signal n272 : unsigned(0 downto 0);
signal n273 : unsigned(0 downto 0);
signal n274 : unsigned(0 downto 0);
signal n275 : unsigned(0 downto 0);
signal n276 : unsigned(0 downto 0);
signal n277 : unsigned(1 downto 0);
signal n278 : unsigned(0 downto 0);
signal n279 : unsigned(0 downto 0);
signal n280 : unsigned(0 downto 0);
signal n281 : unsigned(0 downto 0);
signal n282 : unsigned(0 downto 0);
signal n283 : unsigned(0 downto 0);
signal n284 : unsigned(0 downto 0);
signal n285 : unsigned(0 downto 0);
signal n286 : unsigned(0 downto 0);
signal n287 : unsigned(0 downto 0);
signal n288 : unsigned(0 downto 0);
signal n289 : unsigned(1 downto 0);
signal n290 : unsigned(2 downto 0);
signal n291 : unsigned(1 downto 0);
signal n292 : unsigned(0 downto 0);
signal n293 : unsigned(0 downto 0);
signal n294 : unsigned(0 downto 0);
signal n295 : unsigned(0 downto 0);
signal n296 : unsigned(0 downto 0);
signal n297 : unsigned(0 downto 0);
signal n298 : unsigned(0 downto 0);
signal n299 : unsigned(0 downto 0);
signal n300 : unsigned(0 downto 0);
signal n301 : unsigned(0 downto 0);
signal n302 : unsigned(0 downto 0);
signal n303 : unsigned(0 downto 0) := "0";
signal n304 : unsigned(0 downto 0);
signal n305 : unsigned(0 downto 0);
signal n306 : unsigned(0 downto 0);
signal n307 : unsigned(0 downto 0);
signal n308 : unsigned(0 downto 0) := "0";
signal n309 : unsigned(0 downto 0) := "0";
signal s310_1 : unsigned(3 downto 0);
component cf_rca_16_31 is
port (
i1 : in  unsigned(2 downto 0);
i2 : in  unsigned(3 downto 0);
i3 : in  unsigned(3 downto 0);
i4 : in  unsigned(3 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(3 downto 0);
o1 : out unsigned(3 downto 0));
end component cf_rca_16_31;
begin
n1 <= i6 & i4;
n2 <= "1000";
n3 <= "0100";
n4 <= "0010";
n5 <= "0001";
n6 <= "0000";
n7 <= "000";
n8 <= "1" when n1 = n7 else "0";
n9 <= n6 when n8 = "1" else s310_1;
n10 <= n9(0 downto 0);
process (clock_config_c) begin
  if rising_edge(clock_config_c) then
    if i2 = "1" then
      n11 <= "000000000000000000";
    elsif n10 = "1" then
      n11 <= i3;
    end if;
  end if;
end process;
n12 <= n11(17 downto 17);
n13 <= n11(16 downto 16) &
  n11(15 downto 15) &
  n11(14 downto 14);
n14 <= n11(13 downto 13) &
  n11(12 downto 12) &
  n11(11 downto 11);
n15 <= n11(10 downto 10) &
  n11(9 downto 9) &
  n11(8 downto 8);
n16 <= n11(7 downto 7) &
  n11(6 downto 6) &
  n11(5 downto 5) &
  n11(4 downto 4) &
  n11(3 downto 3) &
  n11(2 downto 2) &
  n11(1 downto 1) &
  n11(0 downto 0);
n17 <= n9(1 downto 1);
process (clock_config_c) begin
  if rising_edge(clock_config_c) then
    if i2 = "1" then
      n18 <= "000000000000000000";
    elsif n17 = "1" then
      n18 <= i3;
    end if;
  end if;
end process;
n19 <= n18(17 downto 17);
n20 <= n18(16 downto 16) &
  n18(15 downto 15) &
  n18(14 downto 14);
n21 <= n18(13 downto 13) &
  n18(12 downto 12) &
  n18(11 downto 11);
n22 <= n18(10 downto 10) &
  n18(9 downto 9) &
  n18(8 downto 8);
n23 <= n18(7 downto 7) &
  n18(6 downto 6) &
  n18(5 downto 5) &
  n18(4 downto 4) &
  n18(3 downto 3) &
  n18(2 downto 2) &
  n18(1 downto 1) &
  n18(0 downto 0);
n24 <= n9(2 downto 2);
process (clock_config_c) begin
  if rising_edge(clock_config_c) then
    if i2 = "1" then
      n25 <= "000000000000000000";
    elsif n24 = "1" then
      n25 <= i3;
    end if;
  end if;
end process;
n26 <= n25(17 downto 17);
n27 <= n25(16 downto 16) &
  n25(15 downto 15) &
  n25(14 downto 14);
n28 <= n25(13 downto 13) &
  n25(12 downto 12) &
  n25(11 downto 11);
n29 <= n25(10 downto 10) &
  n25(9 downto 9) &
  n25(8 downto 8);
n30 <= n25(7 downto 7) &
  n25(6 downto 6) &
  n25(5 downto 5) &
  n25(4 downto 4) &
  n25(3 downto 3) &
  n25(2 downto 2) &
  n25(1 downto 1) &
  n25(0 downto 0);
n31 <= n9(3 downto 3);
process (clock_config_c) begin
  if rising_edge(clock_config_c) then
    if i2 = "1" then
      n32 <= "000000000000000000";
    elsif n31 = "1" then
      n32 <= i3;
    end if;
  end if;
end process;
n33 <= n32(17 downto 17);
n34 <= n32(16 downto 16) &
  n32(15 downto 15) &
  n32(14 downto 14);
n35 <= n32(13 downto 13) &
  n32(12 downto 12) &
  n32(11 downto 11);
n36 <= n32(10 downto 10) &
  n32(9 downto 9) &
  n32(8 downto 8);
n37 <= n32(7 downto 7) &
  n32(6 downto 6) &
  n32(5 downto 5) &
  n32(4 downto 4) &
  n32(3 downto 3) &
  n32(2 downto 2) &
  n32(1 downto 1) &
  n32(0 downto 0);
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n38 <= "0";
    elsif i1 = "1" then
      n38 <= i7;
    end if;
  end if;
end process;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n39 <= "0";
    elsif i1 = "1" then
      n39 <= i5;
    end if;
  end if;
end process;
n40 <= n16(7 downto 7);
n41 <= n16(6 downto 6) &
  n16(5 downto 5) &
  n16(4 downto 4) &
  n16(3 downto 3) &
  n16(2 downto 2) &
  n16(1 downto 1) &
  n16(0 downto 0);
n42 <= n41(6 downto 6);
n43 <= n41(5 downto 5) &
  n41(4 downto 4) &
  n41(3 downto 3) &
  n41(2 downto 2) &
  n41(1 downto 1) &
  n41(0 downto 0);
n44 <= n43(5 downto 5);
n45 <= n43(4 downto 4) &
  n43(3 downto 3) &
  n43(2 downto 2) &
  n43(1 downto 1) &
  n43(0 downto 0);
n46 <= n45(4 downto 4);
n47 <= n45(3 downto 3) &
  n45(2 downto 2) &
  n45(1 downto 1) &
  n45(0 downto 0);
n48 <= n47(3 downto 3);
n49 <= n47(2 downto 2) &
  n47(1 downto 1) &
  n47(0 downto 0);
n50 <= n49(2 downto 2);
n51 <= n49(1 downto 1) &
  n49(0 downto 0);
n52 <= n51(1 downto 1);
n53 <= n51(0 downto 0);
n54 <= n53(0 downto 0);
n55 <= n23(7 downto 7);
n56 <= n23(6 downto 6) &
  n23(5 downto 5) &
  n23(4 downto 4) &
  n23(3 downto 3) &
  n23(2 downto 2) &
  n23(1 downto 1) &
  n23(0 downto 0);
n57 <= n56(6 downto 6);
n58 <= n56(5 downto 5) &
  n56(4 downto 4) &
  n56(3 downto 3) &
  n56(2 downto 2) &
  n56(1 downto 1) &
  n56(0 downto 0);
n59 <= n58(5 downto 5);
n60 <= n58(4 downto 4) &
  n58(3 downto 3) &
  n58(2 downto 2) &
  n58(1 downto 1) &
  n58(0 downto 0);
n61 <= n60(4 downto 4);
n62 <= n60(3 downto 3) &
  n60(2 downto 2) &
  n60(1 downto 1) &
  n60(0 downto 0);
n63 <= n62(3 downto 3);
n64 <= n62(2 downto 2) &
  n62(1 downto 1) &
  n62(0 downto 0);
n65 <= n64(2 downto 2);
n66 <= n64(1 downto 1) &
  n64(0 downto 0);
n67 <= n66(1 downto 1);
n68 <= n66(0 downto 0);
n69 <= n68(0 downto 0);
n70 <= n30(7 downto 7);
n71 <= n30(6 downto 6) &
  n30(5 downto 5) &
  n30(4 downto 4) &
  n30(3 downto 3) &
  n30(2 downto 2) &
  n30(1 downto 1) &
  n30(0 downto 0);
n72 <= n71(6 downto 6);
n73 <= n71(5 downto 5) &
  n71(4 downto 4) &
  n71(3 downto 3) &
  n71(2 downto 2) &
  n71(1 downto 1) &
  n71(0 downto 0);
n74 <= n73(5 downto 5);
n75 <= n73(4 downto 4) &
  n73(3 downto 3) &
  n73(2 downto 2) &
  n73(1 downto 1) &
  n73(0 downto 0);
n76 <= n75(4 downto 4);
n77 <= n75(3 downto 3) &
  n75(2 downto 2) &
  n75(1 downto 1) &
  n75(0 downto 0);
n78 <= n77(3 downto 3);
n79 <= n77(2 downto 2) &
  n77(1 downto 1) &
  n77(0 downto 0);
n80 <= n79(2 downto 2);
n81 <= n79(1 downto 1) &
  n79(0 downto 0);
n82 <= n81(1 downto 1);
n83 <= n81(0 downto 0);
n84 <= n83(0 downto 0);
n85 <= n37(7 downto 7);
n86 <= n37(6 downto 6) &
  n37(5 downto 5) &
  n37(4 downto 4) &
  n37(3 downto 3) &
  n37(2 downto 2) &
  n37(1 downto 1) &
  n37(0 downto 0);
n87 <= n86(6 downto 6);
n88 <= n86(5 downto 5) &
  n86(4 downto 4) &
  n86(3 downto 3) &
  n86(2 downto 2) &
  n86(1 downto 1) &
  n86(0 downto 0);
n89 <= n88(5 downto 5);
n90 <= n88(4 downto 4) &
  n88(3 downto 3) &
  n88(2 downto 2) &
  n88(1 downto 1) &
  n88(0 downto 0);
n91 <= n90(4 downto 4);
n92 <= n90(3 downto 3) &
  n90(2 downto 2) &
  n90(1 downto 1) &
  n90(0 downto 0);
n93 <= n92(3 downto 3);
n94 <= n92(2 downto 2) &
  n92(1 downto 1) &
  n92(0 downto 0);
n95 <= n94(2 downto 2);
n96 <= n94(1 downto 1) &
  n94(0 downto 0);
n97 <= n96(1 downto 1);
n98 <= n96(0 downto 0);
n99 <= n98(0 downto 0);
n100 <= n13(2 downto 2) &
  n13(1 downto 1);
n101 <= n13(0 downto 0);
n102 <= n309 when n101 = "1" else n38;
n103 <= n308 when n101 = "1" else n39;
n104 <= n201 when n101 = "1" else n150;
n105 <= n303 when n101 = "1" else n252;
n106 <= n100(1 downto 1);
n107 <= n100(0 downto 0);
n108 <= n103 when n107 = "1" else n102;
n109 <= n105 when n107 = "1" else n104;
n110 <= n106(0 downto 0);
n111 <= n109 when n110 = "1" else n108;
n112 <= n14(2 downto 2) &
  n14(1 downto 1);
n113 <= n14(0 downto 0);
n114 <= n309 when n113 = "1" else n38;
n115 <= n308 when n113 = "1" else n39;
n116 <= n201 when n113 = "1" else n150;
n117 <= n303 when n113 = "1" else n252;
n118 <= n112(1 downto 1);
n119 <= n112(0 downto 0);
n120 <= n115 when n119 = "1" else n114;
n121 <= n117 when n119 = "1" else n116;
n122 <= n118(0 downto 0);
n123 <= n121 when n122 = "1" else n120;
n124 <= n15(2 downto 2) &
  n15(1 downto 1);
n125 <= n15(0 downto 0);
n126 <= n309 when n125 = "1" else n38;
n127 <= n308 when n125 = "1" else n39;
n128 <= n201 when n125 = "1" else n150;
n129 <= n303 when n125 = "1" else n252;
n130 <= n124(1 downto 1);
n131 <= n124(0 downto 0);
n132 <= n127 when n131 = "1" else n126;
n133 <= n129 when n131 = "1" else n128;
n134 <= n130(0 downto 0);
n135 <= n133 when n134 = "1" else n132;
n136 <= n123 & n135;
n137 <= n111 & n136;
n138 <= n137(2 downto 2) &
  n137(1 downto 1);
n139 <= n137(0 downto 0);
n140 <= n52 when n139 = "1" else n54;
n141 <= n48 when n139 = "1" else n50;
n142 <= n44 when n139 = "1" else n46;
n143 <= n40 when n139 = "1" else n42;
n144 <= n138(1 downto 1);
n145 <= n138(0 downto 0);
n146 <= n141 when n145 = "1" else n140;
n147 <= n143 when n145 = "1" else n142;
n148 <= n144(0 downto 0);
n149 <= n147 when n148 = "1" else n146;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n150 <= "0";
    elsif i1 = "1" then
      n150 <= n149;
    end if;
  end if;
end process;
n151 <= n20(2 downto 2) &
  n20(1 downto 1);
n152 <= n20(0 downto 0);
n153 <= n309 when n152 = "1" else n38;
n154 <= n308 when n152 = "1" else n39;
n155 <= n201 when n152 = "1" else n150;
n156 <= n303 when n152 = "1" else n252;
n157 <= n151(1 downto 1);
n158 <= n151(0 downto 0);
n159 <= n154 when n158 = "1" else n153;
n160 <= n156 when n158 = "1" else n155;
n161 <= n157(0 downto 0);
n162 <= n160 when n161 = "1" else n159;
n163 <= n21(2 downto 2) &
  n21(1 downto 1);
n164 <= n21(0 downto 0);
n165 <= n309 when n164 = "1" else n38;
n166 <= n308 when n164 = "1" else n39;
n167 <= n201 when n164 = "1" else n150;
n168 <= n303 when n164 = "1" else n252;
n169 <= n163(1 downto 1);
n170 <= n163(0 downto 0);
n171 <= n166 when n170 = "1" else n165;
n172 <= n168 when n170 = "1" else n167;
n173 <= n169(0 downto 0);
n174 <= n172 when n173 = "1" else n171;
n175 <= n22(2 downto 2) &
  n22(1 downto 1);
n176 <= n22(0 downto 0);
n177 <= n309 when n176 = "1" else n38;
n178 <= n308 when n176 = "1" else n39;
n179 <= n201 when n176 = "1" else n150;
n180 <= n303 when n176 = "1" else n252;
n181 <= n175(1 downto 1);
n182 <= n175(0 downto 0);
n183 <= n178 when n182 = "1" else n177;
n184 <= n180 when n182 = "1" else n179;
n185 <= n181(0 downto 0);
n186 <= n184 when n185 = "1" else n183;
n187 <= n174 & n186;
n188 <= n162 & n187;
n189 <= n188(2 downto 2) &
  n188(1 downto 1);
n190 <= n188(0 downto 0);
n191 <= n67 when n190 = "1" else n69;
n192 <= n63 when n190 = "1" else n65;
n193 <= n59 when n190 = "1" else n61;
n194 <= n55 when n190 = "1" else n57;
n195 <= n189(1 downto 1);
n196 <= n189(0 downto 0);
n197 <= n192 when n196 = "1" else n191;
n198 <= n194 when n196 = "1" else n193;
n199 <= n195(0 downto 0);
n200 <= n198 when n199 = "1" else n197;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n201 <= "0";
    elsif i1 = "1" then
      n201 <= n200;
    end if;
  end if;
end process;
n202 <= n27(2 downto 2) &
  n27(1 downto 1);
n203 <= n27(0 downto 0);
n204 <= n309 when n203 = "1" else n38;
n205 <= n308 when n203 = "1" else n39;
n206 <= n201 when n203 = "1" else n150;
n207 <= n303 when n203 = "1" else n252;
n208 <= n202(1 downto 1);
n209 <= n202(0 downto 0);
n210 <= n205 when n209 = "1" else n204;
n211 <= n207 when n209 = "1" else n206;
n212 <= n208(0 downto 0);
n213 <= n211 when n212 = "1" else n210;
n214 <= n28(2 downto 2) &
  n28(1 downto 1);
n215 <= n28(0 downto 0);
n216 <= n309 when n215 = "1" else n38;
n217 <= n308 when n215 = "1" else n39;
n218 <= n201 when n215 = "1" else n150;
n219 <= n303 when n215 = "1" else n252;
n220 <= n214(1 downto 1);
n221 <= n214(0 downto 0);
n222 <= n217 when n221 = "1" else n216;
n223 <= n219 when n221 = "1" else n218;
n224 <= n220(0 downto 0);
n225 <= n223 when n224 = "1" else n222;
n226 <= n29(2 downto 2) &
  n29(1 downto 1);
n227 <= n29(0 downto 0);
n228 <= n309 when n227 = "1" else n38;
n229 <= n308 when n227 = "1" else n39;
n230 <= n201 when n227 = "1" else n150;
n231 <= n303 when n227 = "1" else n252;
n232 <= n226(1 downto 1);
n233 <= n226(0 downto 0);
n234 <= n229 when n233 = "1" else n228;
n235 <= n231 when n233 = "1" else n230;
n236 <= n232(0 downto 0);
n237 <= n235 when n236 = "1" else n234;
n238 <= n225 & n237;
n239 <= n213 & n238;
n240 <= n239(2 downto 2) &
  n239(1 downto 1);
n241 <= n239(0 downto 0);
n242 <= n82 when n241 = "1" else n84;
n243 <= n78 when n241 = "1" else n80;
n244 <= n74 when n241 = "1" else n76;
n245 <= n70 when n241 = "1" else n72;
n246 <= n240(1 downto 1);
n247 <= n240(0 downto 0);
n248 <= n243 when n247 = "1" else n242;
n249 <= n245 when n247 = "1" else n244;
n250 <= n246(0 downto 0);
n251 <= n249 when n250 = "1" else n248;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n252 <= "0";
    elsif i1 = "1" then
      n252 <= n251;
    end if;
  end if;
end process;
n253 <= n34(2 downto 2) &
  n34(1 downto 1);
n254 <= n34(0 downto 0);
n255 <= n309 when n254 = "1" else n38;
n256 <= n308 when n254 = "1" else n39;
n257 <= n201 when n254 = "1" else n150;
n258 <= n303 when n254 = "1" else n252;
n259 <= n253(1 downto 1);
n260 <= n253(0 downto 0);
n261 <= n256 when n260 = "1" else n255;
n262 <= n258 when n260 = "1" else n257;
n263 <= n259(0 downto 0);
n264 <= n262 when n263 = "1" else n261;
n265 <= n35(2 downto 2) &
  n35(1 downto 1);
n266 <= n35(0 downto 0);
n267 <= n309 when n266 = "1" else n38;
n268 <= n308 when n266 = "1" else n39;
n269 <= n201 when n266 = "1" else n150;
n270 <= n303 when n266 = "1" else n252;
n271 <= n265(1 downto 1);
n272 <= n265(0 downto 0);
n273 <= n268 when n272 = "1" else n267;
n274 <= n270 when n272 = "1" else n269;
n275 <= n271(0 downto 0);
n276 <= n274 when n275 = "1" else n273;
n277 <= n36(2 downto 2) &
  n36(1 downto 1);
n278 <= n36(0 downto 0);
n279 <= n309 when n278 = "1" else n38;
n280 <= n308 when n278 = "1" else n39;
n281 <= n201 when n278 = "1" else n150;
n282 <= n303 when n278 = "1" else n252;
n283 <= n277(1 downto 1);
n284 <= n277(0 downto 0);
n285 <= n280 when n284 = "1" else n279;
n286 <= n282 when n284 = "1" else n281;
n287 <= n283(0 downto 0);
n288 <= n286 when n287 = "1" else n285;
n289 <= n276 & n288;
n290 <= n264 & n289;
n291 <= n290(2 downto 2) &
  n290(1 downto 1);
n292 <= n290(0 downto 0);
n293 <= n97 when n292 = "1" else n99;
n294 <= n93 when n292 = "1" else n95;
n295 <= n89 when n292 = "1" else n91;
n296 <= n85 when n292 = "1" else n87;
n297 <= n291(1 downto 1);
n298 <= n291(0 downto 0);
n299 <= n294 when n298 = "1" else n293;
n300 <= n296 when n298 = "1" else n295;
n301 <= n297(0 downto 0);
n302 <= n300 when n301 = "1" else n299;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n303 <= "0";
    elsif i1 = "1" then
      n303 <= n302;
    end if;
  end if;
end process;
n304 <= n150 when n12 = "1" else n149;
n305 <= n201 when n19 = "1" else n200;
n306 <= n252 when n26 = "1" else n251;
n307 <= n303 when n33 = "1" else n302;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n308 <= "0";
    elsif i1 = "1" then
      n308 <= i8;
    end if;
  end if;
end process;
process (clock_main_c) begin
  if rising_edge(clock_main_c) then
    if i2 = "1" then
      n309 <= "0";
    elsif i1 = "1" then
      n309 <= i9;
    end if;
  end if;
end process;
s310 : cf_rca_16_31 port map (n1, n2, n3, n4, n5, n6, s310_1);
o4 <= n307;
o3 <= n306;
o2 <= n305;
o1 <= n304;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_28 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(2 downto 0);
i8 : in  unsigned(2 downto 0);
i9 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(2 downto 0);
o4 : out unsigned(2 downto 0));
end entity cf_rca_16_28;
architecture rtl of cf_rca_16_28 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(1 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(1 downto 0);
signal n12 : unsigned(1 downto 0);
signal n13 : unsigned(2 downto 0);
signal n14 : unsigned(2 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(1 downto 0);
signal n17 : unsigned(0 downto 0);
signal n18 : unsigned(0 downto 0);
signal n19 : unsigned(0 downto 0);
signal s20_1 : unsigned(0 downto 0);
signal s20_2 : unsigned(0 downto 0);
signal s20_3 : unsigned(0 downto 0);
signal s20_4 : unsigned(0 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(0 downto 0);
signal s21_4 : unsigned(0 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
component cf_rca_16_30 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_30;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
begin
n1 <= i7(0 downto 0);
n2 <= i8(0 downto 0);
n3 <= i7(2 downto 2) &
  i7(1 downto 1);
n4 <= i8(2 downto 2) &
  i8(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n4(0 downto 0);
n7 <= n3(1 downto 1);
n8 <= n4(1 downto 1);
n9 <= n7(0 downto 0);
n10 <= n8(0 downto 0);
n11 <= s20_1 & s21_1;
n12 <= s20_2 & s21_2;
n13 <= n11 & s22_1;
n14 <= n12 & s22_2;
n15 <= i9(0 downto 0);
n16 <= i9(2 downto 2) &
  i9(1 downto 1);
n17 <= n16(0 downto 0);
n18 <= n16(1 downto 1);
n19 <= n18(0 downto 0);
s20 : cf_rca_16_30 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, s21_4, n9, n10, n19, s20_1, s20_2, s20_3, s20_4);
s21 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, s22_4, n5, n6, s20_3, n17, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i6, n1, n2, s21_3, n15, s22_1, s22_2, s22_3, s22_4);
o4 <= n14;
o3 <= n13;
o2 <= s20_4;
o1 <= s22_3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_27 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(4 downto 0);
i8 : in  unsigned(4 downto 0);
i9 : in  unsigned(4 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(4 downto 0);
o4 : out unsigned(4 downto 0));
end entity cf_rca_16_27;
architecture rtl of cf_rca_16_27 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(3 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(2 downto 0);
signal n9 : unsigned(3 downto 0);
signal n10 : unsigned(3 downto 0);
signal n11 : unsigned(4 downto 0);
signal n12 : unsigned(4 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(3 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(2 downto 0);
signal s17_1 : unsigned(0 downto 0);
signal s17_2 : unsigned(0 downto 0);
signal s17_3 : unsigned(2 downto 0);
signal s17_4 : unsigned(2 downto 0);
signal s18_1 : unsigned(0 downto 0);
signal s18_2 : unsigned(0 downto 0);
signal s18_3 : unsigned(0 downto 0);
signal s18_4 : unsigned(0 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(0 downto 0);
signal s19_4 : unsigned(0 downto 0);
component cf_rca_16_28 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(2 downto 0);
i8 : in  unsigned(2 downto 0);
i9 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(2 downto 0);
o4 : out unsigned(2 downto 0));
end component cf_rca_16_28;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
begin
n1 <= i7(0 downto 0);
n2 <= i8(0 downto 0);
n3 <= i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n4 <= i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n4(0 downto 0);
n7 <= n3(3 downto 3) &
  n3(2 downto 2) &
  n3(1 downto 1);
n8 <= n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1);
n9 <= s17_3 & s18_1;
n10 <= s17_4 & s18_2;
n11 <= n9 & s19_1;
n12 <= n10 & s19_2;
n13 <= i9(0 downto 0);
n14 <= i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n15 <= n14(0 downto 0);
n16 <= n14(3 downto 3) &
  n14(2 downto 2) &
  n14(1 downto 1);
s17 : cf_rca_16_28 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, s18_4, n7, n8, n16, s17_1, s17_2, s17_3, s17_4);
s18 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, s19_4, n5, n6, s17_1, n15, s18_1, s18_2, s18_3, s18_4);
s19 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i6, n1, n2, s18_3, n13, s19_1, s19_2, s19_3, s19_4);
o4 <= n12;
o3 <= n11;
o2 <= s17_2;
o1 <= s19_3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_26 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(6 downto 0);
i8 : in  unsigned(6 downto 0);
i9 : in  unsigned(6 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(6 downto 0);
o4 : out unsigned(6 downto 0));
end entity cf_rca_16_26;
architecture rtl of cf_rca_16_26 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(5 downto 0);
signal n4 : unsigned(5 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(4 downto 0);
signal n8 : unsigned(4 downto 0);
signal n9 : unsigned(5 downto 0);
signal n10 : unsigned(5 downto 0);
signal n11 : unsigned(6 downto 0);
signal n12 : unsigned(6 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(5 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(4 downto 0);
signal s17_1 : unsigned(0 downto 0);
signal s17_2 : unsigned(0 downto 0);
signal s17_3 : unsigned(4 downto 0);
signal s17_4 : unsigned(4 downto 0);
signal s18_1 : unsigned(0 downto 0);
signal s18_2 : unsigned(0 downto 0);
signal s18_3 : unsigned(0 downto 0);
signal s18_4 : unsigned(0 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(0 downto 0);
signal s19_4 : unsigned(0 downto 0);
component cf_rca_16_27 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(4 downto 0);
i8 : in  unsigned(4 downto 0);
i9 : in  unsigned(4 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(4 downto 0);
o4 : out unsigned(4 downto 0));
end component cf_rca_16_27;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
begin
n1 <= i7(0 downto 0);
n2 <= i8(0 downto 0);
n3 <= i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n4 <= i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n4(0 downto 0);
n7 <= n3(5 downto 5) &
  n3(4 downto 4) &
  n3(3 downto 3) &
  n3(2 downto 2) &
  n3(1 downto 1);
n8 <= n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1);
n9 <= s17_3 & s18_1;
n10 <= s17_4 & s18_2;
n11 <= n9 & s19_1;
n12 <= n10 & s19_2;
n13 <= i9(0 downto 0);
n14 <= i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n15 <= n14(0 downto 0);
n16 <= n14(5 downto 5) &
  n14(4 downto 4) &
  n14(3 downto 3) &
  n14(2 downto 2) &
  n14(1 downto 1);
s17 : cf_rca_16_27 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, s18_4, n7, n8, n16, s17_1, s17_2, s17_3, s17_4);
s18 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, s19_4, n5, n6, s17_1, n15, s18_1, s18_2, s18_3, s18_4);
s19 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i6, n1, n2, s18_3, n13, s19_1, s19_2, s19_3, s19_4);
o4 <= n12;
o3 <= n11;
o2 <= s17_2;
o1 <= s19_3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_25 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(8 downto 0);
i8 : in  unsigned(8 downto 0);
i9 : in  unsigned(8 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(8 downto 0);
o4 : out unsigned(8 downto 0));
end entity cf_rca_16_25;
architecture rtl of cf_rca_16_25 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(7 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(6 downto 0);
signal n8 : unsigned(6 downto 0);
signal n9 : unsigned(7 downto 0);
signal n10 : unsigned(7 downto 0);
signal n11 : unsigned(8 downto 0);
signal n12 : unsigned(8 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(7 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(6 downto 0);
signal s17_1 : unsigned(0 downto 0);
signal s17_2 : unsigned(0 downto 0);
signal s17_3 : unsigned(6 downto 0);
signal s17_4 : unsigned(6 downto 0);
signal s18_1 : unsigned(0 downto 0);
signal s18_2 : unsigned(0 downto 0);
signal s18_3 : unsigned(0 downto 0);
signal s18_4 : unsigned(0 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(0 downto 0);
signal s19_4 : unsigned(0 downto 0);
component cf_rca_16_26 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(6 downto 0);
i8 : in  unsigned(6 downto 0);
i9 : in  unsigned(6 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(6 downto 0);
o4 : out unsigned(6 downto 0));
end component cf_rca_16_26;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
begin
n1 <= i7(0 downto 0);
n2 <= i8(0 downto 0);
n3 <= i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n4 <= i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n4(0 downto 0);
n7 <= n3(7 downto 7) &
  n3(6 downto 6) &
  n3(5 downto 5) &
  n3(4 downto 4) &
  n3(3 downto 3) &
  n3(2 downto 2) &
  n3(1 downto 1);
n8 <= n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1);
n9 <= s17_3 & s18_1;
n10 <= s17_4 & s18_2;
n11 <= n9 & s19_1;
n12 <= n10 & s19_2;
n13 <= i9(0 downto 0);
n14 <= i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n15 <= n14(0 downto 0);
n16 <= n14(7 downto 7) &
  n14(6 downto 6) &
  n14(5 downto 5) &
  n14(4 downto 4) &
  n14(3 downto 3) &
  n14(2 downto 2) &
  n14(1 downto 1);
s17 : cf_rca_16_26 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, s18_4, n7, n8, n16, s17_1, s17_2, s17_3, s17_4);
s18 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, s19_4, n5, n6, s17_1, n15, s18_1, s18_2, s18_3, s18_4);
s19 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i6, n1, n2, s18_3, n13, s19_1, s19_2, s19_3, s19_4);
o4 <= n12;
o3 <= n11;
o2 <= s17_2;
o1 <= s19_3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_24 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(10 downto 0);
i8 : in  unsigned(10 downto 0);
i9 : in  unsigned(10 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(10 downto 0);
o4 : out unsigned(10 downto 0));
end entity cf_rca_16_24;
architecture rtl of cf_rca_16_24 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(9 downto 0);
signal n4 : unsigned(9 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0);
signal n9 : unsigned(9 downto 0);
signal n10 : unsigned(9 downto 0);
signal n11 : unsigned(10 downto 0);
signal n12 : unsigned(10 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(9 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(8 downto 0);
signal s17_1 : unsigned(0 downto 0);
signal s17_2 : unsigned(0 downto 0);
signal s17_3 : unsigned(8 downto 0);
signal s17_4 : unsigned(8 downto 0);
signal s18_1 : unsigned(0 downto 0);
signal s18_2 : unsigned(0 downto 0);
signal s18_3 : unsigned(0 downto 0);
signal s18_4 : unsigned(0 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(0 downto 0);
signal s19_4 : unsigned(0 downto 0);
component cf_rca_16_25 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(8 downto 0);
i8 : in  unsigned(8 downto 0);
i9 : in  unsigned(8 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(8 downto 0);
o4 : out unsigned(8 downto 0));
end component cf_rca_16_25;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
begin
n1 <= i7(0 downto 0);
n2 <= i8(0 downto 0);
n3 <= i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n4 <= i8(10 downto 10) &
  i8(9 downto 9) &
  i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n4(0 downto 0);
n7 <= n3(9 downto 9) &
  n3(8 downto 8) &
  n3(7 downto 7) &
  n3(6 downto 6) &
  n3(5 downto 5) &
  n3(4 downto 4) &
  n3(3 downto 3) &
  n3(2 downto 2) &
  n3(1 downto 1);
n8 <= n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1);
n9 <= s17_3 & s18_1;
n10 <= s17_4 & s18_2;
n11 <= n9 & s19_1;
n12 <= n10 & s19_2;
n13 <= i9(0 downto 0);
n14 <= i9(10 downto 10) &
  i9(9 downto 9) &
  i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n15 <= n14(0 downto 0);
n16 <= n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7) &
  n14(6 downto 6) &
  n14(5 downto 5) &
  n14(4 downto 4) &
  n14(3 downto 3) &
  n14(2 downto 2) &
  n14(1 downto 1);
s17 : cf_rca_16_25 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, s18_4, n7, n8, n16, s17_1, s17_2, s17_3, s17_4);
s18 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, s19_4, n5, n6, s17_1, n15, s18_1, s18_2, s18_3, s18_4);
s19 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i6, n1, n2, s18_3, n13, s19_1, s19_2, s19_3, s19_4);
o4 <= n12;
o3 <= n11;
o2 <= s17_2;
o1 <= s19_3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_23 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(12 downto 0);
i8 : in  unsigned(12 downto 0);
i9 : in  unsigned(12 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(12 downto 0);
o4 : out unsigned(12 downto 0));
end entity cf_rca_16_23;
architecture rtl of cf_rca_16_23 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(11 downto 0);
signal n4 : unsigned(11 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(10 downto 0);
signal n8 : unsigned(10 downto 0);
signal n9 : unsigned(11 downto 0);
signal n10 : unsigned(11 downto 0);
signal n11 : unsigned(12 downto 0);
signal n12 : unsigned(12 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(11 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(10 downto 0);
signal s17_1 : unsigned(0 downto 0);
signal s17_2 : unsigned(0 downto 0);
signal s17_3 : unsigned(10 downto 0);
signal s17_4 : unsigned(10 downto 0);
signal s18_1 : unsigned(0 downto 0);
signal s18_2 : unsigned(0 downto 0);
signal s18_3 : unsigned(0 downto 0);
signal s18_4 : unsigned(0 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(0 downto 0);
signal s19_4 : unsigned(0 downto 0);
component cf_rca_16_24 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(10 downto 0);
i8 : in  unsigned(10 downto 0);
i9 : in  unsigned(10 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(10 downto 0);
o4 : out unsigned(10 downto 0));
end component cf_rca_16_24;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
begin
n1 <= i7(0 downto 0);
n2 <= i8(0 downto 0);
n3 <= i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n4 <= i8(12 downto 12) &
  i8(11 downto 11) &
  i8(10 downto 10) &
  i8(9 downto 9) &
  i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n4(0 downto 0);
n7 <= n3(11 downto 11) &
  n3(10 downto 10) &
  n3(9 downto 9) &
  n3(8 downto 8) &
  n3(7 downto 7) &
  n3(6 downto 6) &
  n3(5 downto 5) &
  n3(4 downto 4) &
  n3(3 downto 3) &
  n3(2 downto 2) &
  n3(1 downto 1);
n8 <= n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1);
n9 <= s17_3 & s18_1;
n10 <= s17_4 & s18_2;
n11 <= n9 & s19_1;
n12 <= n10 & s19_2;
n13 <= i9(0 downto 0);
n14 <= i9(12 downto 12) &
  i9(11 downto 11) &
  i9(10 downto 10) &
  i9(9 downto 9) &
  i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n15 <= n14(0 downto 0);
n16 <= n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7) &
  n14(6 downto 6) &
  n14(5 downto 5) &
  n14(4 downto 4) &
  n14(3 downto 3) &
  n14(2 downto 2) &
  n14(1 downto 1);
s17 : cf_rca_16_24 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, s18_4, n7, n8, n16, s17_1, s17_2, s17_3, s17_4);
s18 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, s19_4, n5, n6, s17_1, n15, s18_1, s18_2, s18_3, s18_4);
s19 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i6, n1, n2, s18_3, n13, s19_1, s19_2, s19_3, s19_4);
o4 <= n12;
o3 <= n11;
o2 <= s17_2;
o1 <= s19_3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end entity cf_rca_16_22;
architecture rtl of cf_rca_16_22 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(13 downto 0);
signal n4 : unsigned(13 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(12 downto 0);
signal n8 : unsigned(12 downto 0);
signal n9 : unsigned(13 downto 0);
signal n10 : unsigned(13 downto 0);
signal n11 : unsigned(14 downto 0);
signal n12 : unsigned(14 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(13 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(12 downto 0);
signal s17_1 : unsigned(0 downto 0);
signal s17_2 : unsigned(0 downto 0);
signal s17_3 : unsigned(12 downto 0);
signal s17_4 : unsigned(12 downto 0);
signal s18_1 : unsigned(0 downto 0);
signal s18_2 : unsigned(0 downto 0);
signal s18_3 : unsigned(0 downto 0);
signal s18_4 : unsigned(0 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(0 downto 0);
signal s19_4 : unsigned(0 downto 0);
component cf_rca_16_23 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(12 downto 0);
i8 : in  unsigned(12 downto 0);
i9 : in  unsigned(12 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(12 downto 0);
o4 : out unsigned(12 downto 0));
end component cf_rca_16_23;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
begin
n1 <= i7(0 downto 0);
n2 <= i8(0 downto 0);
n3 <= i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n4 <= i8(14 downto 14) &
  i8(13 downto 13) &
  i8(12 downto 12) &
  i8(11 downto 11) &
  i8(10 downto 10) &
  i8(9 downto 9) &
  i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n4(0 downto 0);
n7 <= n3(13 downto 13) &
  n3(12 downto 12) &
  n3(11 downto 11) &
  n3(10 downto 10) &
  n3(9 downto 9) &
  n3(8 downto 8) &
  n3(7 downto 7) &
  n3(6 downto 6) &
  n3(5 downto 5) &
  n3(4 downto 4) &
  n3(3 downto 3) &
  n3(2 downto 2) &
  n3(1 downto 1);
n8 <= n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1);
n9 <= s17_3 & s18_1;
n10 <= s17_4 & s18_2;
n11 <= n9 & s19_1;
n12 <= n10 & s19_2;
n13 <= i9(0 downto 0);
n14 <= i9(14 downto 14) &
  i9(13 downto 13) &
  i9(12 downto 12) &
  i9(11 downto 11) &
  i9(10 downto 10) &
  i9(9 downto 9) &
  i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n15 <= n14(0 downto 0);
n16 <= n14(13 downto 13) &
  n14(12 downto 12) &
  n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7) &
  n14(6 downto 6) &
  n14(5 downto 5) &
  n14(4 downto 4) &
  n14(3 downto 3) &
  n14(2 downto 2) &
  n14(1 downto 1);
s17 : cf_rca_16_23 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, s18_4, n7, n8, n16, s17_1, s17_2, s17_3, s17_4);
s18 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, s19_4, n5, n6, s17_1, n15, s18_1, s18_2, s18_3, s18_4);
s19 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i6, n1, n2, s18_3, n13, s19_1, s19_2, s19_3, s19_4);
o4 <= n12;
o3 <= n11;
o2 <= s17_2;
o1 <= s19_3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_21 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(8 downto 0);
i8 : in  unsigned(8 downto 0);
i9 : in  unsigned(8 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(8 downto 0);
o4 : out unsigned(8 downto 0));
end entity cf_rca_16_21;
architecture rtl of cf_rca_16_21 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(7 downto 0);
signal n4 : unsigned(7 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(6 downto 0);
signal n8 : unsigned(6 downto 0);
signal n9 : unsigned(7 downto 0);
signal n10 : unsigned(7 downto 0);
signal n11 : unsigned(8 downto 0);
signal n12 : unsigned(8 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(7 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(6 downto 0);
signal s17_1 : unsigned(0 downto 0);
signal s17_2 : unsigned(0 downto 0);
signal s17_3 : unsigned(0 downto 0);
signal s17_4 : unsigned(0 downto 0);
signal s18_1 : unsigned(0 downto 0);
signal s18_2 : unsigned(0 downto 0);
signal s18_3 : unsigned(6 downto 0);
signal s18_4 : unsigned(6 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(0 downto 0);
signal s19_4 : unsigned(0 downto 0);
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_26 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(6 downto 0);
i8 : in  unsigned(6 downto 0);
i9 : in  unsigned(6 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(6 downto 0);
o4 : out unsigned(6 downto 0));
end component cf_rca_16_26;
begin
n1 <= i7(0 downto 0);
n2 <= i8(0 downto 0);
n3 <= i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n4 <= i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n4(0 downto 0);
n7 <= n3(7 downto 7) &
  n3(6 downto 6) &
  n3(5 downto 5) &
  n3(4 downto 4) &
  n3(3 downto 3) &
  n3(2 downto 2) &
  n3(1 downto 1);
n8 <= n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1);
n9 <= s18_3 & s17_1;
n10 <= s18_4 & s17_2;
n11 <= n9 & s19_1;
n12 <= n10 & s19_2;
n13 <= i9(0 downto 0);
n14 <= i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n15 <= n14(0 downto 0);
n16 <= n14(7 downto 7) &
  n14(6 downto 6) &
  n14(5 downto 5) &
  n14(4 downto 4) &
  n14(3 downto 3) &
  n14(2 downto 2) &
  n14(1 downto 1);
s17 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, s19_4, n5, n6, s18_1, n15, s17_1, s17_2, s17_3, s17_4);
s18 : cf_rca_16_26 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, s17_4, n7, n8, n16, s18_1, s18_2, s18_3, s18_4);
s19 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i6, n1, n2, s17_3, n13, s19_1, s19_2, s19_3, s19_4);
o4 <= n12;
o3 <= n11;
o2 <= s18_2;
o1 <= s19_3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_20 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(10 downto 0);
i8 : in  unsigned(10 downto 0);
i9 : in  unsigned(10 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(10 downto 0);
o4 : out unsigned(10 downto 0));
end entity cf_rca_16_20;
architecture rtl of cf_rca_16_20 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(9 downto 0);
signal n4 : unsigned(9 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(8 downto 0);
signal n9 : unsigned(9 downto 0);
signal n10 : unsigned(9 downto 0);
signal n11 : unsigned(10 downto 0);
signal n12 : unsigned(10 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(9 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(8 downto 0);
signal s17_1 : unsigned(0 downto 0);
signal s17_2 : unsigned(0 downto 0);
signal s17_3 : unsigned(0 downto 0);
signal s17_4 : unsigned(0 downto 0);
signal s18_1 : unsigned(0 downto 0);
signal s18_2 : unsigned(0 downto 0);
signal s18_3 : unsigned(8 downto 0);
signal s18_4 : unsigned(8 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(0 downto 0);
signal s19_4 : unsigned(0 downto 0);
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_21 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(8 downto 0);
i8 : in  unsigned(8 downto 0);
i9 : in  unsigned(8 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(8 downto 0);
o4 : out unsigned(8 downto 0));
end component cf_rca_16_21;
begin
n1 <= i7(0 downto 0);
n2 <= i8(0 downto 0);
n3 <= i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n4 <= i8(10 downto 10) &
  i8(9 downto 9) &
  i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n4(0 downto 0);
n7 <= n3(9 downto 9) &
  n3(8 downto 8) &
  n3(7 downto 7) &
  n3(6 downto 6) &
  n3(5 downto 5) &
  n3(4 downto 4) &
  n3(3 downto 3) &
  n3(2 downto 2) &
  n3(1 downto 1);
n8 <= n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1);
n9 <= s18_3 & s17_1;
n10 <= s18_4 & s17_2;
n11 <= n9 & s19_1;
n12 <= n10 & s19_2;
n13 <= i9(0 downto 0);
n14 <= i9(10 downto 10) &
  i9(9 downto 9) &
  i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n15 <= n14(0 downto 0);
n16 <= n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7) &
  n14(6 downto 6) &
  n14(5 downto 5) &
  n14(4 downto 4) &
  n14(3 downto 3) &
  n14(2 downto 2) &
  n14(1 downto 1);
s17 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, s19_4, n5, n6, s18_1, n15, s17_1, s17_2, s17_3, s17_4);
s18 : cf_rca_16_21 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, s17_4, n7, n8, n16, s18_1, s18_2, s18_3, s18_4);
s19 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i6, n1, n2, s17_3, n13, s19_1, s19_2, s19_3, s19_4);
o4 <= n12;
o3 <= n11;
o2 <= s18_2;
o1 <= s19_3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_19 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(12 downto 0);
i8 : in  unsigned(12 downto 0);
i9 : in  unsigned(12 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(12 downto 0);
o4 : out unsigned(12 downto 0));
end entity cf_rca_16_19;
architecture rtl of cf_rca_16_19 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(11 downto 0);
signal n4 : unsigned(11 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(10 downto 0);
signal n8 : unsigned(10 downto 0);
signal n9 : unsigned(11 downto 0);
signal n10 : unsigned(11 downto 0);
signal n11 : unsigned(12 downto 0);
signal n12 : unsigned(12 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(11 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(10 downto 0);
signal s17_1 : unsigned(0 downto 0);
signal s17_2 : unsigned(0 downto 0);
signal s17_3 : unsigned(0 downto 0);
signal s17_4 : unsigned(0 downto 0);
signal s18_1 : unsigned(0 downto 0);
signal s18_2 : unsigned(0 downto 0);
signal s18_3 : unsigned(10 downto 0);
signal s18_4 : unsigned(10 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(0 downto 0);
signal s19_4 : unsigned(0 downto 0);
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_20 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(10 downto 0);
i8 : in  unsigned(10 downto 0);
i9 : in  unsigned(10 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(10 downto 0);
o4 : out unsigned(10 downto 0));
end component cf_rca_16_20;
begin
n1 <= i7(0 downto 0);
n2 <= i8(0 downto 0);
n3 <= i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n4 <= i8(12 downto 12) &
  i8(11 downto 11) &
  i8(10 downto 10) &
  i8(9 downto 9) &
  i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n4(0 downto 0);
n7 <= n3(11 downto 11) &
  n3(10 downto 10) &
  n3(9 downto 9) &
  n3(8 downto 8) &
  n3(7 downto 7) &
  n3(6 downto 6) &
  n3(5 downto 5) &
  n3(4 downto 4) &
  n3(3 downto 3) &
  n3(2 downto 2) &
  n3(1 downto 1);
n8 <= n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1);
n9 <= s18_3 & s17_1;
n10 <= s18_4 & s17_2;
n11 <= n9 & s19_1;
n12 <= n10 & s19_2;
n13 <= i9(0 downto 0);
n14 <= i9(12 downto 12) &
  i9(11 downto 11) &
  i9(10 downto 10) &
  i9(9 downto 9) &
  i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n15 <= n14(0 downto 0);
n16 <= n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7) &
  n14(6 downto 6) &
  n14(5 downto 5) &
  n14(4 downto 4) &
  n14(3 downto 3) &
  n14(2 downto 2) &
  n14(1 downto 1);
s17 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, s19_4, n5, n6, s18_1, n15, s17_1, s17_2, s17_3, s17_4);
s18 : cf_rca_16_20 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, s17_4, n7, n8, n16, s18_1, s18_2, s18_3, s18_4);
s19 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i6, n1, n2, s17_3, n13, s19_1, s19_2, s19_3, s19_4);
o4 <= n12;
o3 <= n11;
o2 <= s18_2;
o1 <= s19_3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_18 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end entity cf_rca_16_18;
architecture rtl of cf_rca_16_18 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(13 downto 0);
signal n4 : unsigned(13 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(12 downto 0);
signal n8 : unsigned(12 downto 0);
signal n9 : unsigned(13 downto 0);
signal n10 : unsigned(13 downto 0);
signal n11 : unsigned(14 downto 0);
signal n12 : unsigned(14 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(13 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(12 downto 0);
signal s17_1 : unsigned(0 downto 0);
signal s17_2 : unsigned(0 downto 0);
signal s17_3 : unsigned(0 downto 0);
signal s17_4 : unsigned(0 downto 0);
signal s18_1 : unsigned(0 downto 0);
signal s18_2 : unsigned(0 downto 0);
signal s18_3 : unsigned(12 downto 0);
signal s18_4 : unsigned(12 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(0 downto 0);
signal s19_4 : unsigned(0 downto 0);
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_19 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(12 downto 0);
i8 : in  unsigned(12 downto 0);
i9 : in  unsigned(12 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(12 downto 0);
o4 : out unsigned(12 downto 0));
end component cf_rca_16_19;
begin
n1 <= i7(0 downto 0);
n2 <= i8(0 downto 0);
n3 <= i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n4 <= i8(14 downto 14) &
  i8(13 downto 13) &
  i8(12 downto 12) &
  i8(11 downto 11) &
  i8(10 downto 10) &
  i8(9 downto 9) &
  i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n4(0 downto 0);
n7 <= n3(13 downto 13) &
  n3(12 downto 12) &
  n3(11 downto 11) &
  n3(10 downto 10) &
  n3(9 downto 9) &
  n3(8 downto 8) &
  n3(7 downto 7) &
  n3(6 downto 6) &
  n3(5 downto 5) &
  n3(4 downto 4) &
  n3(3 downto 3) &
  n3(2 downto 2) &
  n3(1 downto 1);
n8 <= n4(13 downto 13) &
  n4(12 downto 12) &
  n4(11 downto 11) &
  n4(10 downto 10) &
  n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1);
n9 <= s18_3 & s17_1;
n10 <= s18_4 & s17_2;
n11 <= n9 & s19_1;
n12 <= n10 & s19_2;
n13 <= i9(0 downto 0);
n14 <= i9(14 downto 14) &
  i9(13 downto 13) &
  i9(12 downto 12) &
  i9(11 downto 11) &
  i9(10 downto 10) &
  i9(9 downto 9) &
  i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n15 <= n14(0 downto 0);
n16 <= n14(13 downto 13) &
  n14(12 downto 12) &
  n14(11 downto 11) &
  n14(10 downto 10) &
  n14(9 downto 9) &
  n14(8 downto 8) &
  n14(7 downto 7) &
  n14(6 downto 6) &
  n14(5 downto 5) &
  n14(4 downto 4) &
  n14(3 downto 3) &
  n14(2 downto 2) &
  n14(1 downto 1);
s17 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, s19_4, n5, n6, s18_1, n15, s17_1, s17_2, s17_3, s17_4);
s18 : cf_rca_16_19 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, s17_4, n7, n8, n16, s18_1, s18_2, s18_3, s18_4);
s19 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i6, n1, n2, s17_3, n13, s19_1, s19_2, s19_3, s19_4);
o4 <= n12;
o3 <= n11;
o2 <= s18_2;
o1 <= s19_3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_17 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
i10 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0));
end entity cf_rca_16_17;
architecture rtl of cf_rca_16_17 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(14 downto 0);
signal s14_1 : unsigned(15 downto 0);
signal s14_2 : unsigned(15 downto 0);
signal s14_3 : unsigned(15 downto 0);
signal s14_4 : unsigned(15 downto 0);
signal s14_5 : unsigned(15 downto 0);
signal s14_6 : unsigned(15 downto 0);
signal s14_7 : unsigned(15 downto 0);
signal s14_8 : unsigned(15 downto 0);
signal s14_9 : unsigned(15 downto 0);
signal s14_10 : unsigned(15 downto 0);
signal s14_11 : unsigned(15 downto 0);
signal s14_12 : unsigned(15 downto 0);
signal s14_13 : unsigned(15 downto 0);
signal s14_14 : unsigned(15 downto 0);
signal s14_15 : unsigned(15 downto 0);
signal s14_16 : unsigned(15 downto 0);
signal s15_1 : unsigned(15 downto 0);
signal s16_1 : unsigned(0 downto 0);
signal s16_2 : unsigned(0 downto 0);
signal s16_3 : unsigned(14 downto 0);
signal s16_4 : unsigned(14 downto 0);
signal s17_1 : unsigned(0 downto 0);
signal s17_2 : unsigned(0 downto 0);
signal s17_3 : unsigned(0 downto 0);
signal s17_4 : unsigned(0 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s15_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s15_1(15 downto 15) &
  s15_1(14 downto 14) &
  s15_1(13 downto 13) &
  s15_1(12 downto 12) &
  s15_1(11 downto 11) &
  s15_1(10 downto 10) &
  s15_1(9 downto 9) &
  s15_1(8 downto 8) &
  s15_1(7 downto 7) &
  s15_1(6 downto 6) &
  s15_1(5 downto 5) &
  s15_1(4 downto 4) &
  s15_1(3 downto 3) &
  s15_1(2 downto 2) &
  s15_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s16_3 & s17_1;
n11 <= s16_4 & s17_2;
n12 <= i4(0 downto 0);
n13 <= i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5) &
  i4(4 downto 4) &
  i4(3 downto 3) &
  i4(2 downto 2) &
  i4(1 downto 1);
s14 : cf_rca_16_38 port map (s14_1, s14_2, s14_3, s14_4, s14_5, s14_6, s14_7, s14_8, s14_9, s14_10, s14_11, s14_12, s14_13, s14_14, s14_15, s14_16);
s15 : cf_rca_16_32 port map (n2, s14_1, s14_2, s14_3, s14_4, s14_5, s14_6, s14_7, s14_8, s14_9, s14_10, s14_11, s14_12, s14_13, s14_14, s14_15, s14_16, n3, s15_1);
s16 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s17_4, n8, n9, n13, s16_1, s16_2, s16_3, s16_4);
s17 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s16_1, n12, s17_1, s17_2, s17_3, s17_4);
o4 <= n11;
o3 <= n10;
o2 <= s16_2;
o1 <= s17_3;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_16 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(1 downto 0);
i9 : in  unsigned(1 downto 0);
i10 : in  unsigned(1 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(1 downto 0);
o4 : out unsigned(1 downto 0));
end entity cf_rca_16_16;
architecture rtl of cf_rca_16_16 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(0 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(1 downto 0);
signal n18 : unsigned(1 downto 0);
signal s19_1 : unsigned(15 downto 0);
signal s19_2 : unsigned(15 downto 0);
signal s19_3 : unsigned(15 downto 0);
signal s19_4 : unsigned(15 downto 0);
signal s19_5 : unsigned(15 downto 0);
signal s19_6 : unsigned(15 downto 0);
signal s19_7 : unsigned(15 downto 0);
signal s19_8 : unsigned(15 downto 0);
signal s19_9 : unsigned(15 downto 0);
signal s19_10 : unsigned(15 downto 0);
signal s19_11 : unsigned(15 downto 0);
signal s19_12 : unsigned(15 downto 0);
signal s19_13 : unsigned(15 downto 0);
signal s19_14 : unsigned(15 downto 0);
signal s19_15 : unsigned(15 downto 0);
signal s19_16 : unsigned(15 downto 0);
signal s20_1 : unsigned(15 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(14 downto 0);
signal s21_4 : unsigned(14 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
signal s23_1 : unsigned(0 downto 0);
signal s23_2 : unsigned(0 downto 0);
signal s23_3 : unsigned(15 downto 0);
signal s23_4 : unsigned(15 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_17 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
i10 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0));
end component cf_rca_16_17;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s20_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s20_1(15 downto 15) &
  s20_1(14 downto 14) &
  s20_1(13 downto 13) &
  s20_1(12 downto 12) &
  s20_1(11 downto 11) &
  s20_1(10 downto 10) &
  s20_1(9 downto 9) &
  s20_1(8 downto 8) &
  s20_1(7 downto 7) &
  s20_1(6 downto 6) &
  s20_1(5 downto 5) &
  s20_1(4 downto 4) &
  s20_1(3 downto 3) &
  s20_1(2 downto 2) &
  s20_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s21_3 & s22_1;
n11 <= s21_4 & s22_2;
n12 <= i8(1 downto 1);
n13 <= i9(1 downto 1);
n14 <= i10(1 downto 1);
n15 <= s23_3(0 downto 0);
n16 <= s23_3(15 downto 15) &
  s23_3(14 downto 14) &
  s23_3(13 downto 13) &
  s23_3(12 downto 12) &
  s23_3(11 downto 11) &
  s23_3(10 downto 10) &
  s23_3(9 downto 9) &
  s23_3(8 downto 8) &
  s23_3(7 downto 7) &
  s23_3(6 downto 6) &
  s23_3(5 downto 5) &
  s23_3(4 downto 4) &
  s23_3(3 downto 3) &
  s23_3(2 downto 2) &
  s23_3(1 downto 1);
n17 <= s23_1 & s22_3;
n18 <= s23_2 & s21_2;
s19 : cf_rca_16_38 port map (s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16);
s20 : cf_rca_16_32 port map (n2, s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16, n3, s20_1);
s21 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s22_4, n8, n9, n16, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s21_1, n15, s22_1, s22_2, s22_3, s22_4);
s23 : cf_rca_16_17 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_4;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_15 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(2 downto 0);
i9 : in  unsigned(2 downto 0);
i10 : in  unsigned(2 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(2 downto 0);
o4 : out unsigned(2 downto 0));
end entity cf_rca_16_15;
architecture rtl of cf_rca_16_15 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(1 downto 0);
signal n13 : unsigned(1 downto 0);
signal n14 : unsigned(1 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(2 downto 0);
signal n18 : unsigned(2 downto 0);
signal s19_1 : unsigned(15 downto 0);
signal s19_2 : unsigned(15 downto 0);
signal s19_3 : unsigned(15 downto 0);
signal s19_4 : unsigned(15 downto 0);
signal s19_5 : unsigned(15 downto 0);
signal s19_6 : unsigned(15 downto 0);
signal s19_7 : unsigned(15 downto 0);
signal s19_8 : unsigned(15 downto 0);
signal s19_9 : unsigned(15 downto 0);
signal s19_10 : unsigned(15 downto 0);
signal s19_11 : unsigned(15 downto 0);
signal s19_12 : unsigned(15 downto 0);
signal s19_13 : unsigned(15 downto 0);
signal s19_14 : unsigned(15 downto 0);
signal s19_15 : unsigned(15 downto 0);
signal s19_16 : unsigned(15 downto 0);
signal s20_1 : unsigned(15 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(14 downto 0);
signal s21_4 : unsigned(14 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(1 downto 0);
signal s23_4 : unsigned(1 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_16 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(1 downto 0);
i9 : in  unsigned(1 downto 0);
i10 : in  unsigned(1 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(1 downto 0);
o4 : out unsigned(1 downto 0));
end component cf_rca_16_16;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s20_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s20_1(15 downto 15) &
  s20_1(14 downto 14) &
  s20_1(13 downto 13) &
  s20_1(12 downto 12) &
  s20_1(11 downto 11) &
  s20_1(10 downto 10) &
  s20_1(9 downto 9) &
  s20_1(8 downto 8) &
  s20_1(7 downto 7) &
  s20_1(6 downto 6) &
  s20_1(5 downto 5) &
  s20_1(4 downto 4) &
  s20_1(3 downto 3) &
  s20_1(2 downto 2) &
  s20_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s21_3 & s22_1;
n11 <= s21_4 & s22_2;
n12 <= i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s22_3;
n18 <= s23_4 & s21_2;
s19 : cf_rca_16_38 port map (s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16);
s20 : cf_rca_16_32 port map (n2, s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16, n3, s20_1);
s21 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s22_4, n8, n9, n16, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s21_1, n15, s22_1, s22_2, s22_3, s22_4);
s23 : cf_rca_16_16 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_14 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(3 downto 0);
i9 : in  unsigned(3 downto 0);
i10 : in  unsigned(3 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(3 downto 0);
o4 : out unsigned(3 downto 0));
end entity cf_rca_16_14;
architecture rtl of cf_rca_16_14 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(2 downto 0);
signal n13 : unsigned(2 downto 0);
signal n14 : unsigned(2 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(3 downto 0);
signal n18 : unsigned(3 downto 0);
signal s19_1 : unsigned(15 downto 0);
signal s19_2 : unsigned(15 downto 0);
signal s19_3 : unsigned(15 downto 0);
signal s19_4 : unsigned(15 downto 0);
signal s19_5 : unsigned(15 downto 0);
signal s19_6 : unsigned(15 downto 0);
signal s19_7 : unsigned(15 downto 0);
signal s19_8 : unsigned(15 downto 0);
signal s19_9 : unsigned(15 downto 0);
signal s19_10 : unsigned(15 downto 0);
signal s19_11 : unsigned(15 downto 0);
signal s19_12 : unsigned(15 downto 0);
signal s19_13 : unsigned(15 downto 0);
signal s19_14 : unsigned(15 downto 0);
signal s19_15 : unsigned(15 downto 0);
signal s19_16 : unsigned(15 downto 0);
signal s20_1 : unsigned(15 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(14 downto 0);
signal s21_4 : unsigned(14 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(2 downto 0);
signal s23_4 : unsigned(2 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_15 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(2 downto 0);
i9 : in  unsigned(2 downto 0);
i10 : in  unsigned(2 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(2 downto 0);
o4 : out unsigned(2 downto 0));
end component cf_rca_16_15;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s20_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s20_1(15 downto 15) &
  s20_1(14 downto 14) &
  s20_1(13 downto 13) &
  s20_1(12 downto 12) &
  s20_1(11 downto 11) &
  s20_1(10 downto 10) &
  s20_1(9 downto 9) &
  s20_1(8 downto 8) &
  s20_1(7 downto 7) &
  s20_1(6 downto 6) &
  s20_1(5 downto 5) &
  s20_1(4 downto 4) &
  s20_1(3 downto 3) &
  s20_1(2 downto 2) &
  s20_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s21_3 & s22_1;
n11 <= s21_4 & s22_2;
n12 <= i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s22_3;
n18 <= s23_4 & s21_2;
s19 : cf_rca_16_38 port map (s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16);
s20 : cf_rca_16_32 port map (n2, s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16, n3, s20_1);
s21 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s22_4, n8, n9, n16, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s21_1, n15, s22_1, s22_2, s22_3, s22_4);
s23 : cf_rca_16_15 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_13 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(4 downto 0);
i9 : in  unsigned(4 downto 0);
i10 : in  unsigned(4 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(4 downto 0);
o4 : out unsigned(4 downto 0));
end entity cf_rca_16_13;
architecture rtl of cf_rca_16_13 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(3 downto 0);
signal n13 : unsigned(3 downto 0);
signal n14 : unsigned(3 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(4 downto 0);
signal n18 : unsigned(4 downto 0);
signal s19_1 : unsigned(15 downto 0);
signal s19_2 : unsigned(15 downto 0);
signal s19_3 : unsigned(15 downto 0);
signal s19_4 : unsigned(15 downto 0);
signal s19_5 : unsigned(15 downto 0);
signal s19_6 : unsigned(15 downto 0);
signal s19_7 : unsigned(15 downto 0);
signal s19_8 : unsigned(15 downto 0);
signal s19_9 : unsigned(15 downto 0);
signal s19_10 : unsigned(15 downto 0);
signal s19_11 : unsigned(15 downto 0);
signal s19_12 : unsigned(15 downto 0);
signal s19_13 : unsigned(15 downto 0);
signal s19_14 : unsigned(15 downto 0);
signal s19_15 : unsigned(15 downto 0);
signal s19_16 : unsigned(15 downto 0);
signal s20_1 : unsigned(15 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(14 downto 0);
signal s21_4 : unsigned(14 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(3 downto 0);
signal s23_4 : unsigned(3 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_14 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(3 downto 0);
i9 : in  unsigned(3 downto 0);
i10 : in  unsigned(3 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(3 downto 0);
o4 : out unsigned(3 downto 0));
end component cf_rca_16_14;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s20_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s20_1(15 downto 15) &
  s20_1(14 downto 14) &
  s20_1(13 downto 13) &
  s20_1(12 downto 12) &
  s20_1(11 downto 11) &
  s20_1(10 downto 10) &
  s20_1(9 downto 9) &
  s20_1(8 downto 8) &
  s20_1(7 downto 7) &
  s20_1(6 downto 6) &
  s20_1(5 downto 5) &
  s20_1(4 downto 4) &
  s20_1(3 downto 3) &
  s20_1(2 downto 2) &
  s20_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s21_3 & s22_1;
n11 <= s21_4 & s22_2;
n12 <= i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(4 downto 4) &
  i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s22_3;
n18 <= s23_4 & s21_2;
s19 : cf_rca_16_38 port map (s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16);
s20 : cf_rca_16_32 port map (n2, s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16, n3, s20_1);
s21 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s22_4, n8, n9, n16, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s21_1, n15, s22_1, s22_2, s22_3, s22_4);
s23 : cf_rca_16_14 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_12 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(5 downto 0);
i9 : in  unsigned(5 downto 0);
i10 : in  unsigned(5 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(5 downto 0);
o4 : out unsigned(5 downto 0));
end entity cf_rca_16_12;
architecture rtl of cf_rca_16_12 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(4 downto 0);
signal n13 : unsigned(4 downto 0);
signal n14 : unsigned(4 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(5 downto 0);
signal n18 : unsigned(5 downto 0);
signal s19_1 : unsigned(15 downto 0);
signal s19_2 : unsigned(15 downto 0);
signal s19_3 : unsigned(15 downto 0);
signal s19_4 : unsigned(15 downto 0);
signal s19_5 : unsigned(15 downto 0);
signal s19_6 : unsigned(15 downto 0);
signal s19_7 : unsigned(15 downto 0);
signal s19_8 : unsigned(15 downto 0);
signal s19_9 : unsigned(15 downto 0);
signal s19_10 : unsigned(15 downto 0);
signal s19_11 : unsigned(15 downto 0);
signal s19_12 : unsigned(15 downto 0);
signal s19_13 : unsigned(15 downto 0);
signal s19_14 : unsigned(15 downto 0);
signal s19_15 : unsigned(15 downto 0);
signal s19_16 : unsigned(15 downto 0);
signal s20_1 : unsigned(15 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(14 downto 0);
signal s21_4 : unsigned(14 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(4 downto 0);
signal s23_4 : unsigned(4 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_13 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(4 downto 0);
i9 : in  unsigned(4 downto 0);
i10 : in  unsigned(4 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(4 downto 0);
o4 : out unsigned(4 downto 0));
end component cf_rca_16_13;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s20_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s20_1(15 downto 15) &
  s20_1(14 downto 14) &
  s20_1(13 downto 13) &
  s20_1(12 downto 12) &
  s20_1(11 downto 11) &
  s20_1(10 downto 10) &
  s20_1(9 downto 9) &
  s20_1(8 downto 8) &
  s20_1(7 downto 7) &
  s20_1(6 downto 6) &
  s20_1(5 downto 5) &
  s20_1(4 downto 4) &
  s20_1(3 downto 3) &
  s20_1(2 downto 2) &
  s20_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s21_3 & s22_1;
n11 <= s21_4 & s22_2;
n12 <= i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(5 downto 5) &
  i10(4 downto 4) &
  i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s22_3;
n18 <= s23_4 & s21_2;
s19 : cf_rca_16_38 port map (s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16);
s20 : cf_rca_16_32 port map (n2, s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16, n3, s20_1);
s21 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s22_4, n8, n9, n16, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s21_1, n15, s22_1, s22_2, s22_3, s22_4);
s23 : cf_rca_16_13 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_11 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(6 downto 0);
i9 : in  unsigned(6 downto 0);
i10 : in  unsigned(6 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(6 downto 0);
o4 : out unsigned(6 downto 0));
end entity cf_rca_16_11;
architecture rtl of cf_rca_16_11 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(5 downto 0);
signal n13 : unsigned(5 downto 0);
signal n14 : unsigned(5 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(6 downto 0);
signal n18 : unsigned(6 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(0 downto 0);
signal s19_4 : unsigned(0 downto 0);
signal s20_1 : unsigned(0 downto 0);
signal s20_2 : unsigned(0 downto 0);
signal s20_3 : unsigned(14 downto 0);
signal s20_4 : unsigned(14 downto 0);
signal s21_1 : unsigned(15 downto 0);
signal s21_2 : unsigned(15 downto 0);
signal s21_3 : unsigned(15 downto 0);
signal s21_4 : unsigned(15 downto 0);
signal s21_5 : unsigned(15 downto 0);
signal s21_6 : unsigned(15 downto 0);
signal s21_7 : unsigned(15 downto 0);
signal s21_8 : unsigned(15 downto 0);
signal s21_9 : unsigned(15 downto 0);
signal s21_10 : unsigned(15 downto 0);
signal s21_11 : unsigned(15 downto 0);
signal s21_12 : unsigned(15 downto 0);
signal s21_13 : unsigned(15 downto 0);
signal s21_14 : unsigned(15 downto 0);
signal s21_15 : unsigned(15 downto 0);
signal s21_16 : unsigned(15 downto 0);
signal s22_1 : unsigned(15 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(5 downto 0);
signal s23_4 : unsigned(5 downto 0);
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_18 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_18;
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_12 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(5 downto 0);
i9 : in  unsigned(5 downto 0);
i10 : in  unsigned(5 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(5 downto 0);
o4 : out unsigned(5 downto 0));
end component cf_rca_16_12;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s22_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s22_1(15 downto 15) &
  s22_1(14 downto 14) &
  s22_1(13 downto 13) &
  s22_1(12 downto 12) &
  s22_1(11 downto 11) &
  s22_1(10 downto 10) &
  s22_1(9 downto 9) &
  s22_1(8 downto 8) &
  s22_1(7 downto 7) &
  s22_1(6 downto 6) &
  s22_1(5 downto 5) &
  s22_1(4 downto 4) &
  s22_1(3 downto 3) &
  s22_1(2 downto 2) &
  s22_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s20_3 & s19_1;
n11 <= s20_4 & s19_2;
n12 <= i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(6 downto 6) &
  i10(5 downto 5) &
  i10(4 downto 4) &
  i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s19_3;
n18 <= s23_4 & s20_2;
s19 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s20_1, n15, s19_1, s19_2, s19_3, s19_4);
s20 : cf_rca_16_18 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s19_4, n8, n9, n16, s20_1, s20_2, s20_3, s20_4);
s21 : cf_rca_16_38 port map (s21_1, s21_2, s21_3, s21_4, s21_5, s21_6, s21_7, s21_8, s21_9, s21_10, s21_11, s21_12, s21_13, s21_14, s21_15, s21_16);
s22 : cf_rca_16_32 port map (n2, s21_1, s21_2, s21_3, s21_4, s21_5, s21_6, s21_7, s21_8, s21_9, s21_10, s21_11, s21_12, s21_13, s21_14, s21_15, s21_16, n3, s22_1);
s23 : cf_rca_16_12 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_10 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(7 downto 0);
i9 : in  unsigned(7 downto 0);
i10 : in  unsigned(7 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(7 downto 0);
o4 : out unsigned(7 downto 0));
end entity cf_rca_16_10;
architecture rtl of cf_rca_16_10 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(6 downto 0);
signal n13 : unsigned(6 downto 0);
signal n14 : unsigned(6 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(7 downto 0);
signal n18 : unsigned(7 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(14 downto 0);
signal s19_4 : unsigned(14 downto 0);
signal s20_1 : unsigned(0 downto 0);
signal s20_2 : unsigned(0 downto 0);
signal s20_3 : unsigned(0 downto 0);
signal s20_4 : unsigned(0 downto 0);
signal s21_1 : unsigned(15 downto 0);
signal s21_2 : unsigned(15 downto 0);
signal s21_3 : unsigned(15 downto 0);
signal s21_4 : unsigned(15 downto 0);
signal s21_5 : unsigned(15 downto 0);
signal s21_6 : unsigned(15 downto 0);
signal s21_7 : unsigned(15 downto 0);
signal s21_8 : unsigned(15 downto 0);
signal s21_9 : unsigned(15 downto 0);
signal s21_10 : unsigned(15 downto 0);
signal s21_11 : unsigned(15 downto 0);
signal s21_12 : unsigned(15 downto 0);
signal s21_13 : unsigned(15 downto 0);
signal s21_14 : unsigned(15 downto 0);
signal s21_15 : unsigned(15 downto 0);
signal s21_16 : unsigned(15 downto 0);
signal s22_1 : unsigned(15 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(6 downto 0);
signal s23_4 : unsigned(6 downto 0);
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_11 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(6 downto 0);
i9 : in  unsigned(6 downto 0);
i10 : in  unsigned(6 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(6 downto 0);
o4 : out unsigned(6 downto 0));
end component cf_rca_16_11;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s22_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s22_1(15 downto 15) &
  s22_1(14 downto 14) &
  s22_1(13 downto 13) &
  s22_1(12 downto 12) &
  s22_1(11 downto 11) &
  s22_1(10 downto 10) &
  s22_1(9 downto 9) &
  s22_1(8 downto 8) &
  s22_1(7 downto 7) &
  s22_1(6 downto 6) &
  s22_1(5 downto 5) &
  s22_1(4 downto 4) &
  s22_1(3 downto 3) &
  s22_1(2 downto 2) &
  s22_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s19_3 & s20_1;
n11 <= s19_4 & s20_2;
n12 <= i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(7 downto 7) &
  i10(6 downto 6) &
  i10(5 downto 5) &
  i10(4 downto 4) &
  i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s20_3;
n18 <= s23_4 & s19_2;
s19 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s20_4, n8, n9, n16, s19_1, s19_2, s19_3, s19_4);
s20 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s19_1, n15, s20_1, s20_2, s20_3, s20_4);
s21 : cf_rca_16_38 port map (s21_1, s21_2, s21_3, s21_4, s21_5, s21_6, s21_7, s21_8, s21_9, s21_10, s21_11, s21_12, s21_13, s21_14, s21_15, s21_16);
s22 : cf_rca_16_32 port map (n2, s21_1, s21_2, s21_3, s21_4, s21_5, s21_6, s21_7, s21_8, s21_9, s21_10, s21_11, s21_12, s21_13, s21_14, s21_15, s21_16, n3, s22_1);
s23 : cf_rca_16_11 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_9 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(8 downto 0);
i9 : in  unsigned(8 downto 0);
i10 : in  unsigned(8 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(8 downto 0);
o4 : out unsigned(8 downto 0));
end entity cf_rca_16_9;
architecture rtl of cf_rca_16_9 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(7 downto 0);
signal n13 : unsigned(7 downto 0);
signal n14 : unsigned(7 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(8 downto 0);
signal n18 : unsigned(8 downto 0);
signal s19_1 : unsigned(0 downto 0);
signal s19_2 : unsigned(0 downto 0);
signal s19_3 : unsigned(14 downto 0);
signal s19_4 : unsigned(14 downto 0);
signal s20_1 : unsigned(0 downto 0);
signal s20_2 : unsigned(0 downto 0);
signal s20_3 : unsigned(0 downto 0);
signal s20_4 : unsigned(0 downto 0);
signal s21_1 : unsigned(15 downto 0);
signal s21_2 : unsigned(15 downto 0);
signal s21_3 : unsigned(15 downto 0);
signal s21_4 : unsigned(15 downto 0);
signal s21_5 : unsigned(15 downto 0);
signal s21_6 : unsigned(15 downto 0);
signal s21_7 : unsigned(15 downto 0);
signal s21_8 : unsigned(15 downto 0);
signal s21_9 : unsigned(15 downto 0);
signal s21_10 : unsigned(15 downto 0);
signal s21_11 : unsigned(15 downto 0);
signal s21_12 : unsigned(15 downto 0);
signal s21_13 : unsigned(15 downto 0);
signal s21_14 : unsigned(15 downto 0);
signal s21_15 : unsigned(15 downto 0);
signal s21_16 : unsigned(15 downto 0);
signal s22_1 : unsigned(15 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(7 downto 0);
signal s23_4 : unsigned(7 downto 0);
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_10 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(7 downto 0);
i9 : in  unsigned(7 downto 0);
i10 : in  unsigned(7 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(7 downto 0);
o4 : out unsigned(7 downto 0));
end component cf_rca_16_10;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s22_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s22_1(15 downto 15) &
  s22_1(14 downto 14) &
  s22_1(13 downto 13) &
  s22_1(12 downto 12) &
  s22_1(11 downto 11) &
  s22_1(10 downto 10) &
  s22_1(9 downto 9) &
  s22_1(8 downto 8) &
  s22_1(7 downto 7) &
  s22_1(6 downto 6) &
  s22_1(5 downto 5) &
  s22_1(4 downto 4) &
  s22_1(3 downto 3) &
  s22_1(2 downto 2) &
  s22_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s19_3 & s20_1;
n11 <= s19_4 & s20_2;
n12 <= i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(8 downto 8) &
  i10(7 downto 7) &
  i10(6 downto 6) &
  i10(5 downto 5) &
  i10(4 downto 4) &
  i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s20_3;
n18 <= s23_4 & s19_2;
s19 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s20_4, n8, n9, n16, s19_1, s19_2, s19_3, s19_4);
s20 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s19_1, n15, s20_1, s20_2, s20_3, s20_4);
s21 : cf_rca_16_38 port map (s21_1, s21_2, s21_3, s21_4, s21_5, s21_6, s21_7, s21_8, s21_9, s21_10, s21_11, s21_12, s21_13, s21_14, s21_15, s21_16);
s22 : cf_rca_16_32 port map (n2, s21_1, s21_2, s21_3, s21_4, s21_5, s21_6, s21_7, s21_8, s21_9, s21_10, s21_11, s21_12, s21_13, s21_14, s21_15, s21_16, n3, s22_1);
s23 : cf_rca_16_10 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_8 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(9 downto 0);
i9 : in  unsigned(9 downto 0);
i10 : in  unsigned(9 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(9 downto 0);
o4 : out unsigned(9 downto 0));
end entity cf_rca_16_8;
architecture rtl of cf_rca_16_8 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(8 downto 0);
signal n13 : unsigned(8 downto 0);
signal n14 : unsigned(8 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(9 downto 0);
signal n18 : unsigned(9 downto 0);
signal s19_1 : unsigned(15 downto 0);
signal s19_2 : unsigned(15 downto 0);
signal s19_3 : unsigned(15 downto 0);
signal s19_4 : unsigned(15 downto 0);
signal s19_5 : unsigned(15 downto 0);
signal s19_6 : unsigned(15 downto 0);
signal s19_7 : unsigned(15 downto 0);
signal s19_8 : unsigned(15 downto 0);
signal s19_9 : unsigned(15 downto 0);
signal s19_10 : unsigned(15 downto 0);
signal s19_11 : unsigned(15 downto 0);
signal s19_12 : unsigned(15 downto 0);
signal s19_13 : unsigned(15 downto 0);
signal s19_14 : unsigned(15 downto 0);
signal s19_15 : unsigned(15 downto 0);
signal s19_16 : unsigned(15 downto 0);
signal s20_1 : unsigned(15 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(14 downto 0);
signal s21_4 : unsigned(14 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(8 downto 0);
signal s23_4 : unsigned(8 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_9 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(8 downto 0);
i9 : in  unsigned(8 downto 0);
i10 : in  unsigned(8 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(8 downto 0);
o4 : out unsigned(8 downto 0));
end component cf_rca_16_9;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s20_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s20_1(15 downto 15) &
  s20_1(14 downto 14) &
  s20_1(13 downto 13) &
  s20_1(12 downto 12) &
  s20_1(11 downto 11) &
  s20_1(10 downto 10) &
  s20_1(9 downto 9) &
  s20_1(8 downto 8) &
  s20_1(7 downto 7) &
  s20_1(6 downto 6) &
  s20_1(5 downto 5) &
  s20_1(4 downto 4) &
  s20_1(3 downto 3) &
  s20_1(2 downto 2) &
  s20_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s21_3 & s22_1;
n11 <= s21_4 & s22_2;
n12 <= i8(9 downto 9) &
  i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(9 downto 9) &
  i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(9 downto 9) &
  i10(8 downto 8) &
  i10(7 downto 7) &
  i10(6 downto 6) &
  i10(5 downto 5) &
  i10(4 downto 4) &
  i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s22_3;
n18 <= s23_4 & s21_2;
s19 : cf_rca_16_38 port map (s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16);
s20 : cf_rca_16_32 port map (n2, s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16, n3, s20_1);
s21 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s22_4, n8, n9, n16, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s21_1, n15, s22_1, s22_2, s22_3, s22_4);
s23 : cf_rca_16_9 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_7 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(10 downto 0);
i9 : in  unsigned(10 downto 0);
i10 : in  unsigned(10 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(10 downto 0);
o4 : out unsigned(10 downto 0));
end entity cf_rca_16_7;
architecture rtl of cf_rca_16_7 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(9 downto 0);
signal n13 : unsigned(9 downto 0);
signal n14 : unsigned(9 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(10 downto 0);
signal n18 : unsigned(10 downto 0);
signal s19_1 : unsigned(15 downto 0);
signal s19_2 : unsigned(15 downto 0);
signal s19_3 : unsigned(15 downto 0);
signal s19_4 : unsigned(15 downto 0);
signal s19_5 : unsigned(15 downto 0);
signal s19_6 : unsigned(15 downto 0);
signal s19_7 : unsigned(15 downto 0);
signal s19_8 : unsigned(15 downto 0);
signal s19_9 : unsigned(15 downto 0);
signal s19_10 : unsigned(15 downto 0);
signal s19_11 : unsigned(15 downto 0);
signal s19_12 : unsigned(15 downto 0);
signal s19_13 : unsigned(15 downto 0);
signal s19_14 : unsigned(15 downto 0);
signal s19_15 : unsigned(15 downto 0);
signal s19_16 : unsigned(15 downto 0);
signal s20_1 : unsigned(15 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(14 downto 0);
signal s21_4 : unsigned(14 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(9 downto 0);
signal s23_4 : unsigned(9 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_8 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(9 downto 0);
i9 : in  unsigned(9 downto 0);
i10 : in  unsigned(9 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(9 downto 0);
o4 : out unsigned(9 downto 0));
end component cf_rca_16_8;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s20_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s20_1(15 downto 15) &
  s20_1(14 downto 14) &
  s20_1(13 downto 13) &
  s20_1(12 downto 12) &
  s20_1(11 downto 11) &
  s20_1(10 downto 10) &
  s20_1(9 downto 9) &
  s20_1(8 downto 8) &
  s20_1(7 downto 7) &
  s20_1(6 downto 6) &
  s20_1(5 downto 5) &
  s20_1(4 downto 4) &
  s20_1(3 downto 3) &
  s20_1(2 downto 2) &
  s20_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s21_3 & s22_1;
n11 <= s21_4 & s22_2;
n12 <= i8(10 downto 10) &
  i8(9 downto 9) &
  i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(10 downto 10) &
  i9(9 downto 9) &
  i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(10 downto 10) &
  i10(9 downto 9) &
  i10(8 downto 8) &
  i10(7 downto 7) &
  i10(6 downto 6) &
  i10(5 downto 5) &
  i10(4 downto 4) &
  i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s22_3;
n18 <= s23_4 & s21_2;
s19 : cf_rca_16_38 port map (s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16);
s20 : cf_rca_16_32 port map (n2, s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16, n3, s20_1);
s21 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s22_4, n8, n9, n16, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s21_1, n15, s22_1, s22_2, s22_3, s22_4);
s23 : cf_rca_16_8 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_6 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(11 downto 0);
i9 : in  unsigned(11 downto 0);
i10 : in  unsigned(11 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(11 downto 0);
o4 : out unsigned(11 downto 0));
end entity cf_rca_16_6;
architecture rtl of cf_rca_16_6 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(10 downto 0);
signal n13 : unsigned(10 downto 0);
signal n14 : unsigned(10 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(11 downto 0);
signal n18 : unsigned(11 downto 0);
signal s19_1 : unsigned(15 downto 0);
signal s19_2 : unsigned(15 downto 0);
signal s19_3 : unsigned(15 downto 0);
signal s19_4 : unsigned(15 downto 0);
signal s19_5 : unsigned(15 downto 0);
signal s19_6 : unsigned(15 downto 0);
signal s19_7 : unsigned(15 downto 0);
signal s19_8 : unsigned(15 downto 0);
signal s19_9 : unsigned(15 downto 0);
signal s19_10 : unsigned(15 downto 0);
signal s19_11 : unsigned(15 downto 0);
signal s19_12 : unsigned(15 downto 0);
signal s19_13 : unsigned(15 downto 0);
signal s19_14 : unsigned(15 downto 0);
signal s19_15 : unsigned(15 downto 0);
signal s19_16 : unsigned(15 downto 0);
signal s20_1 : unsigned(15 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(14 downto 0);
signal s21_4 : unsigned(14 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(10 downto 0);
signal s23_4 : unsigned(10 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_7 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(10 downto 0);
i9 : in  unsigned(10 downto 0);
i10 : in  unsigned(10 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(10 downto 0);
o4 : out unsigned(10 downto 0));
end component cf_rca_16_7;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s20_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s20_1(15 downto 15) &
  s20_1(14 downto 14) &
  s20_1(13 downto 13) &
  s20_1(12 downto 12) &
  s20_1(11 downto 11) &
  s20_1(10 downto 10) &
  s20_1(9 downto 9) &
  s20_1(8 downto 8) &
  s20_1(7 downto 7) &
  s20_1(6 downto 6) &
  s20_1(5 downto 5) &
  s20_1(4 downto 4) &
  s20_1(3 downto 3) &
  s20_1(2 downto 2) &
  s20_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s21_3 & s22_1;
n11 <= s21_4 & s22_2;
n12 <= i8(11 downto 11) &
  i8(10 downto 10) &
  i8(9 downto 9) &
  i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(11 downto 11) &
  i9(10 downto 10) &
  i9(9 downto 9) &
  i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(11 downto 11) &
  i10(10 downto 10) &
  i10(9 downto 9) &
  i10(8 downto 8) &
  i10(7 downto 7) &
  i10(6 downto 6) &
  i10(5 downto 5) &
  i10(4 downto 4) &
  i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s22_3;
n18 <= s23_4 & s21_2;
s19 : cf_rca_16_38 port map (s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16);
s20 : cf_rca_16_32 port map (n2, s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16, n3, s20_1);
s21 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s22_4, n8, n9, n16, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s21_1, n15, s22_1, s22_2, s22_3, s22_4);
s23 : cf_rca_16_7 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_5 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(12 downto 0);
i9 : in  unsigned(12 downto 0);
i10 : in  unsigned(12 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(12 downto 0);
o4 : out unsigned(12 downto 0));
end entity cf_rca_16_5;
architecture rtl of cf_rca_16_5 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(11 downto 0);
signal n13 : unsigned(11 downto 0);
signal n14 : unsigned(11 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(12 downto 0);
signal n18 : unsigned(12 downto 0);
signal s19_1 : unsigned(15 downto 0);
signal s19_2 : unsigned(15 downto 0);
signal s19_3 : unsigned(15 downto 0);
signal s19_4 : unsigned(15 downto 0);
signal s19_5 : unsigned(15 downto 0);
signal s19_6 : unsigned(15 downto 0);
signal s19_7 : unsigned(15 downto 0);
signal s19_8 : unsigned(15 downto 0);
signal s19_9 : unsigned(15 downto 0);
signal s19_10 : unsigned(15 downto 0);
signal s19_11 : unsigned(15 downto 0);
signal s19_12 : unsigned(15 downto 0);
signal s19_13 : unsigned(15 downto 0);
signal s19_14 : unsigned(15 downto 0);
signal s19_15 : unsigned(15 downto 0);
signal s19_16 : unsigned(15 downto 0);
signal s20_1 : unsigned(15 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(14 downto 0);
signal s21_4 : unsigned(14 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(11 downto 0);
signal s23_4 : unsigned(11 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_6 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(11 downto 0);
i9 : in  unsigned(11 downto 0);
i10 : in  unsigned(11 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(11 downto 0);
o4 : out unsigned(11 downto 0));
end component cf_rca_16_6;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s20_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s20_1(15 downto 15) &
  s20_1(14 downto 14) &
  s20_1(13 downto 13) &
  s20_1(12 downto 12) &
  s20_1(11 downto 11) &
  s20_1(10 downto 10) &
  s20_1(9 downto 9) &
  s20_1(8 downto 8) &
  s20_1(7 downto 7) &
  s20_1(6 downto 6) &
  s20_1(5 downto 5) &
  s20_1(4 downto 4) &
  s20_1(3 downto 3) &
  s20_1(2 downto 2) &
  s20_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s21_3 & s22_1;
n11 <= s21_4 & s22_2;
n12 <= i8(12 downto 12) &
  i8(11 downto 11) &
  i8(10 downto 10) &
  i8(9 downto 9) &
  i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(12 downto 12) &
  i9(11 downto 11) &
  i9(10 downto 10) &
  i9(9 downto 9) &
  i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(12 downto 12) &
  i10(11 downto 11) &
  i10(10 downto 10) &
  i10(9 downto 9) &
  i10(8 downto 8) &
  i10(7 downto 7) &
  i10(6 downto 6) &
  i10(5 downto 5) &
  i10(4 downto 4) &
  i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s22_3;
n18 <= s23_4 & s21_2;
s19 : cf_rca_16_38 port map (s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16);
s20 : cf_rca_16_32 port map (n2, s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16, n3, s20_1);
s21 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s22_4, n8, n9, n16, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s21_1, n15, s22_1, s22_2, s22_3, s22_4);
s23 : cf_rca_16_6 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_4 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(13 downto 0);
i9 : in  unsigned(13 downto 0);
i10 : in  unsigned(13 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(13 downto 0);
o4 : out unsigned(13 downto 0));
end entity cf_rca_16_4;
architecture rtl of cf_rca_16_4 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(12 downto 0);
signal n13 : unsigned(12 downto 0);
signal n14 : unsigned(12 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(13 downto 0);
signal n18 : unsigned(13 downto 0);
signal s19_1 : unsigned(15 downto 0);
signal s19_2 : unsigned(15 downto 0);
signal s19_3 : unsigned(15 downto 0);
signal s19_4 : unsigned(15 downto 0);
signal s19_5 : unsigned(15 downto 0);
signal s19_6 : unsigned(15 downto 0);
signal s19_7 : unsigned(15 downto 0);
signal s19_8 : unsigned(15 downto 0);
signal s19_9 : unsigned(15 downto 0);
signal s19_10 : unsigned(15 downto 0);
signal s19_11 : unsigned(15 downto 0);
signal s19_12 : unsigned(15 downto 0);
signal s19_13 : unsigned(15 downto 0);
signal s19_14 : unsigned(15 downto 0);
signal s19_15 : unsigned(15 downto 0);
signal s19_16 : unsigned(15 downto 0);
signal s20_1 : unsigned(15 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(14 downto 0);
signal s21_4 : unsigned(14 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(12 downto 0);
signal s23_4 : unsigned(12 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_5 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(12 downto 0);
i9 : in  unsigned(12 downto 0);
i10 : in  unsigned(12 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(12 downto 0);
o4 : out unsigned(12 downto 0));
end component cf_rca_16_5;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s20_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s20_1(15 downto 15) &
  s20_1(14 downto 14) &
  s20_1(13 downto 13) &
  s20_1(12 downto 12) &
  s20_1(11 downto 11) &
  s20_1(10 downto 10) &
  s20_1(9 downto 9) &
  s20_1(8 downto 8) &
  s20_1(7 downto 7) &
  s20_1(6 downto 6) &
  s20_1(5 downto 5) &
  s20_1(4 downto 4) &
  s20_1(3 downto 3) &
  s20_1(2 downto 2) &
  s20_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s21_3 & s22_1;
n11 <= s21_4 & s22_2;
n12 <= i8(13 downto 13) &
  i8(12 downto 12) &
  i8(11 downto 11) &
  i8(10 downto 10) &
  i8(9 downto 9) &
  i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(13 downto 13) &
  i9(12 downto 12) &
  i9(11 downto 11) &
  i9(10 downto 10) &
  i9(9 downto 9) &
  i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(13 downto 13) &
  i10(12 downto 12) &
  i10(11 downto 11) &
  i10(10 downto 10) &
  i10(9 downto 9) &
  i10(8 downto 8) &
  i10(7 downto 7) &
  i10(6 downto 6) &
  i10(5 downto 5) &
  i10(4 downto 4) &
  i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s22_3;
n18 <= s23_4 & s21_2;
s19 : cf_rca_16_38 port map (s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16);
s20 : cf_rca_16_32 port map (n2, s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16, n3, s20_1);
s21 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s22_4, n8, n9, n16, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s21_1, n15, s22_1, s22_2, s22_3, s22_4);
s23 : cf_rca_16_5 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_3 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
i10 : in  unsigned(14 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end entity cf_rca_16_3;
architecture rtl of cf_rca_16_3 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(13 downto 0);
signal n13 : unsigned(13 downto 0);
signal n14 : unsigned(13 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(14 downto 0);
signal n18 : unsigned(14 downto 0);
signal s19_1 : unsigned(15 downto 0);
signal s19_2 : unsigned(15 downto 0);
signal s19_3 : unsigned(15 downto 0);
signal s19_4 : unsigned(15 downto 0);
signal s19_5 : unsigned(15 downto 0);
signal s19_6 : unsigned(15 downto 0);
signal s19_7 : unsigned(15 downto 0);
signal s19_8 : unsigned(15 downto 0);
signal s19_9 : unsigned(15 downto 0);
signal s19_10 : unsigned(15 downto 0);
signal s19_11 : unsigned(15 downto 0);
signal s19_12 : unsigned(15 downto 0);
signal s19_13 : unsigned(15 downto 0);
signal s19_14 : unsigned(15 downto 0);
signal s19_15 : unsigned(15 downto 0);
signal s19_16 : unsigned(15 downto 0);
signal s20_1 : unsigned(15 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(14 downto 0);
signal s21_4 : unsigned(14 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(13 downto 0);
signal s23_4 : unsigned(13 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_4 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(13 downto 0);
i9 : in  unsigned(13 downto 0);
i10 : in  unsigned(13 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(13 downto 0);
o4 : out unsigned(13 downto 0));
end component cf_rca_16_4;
begin
n1 <= i8(0 downto 0);
n2 <= n1 & i5;
n3 <= "0000000000000000";
n4 <= i9(0 downto 0);
n5 <= i10(0 downto 0);
n6 <= s20_1(0 downto 0);
n7 <= i7(0 downto 0);
n8 <= s20_1(15 downto 15) &
  s20_1(14 downto 14) &
  s20_1(13 downto 13) &
  s20_1(12 downto 12) &
  s20_1(11 downto 11) &
  s20_1(10 downto 10) &
  s20_1(9 downto 9) &
  s20_1(8 downto 8) &
  s20_1(7 downto 7) &
  s20_1(6 downto 6) &
  s20_1(5 downto 5) &
  s20_1(4 downto 4) &
  s20_1(3 downto 3) &
  s20_1(2 downto 2) &
  s20_1(1 downto 1);
n9 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n10 <= s21_3 & s22_1;
n11 <= s21_4 & s22_2;
n12 <= i8(14 downto 14) &
  i8(13 downto 13) &
  i8(12 downto 12) &
  i8(11 downto 11) &
  i8(10 downto 10) &
  i8(9 downto 9) &
  i8(8 downto 8) &
  i8(7 downto 7) &
  i8(6 downto 6) &
  i8(5 downto 5) &
  i8(4 downto 4) &
  i8(3 downto 3) &
  i8(2 downto 2) &
  i8(1 downto 1);
n13 <= i9(14 downto 14) &
  i9(13 downto 13) &
  i9(12 downto 12) &
  i9(11 downto 11) &
  i9(10 downto 10) &
  i9(9 downto 9) &
  i9(8 downto 8) &
  i9(7 downto 7) &
  i9(6 downto 6) &
  i9(5 downto 5) &
  i9(4 downto 4) &
  i9(3 downto 3) &
  i9(2 downto 2) &
  i9(1 downto 1);
n14 <= i10(14 downto 14) &
  i10(13 downto 13) &
  i10(12 downto 12) &
  i10(11 downto 11) &
  i10(10 downto 10) &
  i10(9 downto 9) &
  i10(8 downto 8) &
  i10(7 downto 7) &
  i10(6 downto 6) &
  i10(5 downto 5) &
  i10(4 downto 4) &
  i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s22_3;
n18 <= s23_4 & s21_2;
s19 : cf_rca_16_38 port map (s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16);
s20 : cf_rca_16_32 port map (n2, s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16, n3, s20_1);
s21 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n5, s22_4, n8, n9, n16, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i6, n4, n6, n7, s21_1, n15, s22_1, s22_2, s22_3, s22_4);
s23 : cf_rca_16_4 port map (clock_config_c, clock_main_c, i1, i2, i3, i4, i5, i6, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_2 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(3 downto 0);
i9 : in  unsigned(1 downto 0);
i10 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0));
end entity cf_rca_16_2;
architecture rtl of cf_rca_16_2 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(4 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(14 downto 0);
signal n9 : unsigned(14 downto 0);
signal n10 : unsigned(15 downto 0);
signal n11 : unsigned(15 downto 0);
signal n12 : unsigned(14 downto 0);
signal n13 : unsigned(14 downto 0);
signal n14 : unsigned(14 downto 0);
signal n15 : unsigned(0 downto 0);
signal n16 : unsigned(14 downto 0);
signal n17 : unsigned(15 downto 0);
signal n18 : unsigned(15 downto 0);
signal s19_1 : unsigned(15 downto 0);
signal s19_2 : unsigned(15 downto 0);
signal s19_3 : unsigned(15 downto 0);
signal s19_4 : unsigned(15 downto 0);
signal s19_5 : unsigned(15 downto 0);
signal s19_6 : unsigned(15 downto 0);
signal s19_7 : unsigned(15 downto 0);
signal s19_8 : unsigned(15 downto 0);
signal s19_9 : unsigned(15 downto 0);
signal s19_10 : unsigned(15 downto 0);
signal s19_11 : unsigned(15 downto 0);
signal s19_12 : unsigned(15 downto 0);
signal s19_13 : unsigned(15 downto 0);
signal s19_14 : unsigned(15 downto 0);
signal s19_15 : unsigned(15 downto 0);
signal s19_16 : unsigned(15 downto 0);
signal s20_1 : unsigned(15 downto 0);
signal s21_1 : unsigned(0 downto 0);
signal s21_2 : unsigned(0 downto 0);
signal s21_3 : unsigned(14 downto 0);
signal s21_4 : unsigned(14 downto 0);
signal s22_1 : unsigned(0 downto 0);
signal s22_2 : unsigned(0 downto 0);
signal s22_3 : unsigned(0 downto 0);
signal s22_4 : unsigned(0 downto 0);
signal s23_1 : unsigned(15 downto 0);
signal s23_2 : unsigned(15 downto 0);
signal s23_3 : unsigned(14 downto 0);
signal s23_4 : unsigned(14 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_22 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(14 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_22;
component cf_rca_16_29 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(1 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0));
end component cf_rca_16_29;
component cf_rca_16_3 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(3 downto 0);
i6 : in  unsigned(1 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(14 downto 0);
i9 : in  unsigned(14 downto 0);
i10 : in  unsigned(14 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(14 downto 0);
o4 : out unsigned(14 downto 0));
end component cf_rca_16_3;
begin
n1 <= i10(0 downto 0);
n2 <= n1 & i8;
n3 <= "0000000000000000";
n4 <= i7(0 downto 0);
n5 <= i6(0 downto 0);
n6 <= s20_1(0 downto 0);
n7 <= i4(0 downto 0);
n8 <= s20_1(15 downto 15) &
  s20_1(14 downto 14) &
  s20_1(13 downto 13) &
  s20_1(12 downto 12) &
  s20_1(11 downto 11) &
  s20_1(10 downto 10) &
  s20_1(9 downto 9) &
  s20_1(8 downto 8) &
  s20_1(7 downto 7) &
  s20_1(6 downto 6) &
  s20_1(5 downto 5) &
  s20_1(4 downto 4) &
  s20_1(3 downto 3) &
  s20_1(2 downto 2) &
  s20_1(1 downto 1);
n9 <= i4(15 downto 15) &
  i4(14 downto 14) &
  i4(13 downto 13) &
  i4(12 downto 12) &
  i4(11 downto 11) &
  i4(10 downto 10) &
  i4(9 downto 9) &
  i4(8 downto 8) &
  i4(7 downto 7) &
  i4(6 downto 6) &
  i4(5 downto 5) &
  i4(4 downto 4) &
  i4(3 downto 3) &
  i4(2 downto 2) &
  i4(1 downto 1);
n10 <= s21_3 & s22_1;
n11 <= s21_4 & s22_2;
n12 <= i10(15 downto 15) &
  i10(14 downto 14) &
  i10(13 downto 13) &
  i10(12 downto 12) &
  i10(11 downto 11) &
  i10(10 downto 10) &
  i10(9 downto 9) &
  i10(8 downto 8) &
  i10(7 downto 7) &
  i10(6 downto 6) &
  i10(5 downto 5) &
  i10(4 downto 4) &
  i10(3 downto 3) &
  i10(2 downto 2) &
  i10(1 downto 1);
n13 <= i7(15 downto 15) &
  i7(14 downto 14) &
  i7(13 downto 13) &
  i7(12 downto 12) &
  i7(11 downto 11) &
  i7(10 downto 10) &
  i7(9 downto 9) &
  i7(8 downto 8) &
  i7(7 downto 7) &
  i7(6 downto 6) &
  i7(5 downto 5) &
  i7(4 downto 4) &
  i7(3 downto 3) &
  i7(2 downto 2) &
  i7(1 downto 1);
n14 <= i6(15 downto 15) &
  i6(14 downto 14) &
  i6(13 downto 13) &
  i6(12 downto 12) &
  i6(11 downto 11) &
  i6(10 downto 10) &
  i6(9 downto 9) &
  i6(8 downto 8) &
  i6(7 downto 7) &
  i6(6 downto 6) &
  i6(5 downto 5) &
  i6(4 downto 4) &
  i6(3 downto 3) &
  i6(2 downto 2) &
  i6(1 downto 1);
n15 <= s23_1(0 downto 0);
n16 <= s23_1(15 downto 15) &
  s23_1(14 downto 14) &
  s23_1(13 downto 13) &
  s23_1(12 downto 12) &
  s23_1(11 downto 11) &
  s23_1(10 downto 10) &
  s23_1(9 downto 9) &
  s23_1(8 downto 8) &
  s23_1(7 downto 7) &
  s23_1(6 downto 6) &
  s23_1(5 downto 5) &
  s23_1(4 downto 4) &
  s23_1(3 downto 3) &
  s23_1(2 downto 2) &
  s23_1(1 downto 1);
n17 <= s23_3 & s22_3;
n18 <= s23_4 & s21_2;
s19 : cf_rca_16_38 port map (s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16);
s20 : cf_rca_16_32 port map (n2, s19_1, s19_2, s19_3, s19_4, s19_5, s19_6, s19_7, s19_8, s19_9, s19_10, s19_11, s19_12, s19_13, s19_14, s19_15, s19_16, n3, s20_1);
s21 : cf_rca_16_22 port map (clock_config_c, clock_main_c, i1, i2, i3, i9, n5, s22_4, n8, n9, n16, s21_1, s21_2, s21_3, s21_4);
s22 : cf_rca_16_29 port map (clock_config_c, clock_main_c, i1, i2, i3, i9, n4, n6, n7, s21_1, n15, s22_1, s22_2, s22_3, s22_4);
s23 : cf_rca_16_3 port map (clock_config_c, clock_main_c, i1, i2, i3, i5, i8, i9, n11, n12, n13, n14, s23_1, s23_2, s23_3, s23_4);
o4 <= n18;
o3 <= n17;
o2 <= s23_2;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16_1 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(9 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0));
end entity cf_rca_16_1;
architecture rtl of cf_rca_16_1 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(3 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(1 downto 0);
signal n6 : unsigned(4 downto 0);
signal n7 : unsigned(15 downto 0);
signal s8_1 : unsigned(15 downto 0);
signal s8_2 : unsigned(15 downto 0);
signal s8_3 : unsigned(15 downto 0);
signal s8_4 : unsigned(15 downto 0);
signal s8_5 : unsigned(15 downto 0);
signal s8_6 : unsigned(15 downto 0);
signal s8_7 : unsigned(15 downto 0);
signal s8_8 : unsigned(15 downto 0);
signal s8_9 : unsigned(15 downto 0);
signal s8_10 : unsigned(15 downto 0);
signal s8_11 : unsigned(15 downto 0);
signal s8_12 : unsigned(15 downto 0);
signal s8_13 : unsigned(15 downto 0);
signal s8_14 : unsigned(15 downto 0);
signal s8_15 : unsigned(15 downto 0);
signal s8_16 : unsigned(15 downto 0);
signal s9_1 : unsigned(15 downto 0);
signal s10_1 : unsigned(15 downto 0);
signal s10_2 : unsigned(15 downto 0);
signal s10_3 : unsigned(15 downto 0);
signal s10_4 : unsigned(15 downto 0);
component cf_rca_16_38 is
port (
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0);
o5 : out unsigned(15 downto 0);
o6 : out unsigned(15 downto 0);
o7 : out unsigned(15 downto 0);
o8 : out unsigned(15 downto 0);
o9 : out unsigned(15 downto 0);
o10 : out unsigned(15 downto 0);
o11 : out unsigned(15 downto 0);
o12 : out unsigned(15 downto 0);
o13 : out unsigned(15 downto 0);
o14 : out unsigned(15 downto 0);
o15 : out unsigned(15 downto 0);
o16 : out unsigned(15 downto 0));
end component cf_rca_16_38;
component cf_rca_16_32 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(15 downto 0);
i9 : in  unsigned(15 downto 0);
i10 : in  unsigned(15 downto 0);
i11 : in  unsigned(15 downto 0);
i12 : in  unsigned(15 downto 0);
i13 : in  unsigned(15 downto 0);
i14 : in  unsigned(15 downto 0);
i15 : in  unsigned(15 downto 0);
i16 : in  unsigned(15 downto 0);
i17 : in  unsigned(15 downto 0);
i18 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_rca_16_32;
component cf_rca_16_2 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
i8 : in  unsigned(3 downto 0);
i9 : in  unsigned(1 downto 0);
i10 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0));
end component cf_rca_16_2;
begin
n1 <= "1";
n2 <= "0";
n3 <= i2(9 downto 9) &
  i2(8 downto 8) &
  i2(7 downto 7) &
  i2(6 downto 6);
n4 <= i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2);
n5 <= i2(1 downto 1) &
  i2(0 downto 0);
n6 <= i1 & n3;
n7 <= "0000000000000000";
s8 : cf_rca_16_38 port map (s8_1, s8_2, s8_3, s8_4, s8_5, s8_6, s8_7, s8_8, s8_9, s8_10, s8_11, s8_12, s8_13, s8_14, s8_15, s8_16);
s9 : cf_rca_16_32 port map (n6, s8_1, s8_2, s8_3, s8_4, s8_5, s8_6, s8_7, s8_8, s8_9, s8_10, s8_11, s8_12, s8_13, s8_14, s8_15, s8_16, n7, s9_1);
s10 : cf_rca_16_2 port map (clock_config_c, clock_main_c, n1, n2, i3, i4, i5, i6, i7, n4, n5, s9_1, s10_1, s10_2, s10_3, s10_4);
o4 <= s10_4;
o3 <= s10_3;
o2 <= s10_2;
o1 <= s10_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_rca_16 is
port(
signal clock_config_c : in std_logic;
signal clock_main_c : in std_logic;
signal config_write_i : in unsigned(0 downto 0);
signal config_addr_i : in unsigned(9 downto 0);
signal config_data_i : in unsigned(17 downto 0);
signal north_i : in unsigned(15 downto 0);
signal south_i : in unsigned(15 downto 0);
signal west_i : in unsigned(15 downto 0);
signal east_i : in unsigned(15 downto 0);
signal north_o : out unsigned(15 downto 0);
signal south_o : out unsigned(15 downto 0);
signal west_o : out unsigned(15 downto 0);
signal east_o : out unsigned(15 downto 0));
end entity cf_rca_16;
architecture rtl of cf_rca_16 is
component cf_rca_16_1 is
port (
clock_config_c : in std_logic;
clock_main_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(9 downto 0);
i3 : in  unsigned(17 downto 0);
i4 : in  unsigned(15 downto 0);
i5 : in  unsigned(15 downto 0);
i6 : in  unsigned(15 downto 0);
i7 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0);
o3 : out unsigned(15 downto 0);
o4 : out unsigned(15 downto 0));
end component cf_rca_16_1;
signal n1 : unsigned(15 downto 0);
signal n2 : unsigned(15 downto 0);
signal n3 : unsigned(15 downto 0);
signal n4 : unsigned(15 downto 0);
begin
s1 : cf_rca_16_1 port map (clock_config_c, clock_main_c, config_write_i, config_addr_i, config_data_i, north_i, south_i, west_i, east_i, n1, n2, n3, n4);
north_o <= n1;
south_o <= n2;
west_o <= n4;
east_o <= n3;
end architecture rtl;


