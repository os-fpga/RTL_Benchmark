module design14_11_35_top #(parameter WIDTH=32,CHANNEL=11) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	reg [WIDTH-1:0] d_in10;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;
	wire [WIDTH-1:0] d_out10;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH+1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 = tmp[WIDTH-1:0];
		d_in1 = tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 = tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 = tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 = tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 = tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 = tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 = tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 = tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 = tmp[(WIDTH*10)-1:WIDTH*9];
		d_in10 = tmp[(WIDTH*11)-1:WIDTH*10];
	end

	design14_11_35 #(.WIDTH(WIDTH)) design14_11_35_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_in10(d_in10),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.d_out10(d_out10),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9^d_out10;

endmodule

module design14_11_35 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_in10, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, d_out10, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	input [WIDTH-1:0] d_in10; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 
	output [WIDTH-1:0] d_out10; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d0_29;
	wire [WIDTH-1:0] wire_d0_30;
	wire [WIDTH-1:0] wire_d0_31;
	wire [WIDTH-1:0] wire_d0_32;
	wire [WIDTH-1:0] wire_d0_33;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d1_29;
	wire [WIDTH-1:0] wire_d1_30;
	wire [WIDTH-1:0] wire_d1_31;
	wire [WIDTH-1:0] wire_d1_32;
	wire [WIDTH-1:0] wire_d1_33;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d2_29;
	wire [WIDTH-1:0] wire_d2_30;
	wire [WIDTH-1:0] wire_d2_31;
	wire [WIDTH-1:0] wire_d2_32;
	wire [WIDTH-1:0] wire_d2_33;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d3_29;
	wire [WIDTH-1:0] wire_d3_30;
	wire [WIDTH-1:0] wire_d3_31;
	wire [WIDTH-1:0] wire_d3_32;
	wire [WIDTH-1:0] wire_d3_33;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d4_29;
	wire [WIDTH-1:0] wire_d4_30;
	wire [WIDTH-1:0] wire_d4_31;
	wire [WIDTH-1:0] wire_d4_32;
	wire [WIDTH-1:0] wire_d4_33;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d5_29;
	wire [WIDTH-1:0] wire_d5_30;
	wire [WIDTH-1:0] wire_d5_31;
	wire [WIDTH-1:0] wire_d5_32;
	wire [WIDTH-1:0] wire_d5_33;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d6_29;
	wire [WIDTH-1:0] wire_d6_30;
	wire [WIDTH-1:0] wire_d6_31;
	wire [WIDTH-1:0] wire_d6_32;
	wire [WIDTH-1:0] wire_d6_33;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d7_29;
	wire [WIDTH-1:0] wire_d7_30;
	wire [WIDTH-1:0] wire_d7_31;
	wire [WIDTH-1:0] wire_d7_32;
	wire [WIDTH-1:0] wire_d7_33;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d8_29;
	wire [WIDTH-1:0] wire_d8_30;
	wire [WIDTH-1:0] wire_d8_31;
	wire [WIDTH-1:0] wire_d8_32;
	wire [WIDTH-1:0] wire_d8_33;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d9_29;
	wire [WIDTH-1:0] wire_d9_30;
	wire [WIDTH-1:0] wire_d9_31;
	wire [WIDTH-1:0] wire_d9_32;
	wire [WIDTH-1:0] wire_d9_33;
	wire [WIDTH-1:0] wire_d10_0;
	wire [WIDTH-1:0] wire_d10_1;
	wire [WIDTH-1:0] wire_d10_2;
	wire [WIDTH-1:0] wire_d10_3;
	wire [WIDTH-1:0] wire_d10_4;
	wire [WIDTH-1:0] wire_d10_5;
	wire [WIDTH-1:0] wire_d10_6;
	wire [WIDTH-1:0] wire_d10_7;
	wire [WIDTH-1:0] wire_d10_8;
	wire [WIDTH-1:0] wire_d10_9;
	wire [WIDTH-1:0] wire_d10_10;
	wire [WIDTH-1:0] wire_d10_11;
	wire [WIDTH-1:0] wire_d10_12;
	wire [WIDTH-1:0] wire_d10_13;
	wire [WIDTH-1:0] wire_d10_14;
	wire [WIDTH-1:0] wire_d10_15;
	wire [WIDTH-1:0] wire_d10_16;
	wire [WIDTH-1:0] wire_d10_17;
	wire [WIDTH-1:0] wire_d10_18;
	wire [WIDTH-1:0] wire_d10_19;
	wire [WIDTH-1:0] wire_d10_20;
	wire [WIDTH-1:0] wire_d10_21;
	wire [WIDTH-1:0] wire_d10_22;
	wire [WIDTH-1:0] wire_d10_23;
	wire [WIDTH-1:0] wire_d10_24;
	wire [WIDTH-1:0] wire_d10_25;
	wire [WIDTH-1:0] wire_d10_26;
	wire [WIDTH-1:0] wire_d10_27;
	wire [WIDTH-1:0] wire_d10_28;
	wire [WIDTH-1:0] wire_d10_29;
	wire [WIDTH-1:0] wire_d10_30;
	wire [WIDTH-1:0] wire_d10_31;
	wire [WIDTH-1:0] wire_d10_32;
	wire [WIDTH-1:0] wire_d10_33;

	register #(.WIDTH(WIDTH)) register_instance00(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	invertion #(.WIDTH(WIDTH)) invertion_instance01(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance02(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance03(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance04(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance05(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance06(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance07(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance08(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance09(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance029(.data_in(wire_d0_28),.data_out(wire_d0_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance030(.data_in(wire_d0_29),.data_out(wire_d0_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance031(.data_in(wire_d0_30),.data_out(wire_d0_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance032(.data_in(wire_d0_31),.data_out(wire_d0_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance033(.data_in(wire_d0_32),.data_out(wire_d0_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance034(.data_in(wire_d0_33),.data_out(d_out0),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance10(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance15(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance17(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance18(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance19(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance129(.data_in(wire_d1_28),.data_out(wire_d1_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance130(.data_in(wire_d1_29),.data_out(wire_d1_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131(.data_in(wire_d1_30),.data_out(wire_d1_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance132(.data_in(wire_d1_31),.data_out(wire_d1_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance133(.data_in(wire_d1_32),.data_out(wire_d1_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance134(.data_in(wire_d1_33),.data_out(d_out1),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance20(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	invertion #(.WIDTH(WIDTH)) invertion_instance21(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance22(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance23(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance24(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance25(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance26(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance27(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance28(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance29(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance229(.data_in(wire_d2_28),.data_out(wire_d2_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance230(.data_in(wire_d2_29),.data_out(wire_d2_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance231(.data_in(wire_d2_30),.data_out(wire_d2_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232(.data_in(wire_d2_31),.data_out(wire_d2_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance233(.data_in(wire_d2_32),.data_out(wire_d2_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance234(.data_in(wire_d2_33),.data_out(d_out2),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance30(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	invertion #(.WIDTH(WIDTH)) invertion_instance31(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance32(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance33(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance34(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance35(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance36(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance37(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance38(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance39(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance329(.data_in(wire_d3_28),.data_out(wire_d3_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance330(.data_in(wire_d3_29),.data_out(wire_d3_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance331(.data_in(wire_d3_30),.data_out(wire_d3_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance332(.data_in(wire_d3_31),.data_out(wire_d3_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333(.data_in(wire_d3_32),.data_out(wire_d3_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance334(.data_in(wire_d3_33),.data_out(d_out3),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance40(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	register #(.WIDTH(WIDTH)) register_instance41(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance42(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance43(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance44(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance45(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance46(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance47(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance48(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance49(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance429(.data_in(wire_d4_28),.data_out(wire_d4_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance430(.data_in(wire_d4_29),.data_out(wire_d4_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance431(.data_in(wire_d4_30),.data_out(wire_d4_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance432(.data_in(wire_d4_31),.data_out(wire_d4_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance433(.data_in(wire_d4_32),.data_out(wire_d4_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434(.data_in(wire_d4_33),.data_out(d_out4),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance50(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	register #(.WIDTH(WIDTH)) register_instance51(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance52(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance53(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance54(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance55(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance56(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance57(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance58(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance59(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance529(.data_in(wire_d5_28),.data_out(wire_d5_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance530(.data_in(wire_d5_29),.data_out(wire_d5_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance531(.data_in(wire_d5_30),.data_out(wire_d5_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance532(.data_in(wire_d5_31),.data_out(wire_d5_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance533(.data_in(wire_d5_32),.data_out(wire_d5_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance534(.data_in(wire_d5_33),.data_out(d_out5),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance60(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	register #(.WIDTH(WIDTH)) register_instance61(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance62(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance63(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance64(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance65(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance66(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance67(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance68(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance69(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance629(.data_in(wire_d6_28),.data_out(wire_d6_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance630(.data_in(wire_d6_29),.data_out(wire_d6_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance631(.data_in(wire_d6_30),.data_out(wire_d6_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance632(.data_in(wire_d6_31),.data_out(wire_d6_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance633(.data_in(wire_d6_32),.data_out(wire_d6_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance634(.data_in(wire_d6_33),.data_out(d_out6),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance70(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	encoder #(.WIDTH(WIDTH)) encoder_instance71(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance72(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance73(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance74(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance75(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance76(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance77(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance78(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance79(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance729(.data_in(wire_d7_28),.data_out(wire_d7_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance730(.data_in(wire_d7_29),.data_out(wire_d7_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance731(.data_in(wire_d7_30),.data_out(wire_d7_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance732(.data_in(wire_d7_31),.data_out(wire_d7_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance733(.data_in(wire_d7_32),.data_out(wire_d7_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance734(.data_in(wire_d7_33),.data_out(d_out7),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance80(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	encoder #(.WIDTH(WIDTH)) encoder_instance81(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance82(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance83(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance84(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance85(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance86(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance87(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance88(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance89(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance829(.data_in(wire_d8_28),.data_out(wire_d8_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance830(.data_in(wire_d8_29),.data_out(wire_d8_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance831(.data_in(wire_d8_30),.data_out(wire_d8_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance832(.data_in(wire_d8_31),.data_out(wire_d8_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance833(.data_in(wire_d8_32),.data_out(wire_d8_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance834(.data_in(wire_d8_33),.data_out(d_out8),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance90(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	invertion #(.WIDTH(WIDTH)) invertion_instance91(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance92(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance93(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance94(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance95(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance96(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance97(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance98(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance99(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance929(.data_in(wire_d9_28),.data_out(wire_d9_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance930(.data_in(wire_d9_29),.data_out(wire_d9_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance931(.data_in(wire_d9_30),.data_out(wire_d9_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance932(.data_in(wire_d9_31),.data_out(wire_d9_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance933(.data_in(wire_d9_32),.data_out(wire_d9_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance934(.data_in(wire_d9_33),.data_out(d_out9),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance100(.data_in(d_in10),.data_out(wire_d10_0),.clk(clk),.rst(rst));            //channel 11
	invertion #(.WIDTH(WIDTH)) invertion_instance101(.data_in(wire_d10_0),.data_out(wire_d10_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance102(.data_in(wire_d10_1),.data_out(wire_d10_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance103(.data_in(wire_d10_2),.data_out(wire_d10_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance104(.data_in(wire_d10_3),.data_out(wire_d10_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance105(.data_in(wire_d10_4),.data_out(wire_d10_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance106(.data_in(wire_d10_5),.data_out(wire_d10_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance107(.data_in(wire_d10_6),.data_out(wire_d10_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance108(.data_in(wire_d10_7),.data_out(wire_d10_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance109(.data_in(wire_d10_8),.data_out(wire_d10_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1010(.data_in(wire_d10_9),.data_out(wire_d10_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1011(.data_in(wire_d10_10),.data_out(wire_d10_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1012(.data_in(wire_d10_11),.data_out(wire_d10_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1013(.data_in(wire_d10_12),.data_out(wire_d10_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1014(.data_in(wire_d10_13),.data_out(wire_d10_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1015(.data_in(wire_d10_14),.data_out(wire_d10_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1016(.data_in(wire_d10_15),.data_out(wire_d10_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1017(.data_in(wire_d10_16),.data_out(wire_d10_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1018(.data_in(wire_d10_17),.data_out(wire_d10_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1019(.data_in(wire_d10_18),.data_out(wire_d10_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1020(.data_in(wire_d10_19),.data_out(wire_d10_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1021(.data_in(wire_d10_20),.data_out(wire_d10_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1022(.data_in(wire_d10_21),.data_out(wire_d10_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1023(.data_in(wire_d10_22),.data_out(wire_d10_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1024(.data_in(wire_d10_23),.data_out(wire_d10_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1025(.data_in(wire_d10_24),.data_out(wire_d10_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1026(.data_in(wire_d10_25),.data_out(wire_d10_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1027(.data_in(wire_d10_26),.data_out(wire_d10_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1028(.data_in(wire_d10_27),.data_out(wire_d10_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1029(.data_in(wire_d10_28),.data_out(wire_d10_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1030(.data_in(wire_d10_29),.data_out(wire_d10_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1031(.data_in(wire_d10_30),.data_out(wire_d10_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1032(.data_in(wire_d10_31),.data_out(wire_d10_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1033(.data_in(wire_d10_32),.data_out(wire_d10_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1034(.data_in(wire_d10_33),.data_out(d_out10),.clk(clk),.rst(rst));


endmodule