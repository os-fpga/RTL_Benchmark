// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: rca_pkg.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2016-04-18-EP on Tue Mar 19 21:50:30 2019
//=============================================================================
// Description: Package for agent rca
//=============================================================================

package rca_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;


  `include "rca_trans.sv"
  `include "rca_config.sv"
  `include "rca_driver.sv"
  `include "rca_monitor.sv"
  `include "rca_sequencer.sv"
  `include "rca_coverage.sv"
  `include "rca_agent.sv"
  `include "rca_seq_lib.sv"

endpackage : rca_pkg
