//------------------------------------------------------------------------
// Filename     : atcbusdec301_config.vh
// Description  : specify AXI slave configurations
//------------------------------------------------------------------------
`include "config.inc"
`include "ae350_config.vh"
`include "ae350_const.vh"
`ifdef ATCBUSDEC301_CONFIG_VH
`else
`define ATCBUSDEC301_CONFIG_VH

`ifdef NDS_BIU_DATA_WIDTH_256
	`define ATCBUSDEC301_DATA_WIDTH_256
`else
`ifdef NDS_BIU_DATA_WIDTH_128
	`define ATCBUSDEC301_DATA_WIDTH_128
`else
`ifdef NDS_BIU_DATA_WIDTH_64
	`define ATCBUSDEC301_DATA_WIDTH_64
`else
	`define ATCBUSDEC301_DATA_WIDTH_32
`endif // NDS_BIU_DATA_WIDTH_64
`endif // NDS_BIU_DATA_WIDTH_128
`endif // NDS_BIU_DATA_WIDTH_256

//`define ATCBUSDEC301_DATA_WIDTH_256
//`define ATCBUSDEC301_DATA_WIDTH_128
//`define ATCBUSDEC301_DATA_WIDTH_64
`define ATCBUSDEC301_ID_WIDTH (`AE350_AXI_ID_WIDTH + 4)
`define ATCBUSDEC301_OOR_ERR_EN 

`define ATCBUSDEC301_SLV1_SUPPORT	// PLIC
`define ATCBUSDEC301_SLV2_SUPPORT	// PLMT
`ifndef PLATFORM_NO_PLIC_SW
`define ATCBUSDEC301_SLV3_SUPPORT	// PLIC_SW
`endif // PLATFORM_NO_PLIC_SW
`ifdef PLATFORM_DEBUG_SUBSYSTEM
        `define ATCBUSDEC301_SLV4_SUPPORT   // DEBUG
`endif // PLATFORM_DEBUG_SUBSYSTEM

//`define	ATCBUSDEC301_ADDR_DECODE_WIDTH	32
//`define	ATCBUSDEC301_SLV1_OFFSET	`ATCBUSDEC301_ADDR_DECODE_WIDTH'hE400_0000
//`define	ATCBUSDEC301_SLV2_OFFSET	`ATCBUSDEC301_ADDR_DECODE_WIDTH'hE600_0000
//`define	ATCBUSDEC301_SLV3_OFFSET	`ATCBUSDEC301_ADDR_DECODE_WIDTH'hE640_0000
//`define	ATCBUSDEC301_SLV4_OFFSET	`ATCBUSDEC301_ADDR_DECODE_WIDTH'hE680_0000
`define	ATCBUSDEC301_ADDR_DECODE_WIDTH	26
`define	ATCBUSDEC301_SLV1_OFFSET	`ATCBUSDEC301_ADDR_DECODE_WIDTH'h0
`define	ATCBUSDEC301_SLV2_OFFSET	`ATCBUSDEC301_ADDR_DECODE_WIDTH'h2000000
`define	ATCBUSDEC301_SLV3_OFFSET	`ATCBUSDEC301_ADDR_DECODE_WIDTH'h2400000
`define	ATCBUSDEC301_SLV4_OFFSET	`ATCBUSDEC301_ADDR_DECODE_WIDTH'h2800000
`define	ATCBUSDEC301_SLV1_SIZE		3	// PLIC 4 MiB
`define	ATCBUSDEC301_SLV2_SIZE		1	// PLMT	1 MiB
`define	ATCBUSDEC301_SLV3_SIZE		3	// PLIC_SW 4 MiB
`define	ATCBUSDEC301_SLV4_SIZE		1	// DEBUG 1MiB

`endif //ATCBUSDEC301_CONFIG_VH
