-- Xilinx Vhdl netlist produced by netgen application (version G.35)
-- Command       : -sim -ofmt vhdl -rpw 100 -w -s 4 MDCT_out.ncd MDCT_out.vhd 
-- Input file    : MDCT_out.ncd
-- Output file   : MDCT_out.vhd
-- Design name   : MDCT
-- # of Entities : 1
-- Xilinx        : f:/Xilinx
-- Device        : 3s1000ft256-4 (ADVANCED 1.32 2004-06-25)

-- This vhdl netlist is a simulation model and uses simulation 
-- primitives which may not represent the true implementation of the 
-- device, however the netlist is functionally correct and should not 
-- be modified. This file cannot be synthesized and should only be used 
-- with supported simulation tools.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library SIMPRIM;
use SIMPRIM.VCOMPONENTS.ALL;
use SIMPRIM.VPACKAGE.ALL;

entity MDCT is
  port (
    idv : in STD_LOGIC := 'X'; 
    rst : in STD_LOGIC := 'X'; 
    clk : in STD_LOGIC := 'X'; 
    ready : out STD_LOGIC; 
    odv : out STD_LOGIC; 
    odv1 : out STD_LOGIC; 
    dcto1 : out STD_LOGIC_VECTOR ( 11 downto 0 ); 
    dcto : out STD_LOGIC_VECTOR ( 11 downto 0 ); 
    dcti : in STD_LOGIC_VECTOR ( 7 downto 0 ) 
  );
end MDCT;

architecture STRUCTURE of MDCT is
  signal GLOBAL_LOGIC0 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1558 : STD_LOGIC; 
  signal clk_int : STD_LOGIC; 
  signal rst_int : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1421_add_10_ix61816z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1421_add_10_ix63810z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1421_add_10_ix268z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1421_add_10_ix2262z63342_O : STD_LOGIC; 
  signal U_DCT1D_nx2262z1 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1702 : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_0_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_0_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_1_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_1_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1580_add_47_ix61816z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_2_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_2_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_3_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_3_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1580_add_47_ix63810z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_4_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_4_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_5_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_5_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1580_add_47_ix268z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_6_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_6_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_7_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_7_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1580_add_47_ix2262z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_8_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_8_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_10_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_10_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1580_add_47_ix22763z63342_O : STD_LOGIC; 
  signal U_DCT2D_nx22763z1 : STD_LOGIC; 
  signal GLOBAL_LOGIC1 : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_0_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_0_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_1_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_1_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_97_sub_41_ix51546z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_2_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_2_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_3_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_3_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_97_sub_41_ix53540z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_4_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_4_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_5_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_5_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_97_sub_41_ix55534z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_6_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_6_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_7_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_7_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_97_sub_41_ix57528z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_8_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_8_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_10_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_10_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_97_sub_41_ix7189z63342_O : STD_LOGIC; 
  signal U_DCT2D_nx7189z1 : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_0_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_0_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_1_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_1_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_100_sub_44_ix36141z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_2_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_2_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_3_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_3_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_100_sub_44_ix38135z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_4_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_4_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_5_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_5_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_100_sub_44_ix40129z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_6_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_6_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_7_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_7_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_100_sub_44_ix42123z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_8_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_8_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_10_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_10_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_100_sub_44_ix16172z63342_O : STD_LOGIC; 
  signal U_DCT2D_nx16172z1 : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1420_add_9_ix1415z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1420_add_9_ix3409z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1420_add_9_ix5403z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1420_add_9_ix7397z63342_O : STD_LOGIC; 
  signal U_DCT1D_nx7397z1 : STD_LOGIC; 
  signal U_DCT2D_ix65206z64235_O : STD_LOGIC; 
  signal U_DCT2D_ix65206z64227_O : STD_LOGIC; 
  signal U_DCT2D_ix65206z64219_O : STD_LOGIC; 
  signal U_DCT2D_ix65206z64211_O : STD_LOGIC; 
  signal U_DCT2D_ix65206z64203_O : STD_LOGIC; 
  signal U_DCT2D_ix65206z64195_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z571 : STD_LOGIC; 
  signal U_DCT2D_ix65206z64185_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z607 : STD_LOGIC; 
  signal U_DCT2D_nx65206z604 : STD_LOGIC; 
  signal U_DCT2D_ix65206z64179_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z601 : STD_LOGIC; 
  signal U_DCT2D_nx65206z598 : STD_LOGIC; 
  signal U_DCT2D_ix65206z64173_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z595 : STD_LOGIC; 
  signal U_DCT2D_nx65206z592 : STD_LOGIC; 
  signal U_DCT2D_ix65206z64167_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z589 : STD_LOGIC; 
  signal U_DCT2D_nx65206z586 : STD_LOGIC; 
  signal U_DCT2D_ix65206z64161_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z583 : STD_LOGIC; 
  signal U_DCT2D_nx65206z580 : STD_LOGIC; 
  signal U_DCT2D_ix65206z64155_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z573 : STD_LOGIC; 
  signal U_DCT2D_ix65206z64151_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z572 : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_0_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_0_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_1_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_1_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1579_add_46_ix1415z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_2_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_2_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_3_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_3_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1579_add_46_ix3409z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_4_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_4_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_5_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_5_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1579_add_46_ix5403z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_6_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_6_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_7_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_7_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1579_add_46_ix7397z63342_O : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_8_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_8_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_10_Q : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_10_Q : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1579_add_46_ix30550z63342_O : STD_LOGIC; 
  signal U_DCT2D_nx30550z1 : STD_LOGIC; 
  signal U_DCT1D_rtlc5_83_sub_4_ix51546z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_83_sub_4_ix53540z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_83_sub_4_ix55534z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_83_sub_4_ix57528z63342_O : STD_LOGIC; 
  signal U_DCT1D_nx57528z1 : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63482_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63474_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63467_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63460_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63453_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63446_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63439_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z79 : STD_LOGIC; 
  signal U_DCT1D_rtlc5_86_sub_7_ix36141z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_86_sub_7_ix38135z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_86_sub_7_ix40129z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_86_sub_7_ix42123z63342_O : STD_LOGIC; 
  signal U_DCT1D_nx42123z1 : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1578_add_45_ix58986z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1578_add_45_ix56992z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1578_add_45_ix54998z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1578_add_45_ix53004z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1578_add_45_ix38337z63342_O : STD_LOGIC; 
  signal U_DCT2D_nx38337z1 : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63608_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63597_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63587_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63577_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63567_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63556_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63546_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63538_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z78 : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63742_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63735_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63728_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63721_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63714_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63706_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63699_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z253 : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1581_add_48_ix56681z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1581_add_48_ix58675z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1581_add_48_ix60669z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1581_add_48_ix62663z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1581_add_48_ix14976z63342_O : STD_LOGIC; 
  signal U_DCT2D_nx14976z1 : STD_LOGIC; 
  signal U_DCT2D_rtlc_389_add_65_ix65206z63383_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_389_add_65_ix65206z63376_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_389_add_65_ix65206z63369_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_389_add_65_ix65206z63362_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_389_add_65_ix65206z63355_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_389_add_65_ix65206z63348_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z5 : STD_LOGIC; 
  signal U_DCT1D_nx59700z428 : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63916_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z424 : STD_LOGIC; 
  signal U_DCT1D_nx59700z420 : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63904_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z416 : STD_LOGIC; 
  signal U_DCT1D_nx59700z412 : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63892_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z408 : STD_LOGIC; 
  signal U_DCT1D_nx59700z404 : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63880_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z400 : STD_LOGIC; 
  signal U_DCT1D_nx59700z396 : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63868_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z392 : STD_LOGIC; 
  signal U_DCT1D_nx59700z388 : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63856_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z384 : STD_LOGIC; 
  signal U_DCT1D_nx59700z253 : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63846_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_99_sub_43_ix41276z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_99_sub_43_ix43270z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_99_sub_43_ix45264z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_99_sub_43_ix47258z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_99_sub_43_ix8385z63342_O : STD_LOGIC; 
  signal U_DCT2D_nx8385z1 : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1419_add_8_ix58986z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1419_add_8_ix56992z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1419_add_8_ix54998z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1419_add_8_ix53004z63342_O : STD_LOGIC; 
  signal U_DCT1D_nx53004z1 : STD_LOGIC; 
  signal U_DCT1D_rtlc5_84_sub_5_ix46411z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_84_sub_5_ix48405z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_84_sub_5_ix50399z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_84_sub_5_ix52393z63342_O : STD_LOGIC; 
  signal U_DCT1D_nx52393z1 : STD_LOGIC; 
  signal U_DCT2D_rtlc5_98_sub_42_ix46411z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_98_sub_42_ix48405z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_98_sub_42_ix50399z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_98_sub_42_ix52393z63342_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5_98_sub_42_ix64938z63342_O : STD_LOGIC; 
  signal U_DCT2D_nx64938z1 : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1422_add_11_ix56681z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1422_add_11_ix58675z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1422_add_11_ix60669z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1422_add_11_ix62663z63342_O : STD_LOGIC; 
  signal U_DCT1D_nx62663z1 : STD_LOGIC; 
  signal U_DCT2D_rtlc_387_add_64_ix65206z63429_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_387_add_64_ix65206z63422_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_387_add_64_ix65206z63415_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_387_add_64_ix65206z63408_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_387_add_64_ix65206z63401_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_387_add_64_ix65206z63392_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z42 : STD_LOGIC; 
  signal U_DCT2D_rtlc_396_add_68_ix65206z63832_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_396_add_68_ix65206z63825_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_396_add_68_ix65206z63818_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_396_add_68_ix65206z63811_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_396_add_68_ix65206z63804_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_396_add_68_ix65206z63797_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z334 : STD_LOGIC; 
  signal U_DCT1D_rtlc5_85_sub_6_ix41276z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_85_sub_6_ix43270z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_85_sub_6_ix45264z63342_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5_85_sub_6_ix47258z63342_O : STD_LOGIC; 
  signal U_DCT1D_nx47258z1 : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63531_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63524_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63517_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63510_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63503_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63496_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63489_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z121 : STD_LOGIC; 
  signal U_DCT2D_nx65206z570 : STD_LOGIC; 
  signal U_DCT2D_nx65206z567 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64139_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z564 : STD_LOGIC; 
  signal U_DCT2D_nx65206z561 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64131_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z557 : STD_LOGIC; 
  signal U_DCT2D_nx65206z553 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64119_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z549 : STD_LOGIC; 
  signal U_DCT2D_nx65206z545 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64108_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z541 : STD_LOGIC; 
  signal U_DCT2D_nx65206z537 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64097_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z533 : STD_LOGIC; 
  signal U_DCT2D_nx65206z529 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64087_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z525 : STD_LOGIC; 
  signal U_DCT2D_nx65206z521 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64077_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z3 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64069_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64060_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64310_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64302_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64290_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64280_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64270_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64260_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64248_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z1 : STD_LOGIC; 
  signal U_DCT1D_nx59700z493 : STD_LOGIC; 
  signal U_DCT1D_nx59700z490 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z64000_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z487 : STD_LOGIC; 
  signal U_DCT1D_nx59700z484 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63992_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z480 : STD_LOGIC; 
  signal U_DCT1D_nx59700z476 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63980_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z472 : STD_LOGIC; 
  signal U_DCT1D_nx59700z468 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63968_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z464 : STD_LOGIC; 
  signal U_DCT1D_nx59700z460 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63957_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z456 : STD_LOGIC; 
  signal U_DCT1D_nx59700z452 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63947_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z448 : STD_LOGIC; 
  signal U_DCT1D_nx59700z444 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63937_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z3 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63929_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_512_add_28_ix59700z63383_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_512_add_28_ix59700z63376_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_512_add_28_ix59700z63369_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_512_add_28_ix59700z63362_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_512_add_28_ix59700z63355_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_512_add_28_ix59700z63348_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z5 : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z64046_O : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z64034_O : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z64022_O : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z64010_O : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z63998_O : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z63986_O : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z63975_O : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z63966_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z252 : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63742_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63735_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63728_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63721_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63714_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63707_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63700_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z255 : STD_LOGIC; 
  signal U_DCT1D_nx59700z330 : STD_LOGIC; 
  signal U_DCT1D_nx59700z333 : STD_LOGIC; 
  signal U_DCT1D_nx59700z332 : STD_LOGIC; 
  signal U_DCT1D_ix740_modgen_add_290_ix59700z63789_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z327 : STD_LOGIC; 
  signal U_DCT1D_nx59700z324 : STD_LOGIC; 
  signal U_DCT1D_ix740_modgen_add_290_ix59700z63781_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z321 : STD_LOGIC; 
  signal U_DCT1D_nx59700z318 : STD_LOGIC; 
  signal U_DCT1D_ix740_modgen_add_290_ix59700z63773_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z315 : STD_LOGIC; 
  signal U_DCT1D_nx59700z312 : STD_LOGIC; 
  signal U_DCT1D_ix740_modgen_add_290_ix59700z63765_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z309 : STD_LOGIC; 
  signal U_DCT1D_nx59700z306 : STD_LOGIC; 
  signal U_DCT1D_ix740_modgen_add_290_ix59700z63757_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z303 : STD_LOGIC; 
  signal U_DCT1D_nx59700z300 : STD_LOGIC; 
  signal U_DCT1D_ix740_modgen_add_290_ix59700z63749_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z254 : STD_LOGIC; 
  signal U_DCT2D_rtlc_394_add_67_ix65206z63788_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_394_add_67_ix65206z63781_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_394_add_67_ix65206z63774_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_394_add_67_ix65206z63767_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_394_add_67_ix65206z63760_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_394_add_67_ix65206z63753_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z297 : STD_LOGIC; 
  signal U_DCT2D_nx65206z248 : STD_LOGIC; 
  signal U_DCT2D_nx65206z251 : STD_LOGIC; 
  signal U_DCT2D_nx65206z250 : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63683_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z245 : STD_LOGIC; 
  signal U_DCT2D_nx65206z242 : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63671_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z239 : STD_LOGIC; 
  signal U_DCT2D_nx65206z236 : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63659_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z233 : STD_LOGIC; 
  signal U_DCT2D_nx65206z230 : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63647_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z227 : STD_LOGIC; 
  signal U_DCT2D_nx65206z224 : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63635_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z221 : STD_LOGIC; 
  signal U_DCT2D_nx65206z218 : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63624_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z215 : STD_LOGIC; 
  signal U_DCT2D_nx65206z212 : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63615_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z4 : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63482_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63474_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63467_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63460_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63453_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63446_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63439_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z79 : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63531_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63524_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63517_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63510_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63503_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63496_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63489_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z121 : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63904_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63892_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63880_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63868_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63856_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63847_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63839_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z296 : STD_LOGIC; 
  signal U_DCT1D_rtlc_510_add_27_ix59700z63429_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_510_add_27_ix59700z63422_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_510_add_27_ix59700z63415_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_510_add_27_ix59700z63408_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_510_add_27_ix59700z63401_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_510_add_27_ix59700z63392_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z42 : STD_LOGIC; 
  signal U_DCT1D_nx59700z248 : STD_LOGIC; 
  signal U_DCT1D_nx59700z251 : STD_LOGIC; 
  signal U_DCT1D_nx59700z250 : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63683_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z245 : STD_LOGIC; 
  signal U_DCT1D_nx59700z242 : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63671_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z239 : STD_LOGIC; 
  signal U_DCT1D_nx59700z236 : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63659_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z233 : STD_LOGIC; 
  signal U_DCT1D_nx59700z230 : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63647_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z227 : STD_LOGIC; 
  signal U_DCT1D_nx59700z224 : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63635_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z221 : STD_LOGIC; 
  signal U_DCT1D_nx59700z218 : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63624_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z215 : STD_LOGIC; 
  signal U_DCT1D_nx59700z212 : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63615_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z4 : STD_LOGIC; 
  signal U_DCT1D_ix59700z64053_O : STD_LOGIC; 
  signal U_DCT1D_ix59700z64047_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n2660 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n2659 : STD_LOGIC; 
  signal U_DCT1D_ix59700z64038_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n2658 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n2657 : STD_LOGIC; 
  signal U_DCT1D_ix59700z64029_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n2656 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n2655 : STD_LOGIC; 
  signal U_DCT1D_ix59700z64020_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n2654 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n2653 : STD_LOGIC; 
  signal U_DCT1D_ix59700z64012_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z1 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n2652 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n2651 : STD_LOGIC; 
  signal U_DCT1D_ix59700z63834_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z369 : STD_LOGIC; 
  signal U_DCT1D_nx59700z366 : STD_LOGIC; 
  signal U_DCT1D_ix59700z63828_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z363 : STD_LOGIC; 
  signal U_DCT1D_nx59700z360 : STD_LOGIC; 
  signal U_DCT1D_ix59700z63822_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z357 : STD_LOGIC; 
  signal U_DCT1D_nx59700z354 : STD_LOGIC; 
  signal U_DCT1D_ix59700z63816_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z351 : STD_LOGIC; 
  signal U_DCT1D_nx59700z348 : STD_LOGIC; 
  signal U_DCT1D_ix59700z63810_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z345 : STD_LOGIC; 
  signal U_DCT1D_nx59700z342 : STD_LOGIC; 
  signal U_DCT1D_ix59700z63804_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z335 : STD_LOGIC; 
  signal U_DCT1D_ix59700z63800_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z334 : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63608_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63597_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63587_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63577_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63567_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63556_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63546_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63538_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z78 : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63959_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63952_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63945_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63938_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63931_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63924_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63917_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z413 : STD_LOGIC; 
  signal nx53675z21 : STD_LOGIC; 
  signal nx53675z18 : STD_LOGIC; 
  signal nx53675z27 : STD_LOGIC; 
  signal nx53675z24 : STD_LOGIC; 
  signal nx53675z587 : STD_LOGIC; 
  signal nx53675z585 : STD_LOGIC; 
  signal U2_ROME8_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROME8_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z658 : STD_LOGIC; 
  signal nx53675z655 : STD_LOGIC; 
  signal nx53675z664 : STD_LOGIC; 
  signal nx53675z661 : STD_LOGIC; 
  signal nx53675z162 : STD_LOGIC; 
  signal nx53675z159 : STD_LOGIC; 
  signal nx53675z97 : STD_LOGIC; 
  signal nx53675z94 : STD_LOGIC; 
  signal nx53675z103 : STD_LOGIC; 
  signal nx53675z100 : STD_LOGIC; 
  signal nx53675z109 : STD_LOGIC; 
  signal nx53675z106 : STD_LOGIC; 
  signal nx53675z115 : STD_LOGIC; 
  signal nx53675z112 : STD_LOGIC; 
  signal nx53675z33 : STD_LOGIC; 
  signal nx53675z30 : STD_LOGIC; 
  signal nx53675z39 : STD_LOGIC; 
  signal nx53675z36 : STD_LOGIC; 
  signal nx53675z45 : STD_LOGIC; 
  signal nx53675z42 : STD_LOGIC; 
  signal nx53675z51 : STD_LOGIC; 
  signal nx53675z48 : STD_LOGIC; 
  signal nx53675z57 : STD_LOGIC; 
  signal nx53675z54 : STD_LOGIC; 
  signal nx53675z593 : STD_LOGIC; 
  signal nx53675z590 : STD_LOGIC; 
  signal nx53675z599 : STD_LOGIC; 
  signal nx53675z596 : STD_LOGIC; 
  signal nx53675z605 : STD_LOGIC; 
  signal nx53675z602 : STD_LOGIC; 
  signal nx53675z611 : STD_LOGIC; 
  signal nx53675z608 : STD_LOGIC; 
  signal nx53675z617 : STD_LOGIC; 
  signal nx53675z614 : STD_LOGIC; 
  signal nx53675z794 : STD_LOGIC; 
  signal nx53675z792 : STD_LOGIC; 
  signal nx53675z723 : STD_LOGIC; 
  signal nx53675z720 : STD_LOGIC; 
  signal nx53675z729 : STD_LOGIC; 
  signal nx53675z726 : STD_LOGIC; 
  signal nx53675z735 : STD_LOGIC; 
  signal nx53675z732 : STD_LOGIC; 
  signal nx53675z1292 : STD_LOGIC; 
  signal nx53675z1289 : STD_LOGIC; 
  signal nx53675z1298 : STD_LOGIC; 
  signal nx53675z1295 : STD_LOGIC; 
  signal nx53675z1304 : STD_LOGIC; 
  signal nx53675z1301 : STD_LOGIC; 
  signal nx53675z1310 : STD_LOGIC; 
  signal nx53675z1307 : STD_LOGIC; 
  signal nx53675z1359 : STD_LOGIC; 
  signal nx53675z1356 : STD_LOGIC; 
  signal nx53675z1365 : STD_LOGIC; 
  signal nx53675z1362 : STD_LOGIC; 
  signal nx53675z670 : STD_LOGIC; 
  signal nx53675z667 : STD_LOGIC; 
  signal nx53675z676 : STD_LOGIC; 
  signal nx53675z673 : STD_LOGIC; 
  signal nx53675z682 : STD_LOGIC; 
  signal nx53675z679 : STD_LOGIC; 
  signal nx53675z688 : STD_LOGIC; 
  signal nx53675z685 : STD_LOGIC; 
  signal nx53675z694 : STD_LOGIC; 
  signal nx53675z691 : STD_LOGIC; 
  signal nx53675z168 : STD_LOGIC; 
  signal nx53675z165 : STD_LOGIC; 
  signal nx53675z174 : STD_LOGIC; 
  signal nx53675z171 : STD_LOGIC; 
  signal nx53675z180 : STD_LOGIC; 
  signal nx53675z177 : STD_LOGIC; 
  signal nx53675z186 : STD_LOGIC; 
  signal nx53675z183 : STD_LOGIC; 
  signal nx53675z191 : STD_LOGIC; 
  signal nx53675z189 : STD_LOGIC; 
  signal nx53675z132 : STD_LOGIC; 
  signal nx53675z130 : STD_LOGIC; 
  signal nx53675z73 : STD_LOGIC; 
  signal nx53675z70 : STD_LOGIC; 
  signal nx53675z1426 : STD_LOGIC; 
  signal nx53675z1424 : STD_LOGIC; 
  signal nx53675z652 : STD_LOGIC; 
  signal nx53675z650 : STD_LOGIC; 
  signal nx53675z304 : STD_LOGIC; 
  signal nx53675z301 : STD_LOGIC; 
  signal nx53675z310 : STD_LOGIC; 
  signal nx53675z307 : STD_LOGIC; 
  signal nx53675z67 : STD_LOGIC; 
  signal nx53675z65 : STD_LOGIC; 
  signal nx53675z79 : STD_LOGIC; 
  signal nx53675z76 : STD_LOGIC; 
  signal nx53675z85 : STD_LOGIC; 
  signal nx53675z82 : STD_LOGIC; 
  signal nx53675z121 : STD_LOGIC; 
  signal nx53675z118 : STD_LOGIC; 
  signal nx53675z126 : STD_LOGIC; 
  signal nx53675z124 : STD_LOGIC; 
  signal U2_ROME1_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROME1_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z9 : STD_LOGIC; 
  signal nx53675z6 : STD_LOGIC; 
  signal nx53675z15 : STD_LOGIC; 
  signal nx53675z12 : STD_LOGIC; 
  signal nx53675z62 : STD_LOGIC; 
  signal nx53675z60 : STD_LOGIC; 
  signal nx53675z623 : STD_LOGIC; 
  signal nx53675z620 : STD_LOGIC; 
  signal nx53675z629 : STD_LOGIC; 
  signal nx53675z626 : STD_LOGIC; 
  signal nx53675z635 : STD_LOGIC; 
  signal nx53675z632 : STD_LOGIC; 
  signal nx53675z641 : STD_LOGIC; 
  signal nx53675z638 : STD_LOGIC; 
  signal nx53675z646 : STD_LOGIC; 
  signal nx53675z644 : STD_LOGIC; 
  signal nx53675z3 : STD_LOGIC; 
  signal nx53675z1 : STD_LOGIC; 
  signal nx53675z873 : STD_LOGIC; 
  signal nx53675z871 : STD_LOGIC; 
  signal nx53675z939 : STD_LOGIC; 
  signal nx53675z936 : STD_LOGIC; 
  signal nx53675z800 : STD_LOGIC; 
  signal nx53675z797 : STD_LOGIC; 
  signal nx53675z806 : STD_LOGIC; 
  signal nx53675z803 : STD_LOGIC; 
  signal nx53675z812 : STD_LOGIC; 
  signal nx53675z809 : STD_LOGIC; 
  signal nx53675z818 : STD_LOGIC; 
  signal nx53675z815 : STD_LOGIC; 
  signal nx53675z824 : STD_LOGIC; 
  signal nx53675z821 : STD_LOGIC; 
  signal U2_ROMO1_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROMO1_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z741 : STD_LOGIC; 
  signal nx53675z738 : STD_LOGIC; 
  signal nx53675z747 : STD_LOGIC; 
  signal nx53675z744 : STD_LOGIC; 
  signal nx53675z753 : STD_LOGIC; 
  signal nx53675z750 : STD_LOGIC; 
  signal nx53675z759 : STD_LOGIC; 
  signal nx53675z756 : STD_LOGIC; 
  signal nx53675z765 : STD_LOGIC; 
  signal nx53675z762 : STD_LOGIC; 
  signal nx53675z203 : STD_LOGIC; 
  signal nx53675z200 : STD_LOGIC; 
  signal nx53675z239 : STD_LOGIC; 
  signal nx53675z236 : STD_LOGIC; 
  signal nx53675z251 : STD_LOGIC; 
  signal nx53675z248 : STD_LOGIC; 
  signal U2_ROME3_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROME3_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z1012 : STD_LOGIC; 
  signal nx53675z1009 : STD_LOGIC; 
  signal nx53675z197 : STD_LOGIC; 
  signal nx53675z195 : STD_LOGIC; 
  signal nx53675z1371 : STD_LOGIC; 
  signal nx53675z1368 : STD_LOGIC; 
  signal nx53675z1377 : STD_LOGIC; 
  signal nx53675z1374 : STD_LOGIC; 
  signal nx53675z1383 : STD_LOGIC; 
  signal nx53675z1380 : STD_LOGIC; 
  signal nx53675z1389 : STD_LOGIC; 
  signal nx53675z1386 : STD_LOGIC; 
  signal nx53675z1395 : STD_LOGIC; 
  signal nx53675z1392 : STD_LOGIC; 
  signal nx53675z1316 : STD_LOGIC; 
  signal nx53675z1313 : STD_LOGIC; 
  signal nx53675z1322 : STD_LOGIC; 
  signal nx53675z1319 : STD_LOGIC; 
  signal nx53675z1328 : STD_LOGIC; 
  signal nx53675z1325 : STD_LOGIC; 
  signal nx53675z1334 : STD_LOGIC; 
  signal nx53675z1331 : STD_LOGIC; 
  signal nx53675z1340 : STD_LOGIC; 
  signal nx53675z1337 : STD_LOGIC; 
  signal nx53675z375 : STD_LOGIC; 
  signal nx53675z372 : STD_LOGIC; 
  signal nx53675z381 : STD_LOGIC; 
  signal nx53675z378 : STD_LOGIC; 
  signal U2_ROMO7_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROMO7_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z700 : STD_LOGIC; 
  signal nx53675z697 : STD_LOGIC; 
  signal nx53675z706 : STD_LOGIC; 
  signal nx53675z703 : STD_LOGIC; 
  signal nx53675z711 : STD_LOGIC; 
  signal nx53675z709 : STD_LOGIC; 
  signal U2_ROME10_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROME10_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z327 : STD_LOGIC; 
  signal nx53675z325 : STD_LOGIC; 
  signal nx53675z138 : STD_LOGIC; 
  signal nx53675z135 : STD_LOGIC; 
  signal nx53675z144 : STD_LOGIC; 
  signal nx53675z141 : STD_LOGIC; 
  signal nx53675z150 : STD_LOGIC; 
  signal nx53675z147 : STD_LOGIC; 
  signal nx53675z156 : STD_LOGIC; 
  signal nx53675z153 : STD_LOGIC; 
  signal U2_ROME2_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROME2_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z1438 : STD_LOGIC; 
  signal nx53675z1435 : STD_LOGIC; 
  signal nx53675z1444 : STD_LOGIC; 
  signal nx53675z1441 : STD_LOGIC; 
  signal nx53675z1450 : STD_LOGIC; 
  signal nx53675z1447 : STD_LOGIC; 
  signal nx53675z1456 : STD_LOGIC; 
  signal nx53675z1453 : STD_LOGIC; 
  signal nx53675z1462 : STD_LOGIC; 
  signal nx53675z1459 : STD_LOGIC; 
  signal nx53675z392 : STD_LOGIC; 
  signal nx53675z390 : STD_LOGIC; 
  signal nx53675z268 : STD_LOGIC; 
  signal nx53675z265 : STD_LOGIC; 
  signal nx53675z274 : STD_LOGIC; 
  signal nx53675z271 : STD_LOGIC; 
  signal nx53675z280 : STD_LOGIC; 
  signal nx53675z277 : STD_LOGIC; 
  signal nx53675z316 : STD_LOGIC; 
  signal nx53675z313 : STD_LOGIC; 
  signal nx53675z321 : STD_LOGIC; 
  signal nx53675z319 : STD_LOGIC; 
  signal U2_ROME4_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROME4_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z91 : STD_LOGIC; 
  signal nx53675z88 : STD_LOGIC; 
  signal nx53675z1511 : STD_LOGIC; 
  signal nx53675z1508 : STD_LOGIC; 
  signal nx53675z958 : STD_LOGIC; 
  signal nx53675z955 : STD_LOGIC; 
  signal nx53675z1018 : STD_LOGIC; 
  signal nx53675z1015 : STD_LOGIC; 
  signal nx53675z879 : STD_LOGIC; 
  signal nx53675z876 : STD_LOGIC; 
  signal nx53675z885 : STD_LOGIC; 
  signal nx53675z882 : STD_LOGIC; 
  signal nx53675z891 : STD_LOGIC; 
  signal nx53675z888 : STD_LOGIC; 
  signal nx53675z897 : STD_LOGIC; 
  signal nx53675z894 : STD_LOGIC; 
  signal nx53675z903 : STD_LOGIC; 
  signal nx53675z900 : STD_LOGIC; 
  signal U2_ROME9_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROME9_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z1505 : STD_LOGIC; 
  signal nx53675z1503 : STD_LOGIC; 
  signal nx53675z1523 : STD_LOGIC; 
  signal nx53675z1520 : STD_LOGIC; 
  signal nx53675z1571 : STD_LOGIC; 
  signal nx53675z1568 : STD_LOGIC; 
  signal nx53675z1577 : STD_LOGIC; 
  signal nx53675z1574 : STD_LOGIC; 
  signal U2_ROMO10_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROMO10_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal U2_ROMO9_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROMO9_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z1079 : STD_LOGIC; 
  signal nx53675z1076 : STD_LOGIC; 
  signal nx53675z952 : STD_LOGIC; 
  signal nx53675z950 : STD_LOGIC; 
  signal nx53675z945 : STD_LOGIC; 
  signal nx53675z942 : STD_LOGIC; 
  signal U2_ROMO2_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROMO2_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z830 : STD_LOGIC; 
  signal nx53675z827 : STD_LOGIC; 
  signal nx53675z836 : STD_LOGIC; 
  signal nx53675z833 : STD_LOGIC; 
  signal nx53675z842 : STD_LOGIC; 
  signal nx53675z839 : STD_LOGIC; 
  signal nx53675z848 : STD_LOGIC; 
  signal nx53675z845 : STD_LOGIC; 
  signal nx53675z854 : STD_LOGIC; 
  signal nx53675z851 : STD_LOGIC; 
  signal nx53675z398 : STD_LOGIC; 
  signal nx53675z395 : STD_LOGIC; 
  signal nx53675z446 : STD_LOGIC; 
  signal nx53675z443 : STD_LOGIC; 
  signal nx53675z451 : STD_LOGIC; 
  signal nx53675z449 : STD_LOGIC; 
  signal U2_ROME6_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROME6_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z771 : STD_LOGIC; 
  signal nx53675z768 : STD_LOGIC; 
  signal nx53675z777 : STD_LOGIC; 
  signal nx53675z774 : STD_LOGIC; 
  signal nx53675z783 : STD_LOGIC; 
  signal nx53675z780 : STD_LOGIC; 
  signal nx53675z789 : STD_LOGIC; 
  signal nx53675z786 : STD_LOGIC; 
  signal nx53675z215 : STD_LOGIC; 
  signal nx53675z212 : STD_LOGIC; 
  signal nx53675z227 : STD_LOGIC; 
  signal nx53675z224 : STD_LOGIC; 
  signal nx53675z1043 : STD_LOGIC; 
  signal nx53675z1040 : STD_LOGIC; 
  signal nx53675z1024 : STD_LOGIC; 
  signal nx53675z1021 : STD_LOGIC; 
  signal nx53675z717 : STD_LOGIC; 
  signal nx53675z715 : STD_LOGIC; 
  signal nx53675z1353 : STD_LOGIC; 
  signal nx53675z1350 : STD_LOGIC; 
  signal nx53675z1401 : STD_LOGIC; 
  signal nx53675z1398 : STD_LOGIC; 
  signal nx53675z1407 : STD_LOGIC; 
  signal nx53675z1404 : STD_LOGIC; 
  signal nx53675z1413 : STD_LOGIC; 
  signal nx53675z1410 : STD_LOGIC; 
  signal nx53675z333 : STD_LOGIC; 
  signal nx53675z330 : STD_LOGIC; 
  signal nx53675z339 : STD_LOGIC; 
  signal nx53675z336 : STD_LOGIC; 
  signal nx53675z345 : STD_LOGIC; 
  signal nx53675z342 : STD_LOGIC; 
  signal nx53675z351 : STD_LOGIC; 
  signal nx53675z348 : STD_LOGIC; 
  signal nx53675z386 : STD_LOGIC; 
  signal nx53675z384 : STD_LOGIC; 
  signal U2_ROME5_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROME5_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z1347 : STD_LOGIC; 
  signal nx53675z1345 : STD_LOGIC; 
  signal nx53675z1419 : STD_LOGIC; 
  signal nx53675z1416 : STD_LOGIC; 
  signal nx53675z463 : STD_LOGIC; 
  signal nx53675z460 : STD_LOGIC; 
  signal nx53675z469 : STD_LOGIC; 
  signal nx53675z466 : STD_LOGIC; 
  signal nx53675z516 : STD_LOGIC; 
  signal nx53675z514 : STD_LOGIC; 
  signal U2_ROME7_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROME7_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z1468 : STD_LOGIC; 
  signal nx53675z1465 : STD_LOGIC; 
  signal nx53675z1474 : STD_LOGIC; 
  signal nx53675z1471 : STD_LOGIC; 
  signal nx53675z1480 : STD_LOGIC; 
  signal nx53675z1477 : STD_LOGIC; 
  signal nx53675z1486 : STD_LOGIC; 
  signal nx53675z1483 : STD_LOGIC; 
  signal U2_ROMO8_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROMO8_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z1085 : STD_LOGIC; 
  signal nx53675z1082 : STD_LOGIC; 
  signal nx53675z286 : STD_LOGIC; 
  signal nx53675z283 : STD_LOGIC; 
  signal nx53675z292 : STD_LOGIC; 
  signal nx53675z289 : STD_LOGIC; 
  signal nx53675z298 : STD_LOGIC; 
  signal nx53675z295 : STD_LOGIC; 
  signal nx53675z209 : STD_LOGIC; 
  signal nx53675z206 : STD_LOGIC; 
  signal nx53675z233 : STD_LOGIC; 
  signal nx53675z230 : STD_LOGIC; 
  signal nx53675z1492 : STD_LOGIC; 
  signal nx53675z1489 : STD_LOGIC; 
  signal nx53675z1037 : STD_LOGIC; 
  signal nx53675z1034 : STD_LOGIC; 
  signal nx53675z970 : STD_LOGIC; 
  signal nx53675z967 : STD_LOGIC; 
  signal nx53675z982 : STD_LOGIC; 
  signal nx53675z979 : STD_LOGIC; 
  signal U2_ROMO3_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROMO3_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z909 : STD_LOGIC; 
  signal nx53675z906 : STD_LOGIC; 
  signal nx53675z915 : STD_LOGIC; 
  signal nx53675z912 : STD_LOGIC; 
  signal nx53675z921 : STD_LOGIC; 
  signal nx53675z918 : STD_LOGIC; 
  signal nx53675z927 : STD_LOGIC; 
  signal nx53675z924 : STD_LOGIC; 
  signal nx53675z1529 : STD_LOGIC; 
  signal nx53675z1526 : STD_LOGIC; 
  signal nx53675z1535 : STD_LOGIC; 
  signal nx53675z1532 : STD_LOGIC; 
  signal nx53675z1541 : STD_LOGIC; 
  signal nx53675z1538 : STD_LOGIC; 
  signal nx53675z1547 : STD_LOGIC; 
  signal nx53675z1544 : STD_LOGIC; 
  signal nx53675z1553 : STD_LOGIC; 
  signal nx53675z1550 : STD_LOGIC; 
  signal nx53675z1031 : STD_LOGIC; 
  signal nx53675z1029 : STD_LOGIC; 
  signal nx53675z860 : STD_LOGIC; 
  signal nx53675z857 : STD_LOGIC; 
  signal nx53675z866 : STD_LOGIC; 
  signal nx53675z863 : STD_LOGIC; 
  signal nx53675z457 : STD_LOGIC; 
  signal nx53675z455 : STD_LOGIC; 
  signal nx53675z404 : STD_LOGIC; 
  signal nx53675z401 : STD_LOGIC; 
  signal nx53675z410 : STD_LOGIC; 
  signal nx53675z407 : STD_LOGIC; 
  signal nx53675z416 : STD_LOGIC; 
  signal nx53675z413 : STD_LOGIC; 
  signal nx53675z422 : STD_LOGIC; 
  signal nx53675z419 : STD_LOGIC; 
  signal nx53675z428 : STD_LOGIC; 
  signal nx53675z425 : STD_LOGIC; 
  signal nx53675z1091 : STD_LOGIC; 
  signal nx53675z1088 : STD_LOGIC; 
  signal nx53675z1103 : STD_LOGIC; 
  signal nx53675z1100 : STD_LOGIC; 
  signal nx53675z1219 : STD_LOGIC; 
  signal nx53675z1216 : STD_LOGIC; 
  signal nx53675z1225 : STD_LOGIC; 
  signal nx53675z1222 : STD_LOGIC; 
  signal nx53675z1110 : STD_LOGIC; 
  signal nx53675z1108 : STD_LOGIC; 
  signal nx53675z1152 : STD_LOGIC; 
  signal nx53675z1149 : STD_LOGIC; 
  signal nx53675z1158 : STD_LOGIC; 
  signal nx53675z1155 : STD_LOGIC; 
  signal nx53675z1164 : STD_LOGIC; 
  signal nx53675z1161 : STD_LOGIC; 
  signal nx53675z1170 : STD_LOGIC; 
  signal nx53675z1167 : STD_LOGIC; 
  signal U2_ROMO4_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROMO4_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z528 : STD_LOGIC; 
  signal nx53675z525 : STD_LOGIC; 
  signal nx53675z534 : STD_LOGIC; 
  signal nx53675z531 : STD_LOGIC; 
  signal nx53675z540 : STD_LOGIC; 
  signal nx53675z537 : STD_LOGIC; 
  signal nx53675z546 : STD_LOGIC; 
  signal nx53675z543 : STD_LOGIC; 
  signal nx53675z262 : STD_LOGIC; 
  signal nx53675z260 : STD_LOGIC; 
  signal nx53675z522 : STD_LOGIC; 
  signal nx53675z520 : STD_LOGIC; 
  signal nx53675z357 : STD_LOGIC; 
  signal nx53675z354 : STD_LOGIC; 
  signal nx53675z363 : STD_LOGIC; 
  signal nx53675z360 : STD_LOGIC; 
  signal nx53675z369 : STD_LOGIC; 
  signal nx53675z366 : STD_LOGIC; 
  signal nx53675z475 : STD_LOGIC; 
  signal nx53675z472 : STD_LOGIC; 
  signal nx53675z481 : STD_LOGIC; 
  signal nx53675z478 : STD_LOGIC; 
  signal nx53675z487 : STD_LOGIC; 
  signal nx53675z484 : STD_LOGIC; 
  signal nx53675z493 : STD_LOGIC; 
  signal nx53675z490 : STD_LOGIC; 
  signal nx53675z499 : STD_LOGIC; 
  signal nx53675z496 : STD_LOGIC; 
  signal nx53675z1432 : STD_LOGIC; 
  signal nx53675z1429 : STD_LOGIC; 
  signal nx53675z1116 : STD_LOGIC; 
  signal nx53675z1113 : STD_LOGIC; 
  signal nx53675z1097 : STD_LOGIC; 
  signal nx53675z1094 : STD_LOGIC; 
  signal nx53675z221 : STD_LOGIC; 
  signal nx53675z218 : STD_LOGIC; 
  signal nx53675z245 : STD_LOGIC; 
  signal nx53675z242 : STD_LOGIC; 
  signal nx53675z256 : STD_LOGIC; 
  signal nx53675z254 : STD_LOGIC; 
  signal nx53675z1049 : STD_LOGIC; 
  signal nx53675z1046 : STD_LOGIC; 
  signal nx53675z994 : STD_LOGIC; 
  signal nx53675z991 : STD_LOGIC; 
  signal nx53675z1006 : STD_LOGIC; 
  signal nx53675z1003 : STD_LOGIC; 
  signal nx53675z1559 : STD_LOGIC; 
  signal nx53675z1556 : STD_LOGIC; 
  signal nx53675z1565 : STD_LOGIC; 
  signal nx53675z1562 : STD_LOGIC; 
  signal nx53675z1055 : STD_LOGIC; 
  signal nx53675z1052 : STD_LOGIC; 
  signal nx53675z1061 : STD_LOGIC; 
  signal nx53675z1058 : STD_LOGIC; 
  signal nx53675z1067 : STD_LOGIC; 
  signal nx53675z1064 : STD_LOGIC; 
  signal nx53675z1073 : STD_LOGIC; 
  signal nx53675z1070 : STD_LOGIC; 
  signal nx53675z434 : STD_LOGIC; 
  signal nx53675z431 : STD_LOGIC; 
  signal nx53675z440 : STD_LOGIC; 
  signal nx53675z437 : STD_LOGIC; 
  signal nx53675z1122 : STD_LOGIC; 
  signal nx53675z1119 : STD_LOGIC; 
  signal nx53675z1498 : STD_LOGIC; 
  signal nx53675z1495 : STD_LOGIC; 
  signal nx53675z1189 : STD_LOGIC; 
  signal nx53675z1187 : STD_LOGIC; 
  signal nx53675z1231 : STD_LOGIC; 
  signal nx53675z1228 : STD_LOGIC; 
  signal nx53675z1237 : STD_LOGIC; 
  signal nx53675z1234 : STD_LOGIC; 
  signal nx53675z1243 : STD_LOGIC; 
  signal nx53675z1240 : STD_LOGIC; 
  signal nx53675z1249 : STD_LOGIC; 
  signal nx53675z1246 : STD_LOGIC; 
  signal nx53675z1255 : STD_LOGIC; 
  signal nx53675z1252 : STD_LOGIC; 
  signal nx53675z1128 : STD_LOGIC; 
  signal nx53675z1125 : STD_LOGIC; 
  signal nx53675z1134 : STD_LOGIC; 
  signal nx53675z1131 : STD_LOGIC; 
  signal nx53675z1140 : STD_LOGIC; 
  signal nx53675z1137 : STD_LOGIC; 
  signal nx53675z1176 : STD_LOGIC; 
  signal nx53675z1173 : STD_LOGIC; 
  signal nx53675z1182 : STD_LOGIC; 
  signal nx53675z1179 : STD_LOGIC; 
  signal U2_ROMO5_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROMO5_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z964 : STD_LOGIC; 
  signal nx53675z961 : STD_LOGIC; 
  signal nx53675z933 : STD_LOGIC; 
  signal nx53675z930 : STD_LOGIC; 
  signal nx53675z552 : STD_LOGIC; 
  signal nx53675z549 : STD_LOGIC; 
  signal nx53675z558 : STD_LOGIC; 
  signal nx53675z555 : STD_LOGIC; 
  signal nx53675z564 : STD_LOGIC; 
  signal nx53675z561 : STD_LOGIC; 
  signal nx53675z570 : STD_LOGIC; 
  signal nx53675z567 : STD_LOGIC; 
  signal nx53675z576 : STD_LOGIC; 
  signal nx53675z573 : STD_LOGIC; 
  signal nx53675z505 : STD_LOGIC; 
  signal nx53675z502 : STD_LOGIC; 
  signal nx53675z511 : STD_LOGIC; 
  signal nx53675z508 : STD_LOGIC; 
  signal nx53675z1195 : STD_LOGIC; 
  signal nx53675z1192 : STD_LOGIC; 
  signal nx53675z1274 : STD_LOGIC; 
  signal nx53675z1271 : STD_LOGIC; 
  signal nx53675z1280 : STD_LOGIC; 
  signal nx53675z1277 : STD_LOGIC; 
  signal nx53675z1201 : STD_LOGIC; 
  signal nx53675z1198 : STD_LOGIC; 
  signal nx53675z1207 : STD_LOGIC; 
  signal nx53675z1204 : STD_LOGIC; 
  signal nx53675z1213 : STD_LOGIC; 
  signal nx53675z1210 : STD_LOGIC; 
  signal nx53675z1261 : STD_LOGIC; 
  signal nx53675z1258 : STD_LOGIC; 
  signal nx53675z1146 : STD_LOGIC; 
  signal nx53675z1143 : STD_LOGIC; 
  signal nx53675z976 : STD_LOGIC; 
  signal nx53675z973 : STD_LOGIC; 
  signal nx53675z581 : STD_LOGIC; 
  signal nx53675z579 : STD_LOGIC; 
  signal U2_ROMO6_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U2_ROMO6_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx53675z1517 : STD_LOGIC; 
  signal nx53675z1514 : STD_LOGIC; 
  signal nx53675z1268 : STD_LOGIC; 
  signal nx53675z1266 : STD_LOGIC; 
  signal nx53675z1286 : STD_LOGIC; 
  signal nx53675z1283 : STD_LOGIC; 
  signal nx53675z988 : STD_LOGIC; 
  signal nx53675z985 : STD_LOGIC; 
  signal nx53675z1000 : STD_LOGIC; 
  signal nx53675z997 : STD_LOGIC; 
  signal nx54672z21 : STD_LOGIC; 
  signal nx54672z18 : STD_LOGIC; 
  signal nx54672z27 : STD_LOGIC; 
  signal nx54672z24 : STD_LOGIC; 
  signal nx54672z587 : STD_LOGIC; 
  signal nx54672z585 : STD_LOGIC; 
  signal U1_ROME8_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROME8_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z162 : STD_LOGIC; 
  signal nx54672z159 : STD_LOGIC; 
  signal nx54672z670 : STD_LOGIC; 
  signal nx54672z667 : STD_LOGIC; 
  signal nx54672z676 : STD_LOGIC; 
  signal nx54672z673 : STD_LOGIC; 
  signal nx54672z730 : STD_LOGIC; 
  signal nx54672z727 : STD_LOGIC; 
  signal nx54672z736 : STD_LOGIC; 
  signal nx54672z733 : STD_LOGIC; 
  signal nx54672z97 : STD_LOGIC; 
  signal nx54672z94 : STD_LOGIC; 
  signal nx54672z103 : STD_LOGIC; 
  signal nx54672z100 : STD_LOGIC; 
  signal nx54672z109 : STD_LOGIC; 
  signal nx54672z106 : STD_LOGIC; 
  signal nx54672z115 : STD_LOGIC; 
  signal nx54672z112 : STD_LOGIC; 
  signal nx54672z33 : STD_LOGIC; 
  signal nx54672z30 : STD_LOGIC; 
  signal nx54672z39 : STD_LOGIC; 
  signal nx54672z36 : STD_LOGIC; 
  signal nx54672z45 : STD_LOGIC; 
  signal nx54672z42 : STD_LOGIC; 
  signal nx54672z51 : STD_LOGIC; 
  signal nx54672z48 : STD_LOGIC; 
  signal nx54672z57 : STD_LOGIC; 
  signal nx54672z54 : STD_LOGIC; 
  signal U1_ROMO8_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROMO8_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z664 : STD_LOGIC; 
  signal nx54672z662 : STD_LOGIC; 
  signal nx54672z593 : STD_LOGIC; 
  signal nx54672z590 : STD_LOGIC; 
  signal nx54672z599 : STD_LOGIC; 
  signal nx54672z596 : STD_LOGIC; 
  signal nx54672z605 : STD_LOGIC; 
  signal nx54672z602 : STD_LOGIC; 
  signal nx54672z611 : STD_LOGIC; 
  signal nx54672z608 : STD_LOGIC; 
  signal nx54672z617 : STD_LOGIC; 
  signal nx54672z614 : STD_LOGIC; 
  signal nx54672z659 : STD_LOGIC; 
  signal nx54672z656 : STD_LOGIC; 
  signal nx54672z168 : STD_LOGIC; 
  signal nx54672z165 : STD_LOGIC; 
  signal nx54672z174 : STD_LOGIC; 
  signal nx54672z171 : STD_LOGIC; 
  signal nx54672z180 : STD_LOGIC; 
  signal nx54672z177 : STD_LOGIC; 
  signal nx54672z186 : STD_LOGIC; 
  signal nx54672z183 : STD_LOGIC; 
  signal nx54672z191 : STD_LOGIC; 
  signal nx54672z189 : STD_LOGIC; 
  signal nx54672z749 : STD_LOGIC; 
  signal nx54672z746 : STD_LOGIC; 
  signal nx54672z755 : STD_LOGIC; 
  signal nx54672z752 : STD_LOGIC; 
  signal nx54672z132 : STD_LOGIC; 
  signal nx54672z130 : STD_LOGIC; 
  signal nx54672z73 : STD_LOGIC; 
  signal nx54672z70 : STD_LOGIC; 
  signal nx54672z743 : STD_LOGIC; 
  signal nx54672z741 : STD_LOGIC; 
  signal nx54672z809 : STD_LOGIC; 
  signal nx54672z806 : STD_LOGIC; 
  signal nx54672z815 : STD_LOGIC; 
  signal nx54672z812 : STD_LOGIC; 
  signal U1_ROMO2_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROMO2_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z682 : STD_LOGIC; 
  signal nx54672z679 : STD_LOGIC; 
  signal nx54672z688 : STD_LOGIC; 
  signal nx54672z685 : STD_LOGIC; 
  signal nx54672z694 : STD_LOGIC; 
  signal nx54672z691 : STD_LOGIC; 
  signal nx54672z700 : STD_LOGIC; 
  signal nx54672z697 : STD_LOGIC; 
  signal nx54672z706 : STD_LOGIC; 
  signal nx54672z703 : STD_LOGIC; 
  signal U1_ROMO1_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROMO1_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z304 : STD_LOGIC; 
  signal nx54672z301 : STD_LOGIC; 
  signal nx54672z310 : STD_LOGIC; 
  signal nx54672z307 : STD_LOGIC; 
  signal nx54672z67 : STD_LOGIC; 
  signal nx54672z65 : STD_LOGIC; 
  signal nx54672z79 : STD_LOGIC; 
  signal nx54672z76 : STD_LOGIC; 
  signal nx54672z85 : STD_LOGIC; 
  signal nx54672z82 : STD_LOGIC; 
  signal nx54672z121 : STD_LOGIC; 
  signal nx54672z118 : STD_LOGIC; 
  signal nx54672z126 : STD_LOGIC; 
  signal nx54672z124 : STD_LOGIC; 
  signal U1_ROME1_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROME1_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z9 : STD_LOGIC; 
  signal nx54672z6 : STD_LOGIC; 
  signal nx54672z15 : STD_LOGIC; 
  signal nx54672z12 : STD_LOGIC; 
  signal nx54672z62 : STD_LOGIC; 
  signal nx54672z60 : STD_LOGIC; 
  signal nx54672z623 : STD_LOGIC; 
  signal nx54672z620 : STD_LOGIC; 
  signal nx54672z629 : STD_LOGIC; 
  signal nx54672z626 : STD_LOGIC; 
  signal nx54672z635 : STD_LOGIC; 
  signal nx54672z632 : STD_LOGIC; 
  signal nx54672z641 : STD_LOGIC; 
  signal nx54672z638 : STD_LOGIC; 
  signal nx54672z647 : STD_LOGIC; 
  signal nx54672z644 : STD_LOGIC; 
  signal nx54672z3 : STD_LOGIC; 
  signal nx54672z1 : STD_LOGIC; 
  signal nx54672z203 : STD_LOGIC; 
  signal nx54672z200 : STD_LOGIC; 
  signal nx54672z239 : STD_LOGIC; 
  signal nx54672z236 : STD_LOGIC; 
  signal nx54672z251 : STD_LOGIC; 
  signal nx54672z248 : STD_LOGIC; 
  signal U1_ROME3_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROME3_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z197 : STD_LOGIC; 
  signal nx54672z195 : STD_LOGIC; 
  signal nx54672z375 : STD_LOGIC; 
  signal nx54672z372 : STD_LOGIC; 
  signal nx54672z381 : STD_LOGIC; 
  signal nx54672z378 : STD_LOGIC; 
  signal nx54672z1010 : STD_LOGIC; 
  signal nx54672z1007 : STD_LOGIC; 
  signal nx54672z327 : STD_LOGIC; 
  signal nx54672z325 : STD_LOGIC; 
  signal nx54672z138 : STD_LOGIC; 
  signal nx54672z135 : STD_LOGIC; 
  signal nx54672z144 : STD_LOGIC; 
  signal nx54672z141 : STD_LOGIC; 
  signal nx54672z150 : STD_LOGIC; 
  signal nx54672z147 : STD_LOGIC; 
  signal nx54672z156 : STD_LOGIC; 
  signal nx54672z153 : STD_LOGIC; 
  signal U1_ROME2_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROME2_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z943 : STD_LOGIC; 
  signal nx54672z940 : STD_LOGIC; 
  signal nx54672z949 : STD_LOGIC; 
  signal nx54672z946 : STD_LOGIC; 
  signal nx54672z955 : STD_LOGIC; 
  signal nx54672z952 : STD_LOGIC; 
  signal nx54672z828 : STD_LOGIC; 
  signal nx54672z825 : STD_LOGIC; 
  signal nx54672z840 : STD_LOGIC; 
  signal nx54672z837 : STD_LOGIC; 
  signal nx54672z876 : STD_LOGIC; 
  signal nx54672z873 : STD_LOGIC; 
  signal nx54672z888 : STD_LOGIC; 
  signal nx54672z885 : STD_LOGIC; 
  signal U1_ROMO3_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROMO3_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z761 : STD_LOGIC; 
  signal nx54672z758 : STD_LOGIC; 
  signal nx54672z767 : STD_LOGIC; 
  signal nx54672z764 : STD_LOGIC; 
  signal nx54672z773 : STD_LOGIC; 
  signal nx54672z770 : STD_LOGIC; 
  signal nx54672z779 : STD_LOGIC; 
  signal nx54672z776 : STD_LOGIC; 
  signal nx54672z785 : STD_LOGIC; 
  signal nx54672z782 : STD_LOGIC; 
  signal nx54672z901 : STD_LOGIC; 
  signal nx54672z899 : STD_LOGIC; 
  signal nx54672z822 : STD_LOGIC; 
  signal nx54672z820 : STD_LOGIC; 
  signal nx54672z712 : STD_LOGIC; 
  signal nx54672z709 : STD_LOGIC; 
  signal nx54672z718 : STD_LOGIC; 
  signal nx54672z715 : STD_LOGIC; 
  signal nx54672z724 : STD_LOGIC; 
  signal nx54672z721 : STD_LOGIC; 
  signal nx54672z392 : STD_LOGIC; 
  signal nx54672z390 : STD_LOGIC; 
  signal nx54672z268 : STD_LOGIC; 
  signal nx54672z265 : STD_LOGIC; 
  signal nx54672z274 : STD_LOGIC; 
  signal nx54672z271 : STD_LOGIC; 
  signal nx54672z280 : STD_LOGIC; 
  signal nx54672z277 : STD_LOGIC; 
  signal nx54672z316 : STD_LOGIC; 
  signal nx54672z313 : STD_LOGIC; 
  signal nx54672z321 : STD_LOGIC; 
  signal nx54672z319 : STD_LOGIC; 
  signal U1_ROME4_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROME4_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z91 : STD_LOGIC; 
  signal nx54672z88 : STD_LOGIC; 
  signal nx54672z653 : STD_LOGIC; 
  signal nx54672z650 : STD_LOGIC; 
  signal nx54672z398 : STD_LOGIC; 
  signal nx54672z395 : STD_LOGIC; 
  signal nx54672z446 : STD_LOGIC; 
  signal nx54672z443 : STD_LOGIC; 
  signal nx54672z451 : STD_LOGIC; 
  signal nx54672z449 : STD_LOGIC; 
  signal U1_ROME6_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROME6_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z215 : STD_LOGIC; 
  signal nx54672z212 : STD_LOGIC; 
  signal nx54672z227 : STD_LOGIC; 
  signal nx54672z224 : STD_LOGIC; 
  signal nx54672z333 : STD_LOGIC; 
  signal nx54672z330 : STD_LOGIC; 
  signal nx54672z339 : STD_LOGIC; 
  signal nx54672z336 : STD_LOGIC; 
  signal nx54672z345 : STD_LOGIC; 
  signal nx54672z342 : STD_LOGIC; 
  signal nx54672z351 : STD_LOGIC; 
  signal nx54672z348 : STD_LOGIC; 
  signal nx54672z386 : STD_LOGIC; 
  signal nx54672z384 : STD_LOGIC; 
  signal U1_ROME5_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROME5_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z1083 : STD_LOGIC; 
  signal nx54672z1080 : STD_LOGIC; 
  signal nx54672z1089 : STD_LOGIC; 
  signal nx54672z1086 : STD_LOGIC; 
  signal nx54672z1095 : STD_LOGIC; 
  signal nx54672z1092 : STD_LOGIC; 
  signal nx54672z1016 : STD_LOGIC; 
  signal nx54672z1013 : STD_LOGIC; 
  signal nx54672z1022 : STD_LOGIC; 
  signal nx54672z1019 : STD_LOGIC; 
  signal nx54672z1028 : STD_LOGIC; 
  signal nx54672z1025 : STD_LOGIC; 
  signal nx54672z1034 : STD_LOGIC; 
  signal nx54672z1031 : STD_LOGIC; 
  signal nx54672z1040 : STD_LOGIC; 
  signal nx54672z1037 : STD_LOGIC; 
  signal nx54672z980 : STD_LOGIC; 
  signal nx54672z978 : STD_LOGIC; 
  signal nx54672z907 : STD_LOGIC; 
  signal nx54672z904 : STD_LOGIC; 
  signal nx54672z919 : STD_LOGIC; 
  signal nx54672z916 : STD_LOGIC; 
  signal nx54672z925 : STD_LOGIC; 
  signal nx54672z922 : STD_LOGIC; 
  signal nx54672z961 : STD_LOGIC; 
  signal nx54672z958 : STD_LOGIC; 
  signal nx54672z967 : STD_LOGIC; 
  signal nx54672z964 : STD_LOGIC; 
  signal nx54672z973 : STD_LOGIC; 
  signal nx54672z970 : STD_LOGIC; 
  signal U1_ROMO4_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROMO4_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z852 : STD_LOGIC; 
  signal nx54672z849 : STD_LOGIC; 
  signal nx54672z864 : STD_LOGIC; 
  signal nx54672z861 : STD_LOGIC; 
  signal nx54672z791 : STD_LOGIC; 
  signal nx54672z788 : STD_LOGIC; 
  signal nx54672z797 : STD_LOGIC; 
  signal nx54672z794 : STD_LOGIC; 
  signal nx54672z463 : STD_LOGIC; 
  signal nx54672z460 : STD_LOGIC; 
  signal nx54672z469 : STD_LOGIC; 
  signal nx54672z466 : STD_LOGIC; 
  signal nx54672z516 : STD_LOGIC; 
  signal nx54672z514 : STD_LOGIC; 
  signal U1_ROME7_modgen_rom_ix2_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROME7_modgen_rom_ix2_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z1150 : STD_LOGIC; 
  signal nx54672z1147 : STD_LOGIC; 
  signal nx54672z1156 : STD_LOGIC; 
  signal nx54672z1153 : STD_LOGIC; 
  signal nx54672z834 : STD_LOGIC; 
  signal nx54672z831 : STD_LOGIC; 
  signal nx54672z803 : STD_LOGIC; 
  signal nx54672z800 : STD_LOGIC; 
  signal nx54672z286 : STD_LOGIC; 
  signal nx54672z283 : STD_LOGIC; 
  signal nx54672z292 : STD_LOGIC; 
  signal nx54672z289 : STD_LOGIC; 
  signal nx54672z298 : STD_LOGIC; 
  signal nx54672z295 : STD_LOGIC; 
  signal nx54672z209 : STD_LOGIC; 
  signal nx54672z206 : STD_LOGIC; 
  signal nx54672z233 : STD_LOGIC; 
  signal nx54672z230 : STD_LOGIC; 
  signal nx54672z457 : STD_LOGIC; 
  signal nx54672z455 : STD_LOGIC; 
  signal nx54672z404 : STD_LOGIC; 
  signal nx54672z401 : STD_LOGIC; 
  signal nx54672z410 : STD_LOGIC; 
  signal nx54672z407 : STD_LOGIC; 
  signal nx54672z416 : STD_LOGIC; 
  signal nx54672z413 : STD_LOGIC; 
  signal nx54672z422 : STD_LOGIC; 
  signal nx54672z419 : STD_LOGIC; 
  signal nx54672z428 : STD_LOGIC; 
  signal nx54672z425 : STD_LOGIC; 
  signal nx54672z528 : STD_LOGIC; 
  signal nx54672z525 : STD_LOGIC; 
  signal nx54672z534 : STD_LOGIC; 
  signal nx54672z531 : STD_LOGIC; 
  signal nx54672z540 : STD_LOGIC; 
  signal nx54672z537 : STD_LOGIC; 
  signal nx54672z546 : STD_LOGIC; 
  signal nx54672z543 : STD_LOGIC; 
  signal nx54672z262 : STD_LOGIC; 
  signal nx54672z260 : STD_LOGIC; 
  signal nx54672z522 : STD_LOGIC; 
  signal nx54672z520 : STD_LOGIC; 
  signal nx54672z357 : STD_LOGIC; 
  signal nx54672z354 : STD_LOGIC; 
  signal nx54672z363 : STD_LOGIC; 
  signal nx54672z360 : STD_LOGIC; 
  signal nx54672z369 : STD_LOGIC; 
  signal nx54672z366 : STD_LOGIC; 
  signal nx54672z1065 : STD_LOGIC; 
  signal nx54672z1062 : STD_LOGIC; 
  signal nx54672z1101 : STD_LOGIC; 
  signal nx54672z1098 : STD_LOGIC; 
  signal nx54672z1107 : STD_LOGIC; 
  signal nx54672z1104 : STD_LOGIC; 
  signal nx54672z1113 : STD_LOGIC; 
  signal nx54672z1110 : STD_LOGIC; 
  signal nx54672z1119 : STD_LOGIC; 
  signal nx54672z1116 : STD_LOGIC; 
  signal nx54672z1125 : STD_LOGIC; 
  signal nx54672z1122 : STD_LOGIC; 
  signal nx54672z986 : STD_LOGIC; 
  signal nx54672z983 : STD_LOGIC; 
  signal nx54672z992 : STD_LOGIC; 
  signal nx54672z989 : STD_LOGIC; 
  signal nx54672z998 : STD_LOGIC; 
  signal nx54672z995 : STD_LOGIC; 
  signal nx54672z1004 : STD_LOGIC; 
  signal nx54672z1001 : STD_LOGIC; 
  signal nx54672z1046 : STD_LOGIC; 
  signal nx54672z1043 : STD_LOGIC; 
  signal nx54672z1052 : STD_LOGIC; 
  signal nx54672z1049 : STD_LOGIC; 
  signal nx54672z1223 : STD_LOGIC; 
  signal nx54672z1220 : STD_LOGIC; 
  signal nx54672z1229 : STD_LOGIC; 
  signal nx54672z1226 : STD_LOGIC; 
  signal nx54672z1059 : STD_LOGIC; 
  signal nx54672z1057 : STD_LOGIC; 
  signal U1_ROMO5_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROMO5_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z931 : STD_LOGIC; 
  signal nx54672z928 : STD_LOGIC; 
  signal nx54672z937 : STD_LOGIC; 
  signal nx54672z934 : STD_LOGIC; 
  signal nx54672z475 : STD_LOGIC; 
  signal nx54672z472 : STD_LOGIC; 
  signal nx54672z481 : STD_LOGIC; 
  signal nx54672z478 : STD_LOGIC; 
  signal nx54672z487 : STD_LOGIC; 
  signal nx54672z484 : STD_LOGIC; 
  signal nx54672z493 : STD_LOGIC; 
  signal nx54672z490 : STD_LOGIC; 
  signal nx54672z499 : STD_LOGIC; 
  signal nx54672z496 : STD_LOGIC; 
  signal nx54672z1235 : STD_LOGIC; 
  signal nx54672z1232 : STD_LOGIC; 
  signal nx54672z1241 : STD_LOGIC; 
  signal nx54672z1238 : STD_LOGIC; 
  signal nx54672z1162 : STD_LOGIC; 
  signal nx54672z1159 : STD_LOGIC; 
  signal nx54672z1168 : STD_LOGIC; 
  signal nx54672z1165 : STD_LOGIC; 
  signal nx54672z1174 : STD_LOGIC; 
  signal nx54672z1171 : STD_LOGIC; 
  signal nx54672z1180 : STD_LOGIC; 
  signal nx54672z1177 : STD_LOGIC; 
  signal nx54672z1186 : STD_LOGIC; 
  signal nx54672z1183 : STD_LOGIC; 
  signal nx54672z846 : STD_LOGIC; 
  signal nx54672z843 : STD_LOGIC; 
  signal nx54672z870 : STD_LOGIC; 
  signal nx54672z867 : STD_LOGIC; 
  signal nx54672z221 : STD_LOGIC; 
  signal nx54672z218 : STD_LOGIC; 
  signal nx54672z245 : STD_LOGIC; 
  signal nx54672z242 : STD_LOGIC; 
  signal nx54672z256 : STD_LOGIC; 
  signal nx54672z254 : STD_LOGIC; 
  signal nx54672z434 : STD_LOGIC; 
  signal nx54672z431 : STD_LOGIC; 
  signal nx54672z440 : STD_LOGIC; 
  signal nx54672z437 : STD_LOGIC; 
  signal nx54672z552 : STD_LOGIC; 
  signal nx54672z549 : STD_LOGIC; 
  signal nx54672z558 : STD_LOGIC; 
  signal nx54672z555 : STD_LOGIC; 
  signal nx54672z564 : STD_LOGIC; 
  signal nx54672z561 : STD_LOGIC; 
  signal nx54672z570 : STD_LOGIC; 
  signal nx54672z567 : STD_LOGIC; 
  signal nx54672z576 : STD_LOGIC; 
  signal nx54672z573 : STD_LOGIC; 
  signal nx54672z1071 : STD_LOGIC; 
  signal nx54672z1068 : STD_LOGIC; 
  signal nx54672z1077 : STD_LOGIC; 
  signal nx54672z1074 : STD_LOGIC; 
  signal nx54672z1131 : STD_LOGIC; 
  signal nx54672z1128 : STD_LOGIC; 
  signal nx54672z505 : STD_LOGIC; 
  signal nx54672z502 : STD_LOGIC; 
  signal nx54672z511 : STD_LOGIC; 
  signal nx54672z508 : STD_LOGIC; 
  signal nx54672z1247 : STD_LOGIC; 
  signal nx54672z1244 : STD_LOGIC; 
  signal nx54672z1253 : STD_LOGIC; 
  signal nx54672z1250 : STD_LOGIC; 
  signal nx54672z1259 : STD_LOGIC; 
  signal nx54672z1256 : STD_LOGIC; 
  signal nx54672z1265 : STD_LOGIC; 
  signal nx54672z1262 : STD_LOGIC; 
  signal nx54672z1271 : STD_LOGIC; 
  signal nx54672z1268 : STD_LOGIC; 
  signal nx54672z1138 : STD_LOGIC; 
  signal nx54672z1136 : STD_LOGIC; 
  signal nx54672z1144 : STD_LOGIC; 
  signal nx54672z1141 : STD_LOGIC; 
  signal nx54672z1192 : STD_LOGIC; 
  signal nx54672z1189 : STD_LOGIC; 
  signal nx54672z1198 : STD_LOGIC; 
  signal nx54672z1195 : STD_LOGIC; 
  signal nx54672z1204 : STD_LOGIC; 
  signal nx54672z1201 : STD_LOGIC; 
  signal nx54672z1210 : STD_LOGIC; 
  signal nx54672z1207 : STD_LOGIC; 
  signal U1_ROMO7_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROMO7_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal U1_ROMO6_modgen_rom_ix0_nx_ro64_32_l : STD_LOGIC; 
  signal U1_ROMO6_modgen_rom_ix0_nx_ro64_32_u : STD_LOGIC; 
  signal nx54672z913 : STD_LOGIC; 
  signal nx54672z910 : STD_LOGIC; 
  signal nx54672z858 : STD_LOGIC; 
  signal nx54672z855 : STD_LOGIC; 
  signal nx54672z882 : STD_LOGIC; 
  signal nx54672z879 : STD_LOGIC; 
  signal nx54672z894 : STD_LOGIC; 
  signal nx54672z891 : STD_LOGIC; 
  signal nx54672z581 : STD_LOGIC; 
  signal nx54672z579 : STD_LOGIC; 
  signal nx54672z1217 : STD_LOGIC; 
  signal nx54672z1215 : STD_LOGIC; 
  signal nx54672z1277 : STD_LOGIC; 
  signal nx54672z1274 : STD_LOGIC; 
  signal nx54672z1283 : STD_LOGIC; 
  signal nx54672z1280 : STD_LOGIC; 
  signal nx54672z1289 : STD_LOGIC; 
  signal nx54672z1286 : STD_LOGIC; 
  signal clk_ibuf_IBUFG : STD_LOGIC; 
  signal idv_int : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1854 : STD_LOGIC; 
  signal U_DCT1D_NOT_rtlcs2 : STD_LOGIC; 
  signal U_DCT1D_rtlc2n465 : STD_LOGIC; 
  signal U_DCT1D_rtlcn339 : STD_LOGIC; 
  signal nx1552z1 : STD_LOGIC; 
  signal nx21201z1 : STD_LOGIC; 
  signal U_DBUFCTL_mem1_lock_reg : STD_LOGIC; 
  signal memswitchwr_s : STD_LOGIC; 
  signal releasewr_s : STD_LOGIC; 
  signal U_DBUFCTL_rtlcn38 : STD_LOGIC; 
  signal requestwr_s : STD_LOGIC; 
  signal requestrd_s : STD_LOGIC; 
  signal U_DBUFCTL_mem1_full_reg : STD_LOGIC; 
  signal U_DBUFCTL_rtlc4n377 : STD_LOGIC; 
  signal reqrdfail_s : STD_LOGIC; 
  signal U_DCT2D_NOT_rtlcs2 : STD_LOGIC; 
  signal U_DCT2D_rtlc2n584 : STD_LOGIC; 
  signal U_DCT2D_completed_reg : STD_LOGIC; 
  signal U_DBUFCTL_rtlc4n374 : STD_LOGIC; 
  signal NOT_U_DBUFCTL_rtlc0n25 : STD_LOGIC; 
  signal memswitchrd_s : STD_LOGIC; 
  signal U_DCT2D_rtlc2n446 : STD_LOGIC; 
  signal U_DBUFCTL_rtlc4n373 : STD_LOGIC; 
  signal U_DBUFCTL_mem2_full_reg : STD_LOGIC; 
  signal U_DBUFCTL_mem2_lock_reg : STD_LOGIC; 
  signal U_DBUFCTL_rtlcn1 : STD_LOGIC; 
  signal U_DBUFCTL_rtlc4n202 : STD_LOGIC; 
  signal nx24581z1 : STD_LOGIC; 
  signal releaserd_s : STD_LOGIC; 
  signal ramwe_s : STD_LOGIC; 
  signal nx43562z1 : STD_LOGIC; 
  signal U_DBUFCTL_rtlcn42 : STD_LOGIC; 
  signal U_DBUFCTL_rtlc4n378 : STD_LOGIC; 
  signal U_DCT1D_ready : STD_LOGIC; 
  signal reqwrfail_s : STD_LOGIC; 
  signal U_DCT1D_NOT_rtlcs1 : STD_LOGIC; 
  signal U_DCT1D_rtlcn1047 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1768 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1612 : STD_LOGIC; 
  signal U_DCT2D_NOT_rtlc2n488 : STD_LOGIC; 
  signal U_DCT2D_nx49413z1 : STD_LOGIC; 
  signal U_DCT2D_rtlc2n576 : STD_LOGIC; 
  signal U_DCT2D_nx39898z2 : STD_LOGIC; 
  signal U_DCT2D_nx40895z2 : STD_LOGIC; 
  signal U_DCT1D_rtlc2n471 : STD_LOGIC; 
  signal U_DCT1D_completed_reg : STD_LOGIC; 
  signal U_DCT1D_rtlc2n365 : STD_LOGIC; 
  signal U_DCT1D_rtlc2n469 : STD_LOGIC; 
  signal nx43562z2 : STD_LOGIC; 
  signal nx53675z1582 : STD_LOGIC; 
  signal U_DCT2D_latch_done_reg : STD_LOGIC; 
  signal U_DCT2D_rtlcn1678 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1690 : STD_LOGIC; 
  signal U_DCT1D_NOT_rtlcs7 : STD_LOGIC; 
  signal U_DCT2D_rtlc2n581 : STD_LOGIC; 
  signal U_DCT2D_rtlcs5 : STD_LOGIC; 
  signal U_DCT2D_rtlcn65 : STD_LOGIC; 
  signal U_DCT2D_rtlc2n582 : STD_LOGIC; 
  signal U_DCT2D_nx6411z1 : STD_LOGIC; 
  signal U_DCT2D_rtlc2n580 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1685 : STD_LOGIC; 
  signal U_DCT2D_rtlc2n579 : STD_LOGIC; 
  signal U_DCT2D_nx41892z3 : STD_LOGIC; 
  signal U_DCT2D_nx41892z2 : STD_LOGIC; 
  signal U_DCT2D_NOT_rtlcs7 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1311 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1684 : STD_LOGIC; 
  signal U_DCT1D_rtlc2n293 : STD_LOGIC; 
  signal U_DCT1D_nx7599z1 : STD_LOGIC; 
  signal U_DCT1D_rtlc2n468 : STD_LOGIC; 
  signal U_DCT1D_latch_done_reg : STD_LOGIC; 
  signal U_DCT1D_rtlcs3 : STD_LOGIC; 
  signal U_DCT1D_nx2819z1 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_0 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_1 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_2 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_3 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_4 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_5 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_6 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_7 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_8 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_9 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_10 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_11 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_12 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_13 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_14 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_15 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_16 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_17 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_18 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_19 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_20 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_21 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_22 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_23 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_24 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_25 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_26 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_27 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_28 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_29 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_30 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_31 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_32 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_33 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_34 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_35 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_36 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_37 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_38 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_39 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_40 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_41 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_42 : STD_LOGIC; 
  signal GLOBAL_LOGIC1_43 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_0 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_1 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_2 : STD_LOGIC; 
  signal GLOBAL_LOGIC0_3 : STD_LOGIC; 
  signal GSR : STD_LOGIC; 
  signal GTS : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_CY0F : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59822z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_XORG : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1421_add_10_ix60819z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx60819z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx61816z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1421_add_10_ix62813z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx62813z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx63810z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1421_add_10_ix64807z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx64807z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx268z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1421_add_10_ix1265z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx1265z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_8_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_8_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_8_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx2262z1_rt : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_8_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_CY0F : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx59822z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_XORG : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1580_add_47_ix60819z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx60819z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx61816z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1580_add_47_ix62813z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx62813z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx63810z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1580_add_47_ix64807z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx64807z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx268z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1580_add_47_ix1265z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx1265z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx2262z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1580_add_47_ix3259z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx3259z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_10_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx22763z1_rt : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_10_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_CY0F : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx49552z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_XORG : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_97_sub_41_ix50549z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx50549z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx51546z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_97_sub_41_ix52543z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx52543z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx53540z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_97_sub_41_ix54537z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx54537z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx55534z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_97_sub_41_ix56531z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx56531z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx57528z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_97_sub_41_ix58525z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx58525z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_10_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx7189z1_rt : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_10_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_CY0F : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx34147z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_XORG : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_100_sub_44_ix35144z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx35144z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx36141z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_100_sub_44_ix37138z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx37138z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx38135z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_100_sub_44_ix39132z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx39132z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx40129z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_100_sub_44_ix41126z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx41126z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx42123z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_100_sub_44_ix43120z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx43120z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_10_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx16172z1_rt : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_10_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_CY0F : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx64957z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_XORG : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1420_add_9_ix418z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx418z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx1415z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1420_add_9_ix2412z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx2412z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx3409z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1420_add_9_ix4406z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx4406z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx5403z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1420_add_9_ix6400z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx6400z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_8_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_8_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_8_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx7397z1_rt : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_8_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_10_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_10_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_10_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z651 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_10_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_10_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64239_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_10_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_10_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z648 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_12_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_12_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_12_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z645 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_12_XORG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64231_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_12_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_12_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_12_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_12_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_12_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_12_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_12_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_12_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z642 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_14_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_14_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_14_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z639 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_14_XORG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64223_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_14_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_14_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_14_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_14_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_14_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_14_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_14_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_14_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z636 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_16_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_16_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_16_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z633 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_16_XORG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64215_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_16_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_16_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_16_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_16_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_16_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_16_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_16_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_16_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z630 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_18_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_18_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_18_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z627 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_18_XORG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64207_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_18_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_18_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_18_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_18_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_18_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_18_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_18_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_18_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z624 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_20_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_20_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_20_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z621 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_20_XORG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64199_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_20_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_20_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_20_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_20_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_20_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_20_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_20_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_20_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z618 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_22_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_22_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_22_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_22_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z615 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1501_22_XORG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64191_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z571_rt : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_9_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_9_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_9_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z613 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_9_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z612 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_9_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_9_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_9_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64188_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_9_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z610 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_9_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z609 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_11_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_11_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_11_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z606 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_11_XORG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64182_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_11_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_11_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_11_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_11_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z603 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_0_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_13_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_13_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_13_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z600 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_13_XORG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64176_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_13_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_13_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_13_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_13_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z597 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_15_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_15_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_15_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z594 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_15_XORG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64170_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_15_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_15_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_15_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_15_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_15_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_15_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_15_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_15_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z591 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_17_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_17_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_17_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z588 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_17_XORG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64164_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_17_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_17_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_17_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_17_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_17_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_17_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_17_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_17_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z585 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_19_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_19_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_19_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z582 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_19_XORG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64158_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_19_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_19_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_19_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_19_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_19_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_19_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_19_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_19_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z579 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_21_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_21_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_21_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z577 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_21_XORG : STD_LOGIC; 
  signal U_DCT2D_ix65206z64153_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_21_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_21_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_21_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_21_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_21_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_21_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_21_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_21_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z575 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_23_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1484_23_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z572_rt : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_CY0F : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx64957z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_XORG : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1579_add_46_ix418z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx418z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx1415z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1579_add_46_ix2412z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx2412z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_2_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx3409z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1579_add_46_ix4406z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx4406z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx5403z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1579_add_46_ix6400z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx6400z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_6_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx7397z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1579_add_46_ix8394z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx8394z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_10_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx30550z1_rt : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_10_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_CY0F : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx49552z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_XORG : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_83_sub_4_ix50549z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx50549z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx51546z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_83_sub_4_ix52543z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx52543z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx53540z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_83_sub_4_ix54537z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx54537z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx55534z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_83_sub_4_ix56531z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx56531z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_8_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_8_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_8_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx57528z1_rt : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_8_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_2_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_2_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_2_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z120 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_2_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_2_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_2_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63485_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_2_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_2_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z117 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_3_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_3_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_3_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z114 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_3_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63478_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_3_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_3_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_3_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_3_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_3_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_3_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_3_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_3_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z111 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_5_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_5_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_5_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z108 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_5_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63471_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_5_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_5_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_5_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_5_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_5_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_5_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_5_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_5_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z105 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_7_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_7_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_7_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z102 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_7_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63463_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_7_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_7_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_7_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_7_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_7_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_7_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_7_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_7_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z99 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_9_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_9_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_9_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z96 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_9_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63456_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_9_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_9_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_9_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_9_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z93 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_11_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_11_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_11_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z90 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_11_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63449_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_11_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_11_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_11_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_11_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z87 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_13_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_13_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_13_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z84 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_13_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_331_add_54_ix65206z63442_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_13_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_13_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_13_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_13_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z81 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_15_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1480_15_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z79_rt : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_CY0F : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx34147z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_XORG : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_86_sub_7_ix35144z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx35144z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx36141z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_86_sub_7_ix37138z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx37138z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx38135z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_86_sub_7_ix39132z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx39132z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx40129z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_86_sub_7_ix41126z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx41126z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_8_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_8_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_8_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx42123z1_rt : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_8_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_CY0F : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx60980z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_XORG : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1578_add_45_ix59983z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx59983z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx58986z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1578_add_45_ix57989z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx57989z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx56992z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1578_add_45_ix55995z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx55995z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx54998z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1578_add_45_ix54001z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx54001z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx53004z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1578_add_45_ix52007z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx52007z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_10_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx38337z1_rt : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_10_CEINV : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z209 : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63608_O_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63612_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z207 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_4_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_4_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_4_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z204 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_4_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63603_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_4_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_4_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_4_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_4_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z201 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_6_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_6_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_6_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z198 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_6_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63592_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_6_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_6_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_6_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_6_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z195 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_8_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_8_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_8_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z192 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_8_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63582_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_8_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_8_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_8_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_8_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z189 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_10_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_10_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z186 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_10_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63572_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_10_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_10_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_10_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_10_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_10_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_10_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_10_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_10_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z183 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_12_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_12_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_12_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z180 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_12_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63561_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_12_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_12_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_12_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_12_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_12_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_12_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_12_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_12_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z177 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_14_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_14_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_14_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z174 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_14_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63551_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_14_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_14_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_14_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_14_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_14_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_14_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_14_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_14_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z171 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_16_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_16_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_16_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z168 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_16_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_336_add_56_ix65206z63542_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_16_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_16_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_16_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_16_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_16_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_16_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_16_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_16_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z165 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_18_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1485_18_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z78_rt : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_7_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_7_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_7_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_7_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z294 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_7_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_7_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_7_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63745_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_7_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_7_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z291 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_9_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_9_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_9_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z288 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_9_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63738_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_9_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_9_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_9_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_9_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z285 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_11_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_11_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_11_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z282 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_11_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63731_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_11_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_11_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_11_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_11_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z279 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_13_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_13_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_13_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z276 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_13_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63724_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_13_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_13_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_13_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_13_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z273 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_15_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_15_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_15_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z270 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_15_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63717_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_15_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_15_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_15_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_15_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_15_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_15_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_15_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_15_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z267 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_17_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_17_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_17_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z264 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_17_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63710_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_17_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_17_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_17_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_17_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_17_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_17_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_17_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_17_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z261 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_19_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_19_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_19_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z258 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_19_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_340_add_58_ix65206z63703_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_19_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_19_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_19_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_19_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_19_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_19_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_19_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_19_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z255 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_21_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1483_21_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z253_rt : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_CY0F : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx54687z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_XORG : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1581_add_48_ix55684z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx55684z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx56681z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1581_add_48_ix57678z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx57678z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx58675z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1581_add_48_ix59672z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx59672z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx60669z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1581_add_48_ix61666z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx61666z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx62663z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_1581_add_48_ix63660z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx63660z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_10_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx14976z1_rt : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_10_CEINV : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_5_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_5_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_5_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_5_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z40 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_5_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_5_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_5_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc_389_add_65_ix65206z63386_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_5_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_5_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z37 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_7_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_7_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_7_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z34 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_7_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_389_add_65_ix65206z63379_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_7_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_7_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_7_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_7_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_7_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_7_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_7_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_7_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z31 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_9_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_9_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_9_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z28 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_9_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_389_add_65_ix65206z63372_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_9_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_9_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_9_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_9_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z25 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_11_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_11_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_11_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z22 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_11_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_389_add_65_ix65206z63365_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_11_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_11_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_11_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_11_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z19 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_13_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_13_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_13_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z16 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_13_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_389_add_65_ix65206z63358_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_13_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_13_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_13_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_13_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z13 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_15_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_15_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_15_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z10 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_15_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_389_add_65_ix65206z63351_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_15_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_15_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_15_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_15_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_15_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_15_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_15_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_15_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z7 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_17_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1493_17_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z5_rt : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_6_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_6_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_6_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z432 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_6_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z431 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_6_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_6_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_6_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63921_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_6_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_6_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z427 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_8_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_8_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_8_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z423 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_8_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63910_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_8_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_8_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_8_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_8_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z419 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_10_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_10_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_10_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z415 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_10_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63898_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_10_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_10_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_10_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_10_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_10_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_10_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_10_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_10_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z411 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_12_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_12_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_12_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z407 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_12_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63886_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_12_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_12_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_12_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_12_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_12_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_12_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_12_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_12_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z403 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_14_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_14_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_14_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z399 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_14_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63874_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_14_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_14_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_14_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_14_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_14_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_14_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_14_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_14_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z395 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_16_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_16_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_16_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z391 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_16_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63862_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_16_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_16_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_16_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_16_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_16_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_16_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_16_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_16_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z387 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_18_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_18_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_18_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z383 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_18_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63851_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_18_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_18_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_18_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_18_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_18_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_18_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_18_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_18_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z380 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_20_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_20_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_20_CY0F : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_20_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z377 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1359_20_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_522_add_32_ix59700z63841_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z252 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_2_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_CY0F : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx39282z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_XORG : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_99_sub_43_ix40279z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx40279z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx41276z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_99_sub_43_ix42273z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx42273z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx43270z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_99_sub_43_ix44267z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx44267z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx45264z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_99_sub_43_ix46261z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx46261z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx47258z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_99_sub_43_ix48255z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx48255z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_10_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx8385z1_rt : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_10_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_CY0F : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx60980z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_XORG : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1419_add_8_ix59983z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59983z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx58986z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1419_add_8_ix57989z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx57989z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx56992z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1419_add_8_ix55995z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx55995z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx54998z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1419_add_8_ix54001z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx54001z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_8_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_8_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_8_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx53004z1_rt : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_8_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_8_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_CY0F : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx44417z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_XORG : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_84_sub_5_ix45414z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx45414z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_0_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx46411z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_84_sub_5_ix47408z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx47408z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx48405z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_84_sub_5_ix49402z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx49402z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx50399z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_84_sub_5_ix51396z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx51396z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_8_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_8_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_8_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx52393z1_rt : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_8_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_CY0F : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx44417z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_XORG : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_98_sub_42_ix45414z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx45414z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx46411z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_98_sub_42_ix47408z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx47408z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx48405z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_98_sub_42_ix49402z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx49402z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx50399z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_98_sub_42_ix51396z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx51396z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_CYINIT : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx52393z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_DYMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5_98_sub_42_ix53390z63342_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_CYSELF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_CYAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_CY0G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx53390z1 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_SRINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_10_XORF : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx64938z1_rt : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_10_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_CY0F : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx54687z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_XORG : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1422_add_11_ix55684z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx55684z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx56681z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1422_add_11_ix57678z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx57678z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx58675z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1422_add_11_ix59672z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59672z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx60669z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_1422_add_11_ix61666z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx61666z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_8_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_8_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_8_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx62663z1_rt : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_8_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_8_CEINV : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_4_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_4_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_4_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z77 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_4_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_4_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_4_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc_387_add_64_ix65206z63433_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_4_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_4_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z74 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_5_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_5_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_5_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z71 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_5_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_387_add_64_ix65206z63426_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_5_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_5_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_5_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_5_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_5_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_5_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_5_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_5_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z68 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_7_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_7_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_7_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z65 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_7_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_387_add_64_ix65206z63419_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_7_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_7_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_7_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_7_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_7_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_7_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_7_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_7_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z62 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_9_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_9_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_9_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z59 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_9_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_387_add_64_ix65206z63412_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_9_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_9_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_9_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_9_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z56 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_11_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_11_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_11_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z53 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_11_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_387_add_64_ix65206z63405_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_11_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_11_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_11_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_11_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z50 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_13_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_13_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_13_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z47 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_13_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_387_add_64_ix65206z63398_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_13_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_13_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_13_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_13_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z44 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_15_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1492_15_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z42_rt : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_9_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_9_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_9_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_9_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z369 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_9_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_9_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_9_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc_396_add_68_ix65206z63835_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_9_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_9_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z366 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_11_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_11_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_11_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z363 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_11_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_396_add_68_ix65206z63828_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_11_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_11_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_11_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_11_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z360 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_13_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_13_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_13_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z357 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_13_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_396_add_68_ix65206z63821_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_13_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_13_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_13_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_13_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z354 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_15_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_15_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_15_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z351 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_15_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_396_add_68_ix65206z63814_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_15_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_15_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_15_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_15_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_15_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_15_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_15_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_15_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z348 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_17_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_17_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_17_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z345 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_17_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_396_add_68_ix65206z63807_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_17_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_17_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_17_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_17_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_17_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_17_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_17_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_17_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z342 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_19_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_19_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_19_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z339 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_19_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_396_add_68_ix65206z63800_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_19_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_19_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_19_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_19_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_19_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_19_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_19_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_19_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z336 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_21_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1495_21_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z334_rt : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_CY0F : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx39282z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_XORG : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_85_sub_6_ix40279z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx40279z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx41276z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_85_sub_6_ix42273z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx42273z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx43270z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_85_sub_6_ix44267z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx44267z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_CYINIT : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx45264z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_DYMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5_85_sub_6_ix46261z63342_O : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_CYSELF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_CYAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_CY0G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx46261z1 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_SRINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_8_DXMUX : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_8_XORF : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_8_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx47258z1_rt : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_8_CLKINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_8_CEINV : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_3_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_3_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_3_CY0F : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_3_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z162 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_3_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_3_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_3_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63535_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_3_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_3_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z159 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_5_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_5_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_5_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z156 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_5_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63528_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_5_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_5_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_5_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_5_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_5_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_5_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_5_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_5_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z153 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_7_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_7_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_7_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z150 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_7_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63521_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_7_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_7_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_7_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_7_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_7_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_7_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_7_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_7_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z147 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_9_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_9_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_9_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z144 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_9_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63514_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_9_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_9_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_9_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_9_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z141 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_11_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_11_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_11_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z138 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_11_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63506_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_11_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_11_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_11_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_11_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z135 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_13_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_13_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_13_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z132 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_13_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63499_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_13_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_13_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_13_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_13_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z129 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_15_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_15_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_15_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z126 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_15_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_493_add_21_ix59700z63492_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_15_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_15_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_15_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_15_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_15_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_15_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_15_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_15_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z123 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_17_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1345_17_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z121_rt : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z569 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64139_O_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64143_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z566 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z563 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64131_O_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z560 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_8_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_8_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_8_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z556 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_8_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64124_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_8_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_8_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_8_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_8_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z552 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_10_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_10_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z548 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_10_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64113_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_10_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_10_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_10_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_10_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_10_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_10_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_10_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_10_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z544 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_12_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_12_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_12_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z540 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_12_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64103_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_12_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_12_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_12_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_12_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_12_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_12_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_12_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_12_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z536 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_14_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_14_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_14_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z532 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_14_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64092_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_14_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_14_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_14_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_14_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_14_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_14_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_14_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_14_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z528 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_16_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_16_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_16_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z524 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_16_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64082_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_16_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_16_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_16_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_16_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_16_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_16_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_16_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_16_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z520 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_18_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_18_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_18_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z517 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_18_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64073_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_18_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_18_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_18_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_18_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_18_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_18_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_18_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_18_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z514 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_20_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_20_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_20_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z511 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_20_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64065_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_20_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_20_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_20_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_20_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_20_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_20_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_20_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_20_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z508 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_22_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_22_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_22_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_22_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z505 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1499_22_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_404_add_70_ix65206z64056_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z2 : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z693 : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64310_O_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64314_O : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z691 : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z689 : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64302_O_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z687 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_12_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_12_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_12_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z684 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_12_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64297_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_12_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_12_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_12_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_12_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_12_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_12_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_12_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_12_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z681 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_14_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_14_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_14_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z678 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_14_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64285_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_14_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_14_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_14_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_14_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_14_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_14_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_14_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_14_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z675 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_4_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_16_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_16_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_16_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z672 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_16_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64275_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_16_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_16_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_16_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_16_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_16_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_16_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_16_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_16_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z669 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_18_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_18_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_18_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z666 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_18_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64265_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_18_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_18_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_18_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_18_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_18_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_18_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_18_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_18_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z663 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_20_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_20_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_20_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z660 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_20_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64253_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_20_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_20_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_20_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_20_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_20_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_20_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_20_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_20_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z657 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_22_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_22_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_22_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_22_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z654 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1491_22_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_385_add_63_ix65206z64243_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z1_rt : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CY0F : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z492 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z64000_O_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z64004_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z489 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z486 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63992_O_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z483 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_8_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_8_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_8_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z479 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_8_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63985_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_8_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_8_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_8_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_8_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z475 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_10_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_10_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_10_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z471 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_10_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63973_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_10_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_10_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_10_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_10_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_10_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_10_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_10_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_10_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z467 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_12_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_12_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_12_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z463 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_12_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63962_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_12_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_12_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_12_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_12_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_12_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_12_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_12_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_12_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z459 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_14_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_14_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_14_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z455 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_14_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63952_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_14_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_14_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_14_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_14_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_14_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_14_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_14_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_14_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z451 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_16_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_16_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_16_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z447 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_16_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63942_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_16_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_16_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_16_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_16_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_16_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_16_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_16_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_16_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z443 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_18_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_18_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_18_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z440 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_18_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63933_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_18_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_18_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_18_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_18_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_18_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_18_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_18_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_18_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z437 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_20_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_20_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_20_CY0F : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_20_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z434 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1350_20_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_508_add_26_ix59700z63925_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_5_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_5_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_5_CY0F : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_5_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z40 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_5_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_5_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_5_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc_512_add_28_ix59700z63386_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_5_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_5_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z37 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_7_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_7_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_7_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z34 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_7_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_512_add_28_ix59700z63379_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_7_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_7_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_7_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_7_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_7_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_7_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_7_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_7_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z31 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_9_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_9_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_9_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z28 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_9_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_512_add_28_ix59700z63372_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_9_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_9_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_9_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_9_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z25 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_11_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_11_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_11_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z22 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_11_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_512_add_28_ix59700z63365_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_11_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_11_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_11_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_11_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z19 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_13_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_13_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_13_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z16 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_13_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_512_add_28_ix59700z63358_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_13_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_13_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_13_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_13_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z13 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_15_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_15_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_15_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z10 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_15_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_512_add_28_ix59700z63351_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_15_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_15_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_15_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_15_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_15_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_15_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_15_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_15_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z7 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_17_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1355_17_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z5_rt : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_2_XORF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_2_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_2_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z503 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_2_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z502 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_2_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_2_XORG : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_2_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z64052_O : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_2_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z500 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_2_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z499 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_4_XORF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_4_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_4_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z497 : STD_LOGIC; 
  signal U_DCT2D_nx65206z496 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_4_XORG : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z64040_O : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_4_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_4_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_4_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z494 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_4_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z493 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_6_XORF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_6_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_6_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z491 : STD_LOGIC; 
  signal U_DCT2D_nx65206z490 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_6_XORG : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z64028_O : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_6_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_6_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_6_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z488 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_6_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z487 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_8_XORF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_8_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_8_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z485 : STD_LOGIC; 
  signal U_DCT2D_nx65206z484 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_8_XORG : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z64016_O : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_8_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_8_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_8_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z482 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_8_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z481 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_10_XORF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_10_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z479 : STD_LOGIC; 
  signal U_DCT2D_nx65206z478 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_10_XORG : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z64004_O : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_10_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_10_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_10_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_10_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_10_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_10_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_10_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z476 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_10_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z475 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_12_XORF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_12_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_12_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z473 : STD_LOGIC; 
  signal U_DCT2D_nx65206z472 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_12_XORG : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z63992_O : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_12_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_12_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_12_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_12_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_12_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_12_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_12_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z470 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_12_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z469 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_14_XORF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_14_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_14_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z467 : STD_LOGIC; 
  signal U_DCT2D_nx65206z466 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_14_XORG : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z63980_O : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_14_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_14_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_14_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_14_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_14_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_14_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_14_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z464 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_14_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z463 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_16_XORF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_16_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_16_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z461 : STD_LOGIC; 
  signal U_DCT2D_nx65206z460 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_16_XORG : STD_LOGIC; 
  signal U_DCT2D_ix946_modgen_add_293_ix65206z63970_O : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_16_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_16_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_16_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_16_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_16_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_16_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_16_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z458 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_16_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z457 : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_18_XORF : STD_LOGIC; 
  signal U_DCT2D_nx115_bus_18_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z252_rt : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_5_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_5_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_5_CY0F : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_5_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z296 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_5_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_5_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_5_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63745_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_5_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_5_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z293 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_7_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_7_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_7_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z290 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_7_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63738_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_7_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_7_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_7_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_7_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_7_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_7_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_7_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_7_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z287 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_9_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_9_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_9_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z284 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_9_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63731_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_9_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_9_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_9_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_9_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z281 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_11_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_11_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_11_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z278 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_11_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63724_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_11_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_11_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_11_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_11_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z275 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_13_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_13_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_13_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z272 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_13_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63717_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_13_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_13_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_13_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_13_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z269 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_15_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_15_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_15_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z266 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_15_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63710_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_15_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_15_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_15_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_15_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_15_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_15_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_15_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_15_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z263 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_17_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_17_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_17_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z260 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_17_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_498_add_23_ix59700z63703_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_17_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_17_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_17_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_17_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_17_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_17_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_17_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_17_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z257 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_19_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1346_19_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z255_rt : STD_LOGIC; 
  signal romodatao4_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z945 : STD_LOGIC; 
  signal romodatao4_s_6_BXINV : STD_LOGIC; 
  signal romodatao4_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z944 : STD_LOGIC; 
  signal romodatao4_s_6_BYINV : STD_LOGIC; 
  signal nx54672z940_F5MUX : STD_LOGIC; 
  signal nx54672z942 : STD_LOGIC; 
  signal nx54672z940_BXINV : STD_LOGIC; 
  signal nx54672z941 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_FFY_RST : STD_LOGIC; 
  signal romodatao4_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z951 : STD_LOGIC; 
  signal romodatao4_s_5_BXINV : STD_LOGIC; 
  signal romodatao4_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z950 : STD_LOGIC; 
  signal romodatao4_s_5_BYINV : STD_LOGIC; 
  signal nx54672z946_F5MUX : STD_LOGIC; 
  signal nx54672z948 : STD_LOGIC; 
  signal nx54672z946_BXINV : STD_LOGIC; 
  signal nx54672z947 : STD_LOGIC; 
  signal romodatao4_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z957 : STD_LOGIC; 
  signal romodatao4_s_4_BXINV : STD_LOGIC; 
  signal romodatao4_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z956 : STD_LOGIC; 
  signal romodatao4_s_4_BYINV : STD_LOGIC; 
  signal nx54672z952_F5MUX : STD_LOGIC; 
  signal nx54672z954 : STD_LOGIC; 
  signal nx54672z952_BXINV : STD_LOGIC; 
  signal nx54672z953 : STD_LOGIC; 
  signal romodatao3_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z830 : STD_LOGIC; 
  signal romodatao3_s_12_BXINV : STD_LOGIC; 
  signal romodatao3_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z829 : STD_LOGIC; 
  signal romodatao3_s_12_BYINV : STD_LOGIC; 
  signal nx54672z825_F5MUX : STD_LOGIC; 
  signal nx54672z827 : STD_LOGIC; 
  signal nx54672z825_BXINV : STD_LOGIC; 
  signal nx54672z826 : STD_LOGIC; 
  signal romodatao3_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z842 : STD_LOGIC; 
  signal romodatao3_s_10_BXINV : STD_LOGIC; 
  signal romodatao3_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z841 : STD_LOGIC; 
  signal romodatao3_s_10_BYINV : STD_LOGIC; 
  signal nx54672z837_F5MUX : STD_LOGIC; 
  signal nx54672z839 : STD_LOGIC; 
  signal nx54672z837_BXINV : STD_LOGIC; 
  signal nx54672z838 : STD_LOGIC; 
  signal romodatao3_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z878 : STD_LOGIC; 
  signal romodatao3_s_4_BXINV : STD_LOGIC; 
  signal romodatao3_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z877 : STD_LOGIC; 
  signal romodatao3_s_4_BYINV : STD_LOGIC; 
  signal nx54672z873_F5MUX : STD_LOGIC; 
  signal nx54672z875 : STD_LOGIC; 
  signal nx54672z873_BXINV : STD_LOGIC; 
  signal nx54672z874 : STD_LOGIC; 
  signal romodatao3_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z890 : STD_LOGIC; 
  signal romodatao3_s_2_BXINV : STD_LOGIC; 
  signal romodatao3_s_2_F6MUX : STD_LOGIC; 
  signal nx54672z889 : STD_LOGIC; 
  signal romodatao3_s_2_BYINV : STD_LOGIC; 
  signal nx54672z885_F5MUX : STD_LOGIC; 
  signal nx54672z887 : STD_LOGIC; 
  signal nx54672z885_BXINV : STD_LOGIC; 
  signal nx54672z886 : STD_LOGIC; 
  signal romodatao3_s_0_F5MUX : STD_LOGIC; 
  signal nx54672z898 : STD_LOGIC; 
  signal romodatao3_s_0_BXINV : STD_LOGIC; 
  signal romodatao3_s_0_F6MUX : STD_LOGIC; 
  signal nx54672z897 : STD_LOGIC; 
  signal romodatao3_s_0_BYINV : STD_LOGIC; 
  signal U1_ROMO3_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROMO3_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROMO3_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROMO3_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romodatao2_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z763 : STD_LOGIC; 
  signal romodatao2_s_10_BXINV : STD_LOGIC; 
  signal romodatao2_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z762 : STD_LOGIC; 
  signal romodatao2_s_10_BYINV : STD_LOGIC; 
  signal nx54672z758_F5MUX : STD_LOGIC; 
  signal nx54672z760 : STD_LOGIC; 
  signal nx54672z758_BXINV : STD_LOGIC; 
  signal nx54672z759 : STD_LOGIC; 
  signal romodatao2_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z769 : STD_LOGIC; 
  signal romodatao2_s_9_BXINV : STD_LOGIC; 
  signal romodatao2_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z768 : STD_LOGIC; 
  signal romodatao2_s_9_BYINV : STD_LOGIC; 
  signal nx54672z764_F5MUX : STD_LOGIC; 
  signal nx54672z766 : STD_LOGIC; 
  signal nx54672z764_BXINV : STD_LOGIC; 
  signal nx54672z765 : STD_LOGIC; 
  signal romodatao2_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z775 : STD_LOGIC; 
  signal romodatao2_s_8_BXINV : STD_LOGIC; 
  signal romodatao2_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z774 : STD_LOGIC; 
  signal romodatao2_s_8_BYINV : STD_LOGIC; 
  signal nx54672z770_F5MUX : STD_LOGIC; 
  signal nx54672z772 : STD_LOGIC; 
  signal nx54672z770_BXINV : STD_LOGIC; 
  signal nx54672z771 : STD_LOGIC; 
  signal romodatao2_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z781 : STD_LOGIC; 
  signal romodatao2_s_7_BXINV : STD_LOGIC; 
  signal romodatao2_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z780 : STD_LOGIC; 
  signal romodatao2_s_7_BYINV : STD_LOGIC; 
  signal nx54672z776_F5MUX : STD_LOGIC; 
  signal nx54672z778 : STD_LOGIC; 
  signal nx54672z776_BXINV : STD_LOGIC; 
  signal nx54672z777 : STD_LOGIC; 
  signal romodatao2_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z787 : STD_LOGIC; 
  signal romodatao2_s_6_BXINV : STD_LOGIC; 
  signal romodatao2_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z786 : STD_LOGIC; 
  signal romodatao2_s_6_BYINV : STD_LOGIC; 
  signal nx54672z782_F5MUX : STD_LOGIC; 
  signal nx54672z784 : STD_LOGIC; 
  signal nx54672z782_BXINV : STD_LOGIC; 
  signal nx54672z783 : STD_LOGIC; 
  signal romodatao4_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z903 : STD_LOGIC; 
  signal romodatao4_s_13_BXINV : STD_LOGIC; 
  signal romodatao4_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z902 : STD_LOGIC; 
  signal romodatao4_s_13_BYINV : STD_LOGIC; 
  signal nx54672z899_F5MUX : STD_LOGIC; 
  signal nx54672z900 : STD_LOGIC; 
  signal nx54672z899_BXINV : STD_LOGIC; 
  signal nx54672z899_G : STD_LOGIC; 
  signal romodatao3_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z824 : STD_LOGIC; 
  signal romodatao3_s_13_BXINV : STD_LOGIC; 
  signal romodatao3_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z823 : STD_LOGIC; 
  signal romodatao3_s_13_BYINV : STD_LOGIC; 
  signal nx54672z820_F5MUX : STD_LOGIC; 
  signal nx54672z821 : STD_LOGIC; 
  signal nx54672z820_BXINV : STD_LOGIC; 
  signal nx54672z820_G : STD_LOGIC; 
  signal romodatao1_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z714 : STD_LOGIC; 
  signal romodatao1_s_5_BXINV : STD_LOGIC; 
  signal romodatao1_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z713 : STD_LOGIC; 
  signal romodatao1_s_5_BYINV : STD_LOGIC; 
  signal nx54672z709_F5MUX : STD_LOGIC; 
  signal nx54672z711 : STD_LOGIC; 
  signal nx54672z709_BXINV : STD_LOGIC; 
  signal nx54672z710 : STD_LOGIC; 
  signal romodatao1_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z720 : STD_LOGIC; 
  signal romodatao1_s_4_BXINV : STD_LOGIC; 
  signal romodatao1_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z719 : STD_LOGIC; 
  signal romodatao1_s_4_BYINV : STD_LOGIC; 
  signal nx54672z715_F5MUX : STD_LOGIC; 
  signal nx54672z717 : STD_LOGIC; 
  signal nx54672z715_BXINV : STD_LOGIC; 
  signal nx54672z716 : STD_LOGIC; 
  signal romodatao1_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z726 : STD_LOGIC; 
  signal romodatao1_s_3_BXINV : STD_LOGIC; 
  signal romodatao1_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z725 : STD_LOGIC; 
  signal romodatao1_s_3_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_0_FFX_RST : STD_LOGIC; 
  signal nx54672z721_F5MUX : STD_LOGIC; 
  signal nx54672z723 : STD_LOGIC; 
  signal nx54672z721_BXINV : STD_LOGIC; 
  signal nx54672z722 : STD_LOGIC; 
  signal romedatao6_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z394 : STD_LOGIC; 
  signal romedatao6_s_13_BXINV : STD_LOGIC; 
  signal romedatao6_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z393 : STD_LOGIC; 
  signal romedatao6_s_13_BYINV : STD_LOGIC; 
  signal nx54672z390_F5MUX : STD_LOGIC; 
  signal nx54672z391 : STD_LOGIC; 
  signal nx54672z390_BXINV : STD_LOGIC; 
  signal nx54672z390_G : STD_LOGIC; 
  signal romedatao4_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z270 : STD_LOGIC; 
  signal romedatao4_s_12_BXINV : STD_LOGIC; 
  signal romedatao4_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z269 : STD_LOGIC; 
  signal romedatao4_s_12_BYINV : STD_LOGIC; 
  signal nx54672z265_F5MUX : STD_LOGIC; 
  signal nx54672z267 : STD_LOGIC; 
  signal nx54672z265_BXINV : STD_LOGIC; 
  signal nx54672z266 : STD_LOGIC; 
  signal romedatao4_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z276 : STD_LOGIC; 
  signal romedatao4_s_11_BXINV : STD_LOGIC; 
  signal romedatao4_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z275 : STD_LOGIC; 
  signal romedatao4_s_11_BYINV : STD_LOGIC; 
  signal nx54672z271_F5MUX : STD_LOGIC; 
  signal nx54672z273 : STD_LOGIC; 
  signal nx54672z271_BXINV : STD_LOGIC; 
  signal nx54672z272 : STD_LOGIC; 
  signal romedatao4_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z282 : STD_LOGIC; 
  signal romedatao4_s_10_BXINV : STD_LOGIC; 
  signal romedatao4_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z281 : STD_LOGIC; 
  signal romedatao4_s_10_BYINV : STD_LOGIC; 
  signal nx54672z277_F5MUX : STD_LOGIC; 
  signal nx54672z279 : STD_LOGIC; 
  signal nx54672z277_BXINV : STD_LOGIC; 
  signal nx54672z278 : STD_LOGIC; 
  signal romedatao4_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z318 : STD_LOGIC; 
  signal romedatao4_s_4_BXINV : STD_LOGIC; 
  signal romedatao4_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z317 : STD_LOGIC; 
  signal romedatao4_s_4_BYINV : STD_LOGIC; 
  signal U_DCT1D_nx59700z428_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z428_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z428_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z428_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z428_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z428_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_nx59700z428_XORG : STD_LOGIC; 
  signal U_DCT1D_nx59700z428_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_ix740_modgen_add_290_ix59700z63793_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z428_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z428_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z329 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_nx59700z420_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z420_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z420_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z326 : STD_LOGIC; 
  signal U_DCT1D_nx59700z420_XORG : STD_LOGIC; 
  signal U_DCT1D_ix740_modgen_add_290_ix59700z63785_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z420_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z420_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_nx59700z420_CYAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z420_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_nx59700z420_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z420_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z420_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z420_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z323 : STD_LOGIC; 
  signal U_DCT1D_nx59700z412_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z412_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z412_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z320 : STD_LOGIC; 
  signal U_DCT1D_nx59700z412_XORG : STD_LOGIC; 
  signal U_DCT1D_ix740_modgen_add_290_ix59700z63777_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z412_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z412_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_nx59700z412_CYAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z412_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_nx59700z412_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z412_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z412_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z412_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z317 : STD_LOGIC; 
  signal U_DCT1D_nx59700z404_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z404_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z404_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z314 : STD_LOGIC; 
  signal U_DCT1D_nx59700z404_XORG : STD_LOGIC; 
  signal U_DCT1D_ix740_modgen_add_290_ix59700z63769_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z404_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z404_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_nx59700z404_CYAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z404_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_nx59700z404_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z404_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z404_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z404_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z311 : STD_LOGIC; 
  signal U_DCT1D_nx59700z396_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z396_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z396_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z308 : STD_LOGIC; 
  signal U_DCT1D_nx59700z396_XORG : STD_LOGIC; 
  signal U_DCT1D_ix740_modgen_add_290_ix59700z63761_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z396_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z396_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_nx59700z396_CYAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z396_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_nx59700z396_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z396_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z396_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z396_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z305 : STD_LOGIC; 
  signal U_DCT1D_nx59700z388_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z388_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z388_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z302 : STD_LOGIC; 
  signal U_DCT1D_nx59700z388_XORG : STD_LOGIC; 
  signal U_DCT1D_ix740_modgen_add_290_ix59700z63753_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z388_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z388_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_nx59700z388_CYAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z388_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_nx59700z388_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z388_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z388_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z388_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z299 : STD_LOGIC; 
  signal U_DCT1D_nx59700z253_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z253_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z254_rt : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_7_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_7_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_7_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_7_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z332 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_7_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_7_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_7_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc_394_add_67_ix65206z63792_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_7_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_7_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z329 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_9_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_9_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_9_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z326 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_9_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_394_add_67_ix65206z63784_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_9_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_9_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_9_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_9_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z323 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_11_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_11_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_11_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z320 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_11_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_394_add_67_ix65206z63777_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_11_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_11_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_11_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_11_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z317 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_13_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_13_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_13_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z314 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_13_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_394_add_67_ix65206z63770_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_13_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_13_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_13_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_13_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z311 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_15_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_15_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_15_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z308 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_15_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_394_add_67_ix65206z63763_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_15_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_15_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_15_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_15_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_15_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_15_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_15_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_15_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z305 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_17_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_17_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_17_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z302 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_17_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_394_add_67_ix65206z63756_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_17_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_17_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_17_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_17_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_17_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_17_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_17_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_17_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z299 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_19_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1494_19_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z297_rt : STD_LOGIC; 
  signal U_DCT2D_nx65206z570_XORF : STD_LOGIC; 
  signal U_DCT2D_nx65206z570_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z570_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z570_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z570_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z570_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_nx65206z570_XORG : STD_LOGIC; 
  signal U_DCT2D_nx65206z570_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63689_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z570_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z570_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z247 : STD_LOGIC; 
  signal U_DCT2D_nx65206z564_XORF : STD_LOGIC; 
  signal U_DCT2D_nx65206z564_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z564_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z244 : STD_LOGIC; 
  signal U_DCT2D_nx65206z564_XORG : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63677_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z564_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z564_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx65206z564_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx65206z564_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx65206z564_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx65206z564_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx65206z564_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z564_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z241 : STD_LOGIC; 
  signal U_DCT2D_nx65206z557_XORF : STD_LOGIC; 
  signal U_DCT2D_nx65206z557_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z557_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z238 : STD_LOGIC; 
  signal U_DCT2D_nx65206z557_XORG : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63665_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z557_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z557_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx65206z557_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx65206z557_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx65206z557_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx65206z557_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx65206z557_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z557_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z235 : STD_LOGIC; 
  signal U_DCT2D_nx65206z549_XORF : STD_LOGIC; 
  signal U_DCT2D_nx65206z549_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z549_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z232 : STD_LOGIC; 
  signal U_DCT2D_nx65206z549_XORG : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63653_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z549_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z549_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx65206z549_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx65206z549_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx65206z549_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx65206z549_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx65206z549_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z549_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z229 : STD_LOGIC; 
  signal U_DCT2D_nx65206z541_XORF : STD_LOGIC; 
  signal U_DCT2D_nx65206z541_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z541_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z226 : STD_LOGIC; 
  signal U_DCT2D_nx65206z541_XORG : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63641_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z541_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z541_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx65206z541_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx65206z541_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx65206z541_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx65206z541_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx65206z541_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z541_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z223 : STD_LOGIC; 
  signal U_DCT2D_nx65206z533_XORF : STD_LOGIC; 
  signal U_DCT2D_nx65206z533_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z533_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z220 : STD_LOGIC; 
  signal U_DCT2D_nx65206z533_XORG : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63629_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z533_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z533_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx65206z533_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx65206z533_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx65206z533_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx65206z533_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx65206z533_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z533_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z217 : STD_LOGIC; 
  signal U_DCT2D_nx65206z525_XORF : STD_LOGIC; 
  signal U_DCT2D_nx65206z525_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z525_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z214 : STD_LOGIC; 
  signal U_DCT2D_nx65206z525_XORG : STD_LOGIC; 
  signal U_DCT2D_ix959_modgen_add_291_ix65206z63619_O : STD_LOGIC; 
  signal U_DCT2D_nx65206z525_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z525_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_nx65206z525_CYAND : STD_LOGIC; 
  signal U_DCT2D_nx65206z525_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_nx65206z525_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_nx65206z525_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_nx65206z525_CY0G : STD_LOGIC; 
  signal U_DCT2D_nx65206z525_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z211 : STD_LOGIC; 
  signal U_DCT2D_nx65206z3_XORF : STD_LOGIC; 
  signal U_DCT2D_nx65206z3_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z4_rt : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_2_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_2_CY0F : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_2_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z120 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_2_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_2_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_2_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63485_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_2_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_2_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z117 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_3_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_3_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_3_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z114 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_3_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63478_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_3_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_3_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_3_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_3_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_3_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_3_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_3_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_3_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z111 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_5_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_5_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_5_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z108 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_5_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63471_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_5_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_5_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_5_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_5_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_5_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_5_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_5_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_5_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z105 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_7_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_7_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_7_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z102 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_7_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63463_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_7_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_7_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_7_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_7_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_7_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_7_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_7_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_7_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z99 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_9_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_9_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_9_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z96 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_9_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63456_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_9_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_9_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_9_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_9_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z93 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_11_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_11_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_11_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z90 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_11_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63449_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_11_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_11_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_11_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_11_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z87 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_13_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_13_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_13_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z84 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_13_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_491_add_20_ix59700z63442_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_13_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_13_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_13_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_13_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z81 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_15_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1344_15_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z79_rt : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_3_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_3_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_3_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_3_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z162 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_3_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_3_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_3_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63535_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_3_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_3_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z159 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_6_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_5_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_5_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_5_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z156 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_5_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63528_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_5_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_5_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_5_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_5_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_5_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_5_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_5_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_5_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z153 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_7_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_7_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_7_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z150 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_7_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63521_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_7_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_7_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_7_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_7_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_7_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_7_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_7_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_7_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z147 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_9_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_9_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_9_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z144 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_9_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63514_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_9_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_9_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_9_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_9_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z141 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_11_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_11_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_11_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z138 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_11_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63506_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_11_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_11_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_11_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_11_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z135 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_13_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_13_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_13_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z132 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_13_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63499_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_13_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_13_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_13_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_13_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z129 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_15_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_15_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_15_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z126 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_15_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_333_add_55_ix65206z63492_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_15_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_15_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_15_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_15_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_15_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_15_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_15_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_15_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z123 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_17_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1481_17_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z121_rt : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_8_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_8_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_8_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_8_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z411 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_8_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_8_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_8_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63910_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_8_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_8_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z408 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_10_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_10_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_10_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z405 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_10_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63898_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_10_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_10_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_10_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_10_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_10_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_10_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_10_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_10_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z402 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_12_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_12_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_12_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z399 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_12_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63886_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_12_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_12_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_12_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_12_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_12_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_12_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_12_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_12_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z396 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_14_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_14_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_14_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z393 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_14_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63874_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_14_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_14_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_14_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_14_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_14_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_14_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_14_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_14_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z390 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_16_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_16_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_16_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z387 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_16_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63862_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_16_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_16_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_16_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_16_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_16_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_16_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_16_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_16_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z384 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_18_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_18_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_18_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z381 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_18_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63851_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_18_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_18_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_18_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_18_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_18_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_18_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_18_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_18_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z378 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_20_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_20_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_20_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z375 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_20_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_399_add_69_ix65206z63843_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_20_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_20_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_20_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_20_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_20_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_20_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_20_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_20_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z372 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_22_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1498_22_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z296_rt : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_4_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_4_CY0F : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_4_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z77 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_4_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_4_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_4_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc_510_add_27_ix59700z63433_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_4_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_4_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z74 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_5_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_5_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_5_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z71 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_5_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_510_add_27_ix59700z63426_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_5_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_5_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_5_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_5_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_5_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_5_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_5_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_5_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z68 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_7_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_7_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_7_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z65 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_7_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_510_add_27_ix59700z63419_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_7_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_7_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_7_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_7_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_7_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_7_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_7_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_7_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z62 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_9_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_9_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_9_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z59 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_9_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_510_add_27_ix59700z63412_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_9_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_9_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_9_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_9_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z56 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_11_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_11_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_11_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z53 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_11_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_510_add_27_ix59700z63405_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_11_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_11_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_11_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_11_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z50 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_13_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_13_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_13_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z47 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_13_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_510_add_27_ix59700z63398_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_13_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_13_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_13_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_13_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z44 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_15_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1354_15_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z42_rt : STD_LOGIC; 
  signal U_DCT1D_nx59700z493_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z493_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z493_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z493_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z493_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z493_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_nx59700z493_XORG : STD_LOGIC; 
  signal U_DCT1D_nx59700z493_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63689_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z493_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z493_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z247 : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_8_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_2_8_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z487_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z487_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z487_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z244 : STD_LOGIC; 
  signal U_DCT1D_nx59700z487_XORG : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63677_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z487_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z487_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_nx59700z487_CYAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z487_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_nx59700z487_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z487_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z487_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z487_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z241 : STD_LOGIC; 
  signal U_DCT1D_nx59700z480_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z480_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z480_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z238 : STD_LOGIC; 
  signal U_DCT1D_nx59700z480_XORG : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63665_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z480_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z480_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_nx59700z480_CYAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z480_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_nx59700z480_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z480_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z480_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z480_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z235 : STD_LOGIC; 
  signal U_DCT1D_nx59700z472_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z472_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z472_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z232 : STD_LOGIC; 
  signal U_DCT1D_nx59700z472_XORG : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63653_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z472_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z472_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_nx59700z472_CYAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z472_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_nx59700z472_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z472_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z472_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z472_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z229 : STD_LOGIC; 
  signal U_DCT1D_nx59700z464_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z464_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z464_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z226 : STD_LOGIC; 
  signal U_DCT1D_nx59700z464_XORG : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63641_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z464_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z464_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_nx59700z464_CYAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z464_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_nx59700z464_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z464_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z464_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z464_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z223 : STD_LOGIC; 
  signal U_DCT1D_nx59700z456_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z456_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z456_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z220 : STD_LOGIC; 
  signal U_DCT1D_nx59700z456_XORG : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63629_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z456_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z456_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_nx59700z456_CYAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z456_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_nx59700z456_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z456_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z456_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z456_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z217 : STD_LOGIC; 
  signal U_DCT1D_nx59700z448_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z448_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z448_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z214 : STD_LOGIC; 
  signal U_DCT1D_nx59700z448_XORG : STD_LOGIC; 
  signal U_DCT1D_ix773_modgen_add_291_ix59700z63619_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z448_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z448_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_nx59700z448_CYAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z448_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_nx59700z448_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z448_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_nx59700z448_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z448_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z211 : STD_LOGIC; 
  signal U_DCT1D_nx59700z3_XORF : STD_LOGIC; 
  signal U_DCT1D_nx59700z3_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z4_rt : STD_LOGIC; 
  signal U_DCT1D_ix59700z64053_O_CYINIT : STD_LOGIC; 
  signal U_DCT1D_ix59700z64053_O_CY0F : STD_LOGIC; 
  signal U_DCT1D_ix59700z64053_O_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z528 : STD_LOGIC; 
  signal U_DCT1D_ix59700z64053_O_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_ix59700z64056_O : STD_LOGIC; 
  signal U_DCT1D_ix59700z64053_O_CY0G : STD_LOGIC; 
  signal U_DCT1D_ix59700z64053_O_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z526 : STD_LOGIC; 
  signal U_DCT1D_ix59700z64047_O_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z524 : STD_LOGIC; 
  signal U_DCT1D_ix59700z64047_O_CYSELF : STD_LOGIC; 
  signal U_DCT1D_ix59700z64047_O_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_ix59700z64047_O_CYAND : STD_LOGIC; 
  signal U_DCT1D_ix59700z64047_O_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_ix59700z64047_O_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_ix59700z64047_O_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_ix59700z64047_O_CY0G : STD_LOGIC; 
  signal U_DCT1D_ix59700z64047_O_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z522 : STD_LOGIC; 
  signal ramdatai_s_0_DXMUX : STD_LOGIC; 
  signal ramdatai_s_0_FXMUX : STD_LOGIC; 
  signal ramdatai_s_0_XORF : STD_LOGIC; 
  signal ramdatai_s_0_CYINIT : STD_LOGIC; 
  signal ramdatai_s_0_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z519 : STD_LOGIC; 
  signal ramdatai_s_0_DYMUX : STD_LOGIC; 
  signal ramdatai_s_0_GYMUX : STD_LOGIC; 
  signal ramdatai_s_0_XORG : STD_LOGIC; 
  signal U_DCT1D_ix59700z64042_O : STD_LOGIC; 
  signal ramdatai_s_0_CYSELF : STD_LOGIC; 
  signal ramdatai_s_0_CYMUXFAST : STD_LOGIC; 
  signal ramdatai_s_0_CYAND : STD_LOGIC; 
  signal ramdatai_s_0_FASTCARRY : STD_LOGIC; 
  signal ramdatai_s_0_CYMUXG2 : STD_LOGIC; 
  signal ramdatai_s_0_CYMUXF2 : STD_LOGIC; 
  signal ramdatai_s_0_CY0G : STD_LOGIC; 
  signal ramdatai_s_0_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z516 : STD_LOGIC; 
  signal ramdatai_s_0_SRINV : STD_LOGIC; 
  signal ramdatai_s_0_CLKINV : STD_LOGIC; 
  signal ramdatai_s_0_CEINV : STD_LOGIC; 
  signal ramdatai_s_2_DXMUX : STD_LOGIC; 
  signal ramdatai_s_2_FXMUX : STD_LOGIC; 
  signal ramdatai_s_2_XORF : STD_LOGIC; 
  signal ramdatai_s_2_CYINIT : STD_LOGIC; 
  signal ramdatai_s_2_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z513 : STD_LOGIC; 
  signal ramdatai_s_2_DYMUX : STD_LOGIC; 
  signal ramdatai_s_2_GYMUX : STD_LOGIC; 
  signal ramdatai_s_2_XORG : STD_LOGIC; 
  signal U_DCT1D_ix59700z64033_O : STD_LOGIC; 
  signal ramdatai_s_2_CYSELF : STD_LOGIC; 
  signal ramdatai_s_2_CYMUXFAST : STD_LOGIC; 
  signal ramdatai_s_2_CYAND : STD_LOGIC; 
  signal ramdatai_s_2_FASTCARRY : STD_LOGIC; 
  signal ramdatai_s_2_CYMUXG2 : STD_LOGIC; 
  signal ramdatai_s_2_CYMUXF2 : STD_LOGIC; 
  signal ramdatai_s_2_CY0G : STD_LOGIC; 
  signal ramdatai_s_2_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z510 : STD_LOGIC; 
  signal ramdatai_s_2_SRINV : STD_LOGIC; 
  signal ramdatai_s_2_CLKINV : STD_LOGIC; 
  signal ramdatai_s_2_CEINV : STD_LOGIC; 
  signal ramdatai_s_4_DXMUX : STD_LOGIC; 
  signal ramdatai_s_4_FXMUX : STD_LOGIC; 
  signal ramdatai_s_4_XORF : STD_LOGIC; 
  signal ramdatai_s_4_CYINIT : STD_LOGIC; 
  signal ramdatai_s_4_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z507 : STD_LOGIC; 
  signal ramdatai_s_4_DYMUX : STD_LOGIC; 
  signal ramdatai_s_4_GYMUX : STD_LOGIC; 
  signal ramdatai_s_4_XORG : STD_LOGIC; 
  signal U_DCT1D_ix59700z64025_O : STD_LOGIC; 
  signal ramdatai_s_4_CYSELF : STD_LOGIC; 
  signal ramdatai_s_4_CYMUXFAST : STD_LOGIC; 
  signal ramdatai_s_4_CYAND : STD_LOGIC; 
  signal ramdatai_s_4_FASTCARRY : STD_LOGIC; 
  signal ramdatai_s_4_CYMUXG2 : STD_LOGIC; 
  signal ramdatai_s_4_CYMUXF2 : STD_LOGIC; 
  signal ramdatai_s_4_CY0G : STD_LOGIC; 
  signal ramdatai_s_4_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z504 : STD_LOGIC; 
  signal ramdatai_s_4_SRINV : STD_LOGIC; 
  signal ramdatai_s_4_CLKINV : STD_LOGIC; 
  signal ramdatai_s_4_CEINV : STD_LOGIC; 
  signal ramdatai_s_6_DXMUX : STD_LOGIC; 
  signal ramdatai_s_6_FXMUX : STD_LOGIC; 
  signal ramdatai_s_6_XORF : STD_LOGIC; 
  signal ramdatai_s_6_CYINIT : STD_LOGIC; 
  signal ramdatai_s_6_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z501 : STD_LOGIC; 
  signal ramdatai_s_6_DYMUX : STD_LOGIC; 
  signal ramdatai_s_6_GYMUX : STD_LOGIC; 
  signal ramdatai_s_6_XORG : STD_LOGIC; 
  signal U_DCT1D_ix59700z64016_O : STD_LOGIC; 
  signal ramdatai_s_6_CYSELF : STD_LOGIC; 
  signal ramdatai_s_6_CYMUXFAST : STD_LOGIC; 
  signal ramdatai_s_6_CYAND : STD_LOGIC; 
  signal ramdatai_s_6_FASTCARRY : STD_LOGIC; 
  signal ramdatai_s_6_CYMUXG2 : STD_LOGIC; 
  signal ramdatai_s_6_CYMUXF2 : STD_LOGIC; 
  signal ramdatai_s_6_CY0G : STD_LOGIC; 
  signal ramdatai_s_6_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z498 : STD_LOGIC; 
  signal ramdatai_s_6_SRINV : STD_LOGIC; 
  signal ramdatai_s_6_CLKINV : STD_LOGIC; 
  signal ramdatai_s_6_CEINV : STD_LOGIC; 
  signal ramdatai_s_8_DXMUX : STD_LOGIC; 
  signal ramdatai_s_8_FXMUX : STD_LOGIC; 
  signal ramdatai_s_8_XORF : STD_LOGIC; 
  signal ramdatai_s_8_CYINIT : STD_LOGIC; 
  signal ramdatai_s_8_CY0F : STD_LOGIC; 
  signal ramdatai_s_8_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z495 : STD_LOGIC; 
  signal ramdatai_s_8_DYMUX : STD_LOGIC; 
  signal ramdatai_s_8_GYMUX : STD_LOGIC; 
  signal ramdatai_s_8_XORG : STD_LOGIC; 
  signal U_DCT1D_ix59700z64007_O : STD_LOGIC; 
  signal U_DCT1D_nx59700z1_rt : STD_LOGIC; 
  signal ramdatai_s_8_SRINV : STD_LOGIC; 
  signal ramdatai_s_8_CLKINV : STD_LOGIC; 
  signal ramdatai_s_8_CEINV : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_7_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_7_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_7_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z375 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_7_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z374 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_7_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_7_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_7_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_ix59700z63837_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_7_CY0G : STD_LOGIC; 
  signal U_DCT1D_nx59700z372 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_7_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z371 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_9_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_9_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_9_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z368 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_9_XORG : STD_LOGIC; 
  signal U_DCT1D_ix59700z63831_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_9_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_9_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_9_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_9_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z365 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_11_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_11_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_11_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z362 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_11_XORG : STD_LOGIC; 
  signal U_DCT1D_ix59700z63825_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_11_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_11_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_11_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_11_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z359 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_13_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_13_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_13_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z356 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_13_XORG : STD_LOGIC; 
  signal U_DCT1D_ix59700z63819_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_13_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_13_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_13_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_13_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z353 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_15_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_15_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_15_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z350 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_15_XORG : STD_LOGIC; 
  signal U_DCT1D_ix59700z63813_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_15_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_15_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_15_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_15_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_15_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_15_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_15_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_15_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z347 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_17_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_17_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_17_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z344 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_17_XORG : STD_LOGIC; 
  signal U_DCT1D_ix59700z63807_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_17_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_17_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_17_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_17_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_17_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_17_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_17_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_17_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z341 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_19_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_19_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_19_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z339 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_19_XORG : STD_LOGIC; 
  signal U_DCT1D_ix59700z63802_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_19_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_19_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_19_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_19_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_19_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_19_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_19_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_19_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z337 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_21_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1347_21_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z334_rt : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CY0F : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYSELF : STD_LOGIC; 
  signal U_DCT1D_nx59700z209 : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63608_O_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYMUXG : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63612_O : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z207 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_4_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_4_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_4_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z204 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_4_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63603_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_4_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_4_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_4_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_4_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_4_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_4_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_4_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_4_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z201 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_6_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_6_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_6_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z198 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_6_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63592_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_6_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_6_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_6_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_6_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_6_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_6_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_6_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_6_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z195 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_8_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_8_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_8_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z192 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_8_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63582_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_8_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_8_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_8_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_8_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_8_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_8_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_8_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_8_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z189 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_10_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_10_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_10_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z186 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_10_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63572_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_10_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_10_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_10_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_10_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_10_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_10_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_10_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_10_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z183 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_12_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_12_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_12_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z180 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_12_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63561_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_12_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_12_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_12_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_12_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_12_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_12_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_12_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_12_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z177 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_14_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_14_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_14_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z174 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_14_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63551_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_14_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_14_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_14_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_14_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_14_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_14_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_14_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_14_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z171 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_16_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_16_CYINIT : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_16_CY0F : STD_LOGIC; 
  signal U_DCT1D_nx59700z168 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_16_XORG : STD_LOGIC; 
  signal U_DCT1D_rtlc_496_add_22_ix59700z63542_O : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_16_CYSELF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_16_CYMUXFAST : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_16_CYAND : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_16_FASTCARRY : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_16_CYMUXG2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_16_CYMUXF2 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_16_CY0G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_16_CYSELG : STD_LOGIC; 
  signal U_DCT1D_nx59700z165 : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_18_XORF : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1348_18_CYINIT : STD_LOGIC; 
  signal U_DCT1D_nx59700z78_rt : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_5_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_5_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_5_CY0F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_5_CYSELF : STD_LOGIC; 
  signal U_DCT2D_nx65206z454 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_5_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_5_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_5_CYMUXG : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63963_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_5_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_5_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z451 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_7_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_7_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_7_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z448 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_7_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63956_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_7_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_7_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_7_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_7_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_7_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_7_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_7_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_7_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z445 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_9_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_9_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_9_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z442 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_9_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63949_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_9_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_9_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_9_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_9_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_9_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_9_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_9_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_9_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z439 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_11_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_11_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_11_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z436 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_11_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63942_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_11_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_11_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_11_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_11_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_11_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_11_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_11_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_11_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z433 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_13_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_13_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_13_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z430 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_13_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63935_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_13_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_13_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_13_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_13_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_13_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_13_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_13_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_13_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z427 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_15_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_15_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_15_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z424 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_15_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63928_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_15_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_15_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_15_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_15_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_15_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_15_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_15_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_15_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z421 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_17_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_17_CYINIT : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_17_CY0F : STD_LOGIC; 
  signal U_DCT2D_nx65206z418 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_17_XORG : STD_LOGIC; 
  signal U_DCT2D_rtlc_338_add_57_ix65206z63921_O : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_17_CYSELF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_17_CYMUXFAST : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_17_CYAND : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_17_FASTCARRY : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_17_CYMUXG2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_17_CYMUXF2 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_17_CY0G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_17_CYSELG : STD_LOGIC; 
  signal U_DCT2D_nx65206z415 : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_19_XORF : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1482_19_CYINIT : STD_LOGIC; 
  signal U_DCT2D_nx65206z413_rt : STD_LOGIC; 
  signal nx53675z1410_F5MUX : STD_LOGIC; 
  signal nx53675z1412 : STD_LOGIC; 
  signal nx53675z1410_BXINV : STD_LOGIC; 
  signal nx53675z1411 : STD_LOGIC; 
  signal rome2datao5_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z335 : STD_LOGIC; 
  signal rome2datao5_s_12_BXINV : STD_LOGIC; 
  signal rome2datao5_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z334 : STD_LOGIC; 
  signal rome2datao5_s_12_BYINV : STD_LOGIC; 
  signal nx53675z330_F5MUX : STD_LOGIC; 
  signal nx53675z332 : STD_LOGIC; 
  signal nx53675z330_BXINV : STD_LOGIC; 
  signal nx53675z331 : STD_LOGIC; 
  signal rome2datao5_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z341 : STD_LOGIC; 
  signal rome2datao5_s_11_BXINV : STD_LOGIC; 
  signal rome2datao5_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z340 : STD_LOGIC; 
  signal rome2datao5_s_11_BYINV : STD_LOGIC; 
  signal nx53675z336_F5MUX : STD_LOGIC; 
  signal nx53675z338 : STD_LOGIC; 
  signal nx53675z336_BXINV : STD_LOGIC; 
  signal nx53675z337 : STD_LOGIC; 
  signal rome2datao5_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z347 : STD_LOGIC; 
  signal rome2datao5_s_10_BXINV : STD_LOGIC; 
  signal rome2datao5_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z346 : STD_LOGIC; 
  signal rome2datao5_s_10_BYINV : STD_LOGIC; 
  signal nx53675z342_F5MUX : STD_LOGIC; 
  signal nx53675z344 : STD_LOGIC; 
  signal nx53675z342_BXINV : STD_LOGIC; 
  signal nx53675z343 : STD_LOGIC; 
  signal rome2datao5_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z353 : STD_LOGIC; 
  signal rome2datao5_s_9_BXINV : STD_LOGIC; 
  signal rome2datao5_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z352 : STD_LOGIC; 
  signal rome2datao5_s_9_BYINV : STD_LOGIC; 
  signal nx53675z348_F5MUX : STD_LOGIC; 
  signal nx53675z350 : STD_LOGIC; 
  signal nx53675z348_BXINV : STD_LOGIC; 
  signal nx53675z349 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_10_FFX_RSTAND : STD_LOGIC; 
  signal rome2datao5_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z388 : STD_LOGIC; 
  signal rome2datao5_s_3_BXINV : STD_LOGIC; 
  signal rome2datao5_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z387 : STD_LOGIC; 
  signal rome2datao5_s_3_BYINV : STD_LOGIC; 
  signal nx53675z384_F5MUX : STD_LOGIC; 
  signal nx53675z385 : STD_LOGIC; 
  signal nx53675z384_BXINV : STD_LOGIC; 
  signal U2_ROME5_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal rome2datao5_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z389 : STD_LOGIC; 
  signal rome2datao5_s_2_BXINV : STD_LOGIC; 
  signal rome2datao5_s_2_F6MUX : STD_LOGIC; 
  signal rome2datao5_s_2_G : STD_LOGIC; 
  signal rome2datao5_s_2_BYINV : STD_LOGIC; 
  signal U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROME5_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romo2datao8_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z1349 : STD_LOGIC; 
  signal romo2datao8_s_13_BXINV : STD_LOGIC; 
  signal romo2datao8_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z1348 : STD_LOGIC; 
  signal romo2datao8_s_13_BYINV : STD_LOGIC; 
  signal nx53675z1345_F5MUX : STD_LOGIC; 
  signal nx53675z1346 : STD_LOGIC; 
  signal nx53675z1345_BXINV : STD_LOGIC; 
  signal nx53675z1345_G : STD_LOGIC; 
  signal romo2datao8_s_1_F5MUX : STD_LOGIC; 
  signal nx53675z1421 : STD_LOGIC; 
  signal romo2datao8_s_1_BXINV : STD_LOGIC; 
  signal romo2datao8_s_1_F6MUX : STD_LOGIC; 
  signal nx53675z1420 : STD_LOGIC; 
  signal romo2datao8_s_1_BYINV : STD_LOGIC; 
  signal nx53675z1416_F5MUX : STD_LOGIC; 
  signal nx53675z1418 : STD_LOGIC; 
  signal nx53675z1416_BXINV : STD_LOGIC; 
  signal nx53675z1417 : STD_LOGIC; 
  signal rome2datao7_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z465 : STD_LOGIC; 
  signal rome2datao7_s_12_BXINV : STD_LOGIC; 
  signal rome2datao7_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z464 : STD_LOGIC; 
  signal rome2datao7_s_12_BYINV : STD_LOGIC; 
  signal nx53675z460_F5MUX : STD_LOGIC; 
  signal nx53675z462 : STD_LOGIC; 
  signal nx53675z460_BXINV : STD_LOGIC; 
  signal nx53675z461 : STD_LOGIC; 
  signal rome2datao7_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z471 : STD_LOGIC; 
  signal rome2datao7_s_11_BXINV : STD_LOGIC; 
  signal rome2datao7_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z470 : STD_LOGIC; 
  signal rome2datao7_s_11_BYINV : STD_LOGIC; 
  signal nx53675z466_F5MUX : STD_LOGIC; 
  signal nx53675z468 : STD_LOGIC; 
  signal nx53675z466_BXINV : STD_LOGIC; 
  signal nx53675z467 : STD_LOGIC; 
  signal rome2datao7_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z518 : STD_LOGIC; 
  signal rome2datao7_s_3_BXINV : STD_LOGIC; 
  signal rome2datao7_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z517 : STD_LOGIC; 
  signal rome2datao7_s_3_BYINV : STD_LOGIC; 
  signal nx53675z514_F5MUX : STD_LOGIC; 
  signal nx53675z515 : STD_LOGIC; 
  signal nx53675z514_BXINV : STD_LOGIC; 
  signal U2_ROME7_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal rome2datao7_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z519 : STD_LOGIC; 
  signal rome2datao7_s_2_BXINV : STD_LOGIC; 
  signal rome2datao7_s_2_F6MUX : STD_LOGIC; 
  signal rome2datao7_s_2_G : STD_LOGIC; 
  signal rome2datao7_s_2_BYINV : STD_LOGIC; 
  signal U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROME7_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romo2datao9_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z1470 : STD_LOGIC; 
  signal romo2datao9_s_6_BXINV : STD_LOGIC; 
  signal romo2datao9_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z1469 : STD_LOGIC; 
  signal romo2datao9_s_6_BYINV : STD_LOGIC; 
  signal nx53675z1465_F5MUX : STD_LOGIC; 
  signal nx53675z1467 : STD_LOGIC; 
  signal nx53675z1465_BXINV : STD_LOGIC; 
  signal nx53675z1466 : STD_LOGIC; 
  signal romo2datao9_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z1476 : STD_LOGIC; 
  signal romo2datao9_s_5_BXINV : STD_LOGIC; 
  signal romo2datao9_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z1475 : STD_LOGIC; 
  signal romo2datao9_s_5_BYINV : STD_LOGIC; 
  signal nx53675z1471_F5MUX : STD_LOGIC; 
  signal nx53675z1473 : STD_LOGIC; 
  signal nx53675z1471_BXINV : STD_LOGIC; 
  signal nx53675z1472 : STD_LOGIC; 
  signal romo2datao9_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z1482 : STD_LOGIC; 
  signal romo2datao9_s_4_BXINV : STD_LOGIC; 
  signal romo2datao9_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z1481 : STD_LOGIC; 
  signal romo2datao9_s_4_BYINV : STD_LOGIC; 
  signal nx53675z1477_F5MUX : STD_LOGIC; 
  signal nx53675z1479 : STD_LOGIC; 
  signal nx53675z1477_BXINV : STD_LOGIC; 
  signal nx53675z1478 : STD_LOGIC; 
  signal romo2datao9_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z1488 : STD_LOGIC; 
  signal romo2datao9_s_3_BXINV : STD_LOGIC; 
  signal romo2datao9_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z1487 : STD_LOGIC; 
  signal romo2datao9_s_3_BYINV : STD_LOGIC; 
  signal nx53675z1483_F5MUX : STD_LOGIC; 
  signal nx53675z1485 : STD_LOGIC; 
  signal nx53675z1483_BXINV : STD_LOGIC; 
  signal nx53675z1484 : STD_LOGIC; 
  signal romo2datao8_s_0_F5MUX : STD_LOGIC; 
  signal nx53675z1423 : STD_LOGIC; 
  signal romo2datao8_s_0_BXINV : STD_LOGIC; 
  signal romo2datao8_s_0_F6MUX : STD_LOGIC; 
  signal nx53675z1422 : STD_LOGIC; 
  signal romo2datao8_s_0_BYINV : STD_LOGIC; 
  signal U2_ROMO8_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROMO8_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROMO8_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROMO8_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romo2datao4_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z1087 : STD_LOGIC; 
  signal romo2datao4_s_4_BXINV : STD_LOGIC; 
  signal romo2datao4_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z1086 : STD_LOGIC; 
  signal romo2datao4_s_4_BYINV : STD_LOGIC; 
  signal nx53675z1082_F5MUX : STD_LOGIC; 
  signal nx53675z1084 : STD_LOGIC; 
  signal nx53675z1082_BXINV : STD_LOGIC; 
  signal nx53675z1083 : STD_LOGIC; 
  signal rome2datao4_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z288 : STD_LOGIC; 
  signal rome2datao4_s_9_BXINV : STD_LOGIC; 
  signal rome2datao4_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z287 : STD_LOGIC; 
  signal rome2datao4_s_9_BYINV : STD_LOGIC; 
  signal nx53675z283_F5MUX : STD_LOGIC; 
  signal nx53675z285 : STD_LOGIC; 
  signal nx53675z283_BXINV : STD_LOGIC; 
  signal nx53675z284 : STD_LOGIC; 
  signal rome2datao4_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z294 : STD_LOGIC; 
  signal rome2datao4_s_8_BXINV : STD_LOGIC; 
  signal rome2datao4_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z293 : STD_LOGIC; 
  signal rome2datao4_s_8_BYINV : STD_LOGIC; 
  signal nx53675z289_F5MUX : STD_LOGIC; 
  signal nx53675z291 : STD_LOGIC; 
  signal nx53675z289_BXINV : STD_LOGIC; 
  signal nx53675z290 : STD_LOGIC; 
  signal rome2datao4_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z300 : STD_LOGIC; 
  signal rome2datao4_s_7_BXINV : STD_LOGIC; 
  signal rome2datao4_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z299 : STD_LOGIC; 
  signal rome2datao4_s_7_BYINV : STD_LOGIC; 
  signal nx53675z295_F5MUX : STD_LOGIC; 
  signal nx53675z297 : STD_LOGIC; 
  signal nx53675z295_BXINV : STD_LOGIC; 
  signal nx53675z296 : STD_LOGIC; 
  signal rome2datao3_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z211 : STD_LOGIC; 
  signal rome2datao3_s_11_BXINV : STD_LOGIC; 
  signal rome2datao3_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z210 : STD_LOGIC; 
  signal rome2datao3_s_11_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_FFY_RST : STD_LOGIC; 
  signal nx53675z206_F5MUX : STD_LOGIC; 
  signal nx53675z208 : STD_LOGIC; 
  signal nx53675z206_BXINV : STD_LOGIC; 
  signal nx53675z207 : STD_LOGIC; 
  signal rome2datao0_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z23 : STD_LOGIC; 
  signal rome2datao0_s_10_BXINV : STD_LOGIC; 
  signal rome2datao0_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z22 : STD_LOGIC; 
  signal rome2datao0_s_10_BYINV : STD_LOGIC; 
  signal nx53675z18_F5MUX : STD_LOGIC; 
  signal nx53675z20 : STD_LOGIC; 
  signal nx53675z18_BXINV : STD_LOGIC; 
  signal nx53675z19 : STD_LOGIC; 
  signal rome2datao0_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z29 : STD_LOGIC; 
  signal rome2datao0_s_9_BXINV : STD_LOGIC; 
  signal rome2datao0_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z28 : STD_LOGIC; 
  signal rome2datao0_s_9_BYINV : STD_LOGIC; 
  signal nx53675z24_F5MUX : STD_LOGIC; 
  signal nx53675z26 : STD_LOGIC; 
  signal nx53675z24_BXINV : STD_LOGIC; 
  signal nx53675z25 : STD_LOGIC; 
  signal rome2datao9_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z589 : STD_LOGIC; 
  signal rome2datao9_s_13_BXINV : STD_LOGIC; 
  signal rome2datao9_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z588 : STD_LOGIC; 
  signal rome2datao9_s_13_BYINV : STD_LOGIC; 
  signal nx53675z585_F5MUX : STD_LOGIC; 
  signal nx53675z586 : STD_LOGIC; 
  signal nx53675z585_BXINV : STD_LOGIC; 
  signal nx53675z585_G : STD_LOGIC; 
  signal rome2datao8_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z584 : STD_LOGIC; 
  signal rome2datao8_s_2_BXINV : STD_LOGIC; 
  signal rome2datao8_s_2_F6MUX : STD_LOGIC; 
  signal rome2datao8_s_2_G : STD_LOGIC; 
  signal rome2datao8_s_2_BYINV : STD_LOGIC; 
  signal U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROME8_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal rome2datao10_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z660 : STD_LOGIC; 
  signal rome2datao10_s_12_BXINV : STD_LOGIC; 
  signal rome2datao10_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z659 : STD_LOGIC; 
  signal rome2datao10_s_12_BYINV : STD_LOGIC; 
  signal nx53675z655_F5MUX : STD_LOGIC; 
  signal nx53675z657 : STD_LOGIC; 
  signal nx53675z655_BXINV : STD_LOGIC; 
  signal nx53675z656 : STD_LOGIC; 
  signal rome2datao10_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z666 : STD_LOGIC; 
  signal rome2datao10_s_11_BXINV : STD_LOGIC; 
  signal rome2datao10_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z665 : STD_LOGIC; 
  signal rome2datao10_s_11_BYINV : STD_LOGIC; 
  signal nx53675z661_F5MUX : STD_LOGIC; 
  signal nx53675z663 : STD_LOGIC; 
  signal nx53675z661_BXINV : STD_LOGIC; 
  signal nx53675z662 : STD_LOGIC; 
  signal rome2datao2_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z164 : STD_LOGIC; 
  signal rome2datao2_s_8_BXINV : STD_LOGIC; 
  signal rome2datao2_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z163 : STD_LOGIC; 
  signal rome2datao2_s_8_BYINV : STD_LOGIC; 
  signal nx53675z159_F5MUX : STD_LOGIC; 
  signal nx53675z161 : STD_LOGIC; 
  signal nx53675z159_BXINV : STD_LOGIC; 
  signal nx53675z160 : STD_LOGIC; 
  signal rome2datao1_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z99 : STD_LOGIC; 
  signal rome2datao1_s_8_BXINV : STD_LOGIC; 
  signal rome2datao1_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z98 : STD_LOGIC; 
  signal rome2datao1_s_8_BYINV : STD_LOGIC; 
  signal nx53675z94_F5MUX : STD_LOGIC; 
  signal nx53675z96 : STD_LOGIC; 
  signal nx53675z94_BXINV : STD_LOGIC; 
  signal nx53675z95 : STD_LOGIC; 
  signal rome2datao1_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z105 : STD_LOGIC; 
  signal rome2datao1_s_7_BXINV : STD_LOGIC; 
  signal rome2datao1_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z104 : STD_LOGIC; 
  signal rome2datao1_s_7_BYINV : STD_LOGIC; 
  signal nx53675z100_F5MUX : STD_LOGIC; 
  signal nx53675z102 : STD_LOGIC; 
  signal nx53675z100_BXINV : STD_LOGIC; 
  signal nx53675z101 : STD_LOGIC; 
  signal rome2datao1_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z111 : STD_LOGIC; 
  signal rome2datao1_s_6_BXINV : STD_LOGIC; 
  signal rome2datao1_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z110 : STD_LOGIC; 
  signal rome2datao1_s_6_BYINV : STD_LOGIC; 
  signal nx53675z106_F5MUX : STD_LOGIC; 
  signal nx53675z108 : STD_LOGIC; 
  signal nx53675z106_BXINV : STD_LOGIC; 
  signal nx53675z107 : STD_LOGIC; 
  signal rome2datao1_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z117 : STD_LOGIC; 
  signal rome2datao1_s_5_BXINV : STD_LOGIC; 
  signal rome2datao1_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z116 : STD_LOGIC; 
  signal rome2datao1_s_5_BYINV : STD_LOGIC; 
  signal nx53675z112_F5MUX : STD_LOGIC; 
  signal nx53675z114 : STD_LOGIC; 
  signal nx53675z112_BXINV : STD_LOGIC; 
  signal nx53675z113 : STD_LOGIC; 
  signal rome2datao0_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z35 : STD_LOGIC; 
  signal rome2datao0_s_8_BXINV : STD_LOGIC; 
  signal rome2datao0_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z34 : STD_LOGIC; 
  signal rome2datao0_s_8_BYINV : STD_LOGIC; 
  signal nx53675z30_F5MUX : STD_LOGIC; 
  signal nx53675z32 : STD_LOGIC; 
  signal nx53675z30_BXINV : STD_LOGIC; 
  signal nx53675z31 : STD_LOGIC; 
  signal rome2datao0_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z41 : STD_LOGIC; 
  signal rome2datao0_s_7_BXINV : STD_LOGIC; 
  signal rome2datao0_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z40 : STD_LOGIC; 
  signal rome2datao0_s_7_BYINV : STD_LOGIC; 
  signal nx53675z36_F5MUX : STD_LOGIC; 
  signal nx53675z38 : STD_LOGIC; 
  signal nx53675z36_BXINV : STD_LOGIC; 
  signal nx53675z37 : STD_LOGIC; 
  signal rome2datao0_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z47 : STD_LOGIC; 
  signal rome2datao0_s_6_BXINV : STD_LOGIC; 
  signal rome2datao0_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z46 : STD_LOGIC; 
  signal rome2datao0_s_6_BYINV : STD_LOGIC; 
  signal nx53675z42_F5MUX : STD_LOGIC; 
  signal nx53675z44 : STD_LOGIC; 
  signal nx53675z42_BXINV : STD_LOGIC; 
  signal nx53675z43 : STD_LOGIC; 
  signal rome2datao0_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z53 : STD_LOGIC; 
  signal rome2datao0_s_5_BXINV : STD_LOGIC; 
  signal rome2datao0_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z52 : STD_LOGIC; 
  signal rome2datao0_s_5_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_0_FFX_RST : STD_LOGIC; 
  signal nx53675z48_F5MUX : STD_LOGIC; 
  signal nx53675z50 : STD_LOGIC; 
  signal nx53675z48_BXINV : STD_LOGIC; 
  signal nx53675z49 : STD_LOGIC; 
  signal rome2datao0_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z59 : STD_LOGIC; 
  signal rome2datao0_s_4_BXINV : STD_LOGIC; 
  signal rome2datao0_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z58 : STD_LOGIC; 
  signal rome2datao0_s_4_BYINV : STD_LOGIC; 
  signal nx53675z54_F5MUX : STD_LOGIC; 
  signal nx53675z56 : STD_LOGIC; 
  signal nx53675z54_BXINV : STD_LOGIC; 
  signal nx53675z55 : STD_LOGIC; 
  signal rome2datao9_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z595 : STD_LOGIC; 
  signal rome2datao9_s_12_BXINV : STD_LOGIC; 
  signal rome2datao9_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z594 : STD_LOGIC; 
  signal rome2datao9_s_12_BYINV : STD_LOGIC; 
  signal nx53675z590_F5MUX : STD_LOGIC; 
  signal nx53675z592 : STD_LOGIC; 
  signal nx53675z590_BXINV : STD_LOGIC; 
  signal nx53675z591 : STD_LOGIC; 
  signal rome2datao9_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z601 : STD_LOGIC; 
  signal rome2datao9_s_11_BXINV : STD_LOGIC; 
  signal rome2datao9_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z600 : STD_LOGIC; 
  signal rome2datao9_s_11_BYINV : STD_LOGIC; 
  signal nx53675z596_F5MUX : STD_LOGIC; 
  signal nx53675z598 : STD_LOGIC; 
  signal nx53675z596_BXINV : STD_LOGIC; 
  signal nx53675z597 : STD_LOGIC; 
  signal rome2datao9_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z607 : STD_LOGIC; 
  signal rome2datao9_s_10_BXINV : STD_LOGIC; 
  signal rome2datao9_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z606 : STD_LOGIC; 
  signal rome2datao9_s_10_BYINV : STD_LOGIC; 
  signal nx53675z602_F5MUX : STD_LOGIC; 
  signal nx53675z604 : STD_LOGIC; 
  signal nx53675z602_BXINV : STD_LOGIC; 
  signal nx53675z603 : STD_LOGIC; 
  signal rome2datao9_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z613 : STD_LOGIC; 
  signal rome2datao9_s_9_BXINV : STD_LOGIC; 
  signal rome2datao9_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z612 : STD_LOGIC; 
  signal rome2datao9_s_9_BYINV : STD_LOGIC; 
  signal nx53675z608_F5MUX : STD_LOGIC; 
  signal nx53675z610 : STD_LOGIC; 
  signal nx53675z608_BXINV : STD_LOGIC; 
  signal nx53675z609 : STD_LOGIC; 
  signal rome2datao9_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z619 : STD_LOGIC; 
  signal rome2datao9_s_8_BXINV : STD_LOGIC; 
  signal rome2datao9_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z618 : STD_LOGIC; 
  signal rome2datao9_s_8_BYINV : STD_LOGIC; 
  signal nx53675z614_F5MUX : STD_LOGIC; 
  signal nx53675z616 : STD_LOGIC; 
  signal nx53675z614_BXINV : STD_LOGIC; 
  signal nx53675z615 : STD_LOGIC; 
  signal romo2datao1_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z796 : STD_LOGIC; 
  signal romo2datao1_s_13_BXINV : STD_LOGIC; 
  signal romo2datao1_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z795 : STD_LOGIC; 
  signal romo2datao1_s_13_BYINV : STD_LOGIC; 
  signal nx53675z792_F5MUX : STD_LOGIC; 
  signal nx53675z793 : STD_LOGIC; 
  signal nx53675z792_BXINV : STD_LOGIC; 
  signal nx53675z792_G : STD_LOGIC; 
  signal romo2datao0_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z725 : STD_LOGIC; 
  signal romo2datao0_s_12_BXINV : STD_LOGIC; 
  signal romo2datao0_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z724 : STD_LOGIC; 
  signal romo2datao0_s_12_BYINV : STD_LOGIC; 
  signal nx53675z720_F5MUX : STD_LOGIC; 
  signal nx53675z722 : STD_LOGIC; 
  signal nx53675z720_BXINV : STD_LOGIC; 
  signal nx53675z721 : STD_LOGIC; 
  signal romo2datao0_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z731 : STD_LOGIC; 
  signal romo2datao0_s_11_BXINV : STD_LOGIC; 
  signal romo2datao0_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z730 : STD_LOGIC; 
  signal romo2datao0_s_11_BYINV : STD_LOGIC; 
  signal nx53675z726_F5MUX : STD_LOGIC; 
  signal nx53675z728 : STD_LOGIC; 
  signal nx53675z726_BXINV : STD_LOGIC; 
  signal nx53675z727 : STD_LOGIC; 
  signal romo2datao0_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z737 : STD_LOGIC; 
  signal romo2datao0_s_10_BXINV : STD_LOGIC; 
  signal romo2datao0_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z736 : STD_LOGIC; 
  signal romo2datao0_s_10_BYINV : STD_LOGIC; 
  signal nx53675z732_F5MUX : STD_LOGIC; 
  signal nx53675z734 : STD_LOGIC; 
  signal nx53675z732_BXINV : STD_LOGIC; 
  signal nx53675z733 : STD_LOGIC; 
  signal romo2datao7_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z1294 : STD_LOGIC; 
  signal romo2datao7_s_9_BXINV : STD_LOGIC; 
  signal romo2datao7_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z1293 : STD_LOGIC; 
  signal romo2datao7_s_9_BYINV : STD_LOGIC; 
  signal nx53675z1289_F5MUX : STD_LOGIC; 
  signal nx53675z1291 : STD_LOGIC; 
  signal nx53675z1289_BXINV : STD_LOGIC; 
  signal nx53675z1290 : STD_LOGIC; 
  signal romo2datao7_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z1300 : STD_LOGIC; 
  signal romo2datao7_s_8_BXINV : STD_LOGIC; 
  signal romo2datao7_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z1299 : STD_LOGIC; 
  signal romo2datao7_s_8_BYINV : STD_LOGIC; 
  signal nx53675z1295_F5MUX : STD_LOGIC; 
  signal nx53675z1297 : STD_LOGIC; 
  signal nx53675z1295_BXINV : STD_LOGIC; 
  signal nx53675z1296 : STD_LOGIC; 
  signal romo2datao7_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z1306 : STD_LOGIC; 
  signal romo2datao7_s_7_BXINV : STD_LOGIC; 
  signal romo2datao7_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z1305 : STD_LOGIC; 
  signal romo2datao7_s_7_BYINV : STD_LOGIC; 
  signal nx53675z1301_F5MUX : STD_LOGIC; 
  signal nx53675z1303 : STD_LOGIC; 
  signal nx53675z1301_BXINV : STD_LOGIC; 
  signal nx53675z1302 : STD_LOGIC; 
  signal romo2datao7_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z1312 : STD_LOGIC; 
  signal romo2datao7_s_6_BXINV : STD_LOGIC; 
  signal romo2datao7_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z1311 : STD_LOGIC; 
  signal romo2datao7_s_6_BYINV : STD_LOGIC; 
  signal nx53675z1307_F5MUX : STD_LOGIC; 
  signal nx53675z1309 : STD_LOGIC; 
  signal nx53675z1307_BXINV : STD_LOGIC; 
  signal nx53675z1308 : STD_LOGIC; 
  signal romo2datao8_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z1361 : STD_LOGIC; 
  signal romo2datao8_s_11_BXINV : STD_LOGIC; 
  signal romo2datao8_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z1360 : STD_LOGIC; 
  signal romo2datao8_s_11_BYINV : STD_LOGIC; 
  signal nx53675z1356_F5MUX : STD_LOGIC; 
  signal nx53675z1358 : STD_LOGIC; 
  signal nx53675z1356_BXINV : STD_LOGIC; 
  signal nx53675z1357 : STD_LOGIC; 
  signal romo2datao8_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z1367 : STD_LOGIC; 
  signal romo2datao8_s_10_BXINV : STD_LOGIC; 
  signal romo2datao8_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z1366 : STD_LOGIC; 
  signal romo2datao8_s_10_BYINV : STD_LOGIC; 
  signal nx53675z1362_F5MUX : STD_LOGIC; 
  signal nx53675z1364 : STD_LOGIC; 
  signal nx53675z1362_BXINV : STD_LOGIC; 
  signal nx53675z1363 : STD_LOGIC; 
  signal rome2datao10_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z672 : STD_LOGIC; 
  signal rome2datao10_s_10_BXINV : STD_LOGIC; 
  signal rome2datao10_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z671 : STD_LOGIC; 
  signal rome2datao10_s_10_BYINV : STD_LOGIC; 
  signal nx53675z667_F5MUX : STD_LOGIC; 
  signal nx53675z669 : STD_LOGIC; 
  signal nx53675z667_BXINV : STD_LOGIC; 
  signal nx53675z668 : STD_LOGIC; 
  signal rome2datao10_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z678 : STD_LOGIC; 
  signal rome2datao10_s_9_BXINV : STD_LOGIC; 
  signal rome2datao10_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z677 : STD_LOGIC; 
  signal rome2datao10_s_9_BYINV : STD_LOGIC; 
  signal nx53675z673_F5MUX : STD_LOGIC; 
  signal nx53675z675 : STD_LOGIC; 
  signal nx53675z673_BXINV : STD_LOGIC; 
  signal nx53675z674 : STD_LOGIC; 
  signal rome2datao10_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z684 : STD_LOGIC; 
  signal rome2datao10_s_8_BXINV : STD_LOGIC; 
  signal rome2datao10_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z683 : STD_LOGIC; 
  signal rome2datao10_s_8_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_FFY_RST : STD_LOGIC; 
  signal nx53675z679_F5MUX : STD_LOGIC; 
  signal nx53675z681 : STD_LOGIC; 
  signal nx53675z679_BXINV : STD_LOGIC; 
  signal nx53675z680 : STD_LOGIC; 
  signal rome2datao10_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z690 : STD_LOGIC; 
  signal rome2datao10_s_7_BXINV : STD_LOGIC; 
  signal rome2datao10_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z689 : STD_LOGIC; 
  signal rome2datao10_s_7_BYINV : STD_LOGIC; 
  signal nx53675z685_F5MUX : STD_LOGIC; 
  signal nx53675z687 : STD_LOGIC; 
  signal nx53675z685_BXINV : STD_LOGIC; 
  signal nx53675z686 : STD_LOGIC; 
  signal rome2datao10_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z696 : STD_LOGIC; 
  signal rome2datao10_s_6_BXINV : STD_LOGIC; 
  signal rome2datao10_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z695 : STD_LOGIC; 
  signal rome2datao10_s_6_BYINV : STD_LOGIC; 
  signal nx53675z691_F5MUX : STD_LOGIC; 
  signal nx53675z693 : STD_LOGIC; 
  signal nx53675z691_BXINV : STD_LOGIC; 
  signal nx53675z692 : STD_LOGIC; 
  signal rome2datao2_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z170 : STD_LOGIC; 
  signal rome2datao2_s_7_BXINV : STD_LOGIC; 
  signal rome2datao2_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z169 : STD_LOGIC; 
  signal rome2datao2_s_7_BYINV : STD_LOGIC; 
  signal nx53675z165_F5MUX : STD_LOGIC; 
  signal nx53675z167 : STD_LOGIC; 
  signal nx53675z165_BXINV : STD_LOGIC; 
  signal nx53675z166 : STD_LOGIC; 
  signal rome2datao2_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z176 : STD_LOGIC; 
  signal rome2datao2_s_6_BXINV : STD_LOGIC; 
  signal rome2datao2_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z175 : STD_LOGIC; 
  signal rome2datao2_s_6_BYINV : STD_LOGIC; 
  signal nx53675z171_F5MUX : STD_LOGIC; 
  signal nx53675z173 : STD_LOGIC; 
  signal nx53675z171_BXINV : STD_LOGIC; 
  signal nx53675z172 : STD_LOGIC; 
  signal rome2datao2_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z182 : STD_LOGIC; 
  signal rome2datao2_s_5_BXINV : STD_LOGIC; 
  signal rome2datao2_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z181 : STD_LOGIC; 
  signal rome2datao2_s_5_BYINV : STD_LOGIC; 
  signal nx53675z177_F5MUX : STD_LOGIC; 
  signal nx53675z179 : STD_LOGIC; 
  signal nx53675z177_BXINV : STD_LOGIC; 
  signal nx53675z178 : STD_LOGIC; 
  signal rome2datao2_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z188 : STD_LOGIC; 
  signal rome2datao2_s_4_BXINV : STD_LOGIC; 
  signal rome2datao2_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z187 : STD_LOGIC; 
  signal rome2datao2_s_4_BYINV : STD_LOGIC; 
  signal nx53675z183_F5MUX : STD_LOGIC; 
  signal nx53675z185 : STD_LOGIC; 
  signal nx53675z183_BXINV : STD_LOGIC; 
  signal nx53675z184 : STD_LOGIC; 
  signal rome2datao2_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z193 : STD_LOGIC; 
  signal rome2datao2_s_3_BXINV : STD_LOGIC; 
  signal rome2datao2_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z192 : STD_LOGIC; 
  signal rome2datao2_s_3_BYINV : STD_LOGIC; 
  signal nx53675z189_F5MUX : STD_LOGIC; 
  signal nx53675z190 : STD_LOGIC; 
  signal nx53675z189_BXINV : STD_LOGIC; 
  signal U2_ROME2_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal rome2datao2_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z134 : STD_LOGIC; 
  signal rome2datao2_s_13_BXINV : STD_LOGIC; 
  signal rome2datao2_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z133 : STD_LOGIC; 
  signal rome2datao2_s_13_BYINV : STD_LOGIC; 
  signal nx53675z130_F5MUX : STD_LOGIC; 
  signal nx53675z131 : STD_LOGIC; 
  signal nx53675z130_BXINV : STD_LOGIC; 
  signal nx53675z130_G : STD_LOGIC; 
  signal rome2datao1_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z75 : STD_LOGIC; 
  signal rome2datao1_s_12_BXINV : STD_LOGIC; 
  signal rome2datao1_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z74 : STD_LOGIC; 
  signal rome2datao1_s_12_BYINV : STD_LOGIC; 
  signal nx53675z70_F5MUX : STD_LOGIC; 
  signal nx53675z72 : STD_LOGIC; 
  signal nx53675z70_BXINV : STD_LOGIC; 
  signal nx53675z71 : STD_LOGIC; 
  signal romo2datao9_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z1428 : STD_LOGIC; 
  signal romo2datao9_s_13_BXINV : STD_LOGIC; 
  signal romo2datao9_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z1427 : STD_LOGIC; 
  signal romo2datao9_s_13_BYINV : STD_LOGIC; 
  signal nx53675z1424_F5MUX : STD_LOGIC; 
  signal nx53675z1425 : STD_LOGIC; 
  signal nx53675z1424_BXINV : STD_LOGIC; 
  signal nx53675z1424_G : STD_LOGIC; 
  signal rome2datao10_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z654 : STD_LOGIC; 
  signal rome2datao10_s_13_BXINV : STD_LOGIC; 
  signal rome2datao10_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z653 : STD_LOGIC; 
  signal rome2datao10_s_13_BYINV : STD_LOGIC; 
  signal nx53675z650_F5MUX : STD_LOGIC; 
  signal nx53675z651 : STD_LOGIC; 
  signal nx53675z650_BXINV : STD_LOGIC; 
  signal nx53675z650_G : STD_LOGIC; 
  signal rome2datao4_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z306 : STD_LOGIC; 
  signal rome2datao4_s_6_BXINV : STD_LOGIC; 
  signal rome2datao4_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z305 : STD_LOGIC; 
  signal rome2datao4_s_6_BYINV : STD_LOGIC; 
  signal nx53675z301_F5MUX : STD_LOGIC; 
  signal nx53675z303 : STD_LOGIC; 
  signal nx53675z301_BXINV : STD_LOGIC; 
  signal nx53675z302 : STD_LOGIC; 
  signal rome2datao4_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z312 : STD_LOGIC; 
  signal rome2datao4_s_5_BXINV : STD_LOGIC; 
  signal rome2datao4_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z311 : STD_LOGIC; 
  signal rome2datao4_s_5_BYINV : STD_LOGIC; 
  signal nx53675z307_F5MUX : STD_LOGIC; 
  signal nx53675z309 : STD_LOGIC; 
  signal nx53675z307_BXINV : STD_LOGIC; 
  signal nx53675z308 : STD_LOGIC; 
  signal rome2datao1_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z69 : STD_LOGIC; 
  signal rome2datao1_s_13_BXINV : STD_LOGIC; 
  signal rome2datao1_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z68 : STD_LOGIC; 
  signal rome2datao1_s_13_BYINV : STD_LOGIC; 
  signal nx53675z65_F5MUX : STD_LOGIC; 
  signal nx53675z66 : STD_LOGIC; 
  signal nx53675z65_BXINV : STD_LOGIC; 
  signal nx53675z65_G : STD_LOGIC; 
  signal rome2datao1_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z81 : STD_LOGIC; 
  signal rome2datao1_s_11_BXINV : STD_LOGIC; 
  signal rome2datao1_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z80 : STD_LOGIC; 
  signal rome2datao1_s_11_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_2_FFX_RST : STD_LOGIC; 
  signal nx53675z76_F5MUX : STD_LOGIC; 
  signal nx53675z78 : STD_LOGIC; 
  signal nx53675z76_BXINV : STD_LOGIC; 
  signal nx53675z77 : STD_LOGIC; 
  signal rome2datao1_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z87 : STD_LOGIC; 
  signal rome2datao1_s_10_BXINV : STD_LOGIC; 
  signal rome2datao1_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z86 : STD_LOGIC; 
  signal rome2datao1_s_10_BYINV : STD_LOGIC; 
  signal nx53675z82_F5MUX : STD_LOGIC; 
  signal nx53675z84 : STD_LOGIC; 
  signal nx53675z82_BXINV : STD_LOGIC; 
  signal nx53675z83 : STD_LOGIC; 
  signal rome2datao1_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z123 : STD_LOGIC; 
  signal rome2datao1_s_4_BXINV : STD_LOGIC; 
  signal rome2datao1_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z122 : STD_LOGIC; 
  signal rome2datao1_s_4_BYINV : STD_LOGIC; 
  signal nx53675z118_F5MUX : STD_LOGIC; 
  signal nx53675z120 : STD_LOGIC; 
  signal nx53675z118_BXINV : STD_LOGIC; 
  signal nx53675z119 : STD_LOGIC; 
  signal rome2datao1_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z128 : STD_LOGIC; 
  signal rome2datao1_s_3_BXINV : STD_LOGIC; 
  signal rome2datao1_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z127 : STD_LOGIC; 
  signal rome2datao1_s_3_BYINV : STD_LOGIC; 
  signal nx53675z124_F5MUX : STD_LOGIC; 
  signal nx53675z125 : STD_LOGIC; 
  signal nx53675z124_BXINV : STD_LOGIC; 
  signal U2_ROME1_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal rome2datao1_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z129 : STD_LOGIC; 
  signal rome2datao1_s_2_BXINV : STD_LOGIC; 
  signal rome2datao1_s_2_F6MUX : STD_LOGIC; 
  signal rome2datao1_s_2_G : STD_LOGIC; 
  signal rome2datao1_s_2_BYINV : STD_LOGIC; 
  signal U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROME1_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal rome2datao0_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z11 : STD_LOGIC; 
  signal rome2datao0_s_12_BXINV : STD_LOGIC; 
  signal rome2datao0_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z10 : STD_LOGIC; 
  signal rome2datao0_s_12_BYINV : STD_LOGIC; 
  signal nx53675z6_F5MUX : STD_LOGIC; 
  signal nx53675z8 : STD_LOGIC; 
  signal nx53675z6_BXINV : STD_LOGIC; 
  signal nx53675z7 : STD_LOGIC; 
  signal rome2datao0_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z17 : STD_LOGIC; 
  signal rome2datao0_s_11_BXINV : STD_LOGIC; 
  signal rome2datao0_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z16 : STD_LOGIC; 
  signal rome2datao0_s_11_BYINV : STD_LOGIC; 
  signal nx53675z12_F5MUX : STD_LOGIC; 
  signal nx53675z14 : STD_LOGIC; 
  signal nx53675z12_BXINV : STD_LOGIC; 
  signal nx53675z13 : STD_LOGIC; 
  signal rome2datao0_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z64 : STD_LOGIC; 
  signal rome2datao0_s_3_BXINV : STD_LOGIC; 
  signal rome2datao0_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z63 : STD_LOGIC; 
  signal rome2datao0_s_3_BYINV : STD_LOGIC; 
  signal nx53675z60_F5MUX : STD_LOGIC; 
  signal nx53675z61 : STD_LOGIC; 
  signal nx53675z60_BXINV : STD_LOGIC; 
  signal U2_ROME0_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal rome2datao9_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z625 : STD_LOGIC; 
  signal rome2datao9_s_7_BXINV : STD_LOGIC; 
  signal rome2datao9_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z624 : STD_LOGIC; 
  signal rome2datao9_s_7_BYINV : STD_LOGIC; 
  signal nx53675z620_F5MUX : STD_LOGIC; 
  signal nx53675z622 : STD_LOGIC; 
  signal nx53675z620_BXINV : STD_LOGIC; 
  signal nx53675z621 : STD_LOGIC; 
  signal rome2datao9_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z631 : STD_LOGIC; 
  signal rome2datao9_s_6_BXINV : STD_LOGIC; 
  signal rome2datao9_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z630 : STD_LOGIC; 
  signal rome2datao9_s_6_BYINV : STD_LOGIC; 
  signal nx53675z626_F5MUX : STD_LOGIC; 
  signal nx53675z628 : STD_LOGIC; 
  signal nx53675z626_BXINV : STD_LOGIC; 
  signal nx53675z627 : STD_LOGIC; 
  signal rome2datao9_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z637 : STD_LOGIC; 
  signal rome2datao9_s_5_BXINV : STD_LOGIC; 
  signal rome2datao9_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z636 : STD_LOGIC; 
  signal rome2datao9_s_5_BYINV : STD_LOGIC; 
  signal nx53675z632_F5MUX : STD_LOGIC; 
  signal nx53675z634 : STD_LOGIC; 
  signal nx53675z632_BXINV : STD_LOGIC; 
  signal nx53675z633 : STD_LOGIC; 
  signal rome2datao9_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z643 : STD_LOGIC; 
  signal rome2datao9_s_4_BXINV : STD_LOGIC; 
  signal rome2datao9_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z642 : STD_LOGIC; 
  signal rome2datao9_s_4_BYINV : STD_LOGIC; 
  signal nx53675z638_F5MUX : STD_LOGIC; 
  signal nx53675z640 : STD_LOGIC; 
  signal nx53675z638_BXINV : STD_LOGIC; 
  signal nx53675z639 : STD_LOGIC; 
  signal rome2datao9_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z648 : STD_LOGIC; 
  signal rome2datao9_s_3_BXINV : STD_LOGIC; 
  signal rome2datao9_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z647 : STD_LOGIC; 
  signal rome2datao9_s_3_BYINV : STD_LOGIC; 
  signal nx53675z644_F5MUX : STD_LOGIC; 
  signal nx53675z645 : STD_LOGIC; 
  signal nx53675z644_BXINV : STD_LOGIC; 
  signal U2_ROME9_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal rome2datao0_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z5 : STD_LOGIC; 
  signal rome2datao0_s_13_BXINV : STD_LOGIC; 
  signal rome2datao0_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z4 : STD_LOGIC; 
  signal rome2datao0_s_13_BYINV : STD_LOGIC; 
  signal nx53675z1_F5MUX : STD_LOGIC; 
  signal nx53675z2 : STD_LOGIC; 
  signal nx53675z1_BXINV : STD_LOGIC; 
  signal nx53675z1_G : STD_LOGIC; 
  signal romo2datao2_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z875 : STD_LOGIC; 
  signal romo2datao2_s_13_BXINV : STD_LOGIC; 
  signal romo2datao2_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z874 : STD_LOGIC; 
  signal romo2datao2_s_13_BYINV : STD_LOGIC; 
  signal nx53675z871_F5MUX : STD_LOGIC; 
  signal nx53675z872 : STD_LOGIC; 
  signal nx53675z871_BXINV : STD_LOGIC; 
  signal nx53675z871_G : STD_LOGIC; 
  signal romo2datao2_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z941 : STD_LOGIC; 
  signal romo2datao2_s_2_BXINV : STD_LOGIC; 
  signal romo2datao2_s_2_F6MUX : STD_LOGIC; 
  signal nx53675z940 : STD_LOGIC; 
  signal romo2datao2_s_2_BYINV : STD_LOGIC; 
  signal nx53675z936_F5MUX : STD_LOGIC; 
  signal nx53675z938 : STD_LOGIC; 
  signal nx53675z936_BXINV : STD_LOGIC; 
  signal nx53675z937 : STD_LOGIC; 
  signal romo2datao1_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z802 : STD_LOGIC; 
  signal romo2datao1_s_12_BXINV : STD_LOGIC; 
  signal romo2datao1_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z801 : STD_LOGIC; 
  signal romo2datao1_s_12_BYINV : STD_LOGIC; 
  signal nx53675z797_F5MUX : STD_LOGIC; 
  signal nx53675z799 : STD_LOGIC; 
  signal nx53675z797_BXINV : STD_LOGIC; 
  signal nx53675z798 : STD_LOGIC; 
  signal romo2datao1_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z808 : STD_LOGIC; 
  signal romo2datao1_s_11_BXINV : STD_LOGIC; 
  signal romo2datao1_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z807 : STD_LOGIC; 
  signal romo2datao1_s_11_BYINV : STD_LOGIC; 
  signal nx53675z803_F5MUX : STD_LOGIC; 
  signal nx53675z805 : STD_LOGIC; 
  signal nx53675z803_BXINV : STD_LOGIC; 
  signal nx53675z804 : STD_LOGIC; 
  signal romo2datao1_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z814 : STD_LOGIC; 
  signal romo2datao1_s_10_BXINV : STD_LOGIC; 
  signal romo2datao1_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z813 : STD_LOGIC; 
  signal romo2datao1_s_10_BYINV : STD_LOGIC; 
  signal nx53675z809_F5MUX : STD_LOGIC; 
  signal nx53675z811 : STD_LOGIC; 
  signal nx53675z809_BXINV : STD_LOGIC; 
  signal nx53675z810 : STD_LOGIC; 
  signal romo2datao1_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z820 : STD_LOGIC; 
  signal romo2datao1_s_9_BXINV : STD_LOGIC; 
  signal romo2datao1_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z819 : STD_LOGIC; 
  signal romo2datao1_s_9_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_FFY_RST : STD_LOGIC; 
  signal nx53675z815_F5MUX : STD_LOGIC; 
  signal nx53675z817 : STD_LOGIC; 
  signal nx53675z815_BXINV : STD_LOGIC; 
  signal nx53675z816 : STD_LOGIC; 
  signal romo2datao1_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z826 : STD_LOGIC; 
  signal romo2datao1_s_8_BXINV : STD_LOGIC; 
  signal romo2datao1_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z825 : STD_LOGIC; 
  signal romo2datao1_s_8_BYINV : STD_LOGIC; 
  signal nx53675z821_F5MUX : STD_LOGIC; 
  signal nx53675z823 : STD_LOGIC; 
  signal nx53675z821_BXINV : STD_LOGIC; 
  signal nx53675z822 : STD_LOGIC; 
  signal romo2datao1_s_0_F5MUX : STD_LOGIC; 
  signal nx53675z870 : STD_LOGIC; 
  signal romo2datao1_s_0_BXINV : STD_LOGIC; 
  signal romo2datao1_s_0_F6MUX : STD_LOGIC; 
  signal nx53675z869 : STD_LOGIC; 
  signal romo2datao1_s_0_BYINV : STD_LOGIC; 
  signal U2_ROMO1_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROMO1_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROMO1_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROMO1_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romo2datao0_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z743 : STD_LOGIC; 
  signal romo2datao0_s_9_BXINV : STD_LOGIC; 
  signal romo2datao0_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z742 : STD_LOGIC; 
  signal romo2datao0_s_9_BYINV : STD_LOGIC; 
  signal nx53675z738_F5MUX : STD_LOGIC; 
  signal nx53675z740 : STD_LOGIC; 
  signal nx53675z738_BXINV : STD_LOGIC; 
  signal nx53675z739 : STD_LOGIC; 
  signal romo2datao0_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z749 : STD_LOGIC; 
  signal romo2datao0_s_8_BXINV : STD_LOGIC; 
  signal romo2datao0_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z748 : STD_LOGIC; 
  signal romo2datao0_s_8_BYINV : STD_LOGIC; 
  signal nx53675z744_F5MUX : STD_LOGIC; 
  signal nx53675z746 : STD_LOGIC; 
  signal nx53675z744_BXINV : STD_LOGIC; 
  signal nx53675z745 : STD_LOGIC; 
  signal romo2datao0_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z755 : STD_LOGIC; 
  signal romo2datao0_s_7_BXINV : STD_LOGIC; 
  signal romo2datao0_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z754 : STD_LOGIC; 
  signal romo2datao0_s_7_BYINV : STD_LOGIC; 
  signal nx53675z750_F5MUX : STD_LOGIC; 
  signal nx53675z752 : STD_LOGIC; 
  signal nx53675z750_BXINV : STD_LOGIC; 
  signal nx53675z751 : STD_LOGIC; 
  signal romo2datao0_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z761 : STD_LOGIC; 
  signal romo2datao0_s_6_BXINV : STD_LOGIC; 
  signal romo2datao0_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z760 : STD_LOGIC; 
  signal romo2datao0_s_6_BYINV : STD_LOGIC; 
  signal nx53675z756_F5MUX : STD_LOGIC; 
  signal nx53675z758 : STD_LOGIC; 
  signal nx53675z756_BXINV : STD_LOGIC; 
  signal nx53675z757 : STD_LOGIC; 
  signal romo2datao0_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z767 : STD_LOGIC; 
  signal romo2datao0_s_5_BXINV : STD_LOGIC; 
  signal romo2datao0_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z766 : STD_LOGIC; 
  signal romo2datao0_s_5_BYINV : STD_LOGIC; 
  signal nx53675z762_F5MUX : STD_LOGIC; 
  signal nx53675z764 : STD_LOGIC; 
  signal nx53675z762_BXINV : STD_LOGIC; 
  signal nx53675z763 : STD_LOGIC; 
  signal rome2datao3_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z205 : STD_LOGIC; 
  signal rome2datao3_s_12_BXINV : STD_LOGIC; 
  signal rome2datao3_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z204 : STD_LOGIC; 
  signal rome2datao3_s_12_BYINV : STD_LOGIC; 
  signal nx53675z200_F5MUX : STD_LOGIC; 
  signal nx53675z202 : STD_LOGIC; 
  signal nx53675z200_BXINV : STD_LOGIC; 
  signal nx53675z201 : STD_LOGIC; 
  signal rome2datao3_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z241 : STD_LOGIC; 
  signal rome2datao3_s_6_BXINV : STD_LOGIC; 
  signal rome2datao3_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z240 : STD_LOGIC; 
  signal rome2datao3_s_6_BYINV : STD_LOGIC; 
  signal nx53675z236_F5MUX : STD_LOGIC; 
  signal nx53675z238 : STD_LOGIC; 
  signal nx53675z236_BXINV : STD_LOGIC; 
  signal nx53675z237 : STD_LOGIC; 
  signal rome2datao3_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z253 : STD_LOGIC; 
  signal rome2datao3_s_4_BXINV : STD_LOGIC; 
  signal rome2datao3_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z252 : STD_LOGIC; 
  signal rome2datao3_s_4_BYINV : STD_LOGIC; 
  signal nx53675z248_F5MUX : STD_LOGIC; 
  signal nx53675z250 : STD_LOGIC; 
  signal nx53675z248_BXINV : STD_LOGIC; 
  signal nx53675z249 : STD_LOGIC; 
  signal rome2datao3_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z259 : STD_LOGIC; 
  signal rome2datao3_s_2_BXINV : STD_LOGIC; 
  signal rome2datao3_s_2_F6MUX : STD_LOGIC; 
  signal rome2datao3_s_2_G : STD_LOGIC; 
  signal rome2datao3_s_2_BYINV : STD_LOGIC; 
  signal U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROME3_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romo2datao3_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z1014 : STD_LOGIC; 
  signal romo2datao3_s_3_BXINV : STD_LOGIC; 
  signal romo2datao3_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z1013 : STD_LOGIC; 
  signal romo2datao3_s_3_BYINV : STD_LOGIC; 
  signal nx53675z1009_F5MUX : STD_LOGIC; 
  signal nx53675z1011 : STD_LOGIC; 
  signal nx53675z1009_BXINV : STD_LOGIC; 
  signal nx53675z1010 : STD_LOGIC; 
  signal rome2datao3_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z199 : STD_LOGIC; 
  signal rome2datao3_s_13_BXINV : STD_LOGIC; 
  signal rome2datao3_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z198 : STD_LOGIC; 
  signal rome2datao3_s_13_BYINV : STD_LOGIC; 
  signal nx53675z195_F5MUX : STD_LOGIC; 
  signal nx53675z196 : STD_LOGIC; 
  signal nx53675z195_BXINV : STD_LOGIC; 
  signal nx53675z195_G : STD_LOGIC; 
  signal romo2datao8_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z1373 : STD_LOGIC; 
  signal romo2datao8_s_9_BXINV : STD_LOGIC; 
  signal romo2datao8_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z1372 : STD_LOGIC; 
  signal romo2datao8_s_9_BYINV : STD_LOGIC; 
  signal nx53675z1368_F5MUX : STD_LOGIC; 
  signal nx53675z1370 : STD_LOGIC; 
  signal nx53675z1368_BXINV : STD_LOGIC; 
  signal nx53675z1369 : STD_LOGIC; 
  signal romo2datao8_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z1379 : STD_LOGIC; 
  signal romo2datao8_s_8_BXINV : STD_LOGIC; 
  signal romo2datao8_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z1378 : STD_LOGIC; 
  signal romo2datao8_s_8_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_4_FFX_RST : STD_LOGIC; 
  signal nx53675z1374_F5MUX : STD_LOGIC; 
  signal nx53675z1376 : STD_LOGIC; 
  signal nx53675z1374_BXINV : STD_LOGIC; 
  signal nx53675z1375 : STD_LOGIC; 
  signal romo2datao8_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z1385 : STD_LOGIC; 
  signal romo2datao8_s_7_BXINV : STD_LOGIC; 
  signal romo2datao8_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z1384 : STD_LOGIC; 
  signal romo2datao8_s_7_BYINV : STD_LOGIC; 
  signal nx53675z1380_F5MUX : STD_LOGIC; 
  signal nx53675z1382 : STD_LOGIC; 
  signal nx53675z1380_BXINV : STD_LOGIC; 
  signal nx53675z1381 : STD_LOGIC; 
  signal romo2datao8_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z1391 : STD_LOGIC; 
  signal romo2datao8_s_6_BXINV : STD_LOGIC; 
  signal romo2datao8_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z1390 : STD_LOGIC; 
  signal romo2datao8_s_6_BYINV : STD_LOGIC; 
  signal nx53675z1386_F5MUX : STD_LOGIC; 
  signal nx53675z1388 : STD_LOGIC; 
  signal nx53675z1386_BXINV : STD_LOGIC; 
  signal nx53675z1387 : STD_LOGIC; 
  signal romo2datao8_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z1397 : STD_LOGIC; 
  signal romo2datao8_s_5_BXINV : STD_LOGIC; 
  signal romo2datao8_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z1396 : STD_LOGIC; 
  signal romo2datao8_s_5_BYINV : STD_LOGIC; 
  signal nx53675z1392_F5MUX : STD_LOGIC; 
  signal nx53675z1394 : STD_LOGIC; 
  signal nx53675z1392_BXINV : STD_LOGIC; 
  signal nx53675z1393 : STD_LOGIC; 
  signal romo2datao7_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z1318 : STD_LOGIC; 
  signal romo2datao7_s_5_BXINV : STD_LOGIC; 
  signal romo2datao7_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z1317 : STD_LOGIC; 
  signal romo2datao7_s_5_BYINV : STD_LOGIC; 
  signal nx53675z1313_F5MUX : STD_LOGIC; 
  signal nx53675z1315 : STD_LOGIC; 
  signal nx53675z1313_BXINV : STD_LOGIC; 
  signal nx53675z1314 : STD_LOGIC; 
  signal romo2datao7_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z1324 : STD_LOGIC; 
  signal romo2datao7_s_4_BXINV : STD_LOGIC; 
  signal romo2datao7_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z1323 : STD_LOGIC; 
  signal romo2datao7_s_4_BYINV : STD_LOGIC; 
  signal nx53675z1319_F5MUX : STD_LOGIC; 
  signal nx53675z1321 : STD_LOGIC; 
  signal nx53675z1319_BXINV : STD_LOGIC; 
  signal nx53675z1320 : STD_LOGIC; 
  signal romo2datao7_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z1330 : STD_LOGIC; 
  signal romo2datao7_s_3_BXINV : STD_LOGIC; 
  signal romo2datao7_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z1329 : STD_LOGIC; 
  signal romo2datao7_s_3_BYINV : STD_LOGIC; 
  signal nx53675z1325_F5MUX : STD_LOGIC; 
  signal nx53675z1327 : STD_LOGIC; 
  signal nx53675z1325_BXINV : STD_LOGIC; 
  signal nx53675z1326 : STD_LOGIC; 
  signal romo2datao7_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z1336 : STD_LOGIC; 
  signal romo2datao7_s_2_BXINV : STD_LOGIC; 
  signal romo2datao7_s_2_F6MUX : STD_LOGIC; 
  signal nx53675z1335 : STD_LOGIC; 
  signal romo2datao7_s_2_BYINV : STD_LOGIC; 
  signal nx53675z1331_F5MUX : STD_LOGIC; 
  signal nx53675z1333 : STD_LOGIC; 
  signal nx53675z1331_BXINV : STD_LOGIC; 
  signal nx53675z1332 : STD_LOGIC; 
  signal romo2datao7_s_1_F5MUX : STD_LOGIC; 
  signal nx53675z1342 : STD_LOGIC; 
  signal romo2datao7_s_1_BXINV : STD_LOGIC; 
  signal romo2datao7_s_1_F6MUX : STD_LOGIC; 
  signal nx53675z1341 : STD_LOGIC; 
  signal romo2datao7_s_1_BYINV : STD_LOGIC; 
  signal nx53675z1337_F5MUX : STD_LOGIC; 
  signal nx53675z1339 : STD_LOGIC; 
  signal nx53675z1337_BXINV : STD_LOGIC; 
  signal nx53675z1338 : STD_LOGIC; 
  signal rome2datao5_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z377 : STD_LOGIC; 
  signal rome2datao5_s_5_BXINV : STD_LOGIC; 
  signal rome2datao5_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z376 : STD_LOGIC; 
  signal rome2datao5_s_5_BYINV : STD_LOGIC; 
  signal nx53675z372_F5MUX : STD_LOGIC; 
  signal nx53675z374 : STD_LOGIC; 
  signal nx53675z372_BXINV : STD_LOGIC; 
  signal nx53675z373 : STD_LOGIC; 
  signal rome2datao5_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z383 : STD_LOGIC; 
  signal rome2datao5_s_4_BXINV : STD_LOGIC; 
  signal rome2datao5_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z382 : STD_LOGIC; 
  signal rome2datao5_s_4_BYINV : STD_LOGIC; 
  signal nx53675z378_F5MUX : STD_LOGIC; 
  signal nx53675z380 : STD_LOGIC; 
  signal nx53675z378_BXINV : STD_LOGIC; 
  signal nx53675z379 : STD_LOGIC; 
  signal romo2datao7_s_0_F5MUX : STD_LOGIC; 
  signal nx53675z1344 : STD_LOGIC; 
  signal romo2datao7_s_0_BXINV : STD_LOGIC; 
  signal romo2datao7_s_0_F6MUX : STD_LOGIC; 
  signal nx53675z1343 : STD_LOGIC; 
  signal romo2datao7_s_0_BYINV : STD_LOGIC; 
  signal U2_ROMO7_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROMO7_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROMO7_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROMO7_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal rome2datao10_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z702 : STD_LOGIC; 
  signal rome2datao10_s_5_BXINV : STD_LOGIC; 
  signal rome2datao10_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z701 : STD_LOGIC; 
  signal rome2datao10_s_5_BYINV : STD_LOGIC; 
  signal nx53675z697_F5MUX : STD_LOGIC; 
  signal nx53675z699 : STD_LOGIC; 
  signal nx53675z697_BXINV : STD_LOGIC; 
  signal nx53675z698 : STD_LOGIC; 
  signal rome2datao10_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z708 : STD_LOGIC; 
  signal rome2datao10_s_4_BXINV : STD_LOGIC; 
  signal rome2datao10_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z707 : STD_LOGIC; 
  signal rome2datao10_s_4_BYINV : STD_LOGIC; 
  signal nx53675z703_F5MUX : STD_LOGIC; 
  signal nx53675z705 : STD_LOGIC; 
  signal nx53675z703_BXINV : STD_LOGIC; 
  signal nx53675z704 : STD_LOGIC; 
  signal rome2datao10_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z713 : STD_LOGIC; 
  signal rome2datao10_s_3_BXINV : STD_LOGIC; 
  signal rome2datao10_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z712 : STD_LOGIC; 
  signal rome2datao10_s_3_BYINV : STD_LOGIC; 
  signal nx53675z709_F5MUX : STD_LOGIC; 
  signal nx53675z710 : STD_LOGIC; 
  signal nx53675z709_BXINV : STD_LOGIC; 
  signal U2_ROME10_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal rome2datao10_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z714 : STD_LOGIC; 
  signal rome2datao10_s_2_BXINV : STD_LOGIC; 
  signal rome2datao10_s_2_F6MUX : STD_LOGIC; 
  signal rome2datao10_s_2_G : STD_LOGIC; 
  signal rome2datao10_s_2_BYINV : STD_LOGIC; 
  signal U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROME10_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal rome2datao5_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z329 : STD_LOGIC; 
  signal rome2datao5_s_13_BXINV : STD_LOGIC; 
  signal rome2datao5_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z328 : STD_LOGIC; 
  signal rome2datao5_s_13_BYINV : STD_LOGIC; 
  signal nx53675z325_F5MUX : STD_LOGIC; 
  signal nx53675z326 : STD_LOGIC; 
  signal nx53675z325_BXINV : STD_LOGIC; 
  signal nx53675z325_G : STD_LOGIC; 
  signal rome2datao2_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z140 : STD_LOGIC; 
  signal rome2datao2_s_12_BXINV : STD_LOGIC; 
  signal rome2datao2_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z139 : STD_LOGIC; 
  signal rome2datao2_s_12_BYINV : STD_LOGIC; 
  signal nx53675z135_F5MUX : STD_LOGIC; 
  signal nx53675z137 : STD_LOGIC; 
  signal nx53675z135_BXINV : STD_LOGIC; 
  signal nx53675z136 : STD_LOGIC; 
  signal rome2datao2_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z146 : STD_LOGIC; 
  signal rome2datao2_s_11_BXINV : STD_LOGIC; 
  signal rome2datao2_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z145 : STD_LOGIC; 
  signal rome2datao2_s_11_BYINV : STD_LOGIC; 
  signal nx53675z141_F5MUX : STD_LOGIC; 
  signal nx53675z143 : STD_LOGIC; 
  signal nx53675z141_BXINV : STD_LOGIC; 
  signal nx53675z142 : STD_LOGIC; 
  signal rome2datao2_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z152 : STD_LOGIC; 
  signal rome2datao2_s_10_BXINV : STD_LOGIC; 
  signal rome2datao2_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z151 : STD_LOGIC; 
  signal rome2datao2_s_10_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_FFY_RST : STD_LOGIC; 
  signal nx53675z147_F5MUX : STD_LOGIC; 
  signal nx53675z149 : STD_LOGIC; 
  signal nx53675z147_BXINV : STD_LOGIC; 
  signal nx53675z148 : STD_LOGIC; 
  signal rome2datao2_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z158 : STD_LOGIC; 
  signal rome2datao2_s_9_BXINV : STD_LOGIC; 
  signal rome2datao2_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z157 : STD_LOGIC; 
  signal rome2datao2_s_9_BYINV : STD_LOGIC; 
  signal nx53675z153_F5MUX : STD_LOGIC; 
  signal nx53675z155 : STD_LOGIC; 
  signal nx53675z153_BXINV : STD_LOGIC; 
  signal nx53675z154 : STD_LOGIC; 
  signal rome2datao2_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z194 : STD_LOGIC; 
  signal rome2datao2_s_2_BXINV : STD_LOGIC; 
  signal rome2datao2_s_2_F6MUX : STD_LOGIC; 
  signal rome2datao2_s_2_G : STD_LOGIC; 
  signal rome2datao2_s_2_BYINV : STD_LOGIC; 
  signal U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROME2_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romo2datao9_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z1440 : STD_LOGIC; 
  signal romo2datao9_s_11_BXINV : STD_LOGIC; 
  signal romo2datao9_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z1439 : STD_LOGIC; 
  signal romo2datao9_s_11_BYINV : STD_LOGIC; 
  signal nx53675z1435_F5MUX : STD_LOGIC; 
  signal nx53675z1437 : STD_LOGIC; 
  signal nx53675z1435_BXINV : STD_LOGIC; 
  signal nx53675z1436 : STD_LOGIC; 
  signal romo2datao9_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z1446 : STD_LOGIC; 
  signal romo2datao9_s_10_BXINV : STD_LOGIC; 
  signal romo2datao9_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z1445 : STD_LOGIC; 
  signal romo2datao9_s_10_BYINV : STD_LOGIC; 
  signal nx53675z1441_F5MUX : STD_LOGIC; 
  signal nx53675z1443 : STD_LOGIC; 
  signal nx53675z1441_BXINV : STD_LOGIC; 
  signal nx53675z1442 : STD_LOGIC; 
  signal romo2datao9_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z1452 : STD_LOGIC; 
  signal romo2datao9_s_9_BXINV : STD_LOGIC; 
  signal romo2datao9_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z1451 : STD_LOGIC; 
  signal romo2datao9_s_9_BYINV : STD_LOGIC; 
  signal nx53675z1447_F5MUX : STD_LOGIC; 
  signal nx53675z1449 : STD_LOGIC; 
  signal nx53675z1447_BXINV : STD_LOGIC; 
  signal nx53675z1448 : STD_LOGIC; 
  signal romo2datao9_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z1458 : STD_LOGIC; 
  signal romo2datao9_s_8_BXINV : STD_LOGIC; 
  signal romo2datao9_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z1457 : STD_LOGIC; 
  signal romo2datao9_s_8_BYINV : STD_LOGIC; 
  signal nx53675z1453_F5MUX : STD_LOGIC; 
  signal nx53675z1455 : STD_LOGIC; 
  signal nx53675z1453_BXINV : STD_LOGIC; 
  signal nx53675z1454 : STD_LOGIC; 
  signal romo2datao9_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z1464 : STD_LOGIC; 
  signal romo2datao9_s_7_BXINV : STD_LOGIC; 
  signal romo2datao9_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z1463 : STD_LOGIC; 
  signal romo2datao9_s_7_BYINV : STD_LOGIC; 
  signal nx53675z1459_F5MUX : STD_LOGIC; 
  signal nx53675z1461 : STD_LOGIC; 
  signal nx53675z1459_BXINV : STD_LOGIC; 
  signal nx53675z1460 : STD_LOGIC; 
  signal rome2datao6_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z394 : STD_LOGIC; 
  signal rome2datao6_s_13_BXINV : STD_LOGIC; 
  signal rome2datao6_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z393 : STD_LOGIC; 
  signal rome2datao6_s_13_BYINV : STD_LOGIC; 
  signal nx53675z390_F5MUX : STD_LOGIC; 
  signal nx53675z391 : STD_LOGIC; 
  signal nx53675z390_BXINV : STD_LOGIC; 
  signal nx53675z390_G : STD_LOGIC; 
  signal rome2datao4_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z270 : STD_LOGIC; 
  signal rome2datao4_s_12_BXINV : STD_LOGIC; 
  signal rome2datao4_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z269 : STD_LOGIC; 
  signal rome2datao4_s_12_BYINV : STD_LOGIC; 
  signal nx53675z265_F5MUX : STD_LOGIC; 
  signal nx53675z267 : STD_LOGIC; 
  signal nx53675z265_BXINV : STD_LOGIC; 
  signal nx53675z266 : STD_LOGIC; 
  signal rome2datao4_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z276 : STD_LOGIC; 
  signal rome2datao4_s_11_BXINV : STD_LOGIC; 
  signal rome2datao4_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z275 : STD_LOGIC; 
  signal rome2datao4_s_11_BYINV : STD_LOGIC; 
  signal nx53675z271_F5MUX : STD_LOGIC; 
  signal nx53675z273 : STD_LOGIC; 
  signal nx53675z271_BXINV : STD_LOGIC; 
  signal nx53675z272 : STD_LOGIC; 
  signal rome2datao4_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z282 : STD_LOGIC; 
  signal rome2datao4_s_10_BXINV : STD_LOGIC; 
  signal rome2datao4_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z281 : STD_LOGIC; 
  signal rome2datao4_s_10_BYINV : STD_LOGIC; 
  signal nx53675z277_F5MUX : STD_LOGIC; 
  signal nx53675z279 : STD_LOGIC; 
  signal nx53675z277_BXINV : STD_LOGIC; 
  signal nx53675z278 : STD_LOGIC; 
  signal rome2datao4_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z318 : STD_LOGIC; 
  signal rome2datao4_s_4_BXINV : STD_LOGIC; 
  signal rome2datao4_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z317 : STD_LOGIC; 
  signal rome2datao4_s_4_BYINV : STD_LOGIC; 
  signal nx53675z313_F5MUX : STD_LOGIC; 
  signal nx53675z315 : STD_LOGIC; 
  signal nx53675z313_BXINV : STD_LOGIC; 
  signal nx53675z314 : STD_LOGIC; 
  signal rome2datao4_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z323 : STD_LOGIC; 
  signal rome2datao4_s_3_BXINV : STD_LOGIC; 
  signal rome2datao4_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z322 : STD_LOGIC; 
  signal rome2datao4_s_3_BYINV : STD_LOGIC; 
  signal nx53675z319_F5MUX : STD_LOGIC; 
  signal nx53675z320 : STD_LOGIC; 
  signal nx53675z319_BXINV : STD_LOGIC; 
  signal U2_ROME4_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal rome2datao4_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z324 : STD_LOGIC; 
  signal rome2datao4_s_2_BXINV : STD_LOGIC; 
  signal rome2datao4_s_2_F6MUX : STD_LOGIC; 
  signal rome2datao4_s_2_G : STD_LOGIC; 
  signal rome2datao4_s_2_BYINV : STD_LOGIC; 
  signal U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROME4_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal rome2datao1_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z93 : STD_LOGIC; 
  signal rome2datao1_s_9_BXINV : STD_LOGIC; 
  signal rome2datao1_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z92 : STD_LOGIC; 
  signal rome2datao1_s_9_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_6_FFX_RST : STD_LOGIC; 
  signal nx53675z88_F5MUX : STD_LOGIC; 
  signal nx53675z90 : STD_LOGIC; 
  signal nx53675z88_BXINV : STD_LOGIC; 
  signal nx53675z89 : STD_LOGIC; 
  signal romo2datao10_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z1513 : STD_LOGIC; 
  signal romo2datao10_s_12_BXINV : STD_LOGIC; 
  signal romo2datao10_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z1512 : STD_LOGIC; 
  signal romo2datao10_s_12_BYINV : STD_LOGIC; 
  signal nx53675z1508_F5MUX : STD_LOGIC; 
  signal nx53675z1510 : STD_LOGIC; 
  signal nx53675z1508_BXINV : STD_LOGIC; 
  signal nx53675z1509 : STD_LOGIC; 
  signal romo2datao3_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z960 : STD_LOGIC; 
  signal romo2datao3_s_12_BXINV : STD_LOGIC; 
  signal romo2datao3_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z959 : STD_LOGIC; 
  signal romo2datao3_s_12_BYINV : STD_LOGIC; 
  signal nx53675z955_F5MUX : STD_LOGIC; 
  signal nx53675z957 : STD_LOGIC; 
  signal nx53675z955_BXINV : STD_LOGIC; 
  signal nx53675z956 : STD_LOGIC; 
  signal romo2datao3_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z1020 : STD_LOGIC; 
  signal romo2datao3_s_2_BXINV : STD_LOGIC; 
  signal romo2datao3_s_2_F6MUX : STD_LOGIC; 
  signal nx53675z1019 : STD_LOGIC; 
  signal romo2datao3_s_2_BYINV : STD_LOGIC; 
  signal nx53675z1015_F5MUX : STD_LOGIC; 
  signal nx53675z1017 : STD_LOGIC; 
  signal nx53675z1015_BXINV : STD_LOGIC; 
  signal nx53675z1016 : STD_LOGIC; 
  signal romo2datao2_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z881 : STD_LOGIC; 
  signal romo2datao2_s_12_BXINV : STD_LOGIC; 
  signal romo2datao2_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z880 : STD_LOGIC; 
  signal romo2datao2_s_12_BYINV : STD_LOGIC; 
  signal nx53675z876_F5MUX : STD_LOGIC; 
  signal nx53675z878 : STD_LOGIC; 
  signal nx53675z876_BXINV : STD_LOGIC; 
  signal nx53675z877 : STD_LOGIC; 
  signal romo2datao2_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z887 : STD_LOGIC; 
  signal romo2datao2_s_11_BXINV : STD_LOGIC; 
  signal romo2datao2_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z886 : STD_LOGIC; 
  signal romo2datao2_s_11_BYINV : STD_LOGIC; 
  signal nx53675z882_F5MUX : STD_LOGIC; 
  signal nx53675z884 : STD_LOGIC; 
  signal nx53675z882_BXINV : STD_LOGIC; 
  signal nx53675z883 : STD_LOGIC; 
  signal romo2datao2_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z893 : STD_LOGIC; 
  signal romo2datao2_s_10_BXINV : STD_LOGIC; 
  signal romo2datao2_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z892 : STD_LOGIC; 
  signal romo2datao2_s_10_BYINV : STD_LOGIC; 
  signal nx53675z888_F5MUX : STD_LOGIC; 
  signal nx53675z890 : STD_LOGIC; 
  signal nx53675z888_BXINV : STD_LOGIC; 
  signal nx53675z889 : STD_LOGIC; 
  signal romo2datao2_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z899 : STD_LOGIC; 
  signal romo2datao2_s_9_BXINV : STD_LOGIC; 
  signal romo2datao2_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z898 : STD_LOGIC; 
  signal romo2datao2_s_9_BYINV : STD_LOGIC; 
  signal nx53675z894_F5MUX : STD_LOGIC; 
  signal nx53675z896 : STD_LOGIC; 
  signal nx53675z894_BXINV : STD_LOGIC; 
  signal nx53675z895 : STD_LOGIC; 
  signal romo2datao2_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z905 : STD_LOGIC; 
  signal romo2datao2_s_8_BXINV : STD_LOGIC; 
  signal romo2datao2_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z904 : STD_LOGIC; 
  signal romo2datao2_s_8_BYINV : STD_LOGIC; 
  signal nx53675z900_F5MUX : STD_LOGIC; 
  signal nx53675z902 : STD_LOGIC; 
  signal nx53675z900_BXINV : STD_LOGIC; 
  signal nx53675z901 : STD_LOGIC; 
  signal rome2datao9_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z649 : STD_LOGIC; 
  signal rome2datao9_s_2_BXINV : STD_LOGIC; 
  signal rome2datao9_s_2_F6MUX : STD_LOGIC; 
  signal rome2datao9_s_2_G : STD_LOGIC; 
  signal rome2datao9_s_2_BYINV : STD_LOGIC; 
  signal U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROME9_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romo2datao10_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z1507 : STD_LOGIC; 
  signal romo2datao10_s_13_BXINV : STD_LOGIC; 
  signal romo2datao10_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z1506 : STD_LOGIC; 
  signal romo2datao10_s_13_BYINV : STD_LOGIC; 
  signal nx53675z1503_F5MUX : STD_LOGIC; 
  signal nx53675z1504 : STD_LOGIC; 
  signal nx53675z1503_BXINV : STD_LOGIC; 
  signal nx53675z1503_G : STD_LOGIC; 
  signal romo2datao10_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z1525 : STD_LOGIC; 
  signal romo2datao10_s_10_BXINV : STD_LOGIC; 
  signal romo2datao10_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z1524 : STD_LOGIC; 
  signal romo2datao10_s_10_BYINV : STD_LOGIC; 
  signal nx53675z1520_F5MUX : STD_LOGIC; 
  signal nx53675z1522 : STD_LOGIC; 
  signal nx53675z1520_BXINV : STD_LOGIC; 
  signal nx53675z1521 : STD_LOGIC; 
  signal romo2datao10_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z1573 : STD_LOGIC; 
  signal romo2datao10_s_2_BXINV : STD_LOGIC; 
  signal romo2datao10_s_2_F6MUX : STD_LOGIC; 
  signal nx53675z1572 : STD_LOGIC; 
  signal romo2datao10_s_2_BYINV : STD_LOGIC; 
  signal nx53675z1568_F5MUX : STD_LOGIC; 
  signal nx53675z1570 : STD_LOGIC; 
  signal nx53675z1568_BXINV : STD_LOGIC; 
  signal nx53675z1569 : STD_LOGIC; 
  signal romo2datao10_s_1_F5MUX : STD_LOGIC; 
  signal nx53675z1579 : STD_LOGIC; 
  signal romo2datao10_s_1_BXINV : STD_LOGIC; 
  signal romo2datao10_s_1_F6MUX : STD_LOGIC; 
  signal nx53675z1578 : STD_LOGIC; 
  signal romo2datao10_s_1_BYINV : STD_LOGIC; 
  signal nx53675z1574_F5MUX : STD_LOGIC; 
  signal nx53675z1576 : STD_LOGIC; 
  signal nx53675z1574_BXINV : STD_LOGIC; 
  signal nx53675z1575 : STD_LOGIC; 
  signal romo2datao10_s_0_F5MUX : STD_LOGIC; 
  signal nx53675z1581 : STD_LOGIC; 
  signal romo2datao10_s_0_BXINV : STD_LOGIC; 
  signal romo2datao10_s_0_F6MUX : STD_LOGIC; 
  signal nx53675z1580 : STD_LOGIC; 
  signal romo2datao10_s_0_BYINV : STD_LOGIC; 
  signal U2_ROMO10_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROMO10_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROMO10_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROMO10_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romo2datao9_s_0_F5MUX : STD_LOGIC; 
  signal nx53675z1502 : STD_LOGIC; 
  signal romo2datao9_s_0_BXINV : STD_LOGIC; 
  signal romo2datao9_s_0_F6MUX : STD_LOGIC; 
  signal nx53675z1501 : STD_LOGIC; 
  signal romo2datao9_s_0_BYINV : STD_LOGIC; 
  signal U2_ROMO9_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROMO9_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROMO9_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROMO9_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romo2datao4_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z1081 : STD_LOGIC; 
  signal romo2datao4_s_5_BXINV : STD_LOGIC; 
  signal romo2datao4_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z1080 : STD_LOGIC; 
  signal romo2datao4_s_5_BYINV : STD_LOGIC; 
  signal nx53675z1076_F5MUX : STD_LOGIC; 
  signal nx53675z1078 : STD_LOGIC; 
  signal nx53675z1076_BXINV : STD_LOGIC; 
  signal nx53675z1077 : STD_LOGIC; 
  signal romo2datao3_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z954 : STD_LOGIC; 
  signal romo2datao3_s_13_BXINV : STD_LOGIC; 
  signal romo2datao3_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z953 : STD_LOGIC; 
  signal romo2datao3_s_13_BYINV : STD_LOGIC; 
  signal nx53675z950_F5MUX : STD_LOGIC; 
  signal nx53675z951 : STD_LOGIC; 
  signal nx53675z950_BXINV : STD_LOGIC; 
  signal nx53675z950_G : STD_LOGIC; 
  signal romo2datao2_s_1_F5MUX : STD_LOGIC; 
  signal nx53675z947 : STD_LOGIC; 
  signal romo2datao2_s_1_BXINV : STD_LOGIC; 
  signal romo2datao2_s_1_F6MUX : STD_LOGIC; 
  signal nx53675z946 : STD_LOGIC; 
  signal romo2datao2_s_1_BYINV : STD_LOGIC; 
  signal nx53675z942_F5MUX : STD_LOGIC; 
  signal nx53675z944 : STD_LOGIC; 
  signal nx53675z942_BXINV : STD_LOGIC; 
  signal nx53675z943 : STD_LOGIC; 
  signal romo2datao2_s_0_F5MUX : STD_LOGIC; 
  signal nx53675z949 : STD_LOGIC; 
  signal romo2datao2_s_0_BXINV : STD_LOGIC; 
  signal romo2datao2_s_0_F6MUX : STD_LOGIC; 
  signal nx53675z948 : STD_LOGIC; 
  signal romo2datao2_s_0_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_FFY_RST : STD_LOGIC; 
  signal U2_ROMO2_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROMO2_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROMO2_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROMO2_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romo2datao1_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z832 : STD_LOGIC; 
  signal romo2datao1_s_7_BXINV : STD_LOGIC; 
  signal romo2datao1_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z831 : STD_LOGIC; 
  signal romo2datao1_s_7_BYINV : STD_LOGIC; 
  signal nx53675z827_F5MUX : STD_LOGIC; 
  signal nx53675z829 : STD_LOGIC; 
  signal nx53675z827_BXINV : STD_LOGIC; 
  signal nx53675z828 : STD_LOGIC; 
  signal romo2datao1_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z838 : STD_LOGIC; 
  signal romo2datao1_s_6_BXINV : STD_LOGIC; 
  signal romo2datao1_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z837 : STD_LOGIC; 
  signal romo2datao1_s_6_BYINV : STD_LOGIC; 
  signal nx53675z833_F5MUX : STD_LOGIC; 
  signal nx53675z835 : STD_LOGIC; 
  signal nx53675z833_BXINV : STD_LOGIC; 
  signal nx53675z834 : STD_LOGIC; 
  signal romo2datao1_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z844 : STD_LOGIC; 
  signal romo2datao1_s_5_BXINV : STD_LOGIC; 
  signal romo2datao1_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z843 : STD_LOGIC; 
  signal romo2datao1_s_5_BYINV : STD_LOGIC; 
  signal nx53675z839_F5MUX : STD_LOGIC; 
  signal nx53675z841 : STD_LOGIC; 
  signal nx53675z839_BXINV : STD_LOGIC; 
  signal nx53675z840 : STD_LOGIC; 
  signal romo2datao1_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z850 : STD_LOGIC; 
  signal romo2datao1_s_4_BXINV : STD_LOGIC; 
  signal romo2datao1_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z849 : STD_LOGIC; 
  signal romo2datao1_s_4_BYINV : STD_LOGIC; 
  signal nx53675z845_F5MUX : STD_LOGIC; 
  signal nx53675z847 : STD_LOGIC; 
  signal nx53675z845_BXINV : STD_LOGIC; 
  signal nx53675z846 : STD_LOGIC; 
  signal romo2datao1_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z856 : STD_LOGIC; 
  signal romo2datao1_s_3_BXINV : STD_LOGIC; 
  signal romo2datao1_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z855 : STD_LOGIC; 
  signal romo2datao1_s_3_BYINV : STD_LOGIC; 
  signal nx53675z851_F5MUX : STD_LOGIC; 
  signal nx53675z853 : STD_LOGIC; 
  signal nx53675z851_BXINV : STD_LOGIC; 
  signal nx53675z852 : STD_LOGIC; 
  signal rome2datao6_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z400 : STD_LOGIC; 
  signal rome2datao6_s_12_BXINV : STD_LOGIC; 
  signal rome2datao6_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z399 : STD_LOGIC; 
  signal rome2datao6_s_12_BYINV : STD_LOGIC; 
  signal nx53675z395_F5MUX : STD_LOGIC; 
  signal nx53675z397 : STD_LOGIC; 
  signal nx53675z395_BXINV : STD_LOGIC; 
  signal nx53675z396 : STD_LOGIC; 
  signal rome2datao6_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z448 : STD_LOGIC; 
  signal rome2datao6_s_4_BXINV : STD_LOGIC; 
  signal rome2datao6_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z447 : STD_LOGIC; 
  signal rome2datao6_s_4_BYINV : STD_LOGIC; 
  signal nx53675z443_F5MUX : STD_LOGIC; 
  signal nx53675z445 : STD_LOGIC; 
  signal nx53675z443_BXINV : STD_LOGIC; 
  signal nx53675z444 : STD_LOGIC; 
  signal rome2datao6_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z453 : STD_LOGIC; 
  signal rome2datao6_s_3_BXINV : STD_LOGIC; 
  signal rome2datao6_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z452 : STD_LOGIC; 
  signal rome2datao6_s_3_BYINV : STD_LOGIC; 
  signal nx53675z449_F5MUX : STD_LOGIC; 
  signal nx53675z450 : STD_LOGIC; 
  signal nx53675z449_BXINV : STD_LOGIC; 
  signal U2_ROME6_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal rome2datao6_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z454 : STD_LOGIC; 
  signal rome2datao6_s_2_BXINV : STD_LOGIC; 
  signal rome2datao6_s_2_F6MUX : STD_LOGIC; 
  signal rome2datao6_s_2_G : STD_LOGIC; 
  signal rome2datao6_s_2_BYINV : STD_LOGIC; 
  signal U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROME6_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romo2datao0_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z773 : STD_LOGIC; 
  signal romo2datao0_s_4_BXINV : STD_LOGIC; 
  signal romo2datao0_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z772 : STD_LOGIC; 
  signal romo2datao0_s_4_BYINV : STD_LOGIC; 
  signal nx53675z768_F5MUX : STD_LOGIC; 
  signal nx53675z770 : STD_LOGIC; 
  signal nx53675z768_BXINV : STD_LOGIC; 
  signal nx53675z769 : STD_LOGIC; 
  signal romo2datao0_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z779 : STD_LOGIC; 
  signal romo2datao0_s_3_BXINV : STD_LOGIC; 
  signal romo2datao0_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z778 : STD_LOGIC; 
  signal romo2datao0_s_3_BYINV : STD_LOGIC; 
  signal nx53675z774_F5MUX : STD_LOGIC; 
  signal nx53675z776 : STD_LOGIC; 
  signal nx53675z774_BXINV : STD_LOGIC; 
  signal nx53675z775 : STD_LOGIC; 
  signal romo2datao0_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z785 : STD_LOGIC; 
  signal romo2datao0_s_2_BXINV : STD_LOGIC; 
  signal romo2datao0_s_2_F6MUX : STD_LOGIC; 
  signal nx53675z784 : STD_LOGIC; 
  signal romo2datao0_s_2_BYINV : STD_LOGIC; 
  signal nx53675z780_F5MUX : STD_LOGIC; 
  signal nx53675z782 : STD_LOGIC; 
  signal nx53675z780_BXINV : STD_LOGIC; 
  signal nx53675z781 : STD_LOGIC; 
  signal romo2datao0_s_1_F5MUX : STD_LOGIC; 
  signal nx53675z791 : STD_LOGIC; 
  signal romo2datao0_s_1_BXINV : STD_LOGIC; 
  signal romo2datao0_s_1_F6MUX : STD_LOGIC; 
  signal nx53675z790 : STD_LOGIC; 
  signal romo2datao0_s_1_BYINV : STD_LOGIC; 
  signal nx53675z786_F5MUX : STD_LOGIC; 
  signal nx53675z788 : STD_LOGIC; 
  signal nx53675z786_BXINV : STD_LOGIC; 
  signal nx53675z787 : STD_LOGIC; 
  signal rome2datao3_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z217 : STD_LOGIC; 
  signal rome2datao3_s_10_BXINV : STD_LOGIC; 
  signal rome2datao3_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z216 : STD_LOGIC; 
  signal rome2datao3_s_10_BYINV : STD_LOGIC; 
  signal nx53675z212_F5MUX : STD_LOGIC; 
  signal nx53675z214 : STD_LOGIC; 
  signal nx53675z212_BXINV : STD_LOGIC; 
  signal nx53675z213 : STD_LOGIC; 
  signal rome2datao3_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z229 : STD_LOGIC; 
  signal rome2datao3_s_8_BXINV : STD_LOGIC; 
  signal rome2datao3_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z228 : STD_LOGIC; 
  signal rome2datao3_s_8_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_2_8_FFX_RST : STD_LOGIC; 
  signal nx53675z224_F5MUX : STD_LOGIC; 
  signal nx53675z226 : STD_LOGIC; 
  signal nx53675z224_BXINV : STD_LOGIC; 
  signal nx53675z225 : STD_LOGIC; 
  signal romo2datao4_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z1045 : STD_LOGIC; 
  signal romo2datao4_s_11_BXINV : STD_LOGIC; 
  signal romo2datao4_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z1044 : STD_LOGIC; 
  signal romo2datao4_s_11_BYINV : STD_LOGIC; 
  signal nx53675z1040_F5MUX : STD_LOGIC; 
  signal nx53675z1042 : STD_LOGIC; 
  signal nx53675z1040_BXINV : STD_LOGIC; 
  signal nx53675z1041 : STD_LOGIC; 
  signal romo2datao3_s_1_F5MUX : STD_LOGIC; 
  signal nx53675z1026 : STD_LOGIC; 
  signal romo2datao3_s_1_BXINV : STD_LOGIC; 
  signal romo2datao3_s_1_F6MUX : STD_LOGIC; 
  signal nx53675z1025 : STD_LOGIC; 
  signal romo2datao3_s_1_BYINV : STD_LOGIC; 
  signal nx53675z1021_F5MUX : STD_LOGIC; 
  signal nx53675z1023 : STD_LOGIC; 
  signal nx53675z1021_BXINV : STD_LOGIC; 
  signal nx53675z1022 : STD_LOGIC; 
  signal romo2datao0_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z719 : STD_LOGIC; 
  signal romo2datao0_s_13_BXINV : STD_LOGIC; 
  signal romo2datao0_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z718 : STD_LOGIC; 
  signal romo2datao0_s_13_BYINV : STD_LOGIC; 
  signal nx53675z715_F5MUX : STD_LOGIC; 
  signal nx53675z716 : STD_LOGIC; 
  signal nx53675z715_BXINV : STD_LOGIC; 
  signal nx53675z715_G : STD_LOGIC; 
  signal romo2datao8_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z1355 : STD_LOGIC; 
  signal romo2datao8_s_12_BXINV : STD_LOGIC; 
  signal romo2datao8_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z1354 : STD_LOGIC; 
  signal romo2datao8_s_12_BYINV : STD_LOGIC; 
  signal nx53675z1350_F5MUX : STD_LOGIC; 
  signal nx53675z1352 : STD_LOGIC; 
  signal nx53675z1350_BXINV : STD_LOGIC; 
  signal nx53675z1351 : STD_LOGIC; 
  signal romo2datao8_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z1403 : STD_LOGIC; 
  signal romo2datao8_s_4_BXINV : STD_LOGIC; 
  signal romo2datao8_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z1402 : STD_LOGIC; 
  signal romo2datao8_s_4_BYINV : STD_LOGIC; 
  signal nx53675z1398_F5MUX : STD_LOGIC; 
  signal nx53675z1400 : STD_LOGIC; 
  signal nx53675z1398_BXINV : STD_LOGIC; 
  signal nx53675z1399 : STD_LOGIC; 
  signal romo2datao8_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z1409 : STD_LOGIC; 
  signal romo2datao8_s_3_BXINV : STD_LOGIC; 
  signal romo2datao8_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z1408 : STD_LOGIC; 
  signal romo2datao8_s_3_BYINV : STD_LOGIC; 
  signal nx53675z1404_F5MUX : STD_LOGIC; 
  signal nx53675z1406 : STD_LOGIC; 
  signal nx53675z1404_BXINV : STD_LOGIC; 
  signal nx53675z1405 : STD_LOGIC; 
  signal romo2datao8_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z1415 : STD_LOGIC; 
  signal romo2datao8_s_2_BXINV : STD_LOGIC; 
  signal romo2datao8_s_2_F6MUX : STD_LOGIC; 
  signal nx53675z1414 : STD_LOGIC; 
  signal romo2datao8_s_2_BYINV : STD_LOGIC; 
  signal rome2datao3_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z235 : STD_LOGIC; 
  signal rome2datao3_s_7_BXINV : STD_LOGIC; 
  signal rome2datao3_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z234 : STD_LOGIC; 
  signal rome2datao3_s_7_BYINV : STD_LOGIC; 
  signal nx53675z230_F5MUX : STD_LOGIC; 
  signal nx53675z232 : STD_LOGIC; 
  signal nx53675z230_BXINV : STD_LOGIC; 
  signal nx53675z231 : STD_LOGIC; 
  signal romo2datao9_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z1494 : STD_LOGIC; 
  signal romo2datao9_s_2_BXINV : STD_LOGIC; 
  signal romo2datao9_s_2_F6MUX : STD_LOGIC; 
  signal nx53675z1493 : STD_LOGIC; 
  signal romo2datao9_s_2_BYINV : STD_LOGIC; 
  signal nx53675z1489_F5MUX : STD_LOGIC; 
  signal nx53675z1491 : STD_LOGIC; 
  signal nx53675z1489_BXINV : STD_LOGIC; 
  signal nx53675z1490 : STD_LOGIC; 
  signal romo2datao4_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z1039 : STD_LOGIC; 
  signal romo2datao4_s_12_BXINV : STD_LOGIC; 
  signal romo2datao4_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z1038 : STD_LOGIC; 
  signal romo2datao4_s_12_BYINV : STD_LOGIC; 
  signal nx53675z1034_F5MUX : STD_LOGIC; 
  signal nx53675z1036 : STD_LOGIC; 
  signal nx53675z1034_BXINV : STD_LOGIC; 
  signal nx53675z1035 : STD_LOGIC; 
  signal romo2datao3_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z972 : STD_LOGIC; 
  signal romo2datao3_s_10_BXINV : STD_LOGIC; 
  signal romo2datao3_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z971 : STD_LOGIC; 
  signal romo2datao3_s_10_BYINV : STD_LOGIC; 
  signal nx53675z967_F5MUX : STD_LOGIC; 
  signal nx53675z969 : STD_LOGIC; 
  signal nx53675z967_BXINV : STD_LOGIC; 
  signal nx53675z968 : STD_LOGIC; 
  signal romo2datao3_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z984 : STD_LOGIC; 
  signal romo2datao3_s_8_BXINV : STD_LOGIC; 
  signal romo2datao3_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z983 : STD_LOGIC; 
  signal romo2datao3_s_8_BYINV : STD_LOGIC; 
  signal nx53675z979_F5MUX : STD_LOGIC; 
  signal nx53675z981 : STD_LOGIC; 
  signal nx53675z979_BXINV : STD_LOGIC; 
  signal nx53675z980 : STD_LOGIC; 
  signal romo2datao3_s_0_F5MUX : STD_LOGIC; 
  signal nx53675z1028 : STD_LOGIC; 
  signal romo2datao3_s_0_BXINV : STD_LOGIC; 
  signal romo2datao3_s_0_F6MUX : STD_LOGIC; 
  signal nx53675z1027 : STD_LOGIC; 
  signal romo2datao3_s_0_BYINV : STD_LOGIC; 
  signal U2_ROMO3_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROMO3_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROMO3_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROMO3_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romo2datao2_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z911 : STD_LOGIC; 
  signal romo2datao2_s_7_BXINV : STD_LOGIC; 
  signal romo2datao2_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z910 : STD_LOGIC; 
  signal romo2datao2_s_7_BYINV : STD_LOGIC; 
  signal nx53675z906_F5MUX : STD_LOGIC; 
  signal nx53675z908 : STD_LOGIC; 
  signal nx53675z906_BXINV : STD_LOGIC; 
  signal nx53675z907 : STD_LOGIC; 
  signal romo2datao2_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z917 : STD_LOGIC; 
  signal romo2datao2_s_6_BXINV : STD_LOGIC; 
  signal romo2datao2_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z916 : STD_LOGIC; 
  signal romo2datao2_s_6_BYINV : STD_LOGIC; 
  signal nx53675z912_F5MUX : STD_LOGIC; 
  signal nx53675z914 : STD_LOGIC; 
  signal nx53675z912_BXINV : STD_LOGIC; 
  signal nx53675z913 : STD_LOGIC; 
  signal romo2datao2_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z923 : STD_LOGIC; 
  signal romo2datao2_s_5_BXINV : STD_LOGIC; 
  signal romo2datao2_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z922 : STD_LOGIC; 
  signal romo2datao2_s_5_BYINV : STD_LOGIC; 
  signal nx53675z918_F5MUX : STD_LOGIC; 
  signal nx53675z920 : STD_LOGIC; 
  signal nx53675z918_BXINV : STD_LOGIC; 
  signal nx53675z919 : STD_LOGIC; 
  signal romo2datao2_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z929 : STD_LOGIC; 
  signal romo2datao2_s_4_BXINV : STD_LOGIC; 
  signal romo2datao2_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z928 : STD_LOGIC; 
  signal romo2datao2_s_4_BYINV : STD_LOGIC; 
  signal nx53675z924_F5MUX : STD_LOGIC; 
  signal nx53675z926 : STD_LOGIC; 
  signal nx53675z924_BXINV : STD_LOGIC; 
  signal nx53675z925 : STD_LOGIC; 
  signal romo2datao10_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z1531 : STD_LOGIC; 
  signal romo2datao10_s_9_BXINV : STD_LOGIC; 
  signal romo2datao10_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z1530 : STD_LOGIC; 
  signal romo2datao10_s_9_BYINV : STD_LOGIC; 
  signal nx53675z1526_F5MUX : STD_LOGIC; 
  signal nx53675z1528 : STD_LOGIC; 
  signal nx53675z1526_BXINV : STD_LOGIC; 
  signal nx53675z1527 : STD_LOGIC; 
  signal romo2datao10_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z1537 : STD_LOGIC; 
  signal romo2datao10_s_8_BXINV : STD_LOGIC; 
  signal romo2datao10_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z1536 : STD_LOGIC; 
  signal romo2datao10_s_8_BYINV : STD_LOGIC; 
  signal nx53675z1532_F5MUX : STD_LOGIC; 
  signal nx53675z1534 : STD_LOGIC; 
  signal nx53675z1532_BXINV : STD_LOGIC; 
  signal nx53675z1533 : STD_LOGIC; 
  signal romo2datao10_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z1543 : STD_LOGIC; 
  signal romo2datao10_s_7_BXINV : STD_LOGIC; 
  signal romo2datao10_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z1542 : STD_LOGIC; 
  signal romo2datao10_s_7_BYINV : STD_LOGIC; 
  signal nx53675z1538_F5MUX : STD_LOGIC; 
  signal nx53675z1540 : STD_LOGIC; 
  signal nx53675z1538_BXINV : STD_LOGIC; 
  signal nx53675z1539 : STD_LOGIC; 
  signal romo2datao10_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z1549 : STD_LOGIC; 
  signal romo2datao10_s_6_BXINV : STD_LOGIC; 
  signal romo2datao10_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z1548 : STD_LOGIC; 
  signal romo2datao10_s_6_BYINV : STD_LOGIC; 
  signal nx53675z1544_F5MUX : STD_LOGIC; 
  signal nx53675z1546 : STD_LOGIC; 
  signal nx53675z1544_BXINV : STD_LOGIC; 
  signal nx53675z1545 : STD_LOGIC; 
  signal romo2datao10_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z1555 : STD_LOGIC; 
  signal romo2datao10_s_5_BXINV : STD_LOGIC; 
  signal romo2datao10_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z1554 : STD_LOGIC; 
  signal romo2datao10_s_5_BYINV : STD_LOGIC; 
  signal nx53675z1550_F5MUX : STD_LOGIC; 
  signal nx53675z1552 : STD_LOGIC; 
  signal nx53675z1550_BXINV : STD_LOGIC; 
  signal nx53675z1551 : STD_LOGIC; 
  signal romo2datao4_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z1033 : STD_LOGIC; 
  signal romo2datao4_s_13_BXINV : STD_LOGIC; 
  signal romo2datao4_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z1032 : STD_LOGIC; 
  signal romo2datao4_s_13_BYINV : STD_LOGIC; 
  signal nx53675z1029_F5MUX : STD_LOGIC; 
  signal nx53675z1030 : STD_LOGIC; 
  signal nx53675z1029_BXINV : STD_LOGIC; 
  signal nx53675z1029_G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_0_FFX_RST : STD_LOGIC; 
  signal romo2datao1_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z862 : STD_LOGIC; 
  signal romo2datao1_s_2_BXINV : STD_LOGIC; 
  signal romo2datao1_s_2_F6MUX : STD_LOGIC; 
  signal nx53675z861 : STD_LOGIC; 
  signal romo2datao1_s_2_BYINV : STD_LOGIC; 
  signal nx53675z857_F5MUX : STD_LOGIC; 
  signal nx53675z859 : STD_LOGIC; 
  signal nx53675z857_BXINV : STD_LOGIC; 
  signal nx53675z858 : STD_LOGIC; 
  signal romo2datao1_s_1_F5MUX : STD_LOGIC; 
  signal nx53675z868 : STD_LOGIC; 
  signal romo2datao1_s_1_BXINV : STD_LOGIC; 
  signal romo2datao1_s_1_F6MUX : STD_LOGIC; 
  signal nx53675z867 : STD_LOGIC; 
  signal romo2datao1_s_1_BYINV : STD_LOGIC; 
  signal nx53675z863_F5MUX : STD_LOGIC; 
  signal nx53675z865 : STD_LOGIC; 
  signal nx53675z863_BXINV : STD_LOGIC; 
  signal nx53675z864 : STD_LOGIC; 
  signal rome2datao7_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z459 : STD_LOGIC; 
  signal rome2datao7_s_13_BXINV : STD_LOGIC; 
  signal rome2datao7_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z458 : STD_LOGIC; 
  signal rome2datao7_s_13_BYINV : STD_LOGIC; 
  signal nx53675z455_F5MUX : STD_LOGIC; 
  signal nx53675z456 : STD_LOGIC; 
  signal nx53675z455_BXINV : STD_LOGIC; 
  signal nx53675z455_G : STD_LOGIC; 
  signal rome2datao6_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z406 : STD_LOGIC; 
  signal rome2datao6_s_11_BXINV : STD_LOGIC; 
  signal rome2datao6_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z405 : STD_LOGIC; 
  signal rome2datao6_s_11_BYINV : STD_LOGIC; 
  signal nx53675z401_F5MUX : STD_LOGIC; 
  signal nx53675z403 : STD_LOGIC; 
  signal nx53675z401_BXINV : STD_LOGIC; 
  signal nx53675z402 : STD_LOGIC; 
  signal rome2datao6_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z412 : STD_LOGIC; 
  signal rome2datao6_s_10_BXINV : STD_LOGIC; 
  signal rome2datao6_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z411 : STD_LOGIC; 
  signal rome2datao6_s_10_BYINV : STD_LOGIC; 
  signal nx53675z407_F5MUX : STD_LOGIC; 
  signal nx53675z409 : STD_LOGIC; 
  signal nx53675z407_BXINV : STD_LOGIC; 
  signal nx53675z408 : STD_LOGIC; 
  signal rome2datao6_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z418 : STD_LOGIC; 
  signal rome2datao6_s_9_BXINV : STD_LOGIC; 
  signal rome2datao6_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z417 : STD_LOGIC; 
  signal rome2datao6_s_9_BYINV : STD_LOGIC; 
  signal nx53675z413_F5MUX : STD_LOGIC; 
  signal nx53675z415 : STD_LOGIC; 
  signal nx53675z413_BXINV : STD_LOGIC; 
  signal nx53675z414 : STD_LOGIC; 
  signal rome2datao6_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z424 : STD_LOGIC; 
  signal rome2datao6_s_8_BXINV : STD_LOGIC; 
  signal rome2datao6_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z423 : STD_LOGIC; 
  signal rome2datao6_s_8_BYINV : STD_LOGIC; 
  signal nx53675z419_F5MUX : STD_LOGIC; 
  signal nx53675z421 : STD_LOGIC; 
  signal nx53675z419_BXINV : STD_LOGIC; 
  signal nx53675z420 : STD_LOGIC; 
  signal rome2datao6_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z430 : STD_LOGIC; 
  signal rome2datao6_s_7_BXINV : STD_LOGIC; 
  signal rome2datao6_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z429 : STD_LOGIC; 
  signal rome2datao6_s_7_BYINV : STD_LOGIC; 
  signal nx53675z425_F5MUX : STD_LOGIC; 
  signal nx53675z427 : STD_LOGIC; 
  signal nx53675z425_BXINV : STD_LOGIC; 
  signal nx53675z426 : STD_LOGIC; 
  signal romo2datao4_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z1093 : STD_LOGIC; 
  signal romo2datao4_s_3_BXINV : STD_LOGIC; 
  signal romo2datao4_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z1092 : STD_LOGIC; 
  signal romo2datao4_s_3_BYINV : STD_LOGIC; 
  signal nx53675z1088_F5MUX : STD_LOGIC; 
  signal nx53675z1090 : STD_LOGIC; 
  signal nx53675z1088_BXINV : STD_LOGIC; 
  signal nx53675z1089 : STD_LOGIC; 
  signal romo2datao4_s_1_F5MUX : STD_LOGIC; 
  signal nx53675z1105 : STD_LOGIC; 
  signal romo2datao4_s_1_BXINV : STD_LOGIC; 
  signal romo2datao4_s_1_F6MUX : STD_LOGIC; 
  signal nx53675z1104 : STD_LOGIC; 
  signal romo2datao4_s_1_BYINV : STD_LOGIC; 
  signal nx53675z1100_F5MUX : STD_LOGIC; 
  signal nx53675z1102 : STD_LOGIC; 
  signal nx53675z1100_BXINV : STD_LOGIC; 
  signal nx53675z1101 : STD_LOGIC; 
  signal romo2datao6_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z1221 : STD_LOGIC; 
  signal romo2datao6_s_8_BXINV : STD_LOGIC; 
  signal romo2datao6_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z1220 : STD_LOGIC; 
  signal romo2datao6_s_8_BYINV : STD_LOGIC; 
  signal nx53675z1216_F5MUX : STD_LOGIC; 
  signal nx53675z1218 : STD_LOGIC; 
  signal nx53675z1216_BXINV : STD_LOGIC; 
  signal nx53675z1217 : STD_LOGIC; 
  signal romo2datao6_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z1227 : STD_LOGIC; 
  signal romo2datao6_s_7_BXINV : STD_LOGIC; 
  signal romo2datao6_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z1226 : STD_LOGIC; 
  signal romo2datao6_s_7_BYINV : STD_LOGIC; 
  signal nx53675z1222_F5MUX : STD_LOGIC; 
  signal nx53675z1224 : STD_LOGIC; 
  signal nx53675z1222_BXINV : STD_LOGIC; 
  signal nx53675z1223 : STD_LOGIC; 
  signal romo2datao5_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z1112 : STD_LOGIC; 
  signal romo2datao5_s_13_BXINV : STD_LOGIC; 
  signal romo2datao5_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z1111 : STD_LOGIC; 
  signal romo2datao5_s_13_BYINV : STD_LOGIC; 
  signal nx53675z1108_F5MUX : STD_LOGIC; 
  signal nx53675z1109 : STD_LOGIC; 
  signal nx53675z1108_BXINV : STD_LOGIC; 
  signal nx53675z1108_G : STD_LOGIC; 
  signal romo2datao5_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z1154 : STD_LOGIC; 
  signal romo2datao5_s_6_BXINV : STD_LOGIC; 
  signal romo2datao5_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z1153 : STD_LOGIC; 
  signal romo2datao5_s_6_BYINV : STD_LOGIC; 
  signal nx53675z1149_F5MUX : STD_LOGIC; 
  signal nx53675z1151 : STD_LOGIC; 
  signal nx53675z1149_BXINV : STD_LOGIC; 
  signal nx53675z1150 : STD_LOGIC; 
  signal romo2datao5_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z1160 : STD_LOGIC; 
  signal romo2datao5_s_5_BXINV : STD_LOGIC; 
  signal romo2datao5_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z1159 : STD_LOGIC; 
  signal romo2datao5_s_5_BYINV : STD_LOGIC; 
  signal nx53675z1155_F5MUX : STD_LOGIC; 
  signal nx53675z1157 : STD_LOGIC; 
  signal nx53675z1155_BXINV : STD_LOGIC; 
  signal nx53675z1156 : STD_LOGIC; 
  signal romo2datao5_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z1166 : STD_LOGIC; 
  signal romo2datao5_s_4_BXINV : STD_LOGIC; 
  signal romo2datao5_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z1165 : STD_LOGIC; 
  signal romo2datao5_s_4_BYINV : STD_LOGIC; 
  signal nx53675z1161_F5MUX : STD_LOGIC; 
  signal nx53675z1163 : STD_LOGIC; 
  signal nx53675z1161_BXINV : STD_LOGIC; 
  signal nx53675z1162 : STD_LOGIC; 
  signal romo2datao5_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z1172 : STD_LOGIC; 
  signal romo2datao5_s_3_BXINV : STD_LOGIC; 
  signal romo2datao5_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z1171 : STD_LOGIC; 
  signal romo2datao5_s_3_BYINV : STD_LOGIC; 
  signal nx53675z1167_F5MUX : STD_LOGIC; 
  signal nx53675z1169 : STD_LOGIC; 
  signal nx53675z1167_BXINV : STD_LOGIC; 
  signal nx53675z1168 : STD_LOGIC; 
  signal romo2datao4_s_0_F5MUX : STD_LOGIC; 
  signal nx53675z1107 : STD_LOGIC; 
  signal romo2datao4_s_0_BXINV : STD_LOGIC; 
  signal romo2datao4_s_0_F6MUX : STD_LOGIC; 
  signal nx53675z1106 : STD_LOGIC; 
  signal romo2datao4_s_0_BYINV : STD_LOGIC; 
  signal U2_ROMO4_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROMO4_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROMO4_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROMO4_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal rome2datao8_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z530 : STD_LOGIC; 
  signal rome2datao8_s_12_BXINV : STD_LOGIC; 
  signal rome2datao8_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z529 : STD_LOGIC; 
  signal rome2datao8_s_12_BYINV : STD_LOGIC; 
  signal nx53675z525_F5MUX : STD_LOGIC; 
  signal nx53675z527 : STD_LOGIC; 
  signal nx53675z525_BXINV : STD_LOGIC; 
  signal nx53675z526 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_FFY_RST : STD_LOGIC; 
  signal rome2datao8_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z536 : STD_LOGIC; 
  signal rome2datao8_s_11_BXINV : STD_LOGIC; 
  signal rome2datao8_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z535 : STD_LOGIC; 
  signal rome2datao8_s_11_BYINV : STD_LOGIC; 
  signal nx53675z531_F5MUX : STD_LOGIC; 
  signal nx53675z533 : STD_LOGIC; 
  signal nx53675z531_BXINV : STD_LOGIC; 
  signal nx53675z532 : STD_LOGIC; 
  signal rome2datao8_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z542 : STD_LOGIC; 
  signal rome2datao8_s_10_BXINV : STD_LOGIC; 
  signal rome2datao8_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z541 : STD_LOGIC; 
  signal rome2datao8_s_10_BYINV : STD_LOGIC; 
  signal nx53675z537_F5MUX : STD_LOGIC; 
  signal nx53675z539 : STD_LOGIC; 
  signal nx53675z537_BXINV : STD_LOGIC; 
  signal nx53675z538 : STD_LOGIC; 
  signal rome2datao8_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z548 : STD_LOGIC; 
  signal rome2datao8_s_9_BXINV : STD_LOGIC; 
  signal rome2datao8_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z547 : STD_LOGIC; 
  signal rome2datao8_s_9_BYINV : STD_LOGIC; 
  signal nx53675z543_F5MUX : STD_LOGIC; 
  signal nx53675z545 : STD_LOGIC; 
  signal nx53675z543_BXINV : STD_LOGIC; 
  signal nx53675z544 : STD_LOGIC; 
  signal rome2datao4_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z264 : STD_LOGIC; 
  signal rome2datao4_s_13_BXINV : STD_LOGIC; 
  signal rome2datao4_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z263 : STD_LOGIC; 
  signal rome2datao4_s_13_BYINV : STD_LOGIC; 
  signal nx53675z260_F5MUX : STD_LOGIC; 
  signal nx53675z261 : STD_LOGIC; 
  signal nx53675z260_BXINV : STD_LOGIC; 
  signal nx53675z260_G : STD_LOGIC; 
  signal rome2datao8_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z524 : STD_LOGIC; 
  signal rome2datao8_s_13_BXINV : STD_LOGIC; 
  signal rome2datao8_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z523 : STD_LOGIC; 
  signal rome2datao8_s_13_BYINV : STD_LOGIC; 
  signal nx53675z520_F5MUX : STD_LOGIC; 
  signal nx53675z521 : STD_LOGIC; 
  signal nx53675z520_BXINV : STD_LOGIC; 
  signal nx53675z520_G : STD_LOGIC; 
  signal rome2datao5_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z359 : STD_LOGIC; 
  signal rome2datao5_s_8_BXINV : STD_LOGIC; 
  signal rome2datao5_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z358 : STD_LOGIC; 
  signal rome2datao5_s_8_BYINV : STD_LOGIC; 
  signal nx53675z354_F5MUX : STD_LOGIC; 
  signal nx53675z356 : STD_LOGIC; 
  signal nx53675z354_BXINV : STD_LOGIC; 
  signal nx53675z355 : STD_LOGIC; 
  signal rome2datao5_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z365 : STD_LOGIC; 
  signal rome2datao5_s_7_BXINV : STD_LOGIC; 
  signal rome2datao5_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z364 : STD_LOGIC; 
  signal rome2datao5_s_7_BYINV : STD_LOGIC; 
  signal nx53675z360_F5MUX : STD_LOGIC; 
  signal nx53675z362 : STD_LOGIC; 
  signal nx53675z360_BXINV : STD_LOGIC; 
  signal nx53675z361 : STD_LOGIC; 
  signal rome2datao5_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z371 : STD_LOGIC; 
  signal rome2datao5_s_6_BXINV : STD_LOGIC; 
  signal rome2datao5_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z370 : STD_LOGIC; 
  signal rome2datao5_s_6_BYINV : STD_LOGIC; 
  signal nx53675z366_F5MUX : STD_LOGIC; 
  signal nx53675z368 : STD_LOGIC; 
  signal nx53675z366_BXINV : STD_LOGIC; 
  signal nx53675z367 : STD_LOGIC; 
  signal rome2datao7_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z477 : STD_LOGIC; 
  signal rome2datao7_s_10_BXINV : STD_LOGIC; 
  signal rome2datao7_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z476 : STD_LOGIC; 
  signal rome2datao7_s_10_BYINV : STD_LOGIC; 
  signal nx53675z472_F5MUX : STD_LOGIC; 
  signal nx53675z474 : STD_LOGIC; 
  signal nx53675z472_BXINV : STD_LOGIC; 
  signal nx53675z473 : STD_LOGIC; 
  signal rome2datao7_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z483 : STD_LOGIC; 
  signal rome2datao7_s_9_BXINV : STD_LOGIC; 
  signal rome2datao7_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z482 : STD_LOGIC; 
  signal rome2datao7_s_9_BYINV : STD_LOGIC; 
  signal nx53675z478_F5MUX : STD_LOGIC; 
  signal nx53675z480 : STD_LOGIC; 
  signal nx53675z478_BXINV : STD_LOGIC; 
  signal nx53675z479 : STD_LOGIC; 
  signal rome2datao7_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z489 : STD_LOGIC; 
  signal rome2datao7_s_8_BXINV : STD_LOGIC; 
  signal rome2datao7_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z488 : STD_LOGIC; 
  signal rome2datao7_s_8_BYINV : STD_LOGIC; 
  signal nx53675z484_F5MUX : STD_LOGIC; 
  signal nx53675z486 : STD_LOGIC; 
  signal nx53675z484_BXINV : STD_LOGIC; 
  signal nx53675z485 : STD_LOGIC; 
  signal rome2datao7_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z495 : STD_LOGIC; 
  signal rome2datao7_s_7_BXINV : STD_LOGIC; 
  signal rome2datao7_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z494 : STD_LOGIC; 
  signal rome2datao7_s_7_BYINV : STD_LOGIC; 
  signal nx53675z490_F5MUX : STD_LOGIC; 
  signal nx53675z492 : STD_LOGIC; 
  signal nx53675z490_BXINV : STD_LOGIC; 
  signal nx53675z491 : STD_LOGIC; 
  signal rome2datao7_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z501 : STD_LOGIC; 
  signal rome2datao7_s_6_BXINV : STD_LOGIC; 
  signal rome2datao7_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z500 : STD_LOGIC; 
  signal rome2datao7_s_6_BYINV : STD_LOGIC; 
  signal nx53675z496_F5MUX : STD_LOGIC; 
  signal nx53675z498 : STD_LOGIC; 
  signal nx53675z496_BXINV : STD_LOGIC; 
  signal nx53675z497 : STD_LOGIC; 
  signal romo2datao9_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z1434 : STD_LOGIC; 
  signal romo2datao9_s_12_BXINV : STD_LOGIC; 
  signal romo2datao9_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z1433 : STD_LOGIC; 
  signal romo2datao9_s_12_BYINV : STD_LOGIC; 
  signal nx53675z1429_F5MUX : STD_LOGIC; 
  signal nx53675z1431 : STD_LOGIC; 
  signal nx53675z1429_BXINV : STD_LOGIC; 
  signal nx53675z1430 : STD_LOGIC; 
  signal romo2datao5_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z1118 : STD_LOGIC; 
  signal romo2datao5_s_12_BXINV : STD_LOGIC; 
  signal romo2datao5_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z1117 : STD_LOGIC; 
  signal romo2datao5_s_12_BYINV : STD_LOGIC; 
  signal nx53675z1113_F5MUX : STD_LOGIC; 
  signal nx53675z1115 : STD_LOGIC; 
  signal nx53675z1113_BXINV : STD_LOGIC; 
  signal nx53675z1114 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_2_FFX_RST : STD_LOGIC; 
  signal romo2datao4_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z1099 : STD_LOGIC; 
  signal romo2datao4_s_2_BXINV : STD_LOGIC; 
  signal romo2datao4_s_2_F6MUX : STD_LOGIC; 
  signal nx53675z1098 : STD_LOGIC; 
  signal romo2datao4_s_2_BYINV : STD_LOGIC; 
  signal nx53675z1094_F5MUX : STD_LOGIC; 
  signal nx53675z1096 : STD_LOGIC; 
  signal nx53675z1094_BXINV : STD_LOGIC; 
  signal nx53675z1095 : STD_LOGIC; 
  signal rome2datao3_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z223 : STD_LOGIC; 
  signal rome2datao3_s_9_BXINV : STD_LOGIC; 
  signal rome2datao3_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z222 : STD_LOGIC; 
  signal rome2datao3_s_9_BYINV : STD_LOGIC; 
  signal nx53675z218_F5MUX : STD_LOGIC; 
  signal nx53675z220 : STD_LOGIC; 
  signal nx53675z218_BXINV : STD_LOGIC; 
  signal nx53675z219 : STD_LOGIC; 
  signal rome2datao3_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z247 : STD_LOGIC; 
  signal rome2datao3_s_5_BXINV : STD_LOGIC; 
  signal rome2datao3_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z246 : STD_LOGIC; 
  signal rome2datao3_s_5_BYINV : STD_LOGIC; 
  signal nx53675z242_F5MUX : STD_LOGIC; 
  signal nx53675z244 : STD_LOGIC; 
  signal nx53675z242_BXINV : STD_LOGIC; 
  signal nx53675z243 : STD_LOGIC; 
  signal rome2datao3_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z258 : STD_LOGIC; 
  signal rome2datao3_s_3_BXINV : STD_LOGIC; 
  signal rome2datao3_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z257 : STD_LOGIC; 
  signal rome2datao3_s_3_BYINV : STD_LOGIC; 
  signal nx53675z254_F5MUX : STD_LOGIC; 
  signal nx53675z255 : STD_LOGIC; 
  signal nx53675z254_BXINV : STD_LOGIC; 
  signal U2_ROME3_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal romo2datao4_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z1051 : STD_LOGIC; 
  signal romo2datao4_s_10_BXINV : STD_LOGIC; 
  signal romo2datao4_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z1050 : STD_LOGIC; 
  signal romo2datao4_s_10_BYINV : STD_LOGIC; 
  signal nx53675z1046_F5MUX : STD_LOGIC; 
  signal nx53675z1048 : STD_LOGIC; 
  signal nx53675z1046_BXINV : STD_LOGIC; 
  signal nx53675z1047 : STD_LOGIC; 
  signal romo2datao3_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z996 : STD_LOGIC; 
  signal romo2datao3_s_6_BXINV : STD_LOGIC; 
  signal romo2datao3_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z995 : STD_LOGIC; 
  signal romo2datao3_s_6_BYINV : STD_LOGIC; 
  signal nx53675z991_F5MUX : STD_LOGIC; 
  signal nx53675z993 : STD_LOGIC; 
  signal nx53675z991_BXINV : STD_LOGIC; 
  signal nx53675z992 : STD_LOGIC; 
  signal romo2datao3_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z1008 : STD_LOGIC; 
  signal romo2datao3_s_4_BXINV : STD_LOGIC; 
  signal romo2datao3_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z1007 : STD_LOGIC; 
  signal romo2datao3_s_4_BYINV : STD_LOGIC; 
  signal nx53675z1003_F5MUX : STD_LOGIC; 
  signal nx53675z1005 : STD_LOGIC; 
  signal nx53675z1003_BXINV : STD_LOGIC; 
  signal nx53675z1004 : STD_LOGIC; 
  signal romo2datao10_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z1561 : STD_LOGIC; 
  signal romo2datao10_s_4_BXINV : STD_LOGIC; 
  signal romo2datao10_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z1560 : STD_LOGIC; 
  signal romo2datao10_s_4_BYINV : STD_LOGIC; 
  signal nx53675z1556_F5MUX : STD_LOGIC; 
  signal nx53675z1558 : STD_LOGIC; 
  signal nx53675z1556_BXINV : STD_LOGIC; 
  signal nx53675z1557 : STD_LOGIC; 
  signal romo2datao10_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z1567 : STD_LOGIC; 
  signal romo2datao10_s_3_BXINV : STD_LOGIC; 
  signal romo2datao10_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z1566 : STD_LOGIC; 
  signal romo2datao10_s_3_BYINV : STD_LOGIC; 
  signal nx53675z1562_F5MUX : STD_LOGIC; 
  signal nx53675z1564 : STD_LOGIC; 
  signal nx53675z1562_BXINV : STD_LOGIC; 
  signal nx53675z1563 : STD_LOGIC; 
  signal romo2datao4_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z1057 : STD_LOGIC; 
  signal romo2datao4_s_9_BXINV : STD_LOGIC; 
  signal romo2datao4_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z1056 : STD_LOGIC; 
  signal romo2datao4_s_9_BYINV : STD_LOGIC; 
  signal nx53675z1052_F5MUX : STD_LOGIC; 
  signal nx53675z1054 : STD_LOGIC; 
  signal nx53675z1052_BXINV : STD_LOGIC; 
  signal nx53675z1053 : STD_LOGIC; 
  signal romo2datao4_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z1063 : STD_LOGIC; 
  signal romo2datao4_s_8_BXINV : STD_LOGIC; 
  signal romo2datao4_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z1062 : STD_LOGIC; 
  signal romo2datao4_s_8_BYINV : STD_LOGIC; 
  signal nx53675z1058_F5MUX : STD_LOGIC; 
  signal nx53675z1060 : STD_LOGIC; 
  signal nx53675z1058_BXINV : STD_LOGIC; 
  signal nx53675z1059 : STD_LOGIC; 
  signal romo2datao4_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z1069 : STD_LOGIC; 
  signal romo2datao4_s_7_BXINV : STD_LOGIC; 
  signal romo2datao4_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z1068 : STD_LOGIC; 
  signal romo2datao4_s_7_BYINV : STD_LOGIC; 
  signal nx53675z1064_F5MUX : STD_LOGIC; 
  signal nx53675z1066 : STD_LOGIC; 
  signal nx53675z1064_BXINV : STD_LOGIC; 
  signal nx53675z1065 : STD_LOGIC; 
  signal romo2datao4_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z1075 : STD_LOGIC; 
  signal romo2datao4_s_6_BXINV : STD_LOGIC; 
  signal romo2datao4_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z1074 : STD_LOGIC; 
  signal romo2datao4_s_6_BYINV : STD_LOGIC; 
  signal nx53675z1070_F5MUX : STD_LOGIC; 
  signal nx53675z1072 : STD_LOGIC; 
  signal nx53675z1070_BXINV : STD_LOGIC; 
  signal nx53675z1071 : STD_LOGIC; 
  signal rome2datao6_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z436 : STD_LOGIC; 
  signal rome2datao6_s_6_BXINV : STD_LOGIC; 
  signal rome2datao6_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z435 : STD_LOGIC; 
  signal rome2datao6_s_6_BYINV : STD_LOGIC; 
  signal nx53675z431_F5MUX : STD_LOGIC; 
  signal nx53675z433 : STD_LOGIC; 
  signal nx53675z431_BXINV : STD_LOGIC; 
  signal nx53675z432 : STD_LOGIC; 
  signal rome2datao6_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z442 : STD_LOGIC; 
  signal rome2datao6_s_5_BXINV : STD_LOGIC; 
  signal rome2datao6_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z441 : STD_LOGIC; 
  signal rome2datao6_s_5_BYINV : STD_LOGIC; 
  signal nx53675z437_F5MUX : STD_LOGIC; 
  signal nx53675z439 : STD_LOGIC; 
  signal nx53675z437_BXINV : STD_LOGIC; 
  signal nx53675z438 : STD_LOGIC; 
  signal romo2datao5_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z1124 : STD_LOGIC; 
  signal romo2datao5_s_11_BXINV : STD_LOGIC; 
  signal romo2datao5_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z1123 : STD_LOGIC; 
  signal romo2datao5_s_11_BYINV : STD_LOGIC; 
  signal nx53675z1119_F5MUX : STD_LOGIC; 
  signal nx53675z1121 : STD_LOGIC; 
  signal nx53675z1119_BXINV : STD_LOGIC; 
  signal nx53675z1120 : STD_LOGIC; 
  signal romo2datao9_s_1_F5MUX : STD_LOGIC; 
  signal nx53675z1500 : STD_LOGIC; 
  signal romo2datao9_s_1_BXINV : STD_LOGIC; 
  signal romo2datao9_s_1_F6MUX : STD_LOGIC; 
  signal nx53675z1499 : STD_LOGIC; 
  signal romo2datao9_s_1_BYINV : STD_LOGIC; 
  signal nx53675z1495_F5MUX : STD_LOGIC; 
  signal nx53675z1497 : STD_LOGIC; 
  signal nx53675z1495_BXINV : STD_LOGIC; 
  signal nx53675z1496 : STD_LOGIC; 
  signal romo2datao6_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z1191 : STD_LOGIC; 
  signal romo2datao6_s_13_BXINV : STD_LOGIC; 
  signal romo2datao6_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z1190 : STD_LOGIC; 
  signal romo2datao6_s_13_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_4_FFX_RST : STD_LOGIC; 
  signal nx53675z1187_F5MUX : STD_LOGIC; 
  signal nx53675z1188 : STD_LOGIC; 
  signal nx53675z1187_BXINV : STD_LOGIC; 
  signal nx53675z1187_G : STD_LOGIC; 
  signal romo2datao6_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z1233 : STD_LOGIC; 
  signal romo2datao6_s_6_BXINV : STD_LOGIC; 
  signal romo2datao6_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z1232 : STD_LOGIC; 
  signal romo2datao6_s_6_BYINV : STD_LOGIC; 
  signal nx53675z1228_F5MUX : STD_LOGIC; 
  signal nx53675z1230 : STD_LOGIC; 
  signal nx53675z1228_BXINV : STD_LOGIC; 
  signal nx53675z1229 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_FFY_RST : STD_LOGIC; 
  signal romo2datao6_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z1239 : STD_LOGIC; 
  signal romo2datao6_s_5_BXINV : STD_LOGIC; 
  signal romo2datao6_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z1238 : STD_LOGIC; 
  signal romo2datao6_s_5_BYINV : STD_LOGIC; 
  signal nx53675z1234_F5MUX : STD_LOGIC; 
  signal nx53675z1236 : STD_LOGIC; 
  signal nx53675z1234_BXINV : STD_LOGIC; 
  signal nx53675z1235 : STD_LOGIC; 
  signal romo2datao6_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z1245 : STD_LOGIC; 
  signal romo2datao6_s_4_BXINV : STD_LOGIC; 
  signal romo2datao6_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z1244 : STD_LOGIC; 
  signal romo2datao6_s_4_BYINV : STD_LOGIC; 
  signal nx53675z1240_F5MUX : STD_LOGIC; 
  signal nx53675z1242 : STD_LOGIC; 
  signal nx53675z1240_BXINV : STD_LOGIC; 
  signal nx53675z1241 : STD_LOGIC; 
  signal romo2datao6_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z1251 : STD_LOGIC; 
  signal romo2datao6_s_3_BXINV : STD_LOGIC; 
  signal romo2datao6_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z1250 : STD_LOGIC; 
  signal romo2datao6_s_3_BYINV : STD_LOGIC; 
  signal nx53675z1246_F5MUX : STD_LOGIC; 
  signal nx53675z1248 : STD_LOGIC; 
  signal nx53675z1246_BXINV : STD_LOGIC; 
  signal nx53675z1247 : STD_LOGIC; 
  signal romo2datao6_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z1257 : STD_LOGIC; 
  signal romo2datao6_s_2_BXINV : STD_LOGIC; 
  signal romo2datao6_s_2_F6MUX : STD_LOGIC; 
  signal nx53675z1256 : STD_LOGIC; 
  signal romo2datao6_s_2_BYINV : STD_LOGIC; 
  signal nx53675z1252_F5MUX : STD_LOGIC; 
  signal nx53675z1254 : STD_LOGIC; 
  signal nx53675z1252_BXINV : STD_LOGIC; 
  signal nx53675z1253 : STD_LOGIC; 
  signal romo2datao5_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z1130 : STD_LOGIC; 
  signal romo2datao5_s_10_BXINV : STD_LOGIC; 
  signal romo2datao5_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z1129 : STD_LOGIC; 
  signal romo2datao5_s_10_BYINV : STD_LOGIC; 
  signal nx53675z1125_F5MUX : STD_LOGIC; 
  signal nx53675z1127 : STD_LOGIC; 
  signal nx53675z1125_BXINV : STD_LOGIC; 
  signal nx53675z1126 : STD_LOGIC; 
  signal romo2datao5_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z1136 : STD_LOGIC; 
  signal romo2datao5_s_9_BXINV : STD_LOGIC; 
  signal romo2datao5_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z1135 : STD_LOGIC; 
  signal romo2datao5_s_9_BYINV : STD_LOGIC; 
  signal nx53675z1131_F5MUX : STD_LOGIC; 
  signal nx53675z1133 : STD_LOGIC; 
  signal nx53675z1131_BXINV : STD_LOGIC; 
  signal nx53675z1132 : STD_LOGIC; 
  signal romo2datao5_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z1142 : STD_LOGIC; 
  signal romo2datao5_s_8_BXINV : STD_LOGIC; 
  signal romo2datao5_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z1141 : STD_LOGIC; 
  signal romo2datao5_s_8_BYINV : STD_LOGIC; 
  signal nx53675z1137_F5MUX : STD_LOGIC; 
  signal nx53675z1139 : STD_LOGIC; 
  signal nx53675z1137_BXINV : STD_LOGIC; 
  signal nx53675z1138 : STD_LOGIC; 
  signal romo2datao5_s_2_F5MUX : STD_LOGIC; 
  signal nx53675z1178 : STD_LOGIC; 
  signal romo2datao5_s_2_BXINV : STD_LOGIC; 
  signal romo2datao5_s_2_F6MUX : STD_LOGIC; 
  signal nx53675z1177 : STD_LOGIC; 
  signal romo2datao5_s_2_BYINV : STD_LOGIC; 
  signal nx53675z1173_F5MUX : STD_LOGIC; 
  signal nx53675z1175 : STD_LOGIC; 
  signal nx53675z1173_BXINV : STD_LOGIC; 
  signal nx53675z1174 : STD_LOGIC; 
  signal romo2datao5_s_1_F5MUX : STD_LOGIC; 
  signal nx53675z1184 : STD_LOGIC; 
  signal romo2datao5_s_1_BXINV : STD_LOGIC; 
  signal romo2datao5_s_1_F6MUX : STD_LOGIC; 
  signal nx53675z1183 : STD_LOGIC; 
  signal romo2datao5_s_1_BYINV : STD_LOGIC; 
  signal nx53675z1179_F5MUX : STD_LOGIC; 
  signal nx53675z1181 : STD_LOGIC; 
  signal nx53675z1179_BXINV : STD_LOGIC; 
  signal nx53675z1180 : STD_LOGIC; 
  signal romo2datao5_s_0_F5MUX : STD_LOGIC; 
  signal nx53675z1186 : STD_LOGIC; 
  signal romo2datao5_s_0_BXINV : STD_LOGIC; 
  signal romo2datao5_s_0_F6MUX : STD_LOGIC; 
  signal nx53675z1185 : STD_LOGIC; 
  signal romo2datao5_s_0_BYINV : STD_LOGIC; 
  signal U2_ROMO5_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROMO5_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROMO5_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROMO5_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romo2datao3_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z966 : STD_LOGIC; 
  signal romo2datao3_s_11_BXINV : STD_LOGIC; 
  signal romo2datao3_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z965 : STD_LOGIC; 
  signal romo2datao3_s_11_BYINV : STD_LOGIC; 
  signal nx53675z961_F5MUX : STD_LOGIC; 
  signal nx53675z963 : STD_LOGIC; 
  signal nx53675z961_BXINV : STD_LOGIC; 
  signal nx53675z962 : STD_LOGIC; 
  signal romo2datao2_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z935 : STD_LOGIC; 
  signal romo2datao2_s_3_BXINV : STD_LOGIC; 
  signal romo2datao2_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z934 : STD_LOGIC; 
  signal romo2datao2_s_3_BYINV : STD_LOGIC; 
  signal nx53675z930_F5MUX : STD_LOGIC; 
  signal nx53675z932 : STD_LOGIC; 
  signal nx53675z930_BXINV : STD_LOGIC; 
  signal nx53675z931 : STD_LOGIC; 
  signal rome2datao8_s_8_F5MUX : STD_LOGIC; 
  signal nx53675z554 : STD_LOGIC; 
  signal rome2datao8_s_8_BXINV : STD_LOGIC; 
  signal rome2datao8_s_8_F6MUX : STD_LOGIC; 
  signal nx53675z553 : STD_LOGIC; 
  signal rome2datao8_s_8_BYINV : STD_LOGIC; 
  signal nx53675z549_F5MUX : STD_LOGIC; 
  signal nx53675z551 : STD_LOGIC; 
  signal nx53675z549_BXINV : STD_LOGIC; 
  signal nx53675z550 : STD_LOGIC; 
  signal rome2datao8_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z560 : STD_LOGIC; 
  signal rome2datao8_s_7_BXINV : STD_LOGIC; 
  signal rome2datao8_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z559 : STD_LOGIC; 
  signal rome2datao8_s_7_BYINV : STD_LOGIC; 
  signal nx53675z555_F5MUX : STD_LOGIC; 
  signal nx53675z557 : STD_LOGIC; 
  signal nx53675z555_BXINV : STD_LOGIC; 
  signal nx53675z556 : STD_LOGIC; 
  signal rome2datao8_s_6_F5MUX : STD_LOGIC; 
  signal nx53675z566 : STD_LOGIC; 
  signal rome2datao8_s_6_BXINV : STD_LOGIC; 
  signal rome2datao8_s_6_F6MUX : STD_LOGIC; 
  signal nx53675z565 : STD_LOGIC; 
  signal rome2datao8_s_6_BYINV : STD_LOGIC; 
  signal nx53675z561_F5MUX : STD_LOGIC; 
  signal nx53675z563 : STD_LOGIC; 
  signal nx53675z561_BXINV : STD_LOGIC; 
  signal nx53675z562 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_4_FFX_RST : STD_LOGIC; 
  signal rome2datao8_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z572 : STD_LOGIC; 
  signal rome2datao8_s_5_BXINV : STD_LOGIC; 
  signal rome2datao8_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z571 : STD_LOGIC; 
  signal rome2datao8_s_5_BYINV : STD_LOGIC; 
  signal nx53675z567_F5MUX : STD_LOGIC; 
  signal nx53675z569 : STD_LOGIC; 
  signal nx53675z567_BXINV : STD_LOGIC; 
  signal nx53675z568 : STD_LOGIC; 
  signal rome2datao8_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z578 : STD_LOGIC; 
  signal rome2datao8_s_4_BXINV : STD_LOGIC; 
  signal rome2datao8_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z577 : STD_LOGIC; 
  signal rome2datao8_s_4_BYINV : STD_LOGIC; 
  signal nx53675z573_F5MUX : STD_LOGIC; 
  signal nx53675z575 : STD_LOGIC; 
  signal nx53675z573_BXINV : STD_LOGIC; 
  signal nx53675z574 : STD_LOGIC; 
  signal rome2datao7_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z507 : STD_LOGIC; 
  signal rome2datao7_s_5_BXINV : STD_LOGIC; 
  signal rome2datao7_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z506 : STD_LOGIC; 
  signal rome2datao7_s_5_BYINV : STD_LOGIC; 
  signal nx53675z502_F5MUX : STD_LOGIC; 
  signal nx53675z504 : STD_LOGIC; 
  signal nx53675z502_BXINV : STD_LOGIC; 
  signal nx53675z503 : STD_LOGIC; 
  signal rome2datao7_s_4_F5MUX : STD_LOGIC; 
  signal nx53675z513 : STD_LOGIC; 
  signal rome2datao7_s_4_BXINV : STD_LOGIC; 
  signal rome2datao7_s_4_F6MUX : STD_LOGIC; 
  signal nx53675z512 : STD_LOGIC; 
  signal rome2datao7_s_4_BYINV : STD_LOGIC; 
  signal nx53675z508_F5MUX : STD_LOGIC; 
  signal nx53675z510 : STD_LOGIC; 
  signal nx53675z508_BXINV : STD_LOGIC; 
  signal nx53675z509 : STD_LOGIC; 
  signal romo2datao6_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z1197 : STD_LOGIC; 
  signal romo2datao6_s_12_BXINV : STD_LOGIC; 
  signal romo2datao6_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z1196 : STD_LOGIC; 
  signal romo2datao6_s_12_BYINV : STD_LOGIC; 
  signal nx53675z1192_F5MUX : STD_LOGIC; 
  signal nx53675z1194 : STD_LOGIC; 
  signal nx53675z1192_BXINV : STD_LOGIC; 
  signal nx53675z1193 : STD_LOGIC; 
  signal romo2datao7_s_12_F5MUX : STD_LOGIC; 
  signal nx53675z1276 : STD_LOGIC; 
  signal romo2datao7_s_12_BXINV : STD_LOGIC; 
  signal romo2datao7_s_12_F6MUX : STD_LOGIC; 
  signal nx53675z1275 : STD_LOGIC; 
  signal romo2datao7_s_12_BYINV : STD_LOGIC; 
  signal nx53675z1271_F5MUX : STD_LOGIC; 
  signal nx53675z1273 : STD_LOGIC; 
  signal nx53675z1271_BXINV : STD_LOGIC; 
  signal nx53675z1272 : STD_LOGIC; 
  signal romo2datao7_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z1282 : STD_LOGIC; 
  signal romo2datao7_s_11_BXINV : STD_LOGIC; 
  signal romo2datao7_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z1281 : STD_LOGIC; 
  signal romo2datao7_s_11_BYINV : STD_LOGIC; 
  signal nx53675z1277_F5MUX : STD_LOGIC; 
  signal nx53675z1279 : STD_LOGIC; 
  signal nx53675z1277_BXINV : STD_LOGIC; 
  signal nx53675z1278 : STD_LOGIC; 
  signal romo2datao6_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z1203 : STD_LOGIC; 
  signal romo2datao6_s_11_BXINV : STD_LOGIC; 
  signal romo2datao6_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z1202 : STD_LOGIC; 
  signal romo2datao6_s_11_BYINV : STD_LOGIC; 
  signal nx53675z1198_F5MUX : STD_LOGIC; 
  signal nx53675z1200 : STD_LOGIC; 
  signal nx53675z1198_BXINV : STD_LOGIC; 
  signal nx53675z1199 : STD_LOGIC; 
  signal romo2datao6_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z1209 : STD_LOGIC; 
  signal romo2datao6_s_10_BXINV : STD_LOGIC; 
  signal romo2datao6_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z1208 : STD_LOGIC; 
  signal romo2datao6_s_10_BYINV : STD_LOGIC; 
  signal nx53675z1204_F5MUX : STD_LOGIC; 
  signal nx53675z1206 : STD_LOGIC; 
  signal nx53675z1204_BXINV : STD_LOGIC; 
  signal nx53675z1205 : STD_LOGIC; 
  signal romo2datao6_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z1215 : STD_LOGIC; 
  signal romo2datao6_s_9_BXINV : STD_LOGIC; 
  signal romo2datao6_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z1214 : STD_LOGIC; 
  signal romo2datao6_s_9_BYINV : STD_LOGIC; 
  signal nx53675z1210_F5MUX : STD_LOGIC; 
  signal nx53675z1212 : STD_LOGIC; 
  signal nx53675z1210_BXINV : STD_LOGIC; 
  signal nx53675z1211 : STD_LOGIC; 
  signal romo2datao6_s_1_F5MUX : STD_LOGIC; 
  signal nx53675z1263 : STD_LOGIC; 
  signal romo2datao6_s_1_BXINV : STD_LOGIC; 
  signal romo2datao6_s_1_F6MUX : STD_LOGIC; 
  signal nx53675z1262 : STD_LOGIC; 
  signal romo2datao6_s_1_BYINV : STD_LOGIC; 
  signal nx53675z1258_F5MUX : STD_LOGIC; 
  signal nx53675z1260 : STD_LOGIC; 
  signal nx53675z1258_BXINV : STD_LOGIC; 
  signal nx53675z1259 : STD_LOGIC; 
  signal romo2datao5_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z1148 : STD_LOGIC; 
  signal romo2datao5_s_7_BXINV : STD_LOGIC; 
  signal romo2datao5_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z1147 : STD_LOGIC; 
  signal romo2datao5_s_7_BYINV : STD_LOGIC; 
  signal nx53675z1143_F5MUX : STD_LOGIC; 
  signal nx53675z1145 : STD_LOGIC; 
  signal nx53675z1143_BXINV : STD_LOGIC; 
  signal nx53675z1144 : STD_LOGIC; 
  signal romo2datao3_s_9_F5MUX : STD_LOGIC; 
  signal nx53675z978 : STD_LOGIC; 
  signal romo2datao3_s_9_BXINV : STD_LOGIC; 
  signal romo2datao3_s_9_F6MUX : STD_LOGIC; 
  signal nx53675z977 : STD_LOGIC; 
  signal romo2datao3_s_9_BYINV : STD_LOGIC; 
  signal nx53675z973_F5MUX : STD_LOGIC; 
  signal nx53675z975 : STD_LOGIC; 
  signal nx53675z973_BXINV : STD_LOGIC; 
  signal nx53675z974 : STD_LOGIC; 
  signal rome2datao8_s_3_F5MUX : STD_LOGIC; 
  signal nx53675z583 : STD_LOGIC; 
  signal rome2datao8_s_3_BXINV : STD_LOGIC; 
  signal rome2datao8_s_3_F6MUX : STD_LOGIC; 
  signal nx53675z582 : STD_LOGIC; 
  signal rome2datao8_s_3_BYINV : STD_LOGIC; 
  signal nx53675z579_F5MUX : STD_LOGIC; 
  signal nx53675z580 : STD_LOGIC; 
  signal nx53675z579_BXINV : STD_LOGIC; 
  signal U2_ROME8_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal romo2datao6_s_0_F5MUX : STD_LOGIC; 
  signal nx53675z1265 : STD_LOGIC; 
  signal romo2datao6_s_0_BXINV : STD_LOGIC; 
  signal romo2datao6_s_0_F6MUX : STD_LOGIC; 
  signal nx53675z1264 : STD_LOGIC; 
  signal romo2datao6_s_0_BYINV : STD_LOGIC; 
  signal U2_ROMO6_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U2_ROMO6_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U2_ROMO6_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U2_ROMO6_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romo2datao10_s_11_F5MUX : STD_LOGIC; 
  signal nx53675z1519 : STD_LOGIC; 
  signal romo2datao10_s_11_BXINV : STD_LOGIC; 
  signal romo2datao10_s_11_F6MUX : STD_LOGIC; 
  signal nx53675z1518 : STD_LOGIC; 
  signal romo2datao10_s_11_BYINV : STD_LOGIC; 
  signal nx53675z1514_F5MUX : STD_LOGIC; 
  signal nx53675z1516 : STD_LOGIC; 
  signal nx53675z1514_BXINV : STD_LOGIC; 
  signal nx53675z1515 : STD_LOGIC; 
  signal romo2datao7_s_13_F5MUX : STD_LOGIC; 
  signal nx53675z1270 : STD_LOGIC; 
  signal romo2datao7_s_13_BXINV : STD_LOGIC; 
  signal romo2datao7_s_13_F6MUX : STD_LOGIC; 
  signal nx53675z1269 : STD_LOGIC; 
  signal romo2datao7_s_13_BYINV : STD_LOGIC; 
  signal nx53675z1266_F5MUX : STD_LOGIC; 
  signal nx53675z1267 : STD_LOGIC; 
  signal nx53675z1266_BXINV : STD_LOGIC; 
  signal nx53675z1266_G : STD_LOGIC; 
  signal romo2datao7_s_10_F5MUX : STD_LOGIC; 
  signal nx53675z1288 : STD_LOGIC; 
  signal romo2datao7_s_10_BXINV : STD_LOGIC; 
  signal romo2datao7_s_10_F6MUX : STD_LOGIC; 
  signal nx53675z1287 : STD_LOGIC; 
  signal romo2datao7_s_10_BYINV : STD_LOGIC; 
  signal nx53675z1283_F5MUX : STD_LOGIC; 
  signal nx53675z1285 : STD_LOGIC; 
  signal nx53675z1283_BXINV : STD_LOGIC; 
  signal nx53675z1284 : STD_LOGIC; 
  signal romo2datao3_s_7_F5MUX : STD_LOGIC; 
  signal nx53675z990 : STD_LOGIC; 
  signal romo2datao3_s_7_BXINV : STD_LOGIC; 
  signal romo2datao3_s_7_F6MUX : STD_LOGIC; 
  signal nx53675z989 : STD_LOGIC; 
  signal romo2datao3_s_7_BYINV : STD_LOGIC; 
  signal nx53675z985_F5MUX : STD_LOGIC; 
  signal nx53675z987 : STD_LOGIC; 
  signal nx53675z985_BXINV : STD_LOGIC; 
  signal nx53675z986 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_FFY_RST : STD_LOGIC; 
  signal romo2datao3_s_5_F5MUX : STD_LOGIC; 
  signal nx53675z1002 : STD_LOGIC; 
  signal romo2datao3_s_5_BXINV : STD_LOGIC; 
  signal romo2datao3_s_5_F6MUX : STD_LOGIC; 
  signal nx53675z1001 : STD_LOGIC; 
  signal romo2datao3_s_5_BYINV : STD_LOGIC; 
  signal nx53675z997_F5MUX : STD_LOGIC; 
  signal nx53675z999 : STD_LOGIC; 
  signal nx53675z997_BXINV : STD_LOGIC; 
  signal nx53675z998 : STD_LOGIC; 
  signal romedatao0_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z23 : STD_LOGIC; 
  signal romedatao0_s_10_BXINV : STD_LOGIC; 
  signal romedatao0_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z22 : STD_LOGIC; 
  signal romedatao0_s_10_BYINV : STD_LOGIC; 
  signal nx54672z18_F5MUX : STD_LOGIC; 
  signal nx54672z20 : STD_LOGIC; 
  signal nx54672z18_BXINV : STD_LOGIC; 
  signal nx54672z19 : STD_LOGIC; 
  signal romedatao0_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z29 : STD_LOGIC; 
  signal romedatao0_s_9_BXINV : STD_LOGIC; 
  signal romedatao0_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z28 : STD_LOGIC; 
  signal romedatao0_s_9_BYINV : STD_LOGIC; 
  signal nx54672z24_F5MUX : STD_LOGIC; 
  signal nx54672z26 : STD_LOGIC; 
  signal nx54672z24_BXINV : STD_LOGIC; 
  signal nx54672z25 : STD_LOGIC; 
  signal romodatao0_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z589 : STD_LOGIC; 
  signal romodatao0_s_13_BXINV : STD_LOGIC; 
  signal romodatao0_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z588 : STD_LOGIC; 
  signal romodatao0_s_13_BYINV : STD_LOGIC; 
  signal nx54672z585_F5MUX : STD_LOGIC; 
  signal nx54672z586 : STD_LOGIC; 
  signal nx54672z585_BXINV : STD_LOGIC; 
  signal nx54672z585_G : STD_LOGIC; 
  signal romedatao8_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z584 : STD_LOGIC; 
  signal romedatao8_s_2_BXINV : STD_LOGIC; 
  signal romedatao8_s_2_F6MUX : STD_LOGIC; 
  signal romedatao8_s_2_G : STD_LOGIC; 
  signal romedatao8_s_2_BYINV : STD_LOGIC; 
  signal U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROME8_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romedatao2_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z164 : STD_LOGIC; 
  signal romedatao2_s_8_BXINV : STD_LOGIC; 
  signal romedatao2_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z163 : STD_LOGIC; 
  signal romedatao2_s_8_BYINV : STD_LOGIC; 
  signal nx54672z159_F5MUX : STD_LOGIC; 
  signal nx54672z161 : STD_LOGIC; 
  signal nx54672z159_BXINV : STD_LOGIC; 
  signal nx54672z160 : STD_LOGIC; 
  signal romodatao1_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z672 : STD_LOGIC; 
  signal romodatao1_s_12_BXINV : STD_LOGIC; 
  signal romodatao1_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z671 : STD_LOGIC; 
  signal romodatao1_s_12_BYINV : STD_LOGIC; 
  signal nx54672z667_F5MUX : STD_LOGIC; 
  signal nx54672z669 : STD_LOGIC; 
  signal nx54672z667_BXINV : STD_LOGIC; 
  signal nx54672z668 : STD_LOGIC; 
  signal romodatao1_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z678 : STD_LOGIC; 
  signal romodatao1_s_11_BXINV : STD_LOGIC; 
  signal romodatao1_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z677 : STD_LOGIC; 
  signal romodatao1_s_11_BYINV : STD_LOGIC; 
  signal nx54672z673_F5MUX : STD_LOGIC; 
  signal nx54672z675 : STD_LOGIC; 
  signal nx54672z673_BXINV : STD_LOGIC; 
  signal nx54672z674 : STD_LOGIC; 
  signal romodatao1_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z732 : STD_LOGIC; 
  signal romodatao1_s_2_BXINV : STD_LOGIC; 
  signal romodatao1_s_2_F6MUX : STD_LOGIC; 
  signal nx54672z731 : STD_LOGIC; 
  signal romodatao1_s_2_BYINV : STD_LOGIC; 
  signal nx54672z727_F5MUX : STD_LOGIC; 
  signal nx54672z729 : STD_LOGIC; 
  signal nx54672z727_BXINV : STD_LOGIC; 
  signal nx54672z728 : STD_LOGIC; 
  signal romodatao1_s_1_F5MUX : STD_LOGIC; 
  signal nx54672z738 : STD_LOGIC; 
  signal romodatao1_s_1_BXINV : STD_LOGIC; 
  signal romodatao1_s_1_F6MUX : STD_LOGIC; 
  signal nx54672z737 : STD_LOGIC; 
  signal romodatao1_s_1_BYINV : STD_LOGIC; 
  signal nx54672z733_F5MUX : STD_LOGIC; 
  signal nx54672z735 : STD_LOGIC; 
  signal nx54672z733_BXINV : STD_LOGIC; 
  signal nx54672z734 : STD_LOGIC; 
  signal romedatao1_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z99 : STD_LOGIC; 
  signal romedatao1_s_8_BXINV : STD_LOGIC; 
  signal romedatao1_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z98 : STD_LOGIC; 
  signal romedatao1_s_8_BYINV : STD_LOGIC; 
  signal nx54672z94_F5MUX : STD_LOGIC; 
  signal nx54672z96 : STD_LOGIC; 
  signal nx54672z94_BXINV : STD_LOGIC; 
  signal nx54672z95 : STD_LOGIC; 
  signal romedatao1_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z105 : STD_LOGIC; 
  signal romedatao1_s_7_BXINV : STD_LOGIC; 
  signal romedatao1_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z104 : STD_LOGIC; 
  signal romedatao1_s_7_BYINV : STD_LOGIC; 
  signal nx54672z100_F5MUX : STD_LOGIC; 
  signal nx54672z102 : STD_LOGIC; 
  signal nx54672z100_BXINV : STD_LOGIC; 
  signal nx54672z101 : STD_LOGIC; 
  signal romedatao1_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z111 : STD_LOGIC; 
  signal romedatao1_s_6_BXINV : STD_LOGIC; 
  signal romedatao1_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z110 : STD_LOGIC; 
  signal romedatao1_s_6_BYINV : STD_LOGIC; 
  signal nx54672z106_F5MUX : STD_LOGIC; 
  signal nx54672z108 : STD_LOGIC; 
  signal nx54672z106_BXINV : STD_LOGIC; 
  signal nx54672z107 : STD_LOGIC; 
  signal romedatao1_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z117 : STD_LOGIC; 
  signal romedatao1_s_5_BXINV : STD_LOGIC; 
  signal romedatao1_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z116 : STD_LOGIC; 
  signal romedatao1_s_5_BYINV : STD_LOGIC; 
  signal nx54672z112_F5MUX : STD_LOGIC; 
  signal nx54672z114 : STD_LOGIC; 
  signal nx54672z112_BXINV : STD_LOGIC; 
  signal nx54672z113 : STD_LOGIC; 
  signal romedatao0_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z35 : STD_LOGIC; 
  signal romedatao0_s_8_BXINV : STD_LOGIC; 
  signal romedatao0_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z34 : STD_LOGIC; 
  signal romedatao0_s_8_BYINV : STD_LOGIC; 
  signal nx54672z30_F5MUX : STD_LOGIC; 
  signal nx54672z32 : STD_LOGIC; 
  signal nx54672z30_BXINV : STD_LOGIC; 
  signal nx54672z31 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_6_FFX_RST : STD_LOGIC; 
  signal romedatao0_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z41 : STD_LOGIC; 
  signal romedatao0_s_7_BXINV : STD_LOGIC; 
  signal romedatao0_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z40 : STD_LOGIC; 
  signal romedatao0_s_7_BYINV : STD_LOGIC; 
  signal nx54672z36_F5MUX : STD_LOGIC; 
  signal nx54672z38 : STD_LOGIC; 
  signal nx54672z36_BXINV : STD_LOGIC; 
  signal nx54672z37 : STD_LOGIC; 
  signal romedatao0_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z47 : STD_LOGIC; 
  signal romedatao0_s_6_BXINV : STD_LOGIC; 
  signal romedatao0_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z46 : STD_LOGIC; 
  signal romedatao0_s_6_BYINV : STD_LOGIC; 
  signal nx54672z42_F5MUX : STD_LOGIC; 
  signal nx54672z44 : STD_LOGIC; 
  signal nx54672z42_BXINV : STD_LOGIC; 
  signal nx54672z43 : STD_LOGIC; 
  signal romedatao0_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z53 : STD_LOGIC; 
  signal romedatao0_s_5_BXINV : STD_LOGIC; 
  signal romedatao0_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z52 : STD_LOGIC; 
  signal romedatao0_s_5_BYINV : STD_LOGIC; 
  signal nx54672z48_F5MUX : STD_LOGIC; 
  signal nx54672z50 : STD_LOGIC; 
  signal nx54672z48_BXINV : STD_LOGIC; 
  signal nx54672z49 : STD_LOGIC; 
  signal romedatao0_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z59 : STD_LOGIC; 
  signal romedatao0_s_4_BXINV : STD_LOGIC; 
  signal romedatao0_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z58 : STD_LOGIC; 
  signal romedatao0_s_4_BYINV : STD_LOGIC; 
  signal nx54672z54_F5MUX : STD_LOGIC; 
  signal nx54672z56 : STD_LOGIC; 
  signal nx54672z54_BXINV : STD_LOGIC; 
  signal nx54672z55 : STD_LOGIC; 
  signal romodatao8_s_0_F5MUX : STD_LOGIC; 
  signal nx54672z1293 : STD_LOGIC; 
  signal romodatao8_s_0_BXINV : STD_LOGIC; 
  signal romodatao8_s_0_F6MUX : STD_LOGIC; 
  signal nx54672z1292 : STD_LOGIC; 
  signal romodatao8_s_0_BYINV : STD_LOGIC; 
  signal U1_ROMO8_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROMO8_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROMO8_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROMO8_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romodatao1_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z666 : STD_LOGIC; 
  signal romodatao1_s_13_BXINV : STD_LOGIC; 
  signal romodatao1_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z665 : STD_LOGIC; 
  signal romodatao1_s_13_BYINV : STD_LOGIC; 
  signal nx54672z662_F5MUX : STD_LOGIC; 
  signal nx54672z663 : STD_LOGIC; 
  signal nx54672z662_BXINV : STD_LOGIC; 
  signal nx54672z662_G : STD_LOGIC; 
  signal romodatao0_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z595 : STD_LOGIC; 
  signal romodatao0_s_12_BXINV : STD_LOGIC; 
  signal romodatao0_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z594 : STD_LOGIC; 
  signal romodatao0_s_12_BYINV : STD_LOGIC; 
  signal nx54672z590_F5MUX : STD_LOGIC; 
  signal nx54672z592 : STD_LOGIC; 
  signal nx54672z590_BXINV : STD_LOGIC; 
  signal nx54672z591 : STD_LOGIC; 
  signal romodatao0_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z601 : STD_LOGIC; 
  signal romodatao0_s_11_BXINV : STD_LOGIC; 
  signal romodatao0_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z600 : STD_LOGIC; 
  signal romodatao0_s_11_BYINV : STD_LOGIC; 
  signal nx54672z596_F5MUX : STD_LOGIC; 
  signal nx54672z598 : STD_LOGIC; 
  signal nx54672z596_BXINV : STD_LOGIC; 
  signal nx54672z597 : STD_LOGIC; 
  signal romodatao0_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z607 : STD_LOGIC; 
  signal romodatao0_s_10_BXINV : STD_LOGIC; 
  signal romodatao0_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z606 : STD_LOGIC; 
  signal romodatao0_s_10_BYINV : STD_LOGIC; 
  signal nx54672z602_F5MUX : STD_LOGIC; 
  signal nx54672z604 : STD_LOGIC; 
  signal nx54672z602_BXINV : STD_LOGIC; 
  signal nx54672z603 : STD_LOGIC; 
  signal romodatao0_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z613 : STD_LOGIC; 
  signal romodatao0_s_9_BXINV : STD_LOGIC; 
  signal romodatao0_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z612 : STD_LOGIC; 
  signal romodatao0_s_9_BYINV : STD_LOGIC; 
  signal nx54672z608_F5MUX : STD_LOGIC; 
  signal nx54672z610 : STD_LOGIC; 
  signal nx54672z608_BXINV : STD_LOGIC; 
  signal nx54672z609 : STD_LOGIC; 
  signal romodatao0_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z619 : STD_LOGIC; 
  signal romodatao0_s_8_BXINV : STD_LOGIC; 
  signal romodatao0_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z618 : STD_LOGIC; 
  signal romodatao0_s_8_BYINV : STD_LOGIC; 
  signal nx54672z614_F5MUX : STD_LOGIC; 
  signal nx54672z616 : STD_LOGIC; 
  signal nx54672z614_BXINV : STD_LOGIC; 
  signal nx54672z615 : STD_LOGIC; 
  signal romodatao0_s_1_F5MUX : STD_LOGIC; 
  signal nx54672z661 : STD_LOGIC; 
  signal romodatao0_s_1_BXINV : STD_LOGIC; 
  signal romodatao0_s_1_F6MUX : STD_LOGIC; 
  signal nx54672z660 : STD_LOGIC; 
  signal romodatao0_s_1_BYINV : STD_LOGIC; 
  signal nx54672z656_F5MUX : STD_LOGIC; 
  signal nx54672z658 : STD_LOGIC; 
  signal nx54672z656_BXINV : STD_LOGIC; 
  signal nx54672z657 : STD_LOGIC; 
  signal romedatao2_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z170 : STD_LOGIC; 
  signal romedatao2_s_7_BXINV : STD_LOGIC; 
  signal romedatao2_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z169 : STD_LOGIC; 
  signal romedatao2_s_7_BYINV : STD_LOGIC; 
  signal nx54672z165_F5MUX : STD_LOGIC; 
  signal nx54672z167 : STD_LOGIC; 
  signal nx54672z165_BXINV : STD_LOGIC; 
  signal nx54672z166 : STD_LOGIC; 
  signal romedatao2_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z176 : STD_LOGIC; 
  signal romedatao2_s_6_BXINV : STD_LOGIC; 
  signal romedatao2_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z175 : STD_LOGIC; 
  signal romedatao2_s_6_BYINV : STD_LOGIC; 
  signal nx54672z171_F5MUX : STD_LOGIC; 
  signal nx54672z173 : STD_LOGIC; 
  signal nx54672z171_BXINV : STD_LOGIC; 
  signal nx54672z172 : STD_LOGIC; 
  signal romedatao2_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z182 : STD_LOGIC; 
  signal romedatao2_s_5_BXINV : STD_LOGIC; 
  signal romedatao2_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z181 : STD_LOGIC; 
  signal romedatao2_s_5_BYINV : STD_LOGIC; 
  signal nx54672z177_F5MUX : STD_LOGIC; 
  signal nx54672z179 : STD_LOGIC; 
  signal nx54672z177_BXINV : STD_LOGIC; 
  signal nx54672z178 : STD_LOGIC; 
  signal romedatao2_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z188 : STD_LOGIC; 
  signal romedatao2_s_4_BXINV : STD_LOGIC; 
  signal romedatao2_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z187 : STD_LOGIC; 
  signal romedatao2_s_4_BYINV : STD_LOGIC; 
  signal nx54672z183_F5MUX : STD_LOGIC; 
  signal nx54672z185 : STD_LOGIC; 
  signal nx54672z183_BXINV : STD_LOGIC; 
  signal nx54672z184 : STD_LOGIC; 
  signal romedatao2_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z193 : STD_LOGIC; 
  signal romedatao2_s_3_BXINV : STD_LOGIC; 
  signal romedatao2_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z192 : STD_LOGIC; 
  signal romedatao2_s_3_BYINV : STD_LOGIC; 
  signal nx54672z189_F5MUX : STD_LOGIC; 
  signal nx54672z190 : STD_LOGIC; 
  signal nx54672z189_BXINV : STD_LOGIC; 
  signal U1_ROME2_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal romodatao2_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z751 : STD_LOGIC; 
  signal romodatao2_s_12_BXINV : STD_LOGIC; 
  signal romodatao2_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z750 : STD_LOGIC; 
  signal romodatao2_s_12_BYINV : STD_LOGIC; 
  signal nx54672z746_F5MUX : STD_LOGIC; 
  signal nx54672z748 : STD_LOGIC; 
  signal nx54672z746_BXINV : STD_LOGIC; 
  signal nx54672z747 : STD_LOGIC; 
  signal romodatao2_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z757 : STD_LOGIC; 
  signal romodatao2_s_11_BXINV : STD_LOGIC; 
  signal romodatao2_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z756 : STD_LOGIC; 
  signal romodatao2_s_11_BYINV : STD_LOGIC; 
  signal nx54672z752_F5MUX : STD_LOGIC; 
  signal nx54672z754 : STD_LOGIC; 
  signal nx54672z752_BXINV : STD_LOGIC; 
  signal nx54672z753 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_FFY_RST : STD_LOGIC; 
  signal romedatao2_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z134 : STD_LOGIC; 
  signal romedatao2_s_13_BXINV : STD_LOGIC; 
  signal romedatao2_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z133 : STD_LOGIC; 
  signal romedatao2_s_13_BYINV : STD_LOGIC; 
  signal nx54672z130_F5MUX : STD_LOGIC; 
  signal nx54672z131 : STD_LOGIC; 
  signal nx54672z130_BXINV : STD_LOGIC; 
  signal nx54672z130_G : STD_LOGIC; 
  signal romedatao1_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z75 : STD_LOGIC; 
  signal romedatao1_s_12_BXINV : STD_LOGIC; 
  signal romedatao1_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z74 : STD_LOGIC; 
  signal romedatao1_s_12_BYINV : STD_LOGIC; 
  signal nx54672z70_F5MUX : STD_LOGIC; 
  signal nx54672z72 : STD_LOGIC; 
  signal nx54672z70_BXINV : STD_LOGIC; 
  signal nx54672z71 : STD_LOGIC; 
  signal romodatao2_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z745 : STD_LOGIC; 
  signal romodatao2_s_13_BXINV : STD_LOGIC; 
  signal romodatao2_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z744 : STD_LOGIC; 
  signal romodatao2_s_13_BYINV : STD_LOGIC; 
  signal nx54672z741_F5MUX : STD_LOGIC; 
  signal nx54672z742 : STD_LOGIC; 
  signal nx54672z741_BXINV : STD_LOGIC; 
  signal nx54672z741_G : STD_LOGIC; 
  signal romodatao2_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z811 : STD_LOGIC; 
  signal romodatao2_s_2_BXINV : STD_LOGIC; 
  signal romodatao2_s_2_F6MUX : STD_LOGIC; 
  signal nx54672z810 : STD_LOGIC; 
  signal romodatao2_s_2_BYINV : STD_LOGIC; 
  signal nx54672z806_F5MUX : STD_LOGIC; 
  signal nx54672z808 : STD_LOGIC; 
  signal nx54672z806_BXINV : STD_LOGIC; 
  signal nx54672z807 : STD_LOGIC; 
  signal romodatao2_s_1_F5MUX : STD_LOGIC; 
  signal nx54672z817 : STD_LOGIC; 
  signal romodatao2_s_1_BXINV : STD_LOGIC; 
  signal romodatao2_s_1_F6MUX : STD_LOGIC; 
  signal nx54672z816 : STD_LOGIC; 
  signal romodatao2_s_1_BYINV : STD_LOGIC; 
  signal nx54672z812_F5MUX : STD_LOGIC; 
  signal nx54672z814 : STD_LOGIC; 
  signal nx54672z812_BXINV : STD_LOGIC; 
  signal nx54672z813 : STD_LOGIC; 
  signal romodatao2_s_0_F5MUX : STD_LOGIC; 
  signal nx54672z819 : STD_LOGIC; 
  signal romodatao2_s_0_BXINV : STD_LOGIC; 
  signal romodatao2_s_0_F6MUX : STD_LOGIC; 
  signal nx54672z818 : STD_LOGIC; 
  signal romodatao2_s_0_BYINV : STD_LOGIC; 
  signal U1_ROMO2_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROMO2_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROMO2_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROMO2_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romodatao1_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z684 : STD_LOGIC; 
  signal romodatao1_s_10_BXINV : STD_LOGIC; 
  signal romodatao1_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z683 : STD_LOGIC; 
  signal romodatao1_s_10_BYINV : STD_LOGIC; 
  signal nx54672z679_F5MUX : STD_LOGIC; 
  signal nx54672z681 : STD_LOGIC; 
  signal nx54672z679_BXINV : STD_LOGIC; 
  signal nx54672z680 : STD_LOGIC; 
  signal romodatao1_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z690 : STD_LOGIC; 
  signal romodatao1_s_9_BXINV : STD_LOGIC; 
  signal romodatao1_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z689 : STD_LOGIC; 
  signal romodatao1_s_9_BYINV : STD_LOGIC; 
  signal nx54672z685_F5MUX : STD_LOGIC; 
  signal nx54672z687 : STD_LOGIC; 
  signal nx54672z685_BXINV : STD_LOGIC; 
  signal nx54672z686 : STD_LOGIC; 
  signal romodatao1_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z696 : STD_LOGIC; 
  signal romodatao1_s_8_BXINV : STD_LOGIC; 
  signal romodatao1_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z695 : STD_LOGIC; 
  signal romodatao1_s_8_BYINV : STD_LOGIC; 
  signal nx54672z691_F5MUX : STD_LOGIC; 
  signal nx54672z693 : STD_LOGIC; 
  signal nx54672z691_BXINV : STD_LOGIC; 
  signal nx54672z692 : STD_LOGIC; 
  signal romodatao1_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z702 : STD_LOGIC; 
  signal romodatao1_s_7_BXINV : STD_LOGIC; 
  signal romodatao1_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z701 : STD_LOGIC; 
  signal romodatao1_s_7_BYINV : STD_LOGIC; 
  signal nx54672z697_F5MUX : STD_LOGIC; 
  signal nx54672z699 : STD_LOGIC; 
  signal nx54672z697_BXINV : STD_LOGIC; 
  signal nx54672z698 : STD_LOGIC; 
  signal romodatao1_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z708 : STD_LOGIC; 
  signal romodatao1_s_6_BXINV : STD_LOGIC; 
  signal romodatao1_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z707 : STD_LOGIC; 
  signal romodatao1_s_6_BYINV : STD_LOGIC; 
  signal nx54672z703_F5MUX : STD_LOGIC; 
  signal nx54672z705 : STD_LOGIC; 
  signal nx54672z703_BXINV : STD_LOGIC; 
  signal nx54672z704 : STD_LOGIC; 
  signal romodatao1_s_0_F5MUX : STD_LOGIC; 
  signal nx54672z740 : STD_LOGIC; 
  signal romodatao1_s_0_BXINV : STD_LOGIC; 
  signal romodatao1_s_0_F6MUX : STD_LOGIC; 
  signal nx54672z739 : STD_LOGIC; 
  signal romodatao1_s_0_BYINV : STD_LOGIC; 
  signal U1_ROMO1_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROMO1_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROMO1_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROMO1_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romedatao4_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z306 : STD_LOGIC; 
  signal romedatao4_s_6_BXINV : STD_LOGIC; 
  signal romedatao4_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z305 : STD_LOGIC; 
  signal romedatao4_s_6_BYINV : STD_LOGIC; 
  signal nx54672z301_F5MUX : STD_LOGIC; 
  signal nx54672z303 : STD_LOGIC; 
  signal nx54672z301_BXINV : STD_LOGIC; 
  signal nx54672z302 : STD_LOGIC; 
  signal romedatao4_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z312 : STD_LOGIC; 
  signal romedatao4_s_5_BXINV : STD_LOGIC; 
  signal romedatao4_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z311 : STD_LOGIC; 
  signal romedatao4_s_5_BYINV : STD_LOGIC; 
  signal nx54672z307_F5MUX : STD_LOGIC; 
  signal nx54672z309 : STD_LOGIC; 
  signal nx54672z307_BXINV : STD_LOGIC; 
  signal nx54672z308 : STD_LOGIC; 
  signal romedatao1_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z69 : STD_LOGIC; 
  signal romedatao1_s_13_BXINV : STD_LOGIC; 
  signal romedatao1_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z68 : STD_LOGIC; 
  signal romedatao1_s_13_BYINV : STD_LOGIC; 
  signal nx54672z65_F5MUX : STD_LOGIC; 
  signal nx54672z66 : STD_LOGIC; 
  signal nx54672z65_BXINV : STD_LOGIC; 
  signal nx54672z65_G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_8_FFX_RST : STD_LOGIC; 
  signal romedatao1_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z81 : STD_LOGIC; 
  signal romedatao1_s_11_BXINV : STD_LOGIC; 
  signal romedatao1_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z80 : STD_LOGIC; 
  signal romedatao1_s_11_BYINV : STD_LOGIC; 
  signal nx54672z76_F5MUX : STD_LOGIC; 
  signal nx54672z78 : STD_LOGIC; 
  signal nx54672z76_BXINV : STD_LOGIC; 
  signal nx54672z77 : STD_LOGIC; 
  signal romedatao1_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z87 : STD_LOGIC; 
  signal romedatao1_s_10_BXINV : STD_LOGIC; 
  signal romedatao1_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z86 : STD_LOGIC; 
  signal romedatao1_s_10_BYINV : STD_LOGIC; 
  signal nx54672z82_F5MUX : STD_LOGIC; 
  signal nx54672z84 : STD_LOGIC; 
  signal nx54672z82_BXINV : STD_LOGIC; 
  signal nx54672z83 : STD_LOGIC; 
  signal romedatao1_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z123 : STD_LOGIC; 
  signal romedatao1_s_4_BXINV : STD_LOGIC; 
  signal romedatao1_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z122 : STD_LOGIC; 
  signal romedatao1_s_4_BYINV : STD_LOGIC; 
  signal nx54672z118_F5MUX : STD_LOGIC; 
  signal nx54672z120 : STD_LOGIC; 
  signal nx54672z118_BXINV : STD_LOGIC; 
  signal nx54672z119 : STD_LOGIC; 
  signal romedatao1_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z128 : STD_LOGIC; 
  signal romedatao1_s_3_BXINV : STD_LOGIC; 
  signal romedatao1_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z127 : STD_LOGIC; 
  signal romedatao1_s_3_BYINV : STD_LOGIC; 
  signal nx54672z124_F5MUX : STD_LOGIC; 
  signal nx54672z125 : STD_LOGIC; 
  signal nx54672z124_BXINV : STD_LOGIC; 
  signal U1_ROME1_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal romedatao1_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z129 : STD_LOGIC; 
  signal romedatao1_s_2_BXINV : STD_LOGIC; 
  signal romedatao1_s_2_F6MUX : STD_LOGIC; 
  signal romedatao1_s_2_G : STD_LOGIC; 
  signal romedatao1_s_2_BYINV : STD_LOGIC; 
  signal U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROME1_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romedatao0_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z11 : STD_LOGIC; 
  signal romedatao0_s_12_BXINV : STD_LOGIC; 
  signal romedatao0_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z10 : STD_LOGIC; 
  signal romedatao0_s_12_BYINV : STD_LOGIC; 
  signal nx54672z6_F5MUX : STD_LOGIC; 
  signal nx54672z8 : STD_LOGIC; 
  signal nx54672z6_BXINV : STD_LOGIC; 
  signal nx54672z7 : STD_LOGIC; 
  signal romedatao0_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z17 : STD_LOGIC; 
  signal romedatao0_s_11_BXINV : STD_LOGIC; 
  signal romedatao0_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z16 : STD_LOGIC; 
  signal romedatao0_s_11_BYINV : STD_LOGIC; 
  signal nx54672z12_F5MUX : STD_LOGIC; 
  signal nx54672z14 : STD_LOGIC; 
  signal nx54672z12_BXINV : STD_LOGIC; 
  signal nx54672z13 : STD_LOGIC; 
  signal romedatao0_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z64 : STD_LOGIC; 
  signal romedatao0_s_3_BXINV : STD_LOGIC; 
  signal romedatao0_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z63 : STD_LOGIC; 
  signal romedatao0_s_3_BYINV : STD_LOGIC; 
  signal nx54672z60_F5MUX : STD_LOGIC; 
  signal nx54672z61 : STD_LOGIC; 
  signal nx54672z60_BXINV : STD_LOGIC; 
  signal U1_ROME0_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal romodatao0_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z625 : STD_LOGIC; 
  signal romodatao0_s_7_BXINV : STD_LOGIC; 
  signal romodatao0_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z624 : STD_LOGIC; 
  signal romodatao0_s_7_BYINV : STD_LOGIC; 
  signal nx54672z620_F5MUX : STD_LOGIC; 
  signal nx54672z622 : STD_LOGIC; 
  signal nx54672z620_BXINV : STD_LOGIC; 
  signal nx54672z621 : STD_LOGIC; 
  signal romodatao0_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z631 : STD_LOGIC; 
  signal romodatao0_s_6_BXINV : STD_LOGIC; 
  signal romodatao0_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z630 : STD_LOGIC; 
  signal romodatao0_s_6_BYINV : STD_LOGIC; 
  signal nx54672z626_F5MUX : STD_LOGIC; 
  signal nx54672z628 : STD_LOGIC; 
  signal nx54672z626_BXINV : STD_LOGIC; 
  signal nx54672z627 : STD_LOGIC; 
  signal romodatao0_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z637 : STD_LOGIC; 
  signal romodatao0_s_5_BXINV : STD_LOGIC; 
  signal romodatao0_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z636 : STD_LOGIC; 
  signal romodatao0_s_5_BYINV : STD_LOGIC; 
  signal nx54672z632_F5MUX : STD_LOGIC; 
  signal nx54672z634 : STD_LOGIC; 
  signal nx54672z632_BXINV : STD_LOGIC; 
  signal nx54672z633 : STD_LOGIC; 
  signal romodatao0_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z643 : STD_LOGIC; 
  signal romodatao0_s_4_BXINV : STD_LOGIC; 
  signal romodatao0_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z642 : STD_LOGIC; 
  signal romodatao0_s_4_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_4_10_FFX_RSTAND : STD_LOGIC; 
  signal nx54672z638_F5MUX : STD_LOGIC; 
  signal nx54672z640 : STD_LOGIC; 
  signal nx54672z638_BXINV : STD_LOGIC; 
  signal nx54672z639 : STD_LOGIC; 
  signal romodatao0_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z649 : STD_LOGIC; 
  signal romodatao0_s_3_BXINV : STD_LOGIC; 
  signal romodatao0_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z648 : STD_LOGIC; 
  signal romodatao0_s_3_BYINV : STD_LOGIC; 
  signal nx54672z644_F5MUX : STD_LOGIC; 
  signal nx54672z646 : STD_LOGIC; 
  signal nx54672z644_BXINV : STD_LOGIC; 
  signal nx54672z645 : STD_LOGIC; 
  signal romedatao0_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z5 : STD_LOGIC; 
  signal romedatao0_s_13_BXINV : STD_LOGIC; 
  signal romedatao0_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z4 : STD_LOGIC; 
  signal romedatao0_s_13_BYINV : STD_LOGIC; 
  signal nx54672z1_F5MUX : STD_LOGIC; 
  signal nx54672z2 : STD_LOGIC; 
  signal nx54672z1_BXINV : STD_LOGIC; 
  signal nx54672z1_G : STD_LOGIC; 
  signal romedatao3_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z205 : STD_LOGIC; 
  signal romedatao3_s_12_BXINV : STD_LOGIC; 
  signal romedatao3_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z204 : STD_LOGIC; 
  signal romedatao3_s_12_BYINV : STD_LOGIC; 
  signal nx54672z200_F5MUX : STD_LOGIC; 
  signal nx54672z202 : STD_LOGIC; 
  signal nx54672z200_BXINV : STD_LOGIC; 
  signal nx54672z201 : STD_LOGIC; 
  signal romedatao3_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z241 : STD_LOGIC; 
  signal romedatao3_s_6_BXINV : STD_LOGIC; 
  signal romedatao3_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z240 : STD_LOGIC; 
  signal romedatao3_s_6_BYINV : STD_LOGIC; 
  signal nx54672z236_F5MUX : STD_LOGIC; 
  signal nx54672z238 : STD_LOGIC; 
  signal nx54672z236_BXINV : STD_LOGIC; 
  signal nx54672z237 : STD_LOGIC; 
  signal romedatao3_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z253 : STD_LOGIC; 
  signal romedatao3_s_4_BXINV : STD_LOGIC; 
  signal romedatao3_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z252 : STD_LOGIC; 
  signal romedatao3_s_4_BYINV : STD_LOGIC; 
  signal nx54672z248_F5MUX : STD_LOGIC; 
  signal nx54672z250 : STD_LOGIC; 
  signal nx54672z248_BXINV : STD_LOGIC; 
  signal nx54672z249 : STD_LOGIC; 
  signal romedatao3_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z259 : STD_LOGIC; 
  signal romedatao3_s_2_BXINV : STD_LOGIC; 
  signal romedatao3_s_2_F6MUX : STD_LOGIC; 
  signal romedatao3_s_2_G : STD_LOGIC; 
  signal romedatao3_s_2_BYINV : STD_LOGIC; 
  signal U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROME3_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romedatao3_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z199 : STD_LOGIC; 
  signal romedatao3_s_13_BXINV : STD_LOGIC; 
  signal romedatao3_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z198 : STD_LOGIC; 
  signal romedatao3_s_13_BYINV : STD_LOGIC; 
  signal nx54672z195_F5MUX : STD_LOGIC; 
  signal nx54672z196 : STD_LOGIC; 
  signal nx54672z195_BXINV : STD_LOGIC; 
  signal nx54672z195_G : STD_LOGIC; 
  signal romedatao5_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z377 : STD_LOGIC; 
  signal romedatao5_s_5_BXINV : STD_LOGIC; 
  signal romedatao5_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z376 : STD_LOGIC; 
  signal romedatao5_s_5_BYINV : STD_LOGIC; 
  signal nx54672z372_F5MUX : STD_LOGIC; 
  signal nx54672z374 : STD_LOGIC; 
  signal nx54672z372_BXINV : STD_LOGIC; 
  signal nx54672z373 : STD_LOGIC; 
  signal romedatao5_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z383 : STD_LOGIC; 
  signal romedatao5_s_4_BXINV : STD_LOGIC; 
  signal romedatao5_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z382 : STD_LOGIC; 
  signal romedatao5_s_4_BYINV : STD_LOGIC; 
  signal nx54672z378_F5MUX : STD_LOGIC; 
  signal nx54672z380 : STD_LOGIC; 
  signal nx54672z378_BXINV : STD_LOGIC; 
  signal nx54672z379 : STD_LOGIC; 
  signal romodatao5_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z1012 : STD_LOGIC; 
  signal romodatao5_s_8_BXINV : STD_LOGIC; 
  signal romodatao5_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z1011 : STD_LOGIC; 
  signal romodatao5_s_8_BYINV : STD_LOGIC; 
  signal nx54672z1007_F5MUX : STD_LOGIC; 
  signal nx54672z1009 : STD_LOGIC; 
  signal nx54672z1007_BXINV : STD_LOGIC; 
  signal nx54672z1008 : STD_LOGIC; 
  signal romedatao5_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z329 : STD_LOGIC; 
  signal romedatao5_s_13_BXINV : STD_LOGIC; 
  signal romedatao5_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z328 : STD_LOGIC; 
  signal romedatao5_s_13_BYINV : STD_LOGIC; 
  signal nx54672z325_F5MUX : STD_LOGIC; 
  signal nx54672z326 : STD_LOGIC; 
  signal nx54672z325_BXINV : STD_LOGIC; 
  signal nx54672z325_G : STD_LOGIC; 
  signal romedatao2_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z140 : STD_LOGIC; 
  signal romedatao2_s_12_BXINV : STD_LOGIC; 
  signal romedatao2_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z139 : STD_LOGIC; 
  signal romedatao2_s_12_BYINV : STD_LOGIC; 
  signal nx54672z135_F5MUX : STD_LOGIC; 
  signal nx54672z137 : STD_LOGIC; 
  signal nx54672z135_BXINV : STD_LOGIC; 
  signal nx54672z136 : STD_LOGIC; 
  signal romedatao2_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z146 : STD_LOGIC; 
  signal romedatao2_s_11_BXINV : STD_LOGIC; 
  signal romedatao2_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z145 : STD_LOGIC; 
  signal romedatao2_s_11_BYINV : STD_LOGIC; 
  signal nx54672z141_F5MUX : STD_LOGIC; 
  signal nx54672z143 : STD_LOGIC; 
  signal nx54672z141_BXINV : STD_LOGIC; 
  signal nx54672z142 : STD_LOGIC; 
  signal romedatao2_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z152 : STD_LOGIC; 
  signal romedatao2_s_10_BXINV : STD_LOGIC; 
  signal romedatao2_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z151 : STD_LOGIC; 
  signal romedatao2_s_10_BYINV : STD_LOGIC; 
  signal nx54672z147_F5MUX : STD_LOGIC; 
  signal nx54672z149 : STD_LOGIC; 
  signal nx54672z147_BXINV : STD_LOGIC; 
  signal nx54672z148 : STD_LOGIC; 
  signal romedatao2_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z158 : STD_LOGIC; 
  signal romedatao2_s_9_BXINV : STD_LOGIC; 
  signal romedatao2_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z157 : STD_LOGIC; 
  signal romedatao2_s_9_BYINV : STD_LOGIC; 
  signal nx54672z153_F5MUX : STD_LOGIC; 
  signal nx54672z155 : STD_LOGIC; 
  signal nx54672z153_BXINV : STD_LOGIC; 
  signal nx54672z154 : STD_LOGIC; 
  signal romedatao2_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z194 : STD_LOGIC; 
  signal romedatao2_s_2_BXINV : STD_LOGIC; 
  signal romedatao2_s_2_F6MUX : STD_LOGIC; 
  signal romedatao2_s_2_G : STD_LOGIC; 
  signal romedatao2_s_2_BYINV : STD_LOGIC; 
  signal U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROME2_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal nx54672z313_F5MUX : STD_LOGIC; 
  signal nx54672z315 : STD_LOGIC; 
  signal nx54672z313_BXINV : STD_LOGIC; 
  signal nx54672z314 : STD_LOGIC; 
  signal romedatao4_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z323 : STD_LOGIC; 
  signal romedatao4_s_3_BXINV : STD_LOGIC; 
  signal romedatao4_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z322 : STD_LOGIC; 
  signal romedatao4_s_3_BYINV : STD_LOGIC; 
  signal nx54672z319_F5MUX : STD_LOGIC; 
  signal nx54672z320 : STD_LOGIC; 
  signal nx54672z319_BXINV : STD_LOGIC; 
  signal U1_ROME4_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal romedatao4_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z324 : STD_LOGIC; 
  signal romedatao4_s_2_BXINV : STD_LOGIC; 
  signal romedatao4_s_2_F6MUX : STD_LOGIC; 
  signal romedatao4_s_2_G : STD_LOGIC; 
  signal romedatao4_s_2_BYINV : STD_LOGIC; 
  signal U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROME4_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romedatao1_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z93 : STD_LOGIC; 
  signal romedatao1_s_9_BXINV : STD_LOGIC; 
  signal romedatao1_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z92 : STD_LOGIC; 
  signal romedatao1_s_9_BYINV : STD_LOGIC; 
  signal nx54672z88_F5MUX : STD_LOGIC; 
  signal nx54672z90 : STD_LOGIC; 
  signal nx54672z88_BXINV : STD_LOGIC; 
  signal nx54672z89 : STD_LOGIC; 
  signal romodatao0_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z655 : STD_LOGIC; 
  signal romodatao0_s_2_BXINV : STD_LOGIC; 
  signal romodatao0_s_2_F6MUX : STD_LOGIC; 
  signal nx54672z654 : STD_LOGIC; 
  signal romodatao0_s_2_BYINV : STD_LOGIC; 
  signal nx54672z650_F5MUX : STD_LOGIC; 
  signal nx54672z652 : STD_LOGIC; 
  signal nx54672z650_BXINV : STD_LOGIC; 
  signal nx54672z651 : STD_LOGIC; 
  signal romedatao6_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z400 : STD_LOGIC; 
  signal romedatao6_s_12_BXINV : STD_LOGIC; 
  signal romedatao6_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z399 : STD_LOGIC; 
  signal romedatao6_s_12_BYINV : STD_LOGIC; 
  signal nx54672z395_F5MUX : STD_LOGIC; 
  signal nx54672z397 : STD_LOGIC; 
  signal nx54672z395_BXINV : STD_LOGIC; 
  signal nx54672z396 : STD_LOGIC; 
  signal romedatao6_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z448 : STD_LOGIC; 
  signal romedatao6_s_4_BXINV : STD_LOGIC; 
  signal romedatao6_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z447 : STD_LOGIC; 
  signal romedatao6_s_4_BYINV : STD_LOGIC; 
  signal nx54672z443_F5MUX : STD_LOGIC; 
  signal nx54672z445 : STD_LOGIC; 
  signal nx54672z443_BXINV : STD_LOGIC; 
  signal nx54672z444 : STD_LOGIC; 
  signal romedatao6_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z453 : STD_LOGIC; 
  signal romedatao6_s_3_BXINV : STD_LOGIC; 
  signal romedatao6_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z452 : STD_LOGIC; 
  signal romedatao6_s_3_BYINV : STD_LOGIC; 
  signal nx54672z449_F5MUX : STD_LOGIC; 
  signal nx54672z450 : STD_LOGIC; 
  signal nx54672z449_BXINV : STD_LOGIC; 
  signal U1_ROME6_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal romedatao6_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z454 : STD_LOGIC; 
  signal romedatao6_s_2_BXINV : STD_LOGIC; 
  signal romedatao6_s_2_F6MUX : STD_LOGIC; 
  signal romedatao6_s_2_G : STD_LOGIC; 
  signal romedatao6_s_2_BYINV : STD_LOGIC; 
  signal U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROME6_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romedatao3_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z217 : STD_LOGIC; 
  signal romedatao3_s_10_BXINV : STD_LOGIC; 
  signal romedatao3_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z216 : STD_LOGIC; 
  signal romedatao3_s_10_BYINV : STD_LOGIC; 
  signal nx54672z212_F5MUX : STD_LOGIC; 
  signal nx54672z214 : STD_LOGIC; 
  signal nx54672z212_BXINV : STD_LOGIC; 
  signal nx54672z213 : STD_LOGIC; 
  signal romedatao3_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z229 : STD_LOGIC; 
  signal romedatao3_s_8_BXINV : STD_LOGIC; 
  signal romedatao3_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z228 : STD_LOGIC; 
  signal romedatao3_s_8_BYINV : STD_LOGIC; 
  signal nx54672z224_F5MUX : STD_LOGIC; 
  signal nx54672z226 : STD_LOGIC; 
  signal nx54672z224_BXINV : STD_LOGIC; 
  signal nx54672z225 : STD_LOGIC; 
  signal romedatao5_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z335 : STD_LOGIC; 
  signal romedatao5_s_12_BXINV : STD_LOGIC; 
  signal romedatao5_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z334 : STD_LOGIC; 
  signal romedatao5_s_12_BYINV : STD_LOGIC; 
  signal nx54672z330_F5MUX : STD_LOGIC; 
  signal nx54672z332 : STD_LOGIC; 
  signal nx54672z330_BXINV : STD_LOGIC; 
  signal nx54672z331 : STD_LOGIC; 
  signal romedatao5_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z341 : STD_LOGIC; 
  signal romedatao5_s_11_BXINV : STD_LOGIC; 
  signal romedatao5_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z340 : STD_LOGIC; 
  signal romedatao5_s_11_BYINV : STD_LOGIC; 
  signal nx54672z336_F5MUX : STD_LOGIC; 
  signal nx54672z338 : STD_LOGIC; 
  signal nx54672z336_BXINV : STD_LOGIC; 
  signal nx54672z337 : STD_LOGIC; 
  signal romedatao5_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z347 : STD_LOGIC; 
  signal romedatao5_s_10_BXINV : STD_LOGIC; 
  signal romedatao5_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z346 : STD_LOGIC; 
  signal romedatao5_s_10_BYINV : STD_LOGIC; 
  signal nx54672z342_F5MUX : STD_LOGIC; 
  signal nx54672z344 : STD_LOGIC; 
  signal nx54672z342_BXINV : STD_LOGIC; 
  signal nx54672z343 : STD_LOGIC; 
  signal romedatao5_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z353 : STD_LOGIC; 
  signal romedatao5_s_9_BXINV : STD_LOGIC; 
  signal romedatao5_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z352 : STD_LOGIC; 
  signal romedatao5_s_9_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_FFY_RST : STD_LOGIC; 
  signal nx54672z348_F5MUX : STD_LOGIC; 
  signal nx54672z350 : STD_LOGIC; 
  signal nx54672z348_BXINV : STD_LOGIC; 
  signal nx54672z349 : STD_LOGIC; 
  signal romedatao5_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z388 : STD_LOGIC; 
  signal romedatao5_s_3_BXINV : STD_LOGIC; 
  signal romedatao5_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z387 : STD_LOGIC; 
  signal romedatao5_s_3_BYINV : STD_LOGIC; 
  signal nx54672z384_F5MUX : STD_LOGIC; 
  signal nx54672z385 : STD_LOGIC; 
  signal nx54672z384_BXINV : STD_LOGIC; 
  signal U1_ROME5_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal romedatao5_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z389 : STD_LOGIC; 
  signal romedatao5_s_2_BXINV : STD_LOGIC; 
  signal romedatao5_s_2_F6MUX : STD_LOGIC; 
  signal romedatao5_s_2_G : STD_LOGIC; 
  signal romedatao5_s_2_BYINV : STD_LOGIC; 
  signal U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROME5_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romodatao6_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z1085 : STD_LOGIC; 
  signal romodatao6_s_9_BXINV : STD_LOGIC; 
  signal romodatao6_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z1084 : STD_LOGIC; 
  signal romodatao6_s_9_BYINV : STD_LOGIC; 
  signal nx54672z1080_F5MUX : STD_LOGIC; 
  signal nx54672z1082 : STD_LOGIC; 
  signal nx54672z1080_BXINV : STD_LOGIC; 
  signal nx54672z1081 : STD_LOGIC; 
  signal romodatao6_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z1091 : STD_LOGIC; 
  signal romodatao6_s_8_BXINV : STD_LOGIC; 
  signal romodatao6_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z1090 : STD_LOGIC; 
  signal romodatao6_s_8_BYINV : STD_LOGIC; 
  signal nx54672z1086_F5MUX : STD_LOGIC; 
  signal nx54672z1088 : STD_LOGIC; 
  signal nx54672z1086_BXINV : STD_LOGIC; 
  signal nx54672z1087 : STD_LOGIC; 
  signal romodatao6_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z1097 : STD_LOGIC; 
  signal romodatao6_s_7_BXINV : STD_LOGIC; 
  signal romodatao6_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z1096 : STD_LOGIC; 
  signal romodatao6_s_7_BYINV : STD_LOGIC; 
  signal nx54672z1092_F5MUX : STD_LOGIC; 
  signal nx54672z1094 : STD_LOGIC; 
  signal nx54672z1092_BXINV : STD_LOGIC; 
  signal nx54672z1093 : STD_LOGIC; 
  signal romodatao5_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z1018 : STD_LOGIC; 
  signal romodatao5_s_7_BXINV : STD_LOGIC; 
  signal romodatao5_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z1017 : STD_LOGIC; 
  signal romodatao5_s_7_BYINV : STD_LOGIC; 
  signal nx54672z1013_F5MUX : STD_LOGIC; 
  signal nx54672z1015 : STD_LOGIC; 
  signal nx54672z1013_BXINV : STD_LOGIC; 
  signal nx54672z1014 : STD_LOGIC; 
  signal romodatao5_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z1024 : STD_LOGIC; 
  signal romodatao5_s_6_BXINV : STD_LOGIC; 
  signal romodatao5_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z1023 : STD_LOGIC; 
  signal romodatao5_s_6_BYINV : STD_LOGIC; 
  signal nx54672z1019_F5MUX : STD_LOGIC; 
  signal nx54672z1021 : STD_LOGIC; 
  signal nx54672z1019_BXINV : STD_LOGIC; 
  signal nx54672z1020 : STD_LOGIC; 
  signal romodatao5_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z1030 : STD_LOGIC; 
  signal romodatao5_s_5_BXINV : STD_LOGIC; 
  signal romodatao5_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z1029 : STD_LOGIC; 
  signal romodatao5_s_5_BYINV : STD_LOGIC; 
  signal nx54672z1025_F5MUX : STD_LOGIC; 
  signal nx54672z1027 : STD_LOGIC; 
  signal nx54672z1025_BXINV : STD_LOGIC; 
  signal nx54672z1026 : STD_LOGIC; 
  signal romodatao5_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z1036 : STD_LOGIC; 
  signal romodatao5_s_4_BXINV : STD_LOGIC; 
  signal romodatao5_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z1035 : STD_LOGIC; 
  signal romodatao5_s_4_BYINV : STD_LOGIC; 
  signal nx54672z1031_F5MUX : STD_LOGIC; 
  signal nx54672z1033 : STD_LOGIC; 
  signal nx54672z1031_BXINV : STD_LOGIC; 
  signal nx54672z1032 : STD_LOGIC; 
  signal romodatao5_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z1042 : STD_LOGIC; 
  signal romodatao5_s_3_BXINV : STD_LOGIC; 
  signal romodatao5_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z1041 : STD_LOGIC; 
  signal romodatao5_s_3_BYINV : STD_LOGIC; 
  signal nx54672z1037_F5MUX : STD_LOGIC; 
  signal nx54672z1039 : STD_LOGIC; 
  signal nx54672z1037_BXINV : STD_LOGIC; 
  signal nx54672z1038 : STD_LOGIC; 
  signal romodatao5_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z982 : STD_LOGIC; 
  signal romodatao5_s_13_BXINV : STD_LOGIC; 
  signal romodatao5_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z981 : STD_LOGIC; 
  signal romodatao5_s_13_BYINV : STD_LOGIC; 
  signal nx54672z978_F5MUX : STD_LOGIC; 
  signal nx54672z979 : STD_LOGIC; 
  signal nx54672z978_BXINV : STD_LOGIC; 
  signal nx54672z978_G : STD_LOGIC; 
  signal romodatao4_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z909 : STD_LOGIC; 
  signal romodatao4_s_12_BXINV : STD_LOGIC; 
  signal romodatao4_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z908 : STD_LOGIC; 
  signal romodatao4_s_12_BYINV : STD_LOGIC; 
  signal nx54672z904_F5MUX : STD_LOGIC; 
  signal nx54672z906 : STD_LOGIC; 
  signal nx54672z904_BXINV : STD_LOGIC; 
  signal nx54672z905 : STD_LOGIC; 
  signal romodatao4_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z921 : STD_LOGIC; 
  signal romodatao4_s_10_BXINV : STD_LOGIC; 
  signal romodatao4_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z920 : STD_LOGIC; 
  signal romodatao4_s_10_BYINV : STD_LOGIC; 
  signal nx54672z916_F5MUX : STD_LOGIC; 
  signal nx54672z918 : STD_LOGIC; 
  signal nx54672z916_BXINV : STD_LOGIC; 
  signal nx54672z917 : STD_LOGIC; 
  signal romodatao4_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z927 : STD_LOGIC; 
  signal romodatao4_s_9_BXINV : STD_LOGIC; 
  signal romodatao4_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z926 : STD_LOGIC; 
  signal romodatao4_s_9_BYINV : STD_LOGIC; 
  signal nx54672z922_F5MUX : STD_LOGIC; 
  signal nx54672z924 : STD_LOGIC; 
  signal nx54672z922_BXINV : STD_LOGIC; 
  signal nx54672z923 : STD_LOGIC; 
  signal romodatao4_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z963 : STD_LOGIC; 
  signal romodatao4_s_3_BXINV : STD_LOGIC; 
  signal romodatao4_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z962 : STD_LOGIC; 
  signal romodatao4_s_3_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_2_FFX_RST : STD_LOGIC; 
  signal nx54672z958_F5MUX : STD_LOGIC; 
  signal nx54672z960 : STD_LOGIC; 
  signal nx54672z958_BXINV : STD_LOGIC; 
  signal nx54672z959 : STD_LOGIC; 
  signal romodatao4_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z969 : STD_LOGIC; 
  signal romodatao4_s_2_BXINV : STD_LOGIC; 
  signal romodatao4_s_2_F6MUX : STD_LOGIC; 
  signal nx54672z968 : STD_LOGIC; 
  signal romodatao4_s_2_BYINV : STD_LOGIC; 
  signal nx54672z964_F5MUX : STD_LOGIC; 
  signal nx54672z966 : STD_LOGIC; 
  signal nx54672z964_BXINV : STD_LOGIC; 
  signal nx54672z965 : STD_LOGIC; 
  signal romodatao4_s_1_F5MUX : STD_LOGIC; 
  signal nx54672z975 : STD_LOGIC; 
  signal romodatao4_s_1_BXINV : STD_LOGIC; 
  signal romodatao4_s_1_F6MUX : STD_LOGIC; 
  signal nx54672z974 : STD_LOGIC; 
  signal romodatao4_s_1_BYINV : STD_LOGIC; 
  signal nx54672z970_F5MUX : STD_LOGIC; 
  signal nx54672z972 : STD_LOGIC; 
  signal nx54672z970_BXINV : STD_LOGIC; 
  signal nx54672z971 : STD_LOGIC; 
  signal romodatao4_s_0_F5MUX : STD_LOGIC; 
  signal nx54672z977 : STD_LOGIC; 
  signal romodatao4_s_0_BXINV : STD_LOGIC; 
  signal romodatao4_s_0_F6MUX : STD_LOGIC; 
  signal nx54672z976 : STD_LOGIC; 
  signal romodatao4_s_0_BYINV : STD_LOGIC; 
  signal U1_ROMO4_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROMO4_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROMO4_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROMO4_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romodatao3_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z854 : STD_LOGIC; 
  signal romodatao3_s_8_BXINV : STD_LOGIC; 
  signal romodatao3_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z853 : STD_LOGIC; 
  signal romodatao3_s_8_BYINV : STD_LOGIC; 
  signal nx54672z849_F5MUX : STD_LOGIC; 
  signal nx54672z851 : STD_LOGIC; 
  signal nx54672z849_BXINV : STD_LOGIC; 
  signal nx54672z850 : STD_LOGIC; 
  signal romodatao3_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z866 : STD_LOGIC; 
  signal romodatao3_s_6_BXINV : STD_LOGIC; 
  signal romodatao3_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z865 : STD_LOGIC; 
  signal romodatao3_s_6_BYINV : STD_LOGIC; 
  signal nx54672z861_F5MUX : STD_LOGIC; 
  signal nx54672z863 : STD_LOGIC; 
  signal nx54672z861_BXINV : STD_LOGIC; 
  signal nx54672z862 : STD_LOGIC; 
  signal romodatao2_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z793 : STD_LOGIC; 
  signal romodatao2_s_5_BXINV : STD_LOGIC; 
  signal romodatao2_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z792 : STD_LOGIC; 
  signal romodatao2_s_5_BYINV : STD_LOGIC; 
  signal nx54672z788_F5MUX : STD_LOGIC; 
  signal nx54672z790 : STD_LOGIC; 
  signal nx54672z788_BXINV : STD_LOGIC; 
  signal nx54672z789 : STD_LOGIC; 
  signal romodatao2_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z799 : STD_LOGIC; 
  signal romodatao2_s_4_BXINV : STD_LOGIC; 
  signal romodatao2_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z798 : STD_LOGIC; 
  signal romodatao2_s_4_BYINV : STD_LOGIC; 
  signal nx54672z794_F5MUX : STD_LOGIC; 
  signal nx54672z796 : STD_LOGIC; 
  signal nx54672z794_BXINV : STD_LOGIC; 
  signal nx54672z795 : STD_LOGIC; 
  signal romedatao7_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z465 : STD_LOGIC; 
  signal romedatao7_s_12_BXINV : STD_LOGIC; 
  signal romedatao7_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z464 : STD_LOGIC; 
  signal romedatao7_s_12_BYINV : STD_LOGIC; 
  signal nx54672z460_F5MUX : STD_LOGIC; 
  signal nx54672z462 : STD_LOGIC; 
  signal nx54672z460_BXINV : STD_LOGIC; 
  signal nx54672z461 : STD_LOGIC; 
  signal romedatao7_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z471 : STD_LOGIC; 
  signal romedatao7_s_11_BXINV : STD_LOGIC; 
  signal romedatao7_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z470 : STD_LOGIC; 
  signal romedatao7_s_11_BYINV : STD_LOGIC; 
  signal nx54672z466_F5MUX : STD_LOGIC; 
  signal nx54672z468 : STD_LOGIC; 
  signal nx54672z466_BXINV : STD_LOGIC; 
  signal nx54672z467 : STD_LOGIC; 
  signal romedatao7_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z518 : STD_LOGIC; 
  signal romedatao7_s_3_BXINV : STD_LOGIC; 
  signal romedatao7_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z517 : STD_LOGIC; 
  signal romedatao7_s_3_BYINV : STD_LOGIC; 
  signal nx54672z514_F5MUX : STD_LOGIC; 
  signal nx54672z515 : STD_LOGIC; 
  signal nx54672z514_BXINV : STD_LOGIC; 
  signal U1_ROME7_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal romedatao7_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z519 : STD_LOGIC; 
  signal romedatao7_s_2_BXINV : STD_LOGIC; 
  signal romedatao7_s_2_F6MUX : STD_LOGIC; 
  signal romedatao7_s_2_G : STD_LOGIC; 
  signal romedatao7_s_2_BYINV : STD_LOGIC; 
  signal U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROME7_modgen_rom_ix2_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_G : STD_LOGIC; 
  signal romodatao7_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z1152 : STD_LOGIC; 
  signal romodatao7_s_11_BXINV : STD_LOGIC; 
  signal romodatao7_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z1151 : STD_LOGIC; 
  signal romodatao7_s_11_BYINV : STD_LOGIC; 
  signal nx54672z1147_F5MUX : STD_LOGIC; 
  signal nx54672z1149 : STD_LOGIC; 
  signal nx54672z1147_BXINV : STD_LOGIC; 
  signal nx54672z1148 : STD_LOGIC; 
  signal romodatao7_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z1158 : STD_LOGIC; 
  signal romodatao7_s_10_BXINV : STD_LOGIC; 
  signal romodatao7_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z1157 : STD_LOGIC; 
  signal romodatao7_s_10_BYINV : STD_LOGIC; 
  signal nx54672z1153_F5MUX : STD_LOGIC; 
  signal nx54672z1155 : STD_LOGIC; 
  signal nx54672z1153_BXINV : STD_LOGIC; 
  signal nx54672z1154 : STD_LOGIC; 
  signal romodatao3_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z836 : STD_LOGIC; 
  signal romodatao3_s_11_BXINV : STD_LOGIC; 
  signal romodatao3_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z835 : STD_LOGIC; 
  signal romodatao3_s_11_BYINV : STD_LOGIC; 
  signal nx54672z831_F5MUX : STD_LOGIC; 
  signal nx54672z833 : STD_LOGIC; 
  signal nx54672z831_BXINV : STD_LOGIC; 
  signal nx54672z832 : STD_LOGIC; 
  signal romodatao2_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z805 : STD_LOGIC; 
  signal romodatao2_s_3_BXINV : STD_LOGIC; 
  signal romodatao2_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z804 : STD_LOGIC; 
  signal romodatao2_s_3_BYINV : STD_LOGIC; 
  signal nx54672z800_F5MUX : STD_LOGIC; 
  signal nx54672z802 : STD_LOGIC; 
  signal nx54672z800_BXINV : STD_LOGIC; 
  signal nx54672z801 : STD_LOGIC; 
  signal romedatao4_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z288 : STD_LOGIC; 
  signal romedatao4_s_9_BXINV : STD_LOGIC; 
  signal romedatao4_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z287 : STD_LOGIC; 
  signal romedatao4_s_9_BYINV : STD_LOGIC; 
  signal nx54672z283_F5MUX : STD_LOGIC; 
  signal nx54672z285 : STD_LOGIC; 
  signal nx54672z283_BXINV : STD_LOGIC; 
  signal nx54672z284 : STD_LOGIC; 
  signal romedatao4_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z294 : STD_LOGIC; 
  signal romedatao4_s_8_BXINV : STD_LOGIC; 
  signal romedatao4_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z293 : STD_LOGIC; 
  signal romedatao4_s_8_BYINV : STD_LOGIC; 
  signal nx54672z289_F5MUX : STD_LOGIC; 
  signal nx54672z291 : STD_LOGIC; 
  signal nx54672z289_BXINV : STD_LOGIC; 
  signal nx54672z290 : STD_LOGIC; 
  signal romedatao4_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z300 : STD_LOGIC; 
  signal romedatao4_s_7_BXINV : STD_LOGIC; 
  signal romedatao4_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z299 : STD_LOGIC; 
  signal romedatao4_s_7_BYINV : STD_LOGIC; 
  signal nx54672z295_F5MUX : STD_LOGIC; 
  signal nx54672z297 : STD_LOGIC; 
  signal nx54672z295_BXINV : STD_LOGIC; 
  signal nx54672z296 : STD_LOGIC; 
  signal romedatao3_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z211 : STD_LOGIC; 
  signal romedatao3_s_11_BXINV : STD_LOGIC; 
  signal romedatao3_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z210 : STD_LOGIC; 
  signal romedatao3_s_11_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_FFY_RST : STD_LOGIC; 
  signal nx54672z206_F5MUX : STD_LOGIC; 
  signal nx54672z208 : STD_LOGIC; 
  signal nx54672z206_BXINV : STD_LOGIC; 
  signal nx54672z207 : STD_LOGIC; 
  signal romedatao3_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z235 : STD_LOGIC; 
  signal romedatao3_s_7_BXINV : STD_LOGIC; 
  signal romedatao3_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z234 : STD_LOGIC; 
  signal romedatao3_s_7_BYINV : STD_LOGIC; 
  signal nx54672z230_F5MUX : STD_LOGIC; 
  signal nx54672z232 : STD_LOGIC; 
  signal nx54672z230_BXINV : STD_LOGIC; 
  signal nx54672z231 : STD_LOGIC; 
  signal romedatao7_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z459 : STD_LOGIC; 
  signal romedatao7_s_13_BXINV : STD_LOGIC; 
  signal romedatao7_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z458 : STD_LOGIC; 
  signal romedatao7_s_13_BYINV : STD_LOGIC; 
  signal nx54672z455_F5MUX : STD_LOGIC; 
  signal nx54672z456 : STD_LOGIC; 
  signal nx54672z455_BXINV : STD_LOGIC; 
  signal nx54672z455_G : STD_LOGIC; 
  signal romedatao6_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z406 : STD_LOGIC; 
  signal romedatao6_s_11_BXINV : STD_LOGIC; 
  signal romedatao6_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z405 : STD_LOGIC; 
  signal romedatao6_s_11_BYINV : STD_LOGIC; 
  signal nx54672z401_F5MUX : STD_LOGIC; 
  signal nx54672z403 : STD_LOGIC; 
  signal nx54672z401_BXINV : STD_LOGIC; 
  signal nx54672z402 : STD_LOGIC; 
  signal romedatao6_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z412 : STD_LOGIC; 
  signal romedatao6_s_10_BXINV : STD_LOGIC; 
  signal romedatao6_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z411 : STD_LOGIC; 
  signal romedatao6_s_10_BYINV : STD_LOGIC; 
  signal nx54672z407_F5MUX : STD_LOGIC; 
  signal nx54672z409 : STD_LOGIC; 
  signal nx54672z407_BXINV : STD_LOGIC; 
  signal nx54672z408 : STD_LOGIC; 
  signal romedatao6_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z418 : STD_LOGIC; 
  signal romedatao6_s_9_BXINV : STD_LOGIC; 
  signal romedatao6_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z417 : STD_LOGIC; 
  signal romedatao6_s_9_BYINV : STD_LOGIC; 
  signal nx54672z413_F5MUX : STD_LOGIC; 
  signal nx54672z415 : STD_LOGIC; 
  signal nx54672z413_BXINV : STD_LOGIC; 
  signal nx54672z414 : STD_LOGIC; 
  signal romedatao6_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z424 : STD_LOGIC; 
  signal romedatao6_s_8_BXINV : STD_LOGIC; 
  signal romedatao6_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z423 : STD_LOGIC; 
  signal romedatao6_s_8_BYINV : STD_LOGIC; 
  signal nx54672z419_F5MUX : STD_LOGIC; 
  signal nx54672z421 : STD_LOGIC; 
  signal nx54672z419_BXINV : STD_LOGIC; 
  signal nx54672z420 : STD_LOGIC; 
  signal romedatao6_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z430 : STD_LOGIC; 
  signal romedatao6_s_7_BXINV : STD_LOGIC; 
  signal romedatao6_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z429 : STD_LOGIC; 
  signal romedatao6_s_7_BYINV : STD_LOGIC; 
  signal nx54672z425_F5MUX : STD_LOGIC; 
  signal nx54672z427 : STD_LOGIC; 
  signal nx54672z425_BXINV : STD_LOGIC; 
  signal nx54672z426 : STD_LOGIC; 
  signal romedatao8_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z530 : STD_LOGIC; 
  signal romedatao8_s_12_BXINV : STD_LOGIC; 
  signal romedatao8_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z529 : STD_LOGIC; 
  signal romedatao8_s_12_BYINV : STD_LOGIC; 
  signal nx54672z525_F5MUX : STD_LOGIC; 
  signal nx54672z527 : STD_LOGIC; 
  signal nx54672z525_BXINV : STD_LOGIC; 
  signal nx54672z526 : STD_LOGIC; 
  signal romedatao8_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z536 : STD_LOGIC; 
  signal romedatao8_s_11_BXINV : STD_LOGIC; 
  signal romedatao8_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z535 : STD_LOGIC; 
  signal romedatao8_s_11_BYINV : STD_LOGIC; 
  signal nx54672z531_F5MUX : STD_LOGIC; 
  signal nx54672z533 : STD_LOGIC; 
  signal nx54672z531_BXINV : STD_LOGIC; 
  signal nx54672z532 : STD_LOGIC; 
  signal romedatao8_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z542 : STD_LOGIC; 
  signal romedatao8_s_10_BXINV : STD_LOGIC; 
  signal romedatao8_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z541 : STD_LOGIC; 
  signal romedatao8_s_10_BYINV : STD_LOGIC; 
  signal nx54672z537_F5MUX : STD_LOGIC; 
  signal nx54672z539 : STD_LOGIC; 
  signal nx54672z537_BXINV : STD_LOGIC; 
  signal nx54672z538 : STD_LOGIC; 
  signal romedatao8_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z548 : STD_LOGIC; 
  signal romedatao8_s_9_BXINV : STD_LOGIC; 
  signal romedatao8_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z547 : STD_LOGIC; 
  signal romedatao8_s_9_BYINV : STD_LOGIC; 
  signal nx54672z543_F5MUX : STD_LOGIC; 
  signal nx54672z545 : STD_LOGIC; 
  signal nx54672z543_BXINV : STD_LOGIC; 
  signal nx54672z544 : STD_LOGIC; 
  signal romedatao4_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z264 : STD_LOGIC; 
  signal romedatao4_s_13_BXINV : STD_LOGIC; 
  signal romedatao4_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z263 : STD_LOGIC; 
  signal romedatao4_s_13_BYINV : STD_LOGIC; 
  signal nx54672z260_F5MUX : STD_LOGIC; 
  signal nx54672z261 : STD_LOGIC; 
  signal nx54672z260_BXINV : STD_LOGIC; 
  signal nx54672z260_G : STD_LOGIC; 
  signal romedatao8_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z524 : STD_LOGIC; 
  signal romedatao8_s_13_BXINV : STD_LOGIC; 
  signal romedatao8_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z523 : STD_LOGIC; 
  signal romedatao8_s_13_BYINV : STD_LOGIC; 
  signal nx54672z520_F5MUX : STD_LOGIC; 
  signal nx54672z521 : STD_LOGIC; 
  signal nx54672z520_BXINV : STD_LOGIC; 
  signal nx54672z520_G : STD_LOGIC; 
  signal romedatao5_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z359 : STD_LOGIC; 
  signal romedatao5_s_8_BXINV : STD_LOGIC; 
  signal romedatao5_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z358 : STD_LOGIC; 
  signal romedatao5_s_8_BYINV : STD_LOGIC; 
  signal nx54672z354_F5MUX : STD_LOGIC; 
  signal nx54672z356 : STD_LOGIC; 
  signal nx54672z354_BXINV : STD_LOGIC; 
  signal nx54672z355 : STD_LOGIC; 
  signal romedatao5_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z365 : STD_LOGIC; 
  signal romedatao5_s_7_BXINV : STD_LOGIC; 
  signal romedatao5_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z364 : STD_LOGIC; 
  signal romedatao5_s_7_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_4_FFX_RST : STD_LOGIC; 
  signal nx54672z360_F5MUX : STD_LOGIC; 
  signal nx54672z362 : STD_LOGIC; 
  signal nx54672z360_BXINV : STD_LOGIC; 
  signal nx54672z361 : STD_LOGIC; 
  signal romedatao5_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z371 : STD_LOGIC; 
  signal romedatao5_s_6_BXINV : STD_LOGIC; 
  signal romedatao5_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z370 : STD_LOGIC; 
  signal romedatao5_s_6_BYINV : STD_LOGIC; 
  signal nx54672z366_F5MUX : STD_LOGIC; 
  signal nx54672z368 : STD_LOGIC; 
  signal nx54672z366_BXINV : STD_LOGIC; 
  signal nx54672z367 : STD_LOGIC; 
  signal romodatao6_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z1067 : STD_LOGIC; 
  signal romodatao6_s_12_BXINV : STD_LOGIC; 
  signal romodatao6_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z1066 : STD_LOGIC; 
  signal romodatao6_s_12_BYINV : STD_LOGIC; 
  signal nx54672z1062_F5MUX : STD_LOGIC; 
  signal nx54672z1064 : STD_LOGIC; 
  signal nx54672z1062_BXINV : STD_LOGIC; 
  signal nx54672z1063 : STD_LOGIC; 
  signal romodatao6_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z1103 : STD_LOGIC; 
  signal romodatao6_s_6_BXINV : STD_LOGIC; 
  signal romodatao6_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z1102 : STD_LOGIC; 
  signal romodatao6_s_6_BYINV : STD_LOGIC; 
  signal nx54672z1098_F5MUX : STD_LOGIC; 
  signal nx54672z1100 : STD_LOGIC; 
  signal nx54672z1098_BXINV : STD_LOGIC; 
  signal nx54672z1099 : STD_LOGIC; 
  signal romodatao6_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z1109 : STD_LOGIC; 
  signal romodatao6_s_5_BXINV : STD_LOGIC; 
  signal romodatao6_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z1108 : STD_LOGIC; 
  signal romodatao6_s_5_BYINV : STD_LOGIC; 
  signal nx54672z1104_F5MUX : STD_LOGIC; 
  signal nx54672z1106 : STD_LOGIC; 
  signal nx54672z1104_BXINV : STD_LOGIC; 
  signal nx54672z1105 : STD_LOGIC; 
  signal romodatao6_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z1115 : STD_LOGIC; 
  signal romodatao6_s_4_BXINV : STD_LOGIC; 
  signal romodatao6_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z1114 : STD_LOGIC; 
  signal romodatao6_s_4_BYINV : STD_LOGIC; 
  signal nx54672z1110_F5MUX : STD_LOGIC; 
  signal nx54672z1112 : STD_LOGIC; 
  signal nx54672z1110_BXINV : STD_LOGIC; 
  signal nx54672z1111 : STD_LOGIC; 
  signal romodatao6_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z1121 : STD_LOGIC; 
  signal romodatao6_s_3_BXINV : STD_LOGIC; 
  signal romodatao6_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z1120 : STD_LOGIC; 
  signal romodatao6_s_3_BYINV : STD_LOGIC; 
  signal nx54672z1116_F5MUX : STD_LOGIC; 
  signal nx54672z1118 : STD_LOGIC; 
  signal nx54672z1116_BXINV : STD_LOGIC; 
  signal nx54672z1117 : STD_LOGIC; 
  signal romodatao6_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z1127 : STD_LOGIC; 
  signal romodatao6_s_2_BXINV : STD_LOGIC; 
  signal romodatao6_s_2_F6MUX : STD_LOGIC; 
  signal nx54672z1126 : STD_LOGIC; 
  signal romodatao6_s_2_BYINV : STD_LOGIC; 
  signal nx54672z1122_F5MUX : STD_LOGIC; 
  signal nx54672z1124 : STD_LOGIC; 
  signal nx54672z1122_BXINV : STD_LOGIC; 
  signal nx54672z1123 : STD_LOGIC; 
  signal romodatao5_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z988 : STD_LOGIC; 
  signal romodatao5_s_12_BXINV : STD_LOGIC; 
  signal romodatao5_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z987 : STD_LOGIC; 
  signal romodatao5_s_12_BYINV : STD_LOGIC; 
  signal nx54672z983_F5MUX : STD_LOGIC; 
  signal nx54672z985 : STD_LOGIC; 
  signal nx54672z983_BXINV : STD_LOGIC; 
  signal nx54672z984 : STD_LOGIC; 
  signal romodatao5_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z994 : STD_LOGIC; 
  signal romodatao5_s_11_BXINV : STD_LOGIC; 
  signal romodatao5_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z993 : STD_LOGIC; 
  signal romodatao5_s_11_BYINV : STD_LOGIC; 
  signal nx54672z989_F5MUX : STD_LOGIC; 
  signal nx54672z991 : STD_LOGIC; 
  signal nx54672z989_BXINV : STD_LOGIC; 
  signal nx54672z990 : STD_LOGIC; 
  signal romodatao5_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z1000 : STD_LOGIC; 
  signal romodatao5_s_10_BXINV : STD_LOGIC; 
  signal romodatao5_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z999 : STD_LOGIC; 
  signal romodatao5_s_10_BYINV : STD_LOGIC; 
  signal nx54672z995_F5MUX : STD_LOGIC; 
  signal nx54672z997 : STD_LOGIC; 
  signal nx54672z995_BXINV : STD_LOGIC; 
  signal nx54672z996 : STD_LOGIC; 
  signal romodatao5_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z1006 : STD_LOGIC; 
  signal romodatao5_s_9_BXINV : STD_LOGIC; 
  signal romodatao5_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z1005 : STD_LOGIC; 
  signal romodatao5_s_9_BYINV : STD_LOGIC; 
  signal nx54672z1001_F5MUX : STD_LOGIC; 
  signal nx54672z1003 : STD_LOGIC; 
  signal nx54672z1001_BXINV : STD_LOGIC; 
  signal nx54672z1002 : STD_LOGIC; 
  signal romodatao5_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z1048 : STD_LOGIC; 
  signal romodatao5_s_2_BXINV : STD_LOGIC; 
  signal romodatao5_s_2_F6MUX : STD_LOGIC; 
  signal nx54672z1047 : STD_LOGIC; 
  signal romodatao5_s_2_BYINV : STD_LOGIC; 
  signal nx54672z1043_F5MUX : STD_LOGIC; 
  signal nx54672z1045 : STD_LOGIC; 
  signal nx54672z1043_BXINV : STD_LOGIC; 
  signal nx54672z1044 : STD_LOGIC; 
  signal romodatao5_s_1_F5MUX : STD_LOGIC; 
  signal nx54672z1054 : STD_LOGIC; 
  signal romodatao5_s_1_BXINV : STD_LOGIC; 
  signal romodatao5_s_1_F6MUX : STD_LOGIC; 
  signal nx54672z1053 : STD_LOGIC; 
  signal romodatao5_s_1_BYINV : STD_LOGIC; 
  signal nx54672z1049_F5MUX : STD_LOGIC; 
  signal nx54672z1051 : STD_LOGIC; 
  signal nx54672z1049_BXINV : STD_LOGIC; 
  signal nx54672z1050 : STD_LOGIC; 
  signal romodatao8_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z1225 : STD_LOGIC; 
  signal romodatao8_s_12_BXINV : STD_LOGIC; 
  signal romodatao8_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z1224 : STD_LOGIC; 
  signal romodatao8_s_12_BYINV : STD_LOGIC; 
  signal nx54672z1220_F5MUX : STD_LOGIC; 
  signal nx54672z1222 : STD_LOGIC; 
  signal nx54672z1220_BXINV : STD_LOGIC; 
  signal nx54672z1221 : STD_LOGIC; 
  signal romodatao8_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z1231 : STD_LOGIC; 
  signal romodatao8_s_11_BXINV : STD_LOGIC; 
  signal romodatao8_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z1230 : STD_LOGIC; 
  signal romodatao8_s_11_BYINV : STD_LOGIC; 
  signal nx54672z1226_F5MUX : STD_LOGIC; 
  signal nx54672z1228 : STD_LOGIC; 
  signal nx54672z1226_BXINV : STD_LOGIC; 
  signal nx54672z1227 : STD_LOGIC; 
  signal romodatao6_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z1061 : STD_LOGIC; 
  signal romodatao6_s_13_BXINV : STD_LOGIC; 
  signal romodatao6_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z1060 : STD_LOGIC; 
  signal romodatao6_s_13_BYINV : STD_LOGIC; 
  signal nx54672z1057_F5MUX : STD_LOGIC; 
  signal nx54672z1058 : STD_LOGIC; 
  signal nx54672z1057_BXINV : STD_LOGIC; 
  signal nx54672z1057_G : STD_LOGIC; 
  signal romodatao5_s_0_F5MUX : STD_LOGIC; 
  signal nx54672z1056 : STD_LOGIC; 
  signal romodatao5_s_0_BXINV : STD_LOGIC; 
  signal romodatao5_s_0_F6MUX : STD_LOGIC; 
  signal nx54672z1055 : STD_LOGIC; 
  signal romodatao5_s_0_BYINV : STD_LOGIC; 
  signal U1_ROMO5_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROMO5_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROMO5_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROMO5_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romodatao4_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z933 : STD_LOGIC; 
  signal romodatao4_s_8_BXINV : STD_LOGIC; 
  signal romodatao4_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z932 : STD_LOGIC; 
  signal romodatao4_s_8_BYINV : STD_LOGIC; 
  signal nx54672z928_F5MUX : STD_LOGIC; 
  signal nx54672z930 : STD_LOGIC; 
  signal nx54672z928_BXINV : STD_LOGIC; 
  signal nx54672z929 : STD_LOGIC; 
  signal romodatao4_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z939 : STD_LOGIC; 
  signal romodatao4_s_7_BXINV : STD_LOGIC; 
  signal romodatao4_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z938 : STD_LOGIC; 
  signal romodatao4_s_7_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_FFY_RST : STD_LOGIC; 
  signal nx54672z934_F5MUX : STD_LOGIC; 
  signal nx54672z936 : STD_LOGIC; 
  signal nx54672z934_BXINV : STD_LOGIC; 
  signal nx54672z935 : STD_LOGIC; 
  signal romedatao7_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z477 : STD_LOGIC; 
  signal romedatao7_s_10_BXINV : STD_LOGIC; 
  signal romedatao7_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z476 : STD_LOGIC; 
  signal romedatao7_s_10_BYINV : STD_LOGIC; 
  signal nx54672z472_F5MUX : STD_LOGIC; 
  signal nx54672z474 : STD_LOGIC; 
  signal nx54672z472_BXINV : STD_LOGIC; 
  signal nx54672z473 : STD_LOGIC; 
  signal romedatao7_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z483 : STD_LOGIC; 
  signal romedatao7_s_9_BXINV : STD_LOGIC; 
  signal romedatao7_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z482 : STD_LOGIC; 
  signal romedatao7_s_9_BYINV : STD_LOGIC; 
  signal nx54672z478_F5MUX : STD_LOGIC; 
  signal nx54672z480 : STD_LOGIC; 
  signal nx54672z478_BXINV : STD_LOGIC; 
  signal nx54672z479 : STD_LOGIC; 
  signal romedatao7_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z489 : STD_LOGIC; 
  signal romedatao7_s_8_BXINV : STD_LOGIC; 
  signal romedatao7_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z488 : STD_LOGIC; 
  signal romedatao7_s_8_BYINV : STD_LOGIC; 
  signal nx54672z484_F5MUX : STD_LOGIC; 
  signal nx54672z486 : STD_LOGIC; 
  signal nx54672z484_BXINV : STD_LOGIC; 
  signal nx54672z485 : STD_LOGIC; 
  signal romedatao7_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z495 : STD_LOGIC; 
  signal romedatao7_s_7_BXINV : STD_LOGIC; 
  signal romedatao7_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z494 : STD_LOGIC; 
  signal romedatao7_s_7_BYINV : STD_LOGIC; 
  signal nx54672z490_F5MUX : STD_LOGIC; 
  signal nx54672z492 : STD_LOGIC; 
  signal nx54672z490_BXINV : STD_LOGIC; 
  signal nx54672z491 : STD_LOGIC; 
  signal romedatao7_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z501 : STD_LOGIC; 
  signal romedatao7_s_6_BXINV : STD_LOGIC; 
  signal romedatao7_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z500 : STD_LOGIC; 
  signal romedatao7_s_6_BYINV : STD_LOGIC; 
  signal nx54672z496_F5MUX : STD_LOGIC; 
  signal nx54672z498 : STD_LOGIC; 
  signal nx54672z496_BXINV : STD_LOGIC; 
  signal nx54672z497 : STD_LOGIC; 
  signal romodatao8_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z1237 : STD_LOGIC; 
  signal romodatao8_s_10_BXINV : STD_LOGIC; 
  signal romodatao8_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z1236 : STD_LOGIC; 
  signal romodatao8_s_10_BYINV : STD_LOGIC; 
  signal nx54672z1232_F5MUX : STD_LOGIC; 
  signal nx54672z1234 : STD_LOGIC; 
  signal nx54672z1232_BXINV : STD_LOGIC; 
  signal nx54672z1233 : STD_LOGIC; 
  signal romodatao8_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z1243 : STD_LOGIC; 
  signal romodatao8_s_9_BXINV : STD_LOGIC; 
  signal romodatao8_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z1242 : STD_LOGIC; 
  signal romodatao8_s_9_BYINV : STD_LOGIC; 
  signal nx54672z1238_F5MUX : STD_LOGIC; 
  signal nx54672z1240 : STD_LOGIC; 
  signal nx54672z1238_BXINV : STD_LOGIC; 
  signal nx54672z1239 : STD_LOGIC; 
  signal romodatao7_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z1164 : STD_LOGIC; 
  signal romodatao7_s_9_BXINV : STD_LOGIC; 
  signal romodatao7_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z1163 : STD_LOGIC; 
  signal romodatao7_s_9_BYINV : STD_LOGIC; 
  signal ramdatai_s_0_FFX_RST : STD_LOGIC; 
  signal ramdatai_s_2_FFY_RST : STD_LOGIC; 
  signal ramdatai_s_2_FFX_RST : STD_LOGIC; 
  signal nx54672z1159_F5MUX : STD_LOGIC; 
  signal nx54672z1161 : STD_LOGIC; 
  signal nx54672z1159_BXINV : STD_LOGIC; 
  signal nx54672z1160 : STD_LOGIC; 
  signal romodatao7_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z1170 : STD_LOGIC; 
  signal romodatao7_s_8_BXINV : STD_LOGIC; 
  signal romodatao7_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z1169 : STD_LOGIC; 
  signal romodatao7_s_8_BYINV : STD_LOGIC; 
  signal nx54672z1165_F5MUX : STD_LOGIC; 
  signal nx54672z1167 : STD_LOGIC; 
  signal nx54672z1165_BXINV : STD_LOGIC; 
  signal nx54672z1166 : STD_LOGIC; 
  signal romodatao7_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z1176 : STD_LOGIC; 
  signal romodatao7_s_7_BXINV : STD_LOGIC; 
  signal romodatao7_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z1175 : STD_LOGIC; 
  signal romodatao7_s_7_BYINV : STD_LOGIC; 
  signal nx54672z1171_F5MUX : STD_LOGIC; 
  signal nx54672z1173 : STD_LOGIC; 
  signal nx54672z1171_BXINV : STD_LOGIC; 
  signal nx54672z1172 : STD_LOGIC; 
  signal romodatao7_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z1182 : STD_LOGIC; 
  signal romodatao7_s_6_BXINV : STD_LOGIC; 
  signal romodatao7_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z1181 : STD_LOGIC; 
  signal romodatao7_s_6_BYINV : STD_LOGIC; 
  signal nx54672z1177_F5MUX : STD_LOGIC; 
  signal nx54672z1179 : STD_LOGIC; 
  signal nx54672z1177_BXINV : STD_LOGIC; 
  signal nx54672z1178 : STD_LOGIC; 
  signal romodatao7_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z1188 : STD_LOGIC; 
  signal romodatao7_s_5_BXINV : STD_LOGIC; 
  signal romodatao7_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z1187 : STD_LOGIC; 
  signal romodatao7_s_5_BYINV : STD_LOGIC; 
  signal nx54672z1183_F5MUX : STD_LOGIC; 
  signal nx54672z1185 : STD_LOGIC; 
  signal nx54672z1183_BXINV : STD_LOGIC; 
  signal nx54672z1184 : STD_LOGIC; 
  signal romodatao3_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z848 : STD_LOGIC; 
  signal romodatao3_s_9_BXINV : STD_LOGIC; 
  signal romodatao3_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z847 : STD_LOGIC; 
  signal romodatao3_s_9_BYINV : STD_LOGIC; 
  signal nx54672z843_F5MUX : STD_LOGIC; 
  signal nx54672z845 : STD_LOGIC; 
  signal nx54672z843_BXINV : STD_LOGIC; 
  signal nx54672z844 : STD_LOGIC; 
  signal romodatao3_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z872 : STD_LOGIC; 
  signal romodatao3_s_5_BXINV : STD_LOGIC; 
  signal romodatao3_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z871 : STD_LOGIC; 
  signal romodatao3_s_5_BYINV : STD_LOGIC; 
  signal nx54672z867_F5MUX : STD_LOGIC; 
  signal nx54672z869 : STD_LOGIC; 
  signal nx54672z867_BXINV : STD_LOGIC; 
  signal nx54672z868 : STD_LOGIC; 
  signal romedatao3_s_9_F5MUX : STD_LOGIC; 
  signal nx54672z223 : STD_LOGIC; 
  signal romedatao3_s_9_BXINV : STD_LOGIC; 
  signal romedatao3_s_9_F6MUX : STD_LOGIC; 
  signal nx54672z222 : STD_LOGIC; 
  signal romedatao3_s_9_BYINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_6_FFX_RST : STD_LOGIC; 
  signal nx54672z218_F5MUX : STD_LOGIC; 
  signal nx54672z220 : STD_LOGIC; 
  signal nx54672z218_BXINV : STD_LOGIC; 
  signal nx54672z219 : STD_LOGIC; 
  signal romedatao3_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z247 : STD_LOGIC; 
  signal romedatao3_s_5_BXINV : STD_LOGIC; 
  signal romedatao3_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z246 : STD_LOGIC; 
  signal romedatao3_s_5_BYINV : STD_LOGIC; 
  signal nx54672z242_F5MUX : STD_LOGIC; 
  signal nx54672z244 : STD_LOGIC; 
  signal nx54672z242_BXINV : STD_LOGIC; 
  signal nx54672z243 : STD_LOGIC; 
  signal romedatao3_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z258 : STD_LOGIC; 
  signal romedatao3_s_3_BXINV : STD_LOGIC; 
  signal romedatao3_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z257 : STD_LOGIC; 
  signal romedatao3_s_3_BYINV : STD_LOGIC; 
  signal nx54672z254_F5MUX : STD_LOGIC; 
  signal nx54672z255 : STD_LOGIC; 
  signal nx54672z254_BXINV : STD_LOGIC; 
  signal U1_ROME3_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal romedatao6_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z436 : STD_LOGIC; 
  signal romedatao6_s_6_BXINV : STD_LOGIC; 
  signal romedatao6_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z435 : STD_LOGIC; 
  signal romedatao6_s_6_BYINV : STD_LOGIC; 
  signal nx54672z431_F5MUX : STD_LOGIC; 
  signal nx54672z433 : STD_LOGIC; 
  signal nx54672z431_BXINV : STD_LOGIC; 
  signal nx54672z432 : STD_LOGIC; 
  signal romedatao6_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z442 : STD_LOGIC; 
  signal romedatao6_s_5_BXINV : STD_LOGIC; 
  signal romedatao6_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z441 : STD_LOGIC; 
  signal romedatao6_s_5_BYINV : STD_LOGIC; 
  signal nx54672z437_F5MUX : STD_LOGIC; 
  signal nx54672z439 : STD_LOGIC; 
  signal nx54672z437_BXINV : STD_LOGIC; 
  signal nx54672z438 : STD_LOGIC; 
  signal romedatao8_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z554 : STD_LOGIC; 
  signal romedatao8_s_8_BXINV : STD_LOGIC; 
  signal romedatao8_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z553 : STD_LOGIC; 
  signal romedatao8_s_8_BYINV : STD_LOGIC; 
  signal nx54672z549_F5MUX : STD_LOGIC; 
  signal nx54672z551 : STD_LOGIC; 
  signal nx54672z549_BXINV : STD_LOGIC; 
  signal nx54672z550 : STD_LOGIC; 
  signal romedatao8_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z560 : STD_LOGIC; 
  signal romedatao8_s_7_BXINV : STD_LOGIC; 
  signal romedatao8_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z559 : STD_LOGIC; 
  signal romedatao8_s_7_BYINV : STD_LOGIC; 
  signal nx54672z555_F5MUX : STD_LOGIC; 
  signal nx54672z557 : STD_LOGIC; 
  signal nx54672z555_BXINV : STD_LOGIC; 
  signal nx54672z556 : STD_LOGIC; 
  signal romedatao8_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z566 : STD_LOGIC; 
  signal romedatao8_s_6_BXINV : STD_LOGIC; 
  signal romedatao8_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z565 : STD_LOGIC; 
  signal romedatao8_s_6_BYINV : STD_LOGIC; 
  signal nx54672z561_F5MUX : STD_LOGIC; 
  signal nx54672z563 : STD_LOGIC; 
  signal nx54672z561_BXINV : STD_LOGIC; 
  signal nx54672z562 : STD_LOGIC; 
  signal romedatao8_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z572 : STD_LOGIC; 
  signal romedatao8_s_5_BXINV : STD_LOGIC; 
  signal romedatao8_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z571 : STD_LOGIC; 
  signal romedatao8_s_5_BYINV : STD_LOGIC; 
  signal nx54672z567_F5MUX : STD_LOGIC; 
  signal nx54672z569 : STD_LOGIC; 
  signal nx54672z567_BXINV : STD_LOGIC; 
  signal nx54672z568 : STD_LOGIC; 
  signal romedatao8_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z578 : STD_LOGIC; 
  signal romedatao8_s_4_BXINV : STD_LOGIC; 
  signal romedatao8_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z577 : STD_LOGIC; 
  signal romedatao8_s_4_BYINV : STD_LOGIC; 
  signal nx54672z573_F5MUX : STD_LOGIC; 
  signal nx54672z575 : STD_LOGIC; 
  signal nx54672z573_BXINV : STD_LOGIC; 
  signal nx54672z574 : STD_LOGIC; 
  signal romodatao6_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z1073 : STD_LOGIC; 
  signal romodatao6_s_11_BXINV : STD_LOGIC; 
  signal romodatao6_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z1072 : STD_LOGIC; 
  signal romodatao6_s_11_BYINV : STD_LOGIC; 
  signal nx54672z1068_F5MUX : STD_LOGIC; 
  signal nx54672z1070 : STD_LOGIC; 
  signal nx54672z1068_BXINV : STD_LOGIC; 
  signal nx54672z1069 : STD_LOGIC; 
  signal romodatao6_s_10_F5MUX : STD_LOGIC; 
  signal nx54672z1079 : STD_LOGIC; 
  signal romodatao6_s_10_BXINV : STD_LOGIC; 
  signal romodatao6_s_10_F6MUX : STD_LOGIC; 
  signal nx54672z1078 : STD_LOGIC; 
  signal romodatao6_s_10_BYINV : STD_LOGIC; 
  signal nx54672z1074_F5MUX : STD_LOGIC; 
  signal nx54672z1076 : STD_LOGIC; 
  signal nx54672z1074_BXINV : STD_LOGIC; 
  signal nx54672z1075 : STD_LOGIC; 
  signal romodatao6_s_1_F5MUX : STD_LOGIC; 
  signal nx54672z1133 : STD_LOGIC; 
  signal romodatao6_s_1_BXINV : STD_LOGIC; 
  signal romodatao6_s_1_F6MUX : STD_LOGIC; 
  signal nx54672z1132 : STD_LOGIC; 
  signal romodatao6_s_1_BYINV : STD_LOGIC; 
  signal nx54672z1128_F5MUX : STD_LOGIC; 
  signal nx54672z1130 : STD_LOGIC; 
  signal nx54672z1128_BXINV : STD_LOGIC; 
  signal nx54672z1129 : STD_LOGIC; 
  signal romedatao7_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z507 : STD_LOGIC; 
  signal romedatao7_s_5_BXINV : STD_LOGIC; 
  signal romedatao7_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z506 : STD_LOGIC; 
  signal romedatao7_s_5_BYINV : STD_LOGIC; 
  signal nx54672z502_F5MUX : STD_LOGIC; 
  signal nx54672z504 : STD_LOGIC; 
  signal nx54672z502_BXINV : STD_LOGIC; 
  signal nx54672z503 : STD_LOGIC; 
  signal romedatao7_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z513 : STD_LOGIC; 
  signal romedatao7_s_4_BXINV : STD_LOGIC; 
  signal romedatao7_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z512 : STD_LOGIC; 
  signal romedatao7_s_4_BYINV : STD_LOGIC; 
  signal nx54672z508_F5MUX : STD_LOGIC; 
  signal nx54672z510 : STD_LOGIC; 
  signal nx54672z508_BXINV : STD_LOGIC; 
  signal nx54672z509 : STD_LOGIC; 
  signal romodatao8_s_8_F5MUX : STD_LOGIC; 
  signal nx54672z1249 : STD_LOGIC; 
  signal romodatao8_s_8_BXINV : STD_LOGIC; 
  signal romodatao8_s_8_F6MUX : STD_LOGIC; 
  signal nx54672z1248 : STD_LOGIC; 
  signal romodatao8_s_8_BYINV : STD_LOGIC; 
  signal nx54672z1244_F5MUX : STD_LOGIC; 
  signal nx54672z1246 : STD_LOGIC; 
  signal nx54672z1244_BXINV : STD_LOGIC; 
  signal nx54672z1245 : STD_LOGIC; 
  signal romodatao8_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z1255 : STD_LOGIC; 
  signal romodatao8_s_7_BXINV : STD_LOGIC; 
  signal romodatao8_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z1254 : STD_LOGIC; 
  signal romodatao8_s_7_BYINV : STD_LOGIC; 
  signal nx54672z1250_F5MUX : STD_LOGIC; 
  signal nx54672z1252 : STD_LOGIC; 
  signal nx54672z1250_BXINV : STD_LOGIC; 
  signal nx54672z1251 : STD_LOGIC; 
  signal romodatao8_s_6_F5MUX : STD_LOGIC; 
  signal nx54672z1261 : STD_LOGIC; 
  signal romodatao8_s_6_BXINV : STD_LOGIC; 
  signal romodatao8_s_6_F6MUX : STD_LOGIC; 
  signal nx54672z1260 : STD_LOGIC; 
  signal romodatao8_s_6_BYINV : STD_LOGIC; 
  signal nx54672z1256_F5MUX : STD_LOGIC; 
  signal nx54672z1258 : STD_LOGIC; 
  signal nx54672z1256_BXINV : STD_LOGIC; 
  signal nx54672z1257 : STD_LOGIC; 
  signal romodatao8_s_5_F5MUX : STD_LOGIC; 
  signal nx54672z1267 : STD_LOGIC; 
  signal romodatao8_s_5_BXINV : STD_LOGIC; 
  signal romodatao8_s_5_F6MUX : STD_LOGIC; 
  signal nx54672z1266 : STD_LOGIC; 
  signal romodatao8_s_5_BYINV : STD_LOGIC; 
  signal nx54672z1262_F5MUX : STD_LOGIC; 
  signal nx54672z1264 : STD_LOGIC; 
  signal nx54672z1262_BXINV : STD_LOGIC; 
  signal nx54672z1263 : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_FFY_RST : STD_LOGIC; 
  signal romodatao8_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z1273 : STD_LOGIC; 
  signal romodatao8_s_4_BXINV : STD_LOGIC; 
  signal romodatao8_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z1272 : STD_LOGIC; 
  signal romodatao8_s_4_BYINV : STD_LOGIC; 
  signal nx54672z1268_F5MUX : STD_LOGIC; 
  signal nx54672z1270 : STD_LOGIC; 
  signal nx54672z1268_BXINV : STD_LOGIC; 
  signal nx54672z1269 : STD_LOGIC; 
  signal romodatao7_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z1140 : STD_LOGIC; 
  signal romodatao7_s_13_BXINV : STD_LOGIC; 
  signal romodatao7_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z1139 : STD_LOGIC; 
  signal romodatao7_s_13_BYINV : STD_LOGIC; 
  signal nx54672z1136_F5MUX : STD_LOGIC; 
  signal nx54672z1137 : STD_LOGIC; 
  signal nx54672z1136_BXINV : STD_LOGIC; 
  signal nx54672z1136_G : STD_LOGIC; 
  signal romodatao7_s_12_F5MUX : STD_LOGIC; 
  signal nx54672z1146 : STD_LOGIC; 
  signal romodatao7_s_12_BXINV : STD_LOGIC; 
  signal romodatao7_s_12_F6MUX : STD_LOGIC; 
  signal nx54672z1145 : STD_LOGIC; 
  signal romodatao7_s_12_BYINV : STD_LOGIC; 
  signal nx54672z1141_F5MUX : STD_LOGIC; 
  signal nx54672z1143 : STD_LOGIC; 
  signal nx54672z1141_BXINV : STD_LOGIC; 
  signal nx54672z1142 : STD_LOGIC; 
  signal romodatao7_s_4_F5MUX : STD_LOGIC; 
  signal nx54672z1194 : STD_LOGIC; 
  signal romodatao7_s_4_BXINV : STD_LOGIC; 
  signal romodatao7_s_4_F6MUX : STD_LOGIC; 
  signal nx54672z1193 : STD_LOGIC; 
  signal romodatao7_s_4_BYINV : STD_LOGIC; 
  signal nx54672z1189_F5MUX : STD_LOGIC; 
  signal nx54672z1191 : STD_LOGIC; 
  signal nx54672z1189_BXINV : STD_LOGIC; 
  signal nx54672z1190 : STD_LOGIC; 
  signal romodatao7_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z1200 : STD_LOGIC; 
  signal romodatao7_s_3_BXINV : STD_LOGIC; 
  signal romodatao7_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z1199 : STD_LOGIC; 
  signal romodatao7_s_3_BYINV : STD_LOGIC; 
  signal nx54672z1195_F5MUX : STD_LOGIC; 
  signal nx54672z1197 : STD_LOGIC; 
  signal nx54672z1195_BXINV : STD_LOGIC; 
  signal nx54672z1196 : STD_LOGIC; 
  signal romodatao7_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z1206 : STD_LOGIC; 
  signal romodatao7_s_2_BXINV : STD_LOGIC; 
  signal romodatao7_s_2_F6MUX : STD_LOGIC; 
  signal nx54672z1205 : STD_LOGIC; 
  signal romodatao7_s_2_BYINV : STD_LOGIC; 
  signal nx54672z1201_F5MUX : STD_LOGIC; 
  signal nx54672z1203 : STD_LOGIC; 
  signal nx54672z1201_BXINV : STD_LOGIC; 
  signal nx54672z1202 : STD_LOGIC; 
  signal romodatao7_s_1_F5MUX : STD_LOGIC; 
  signal nx54672z1212 : STD_LOGIC; 
  signal romodatao7_s_1_BXINV : STD_LOGIC; 
  signal romodatao7_s_1_F6MUX : STD_LOGIC; 
  signal nx54672z1211 : STD_LOGIC; 
  signal romodatao7_s_1_BYINV : STD_LOGIC; 
  signal nx54672z1207_F5MUX : STD_LOGIC; 
  signal nx54672z1209 : STD_LOGIC; 
  signal nx54672z1207_BXINV : STD_LOGIC; 
  signal nx54672z1208 : STD_LOGIC; 
  signal romodatao7_s_0_F5MUX : STD_LOGIC; 
  signal nx54672z1214 : STD_LOGIC; 
  signal romodatao7_s_0_BXINV : STD_LOGIC; 
  signal romodatao7_s_0_F6MUX : STD_LOGIC; 
  signal nx54672z1213 : STD_LOGIC; 
  signal romodatao7_s_0_BYINV : STD_LOGIC; 
  signal U1_ROMO7_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROMO7_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROMO7_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROMO7_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romodatao6_s_0_F5MUX : STD_LOGIC; 
  signal nx54672z1135 : STD_LOGIC; 
  signal romodatao6_s_0_BXINV : STD_LOGIC; 
  signal romodatao6_s_0_F6MUX : STD_LOGIC; 
  signal nx54672z1134 : STD_LOGIC; 
  signal romodatao6_s_0_BYINV : STD_LOGIC; 
  signal U1_ROMO6_modgen_rom_ix0_nx_ro64_32_u_F5MUX : STD_LOGIC; 
  signal U1_ROMO6_modgen_rom_ix0_nx_rm64_16_l : STD_LOGIC; 
  signal U1_ROMO6_modgen_rom_ix0_nx_ro64_32_u_BXINV : STD_LOGIC; 
  signal U1_ROMO6_modgen_rom_ix0_nx_rm64_16_u : STD_LOGIC; 
  signal romodatao4_s_11_F5MUX : STD_LOGIC; 
  signal nx54672z915 : STD_LOGIC; 
  signal romodatao4_s_11_BXINV : STD_LOGIC; 
  signal romodatao4_s_11_F6MUX : STD_LOGIC; 
  signal nx54672z914 : STD_LOGIC; 
  signal romodatao4_s_11_BYINV : STD_LOGIC; 
  signal nx54672z910_F5MUX : STD_LOGIC; 
  signal nx54672z912 : STD_LOGIC; 
  signal nx54672z910_BXINV : STD_LOGIC; 
  signal nx54672z911 : STD_LOGIC; 
  signal romodatao3_s_7_F5MUX : STD_LOGIC; 
  signal nx54672z860 : STD_LOGIC; 
  signal romodatao3_s_7_BXINV : STD_LOGIC; 
  signal romodatao3_s_7_F6MUX : STD_LOGIC; 
  signal nx54672z859 : STD_LOGIC; 
  signal romodatao3_s_7_BYINV : STD_LOGIC; 
  signal nx54672z855_F5MUX : STD_LOGIC; 
  signal nx54672z857 : STD_LOGIC; 
  signal nx54672z855_BXINV : STD_LOGIC; 
  signal nx54672z856 : STD_LOGIC; 
  signal romodatao3_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z884 : STD_LOGIC; 
  signal romodatao3_s_3_BXINV : STD_LOGIC; 
  signal romodatao3_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z883 : STD_LOGIC; 
  signal romodatao3_s_3_BYINV : STD_LOGIC; 
  signal nx54672z879_F5MUX : STD_LOGIC; 
  signal nx54672z881 : STD_LOGIC; 
  signal nx54672z879_BXINV : STD_LOGIC; 
  signal nx54672z880 : STD_LOGIC; 
  signal romodatao3_s_1_F5MUX : STD_LOGIC; 
  signal nx54672z896 : STD_LOGIC; 
  signal romodatao3_s_1_BXINV : STD_LOGIC; 
  signal romodatao3_s_1_F6MUX : STD_LOGIC; 
  signal nx54672z895 : STD_LOGIC; 
  signal romodatao3_s_1_BYINV : STD_LOGIC; 
  signal nx54672z891_F5MUX : STD_LOGIC; 
  signal nx54672z893 : STD_LOGIC; 
  signal nx54672z891_BXINV : STD_LOGIC; 
  signal nx54672z892 : STD_LOGIC; 
  signal romedatao8_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z583 : STD_LOGIC; 
  signal romedatao8_s_3_BXINV : STD_LOGIC; 
  signal romedatao8_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z582 : STD_LOGIC; 
  signal romedatao8_s_3_BYINV : STD_LOGIC; 
  signal nx54672z579_F5MUX : STD_LOGIC; 
  signal nx54672z580 : STD_LOGIC; 
  signal nx54672z579_BXINV : STD_LOGIC; 
  signal U1_ROME8_modgen_rom_ix2_nx_rm64_16_u : STD_LOGIC; 
  signal romodatao8_s_13_F5MUX : STD_LOGIC; 
  signal nx54672z1219 : STD_LOGIC; 
  signal romodatao8_s_13_BXINV : STD_LOGIC; 
  signal romodatao8_s_13_F6MUX : STD_LOGIC; 
  signal nx54672z1218 : STD_LOGIC; 
  signal romodatao8_s_13_BYINV : STD_LOGIC; 
  signal nx54672z1215_F5MUX : STD_LOGIC; 
  signal nx54672z1216 : STD_LOGIC; 
  signal nx54672z1215_BXINV : STD_LOGIC; 
  signal nx54672z1215_G : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_8_FFX_RST : STD_LOGIC; 
  signal romodatao8_s_3_F5MUX : STD_LOGIC; 
  signal nx54672z1279 : STD_LOGIC; 
  signal romodatao8_s_3_BXINV : STD_LOGIC; 
  signal romodatao8_s_3_F6MUX : STD_LOGIC; 
  signal nx54672z1278 : STD_LOGIC; 
  signal romodatao8_s_3_BYINV : STD_LOGIC; 
  signal nx54672z1274_F5MUX : STD_LOGIC; 
  signal nx54672z1276 : STD_LOGIC; 
  signal nx54672z1274_BXINV : STD_LOGIC; 
  signal nx54672z1275 : STD_LOGIC; 
  signal romodatao8_s_2_F5MUX : STD_LOGIC; 
  signal nx54672z1285 : STD_LOGIC; 
  signal romodatao8_s_2_BXINV : STD_LOGIC; 
  signal romodatao8_s_2_F6MUX : STD_LOGIC; 
  signal nx54672z1284 : STD_LOGIC; 
  signal romodatao8_s_2_BYINV : STD_LOGIC; 
  signal nx54672z1280_F5MUX : STD_LOGIC; 
  signal nx54672z1282 : STD_LOGIC; 
  signal nx54672z1280_BXINV : STD_LOGIC; 
  signal nx54672z1281 : STD_LOGIC; 
  signal romodatao8_s_1_F5MUX : STD_LOGIC; 
  signal nx54672z1291 : STD_LOGIC; 
  signal romodatao8_s_1_BXINV : STD_LOGIC; 
  signal romodatao8_s_1_F6MUX : STD_LOGIC; 
  signal nx54672z1290 : STD_LOGIC; 
  signal romodatao8_s_1_BYINV : STD_LOGIC; 
  signal nx54672z1286_F5MUX : STD_LOGIC; 
  signal nx54672z1288 : STD_LOGIC; 
  signal nx54672z1286_BXINV : STD_LOGIC; 
  signal nx54672z1287 : STD_LOGIC; 
  signal dcto1_10_ENABLE : STD_LOGIC; 
  signal dcto1_10_GTS_OR_T : STD_LOGIC; 
  signal dcto1_10_O : STD_LOGIC; 
  signal dcto1_11_ENABLE : STD_LOGIC; 
  signal dcto1_11_GTS_OR_T : STD_LOGIC; 
  signal dcto1_11_O : STD_LOGIC; 
  signal clk_INBUF : STD_LOGIC; 
  signal idv_INBUF : STD_LOGIC; 
  signal odv_ENABLE : STD_LOGIC; 
  signal odv_GTS_OR_T : STD_LOGIC; 
  signal odv_O : STD_LOGIC; 
  signal rst_INBUF : STD_LOGIC; 
  signal odv1_ENABLE : STD_LOGIC; 
  signal odv1_GTS_OR_T : STD_LOGIC; 
  signal odv1_O : STD_LOGIC; 
  signal dcti_0_INBUF : STD_LOGIC; 
  signal dcti_1_INBUF : STD_LOGIC; 
  signal dcti_2_INBUF : STD_LOGIC; 
  signal dcti_3_INBUF : STD_LOGIC; 
  signal dcti_4_INBUF : STD_LOGIC; 
  signal dcti_5_INBUF : STD_LOGIC; 
  signal dcti_6_INBUF : STD_LOGIC; 
  signal dcti_7_INBUF : STD_LOGIC; 
  signal dcto_0_ENABLE : STD_LOGIC; 
  signal dcto_0_GTS_OR_T : STD_LOGIC; 
  signal dcto_0_O : STD_LOGIC; 
  signal dcto_1_ENABLE : STD_LOGIC; 
  signal dcto_1_GTS_OR_T : STD_LOGIC; 
  signal dcto_1_O : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_7_10_FFX_RSTAND : STD_LOGIC; 
  signal dcto_2_ENABLE : STD_LOGIC; 
  signal dcto_2_GTS_OR_T : STD_LOGIC; 
  signal dcto_2_O : STD_LOGIC; 
  signal dcto_3_ENABLE : STD_LOGIC; 
  signal dcto_3_GTS_OR_T : STD_LOGIC; 
  signal dcto_3_O : STD_LOGIC; 
  signal dcto_4_ENABLE : STD_LOGIC; 
  signal dcto_4_GTS_OR_T : STD_LOGIC; 
  signal dcto_4_O : STD_LOGIC; 
  signal dcto_5_ENABLE : STD_LOGIC; 
  signal dcto_5_GTS_OR_T : STD_LOGIC; 
  signal dcto_5_O : STD_LOGIC; 
  signal dcto_6_ENABLE : STD_LOGIC; 
  signal dcto_6_GTS_OR_T : STD_LOGIC; 
  signal dcto_6_O : STD_LOGIC; 
  signal dcto_7_ENABLE : STD_LOGIC; 
  signal dcto_7_GTS_OR_T : STD_LOGIC; 
  signal dcto_7_O : STD_LOGIC; 
  signal dcto_8_ENABLE : STD_LOGIC; 
  signal dcto_8_GTS_OR_T : STD_LOGIC; 
  signal dcto_8_O : STD_LOGIC; 
  signal dcto_9_ENABLE : STD_LOGIC; 
  signal dcto_9_GTS_OR_T : STD_LOGIC; 
  signal dcto_9_O : STD_LOGIC; 
  signal ready_ENABLE : STD_LOGIC; 
  signal ready_GTS_OR_T : STD_LOGIC; 
  signal ready_O : STD_LOGIC; 
  signal dcto_10_ENABLE : STD_LOGIC; 
  signal dcto_10_GTS_OR_T : STD_LOGIC; 
  signal dcto_10_O : STD_LOGIC; 
  signal dcto_11_ENABLE : STD_LOGIC; 
  signal dcto_11_GTS_OR_T : STD_LOGIC; 
  signal dcto_11_O : STD_LOGIC; 
  signal dcto1_0_ENABLE : STD_LOGIC; 
  signal dcto1_0_GTS_OR_T : STD_LOGIC; 
  signal dcto1_0_O : STD_LOGIC; 
  signal dcto1_1_ENABLE : STD_LOGIC; 
  signal dcto1_1_GTS_OR_T : STD_LOGIC; 
  signal dcto1_1_O : STD_LOGIC; 
  signal dcto1_2_ENABLE : STD_LOGIC; 
  signal dcto1_2_GTS_OR_T : STD_LOGIC; 
  signal dcto1_2_O : STD_LOGIC; 
  signal dcto1_3_ENABLE : STD_LOGIC; 
  signal dcto1_3_GTS_OR_T : STD_LOGIC; 
  signal dcto1_3_O : STD_LOGIC; 
  signal dcto1_4_ENABLE : STD_LOGIC; 
  signal dcto1_4_GTS_OR_T : STD_LOGIC; 
  signal dcto1_4_O : STD_LOGIC; 
  signal dcto1_5_ENABLE : STD_LOGIC; 
  signal dcto1_5_GTS_OR_T : STD_LOGIC; 
  signal dcto1_5_O : STD_LOGIC; 
  signal dcto1_6_ENABLE : STD_LOGIC; 
  signal dcto1_6_GTS_OR_T : STD_LOGIC; 
  signal dcto1_6_O : STD_LOGIC; 
  signal dcto1_7_ENABLE : STD_LOGIC; 
  signal dcto1_7_GTS_OR_T : STD_LOGIC; 
  signal dcto1_7_O : STD_LOGIC; 
  signal dcto1_8_ENABLE : STD_LOGIC; 
  signal dcto1_8_GTS_OR_T : STD_LOGIC; 
  signal dcto1_8_O : STD_LOGIC; 
  signal dcto1_9_ENABLE : STD_LOGIC; 
  signal dcto1_9_GTS_OR_T : STD_LOGIC; 
  signal dcto1_9_O : STD_LOGIC; 
  signal clk_ibuf_BUFG_S_INVNOT : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOPB3 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOPB2 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOPB1 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOPB0 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB31 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB30 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB29 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB28 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB27 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB26 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB25 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB24 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB23 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB22 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB21 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB20 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB19 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB18 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB17 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB16 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB15 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB14 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB13 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB12 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB11 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOB10 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOPA3 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOPA2 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOPA1 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOPA0 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA31 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA30 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA29 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA28 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA27 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA26 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA25 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA24 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA23 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA22 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA21 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA20 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA19 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA18 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA17 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA16 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA15 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA14 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA13 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA12 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA11 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA10 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA9 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA8 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA7 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA6 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA5 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA4 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA3 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA2 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA1 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DOA0 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIPB3 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIPB2 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIPB1 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIPB0 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB31 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB30 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB29 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB28 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB27 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB26 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB25 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB24 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB23 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB22 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB21 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB20 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB19 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB18 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB17 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB16 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB15 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB14 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB13 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB12 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB11 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB10 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB9 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB8 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB7 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB6 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB5 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB4 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB3 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB2 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB1 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIB0 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIPA3 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIPA2 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA31 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA30 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA29 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA28 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA27 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA26 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA25 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA24 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA23 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA22 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA21 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA20 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA19 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA18 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA17 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_DIA16 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_ADDRB0 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_ADDRB1 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_ADDRB2 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_ADDRB3 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_ADDRA0 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_ADDRA1 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_ADDRA2 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_ADDRA3 : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_WEB_INTNOT : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_SSRB_INTNOT : STD_LOGIC; 
  signal U2_RAM_mem_ix3035z34088_SSRA_INTNOT : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOPB3 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOPB2 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOPB1 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOPB0 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB31 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB30 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB29 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB28 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB27 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB26 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB25 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB24 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB23 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB22 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB21 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB20 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB19 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB18 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB17 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB16 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB15 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB14 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB13 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB12 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB11 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOB10 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOPA3 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOPA2 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOPA1 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOPA0 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA31 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA30 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA29 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA28 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA27 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA26 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA25 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA24 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA23 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA22 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA21 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA20 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA19 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA18 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA17 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA16 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA15 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA14 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA13 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA12 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA11 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA10 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA9 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA8 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA7 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA6 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA5 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA4 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA3 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA2 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA1 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DOA0 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIPB3 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIPB2 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIPB1 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIPB0 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB31 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB30 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB29 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB28 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB27 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB26 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB25 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB24 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB23 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB22 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB21 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB20 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB19 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB18 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB17 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB16 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB15 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB14 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB13 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB12 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB11 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB10 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB9 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB8 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB7 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB6 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB5 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB4 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB3 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB2 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB1 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIB0 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIPA3 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIPA2 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA31 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA30 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA29 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA28 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA27 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA26 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA25 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA24 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA23 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA22 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA21 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA20 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA19 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA18 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA17 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_DIA16 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_ADDRB0 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_ADDRB1 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_ADDRB2 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_ADDRB3 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_ADDRA0 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_ADDRA1 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_ADDRA2 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_ADDRA3 : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_WEB_INTNOT : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_SSRB_INTNOT : STD_LOGIC; 
  signal U1_RAM_mem_ix3035z34088_SSRA_INTNOT : STD_LOGIC; 
  signal U_DBUFCTL_rtlc4n377_F5MUX : STD_LOGIC; 
  signal nx31259z2 : STD_LOGIC; 
  signal U_DBUFCTL_rtlc4n377_BXINV : STD_LOGIC; 
  signal nx31259z1 : STD_LOGIC; 
  signal U_DCT2D_rtlc2n584_F5MUX : STD_LOGIC; 
  signal U_DCT2D_nx1822z2 : STD_LOGIC; 
  signal U_DCT2D_rtlc2n584_BXINV : STD_LOGIC; 
  signal U_DCT2D_nx1822z1 : STD_LOGIC; 
  signal U_DCT2D_istate_reg_1_DXMUX : STD_LOGIC; 
  signal U_DCT2D_rtlcn348 : STD_LOGIC; 
  signal U_DCT2D_istate_reg_1_DYMUX : STD_LOGIC; 
  signal U_DCT2D_istate_reg_1_SRINV : STD_LOGIC; 
  signal U_DCT2D_istate_reg_1_CLKINV : STD_LOGIC; 
  signal U_DCT2D_istate_reg_1_CEINV : STD_LOGIC; 
  signal memswitchrd_s_DXMUX : STD_LOGIC; 
  signal memswitchrd_s_FXMUX : STD_LOGIC; 
  signal memswitchrd_s_F : STD_LOGIC; 
  signal memswitchrd_s_CLKINV : STD_LOGIC; 
  signal memswitchrd_s_CEINV : STD_LOGIC; 
  signal ramraddro_s_5_DXMUX : STD_LOGIC; 
  signal U_DCT2D_nx51407z1 : STD_LOGIC; 
  signal ramraddro_s_5_DYMUX : STD_LOGIC; 
  signal U_DCT2D_nx50410z1 : STD_LOGIC; 
  signal ramraddro_s_5_SRINV : STD_LOGIC; 
  signal ramraddro_s_5_CLKINV : STD_LOGIC; 
  signal ramraddro_s_5_CEINV : STD_LOGIC; 
  signal memswitchwr_s_F : STD_LOGIC; 
  signal memswitchwr_s_DYMUX : STD_LOGIC; 
  signal memswitchwr_s_GYMUX : STD_LOGIC; 
  signal memswitchwr_s_G : STD_LOGIC; 
  signal memswitchwr_s_CLKINV : STD_LOGIC; 
  signal memswitchwr_s_CEINV : STD_LOGIC; 
  signal U_DBUFCTL_mem1_full_reg_F : STD_LOGIC; 
  signal U_DBUFCTL_mem1_full_reg_DYMUX : STD_LOGIC; 
  signal U_DBUFCTL_mem1_full_reg_GYMUX : STD_LOGIC; 
  signal U_DBUFCTL_mem1_full_reg_G : STD_LOGIC; 
  signal U_DBUFCTL_mem1_full_reg_CLKINV : STD_LOGIC; 
  signal U_DBUFCTL_mem1_full_reg_CEINV : STD_LOGIC; 
  signal U_DBUFCTL_mem1_lock_reg_F : STD_LOGIC; 
  signal U_DBUFCTL_mem1_lock_reg_DYMUX : STD_LOGIC; 
  signal U_DBUFCTL_rtlcn35 : STD_LOGIC; 
  signal U_DBUFCTL_mem1_lock_reg_CLKINV : STD_LOGIC; 
  signal U_DBUFCTL_mem1_lock_reg_CEINV : STD_LOGIC; 
  signal U_DBUFCTL_mem2_full_reg_F : STD_LOGIC; 
  signal U_DBUFCTL_mem2_full_reg_DYMUX : STD_LOGIC; 
  signal U_DBUFCTL_mem2_full_reg_GYMUX : STD_LOGIC; 
  signal U_DBUFCTL_mem2_full_reg_G : STD_LOGIC; 
  signal U_DBUFCTL_mem2_full_reg_CLKINV : STD_LOGIC; 
  signal U_DBUFCTL_mem2_full_reg_CEINV : STD_LOGIC; 
  signal U_DBUFCTL_mem2_lock_reg_F : STD_LOGIC; 
  signal U_DBUFCTL_mem2_lock_reg_DYMUX : STD_LOGIC; 
  signal U_DBUFCTL_rtlcn76 : STD_LOGIC; 
  signal U_DBUFCTL_mem2_lock_reg_CLKINV : STD_LOGIC; 
  signal U_DBUFCTL_mem2_lock_reg_CEINV : STD_LOGIC; 
  signal U_DCT2D_col_reg_2_DYMUX : STD_LOGIC; 
  signal U_DCT2D_nx35453z1 : STD_LOGIC; 
  signal U_DCT2D_col_reg_2_CLKINV : STD_LOGIC; 
  signal U_DCT2D_col_reg_2_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_col_reg_2_DYMUX : STD_LOGIC; 
  signal U_DCT1D_nx35453z1 : STD_LOGIC; 
  signal U_DCT1D_col_reg_2_CLKINV : STD_LOGIC; 
  signal U_DCT1D_col_reg_2_CEINV : STD_LOGIC; 
  signal U_DCT1D_ready_F : STD_LOGIC; 
  signal U_DCT1D_ready_DYMUX : STD_LOGIC; 
  signal U_DCT1D_ready_GYMUX : STD_LOGIC; 
  signal U_DCT1D_ready_G : STD_LOGIC; 
  signal U_DCT1D_ready_CLKINV : STD_LOGIC; 
  signal U_DCT1D_ready_CEINV : STD_LOGIC; 
  signal U_DCT1D_row_reg_2_DYMUX : STD_LOGIC; 
  signal U_DCT1D_nx53037z1 : STD_LOGIC; 
  signal U_DCT1D_row_reg_2_CLKINV : STD_LOGIC; 
  signal U_DCT1D_row_reg_2_CEINV : STD_LOGIC; 
  signal rome2addro0_s_5_DXMUX : STD_LOGIC; 
  signal rome2addro0_s_5_DYMUX : STD_LOGIC; 
  signal rome2addro0_s_5_SRINV : STD_LOGIC; 
  signal rome2addro0_s_5_CLKINV : STD_LOGIC; 
  signal rome2addro0_s_5_CEINV : STD_LOGIC; 
  signal romeaddro0_s_5_DXMUX : STD_LOGIC; 
  signal romeaddro0_s_5_DYMUX : STD_LOGIC; 
  signal romeaddro0_s_5_SRINV : STD_LOGIC; 
  signal romeaddro0_s_5_CLKINV : STD_LOGIC; 
  signal romeaddro0_s_5_CEINV : STD_LOGIC; 
  signal ramraddro_s_0_F : STD_LOGIC; 
  signal ramraddro_s_0_DYMUX : STD_LOGIC; 
  signal U_DCT2D_nx38901z1 : STD_LOGIC; 
  signal ramraddro_s_0_CLKINV : STD_LOGIC; 
  signal ramraddro_s_0_CEINV : STD_LOGIC; 
  signal ramraddro_s_1_F : STD_LOGIC; 
  signal ramraddro_s_1_DYMUX : STD_LOGIC; 
  signal U_DCT2D_nx39898z1 : STD_LOGIC; 
  signal ramraddro_s_1_CLKINV : STD_LOGIC; 
  signal ramraddro_s_1_CEINV : STD_LOGIC; 
  signal ramraddro_s_2_DYMUX : STD_LOGIC; 
  signal U_DCT2D_nx40895z1 : STD_LOGIC; 
  signal ramraddro_s_2_CLKINV : STD_LOGIC; 
  signal ramraddro_s_2_CEINV : STD_LOGIC; 
  signal U_DCT1D_istate_reg_1_DXMUX : STD_LOGIC; 
  signal U_DCT1D_rtlcn403 : STD_LOGIC; 
  signal U_DCT1D_istate_reg_1_DYMUX : STD_LOGIC; 
  signal U_DCT1D_rtlcn349 : STD_LOGIC; 
  signal U_DCT1D_istate_reg_1_SRINV : STD_LOGIC; 
  signal U_DCT1D_istate_reg_1_CLKINV : STD_LOGIC; 
  signal U_DCT1D_istate_reg_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_2_DYMUX : STD_LOGIC; 
  signal U_DCT1D_nx59993z1 : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_2_CLKINV : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_2_CEINV : STD_LOGIC; 
  signal reqrdfail_s_F : STD_LOGIC; 
  signal reqrdfail_s_DYMUX : STD_LOGIC; 
  signal U_DBUFCTL_rtlcn7 : STD_LOGIC; 
  signal reqrdfail_s_CLKINV : STD_LOGIC; 
  signal reqrdfail_s_CEINV : STD_LOGIC; 
  signal reqwrfail_s_DYMUX : STD_LOGIC; 
  signal U_DBUFCTL_rtlc4n197 : STD_LOGIC; 
  signal reqwrfail_s_CLKINV : STD_LOGIC; 
  signal reqwrfail_s_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_1_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_1_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_1_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_1_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_1_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_3_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_3_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_3_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_3_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_3_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_5_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_5_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_5_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_5_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_5_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_7_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_7_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_7_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_7_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_7_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_10_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_10_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_10_CEINV : STD_LOGIC; 
  signal U_DCT2D_nx65206z252_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z571_G : STD_LOGIC; 
  signal U_DCT1D_rtlc2n469_F : STD_LOGIC; 
  signal U_DCT1D_rtlc2n469_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z251_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z251_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z218_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z218_G : STD_LOGIC; 
  signal ramraddro_s_3_DYMUX : STD_LOGIC; 
  signal ramraddro_s_3_BYINVNOT : STD_LOGIC; 
  signal ramraddro_s_3_CLKINV : STD_LOGIC; 
  signal ramraddro_s_3_CEINV : STD_LOGIC; 
  signal requestwr_s_DYMUX : STD_LOGIC; 
  signal requestwr_s_BYINVNOT : STD_LOGIC; 
  signal requestwr_s_CLKINV : STD_LOGIC; 
  signal requestwr_s_CEINV : STD_LOGIC; 
  signal U_DBUFCTL_rtlc4n378_F : STD_LOGIC; 
  signal U_DBUFCTL_rtlc4n378_G : STD_LOGIC; 
  signal U_DBUFCTL_rtlc4n374_G : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1702_F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1702_G : STD_LOGIC; 
  signal U_DCT1D_state_reg_1_DXMUX : STD_LOGIC; 
  signal U_DCT1D_state_reg_1_DYMUX : STD_LOGIC; 
  signal U_DCT1D_state_reg_1_G : STD_LOGIC; 
  signal U_DCT1D_state_reg_1_BYINVNOT : STD_LOGIC; 
  signal U_DCT1D_state_reg_1_SRINV : STD_LOGIC; 
  signal U_DCT1D_state_reg_1_CLKINV : STD_LOGIC; 
  signal U_DCT1D_state_reg_1_CEINV : STD_LOGIC; 
  signal U_DCT2D_rtlc2n581_F : STD_LOGIC; 
  signal U_DCT2D_rtlc2n581_G : STD_LOGIC; 
  signal U_DCT2D_nx64938z1_F : STD_LOGIC; 
  signal U_DCT2D_nx64938z1_G : STD_LOGIC; 
  signal U_DCT2D_rtlcs5_F : STD_LOGIC; 
  signal U_DCT2D_rtlcs5_G : STD_LOGIC; 
  signal U_DCT2D_rtlc2n580_F : STD_LOGIC; 
  signal U_DCT2D_rtlc2n580_G : STD_LOGIC; 
  signal U_DCT2D_nx14976z1_F : STD_LOGIC; 
  signal U_DCT2D_nx14976z1_G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_0_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_col_reg_0_DXMUX : STD_LOGIC; 
  signal U_DCT2D_col_reg_0_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_col_reg_0_DYMUX : STD_LOGIC; 
  signal U_DCT2D_nx36450z1 : STD_LOGIC; 
  signal U_DCT2D_col_reg_0_SRINV : STD_LOGIC; 
  signal U_DCT2D_col_reg_0_CLKINV : STD_LOGIC; 
  signal U_DCT2D_col_reg_0_CEINV : STD_LOGIC; 
  signal U_DCT1D_col_reg_0_DXMUX : STD_LOGIC; 
  signal U_DCT1D_col_reg_0_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_col_reg_0_DYMUX : STD_LOGIC; 
  signal U_DCT1D_nx36450z1 : STD_LOGIC; 
  signal U_DCT1D_col_reg_0_SRINV : STD_LOGIC; 
  signal U_DCT1D_col_reg_0_CLKINV : STD_LOGIC; 
  signal U_DCT1D_col_reg_0_CEINV : STD_LOGIC; 
  signal U_DCT2D_nx8385z1_F : STD_LOGIC; 
  signal U_DCT2D_nx8385z1_G : STD_LOGIC; 
  signal U_DCT1D_completed_reg_DYMUX : STD_LOGIC; 
  signal U_DCT1D_completed_reg_CLKINV : STD_LOGIC; 
  signal U_DCT1D_completed_reg_CEINV : STD_LOGIC; 
  signal U_DCT2D_nx38337z1_F : STD_LOGIC; 
  signal U_DCT2D_nx38337z1_G : STD_LOGIC; 
  signal U_DCT1D_nx47258z1_F : STD_LOGIC; 
  signal U_DCT1D_nx47258z1_G : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_1_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_1_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_1_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_1_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_3_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_3_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_3_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_3_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_5_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_5_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_5_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_5_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_5_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_7_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_7_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_7_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_7_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_7_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_1_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_1_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_1_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_1_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_3_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_3_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_3_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_3_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_5_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_5_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_5_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_5_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_5_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_7_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_7_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_7_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_7_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_7_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_1_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_1_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_1_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_1_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_3_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_3_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_3_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_3_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_5_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_5_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_5_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_5_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_5_CEINV : STD_LOGIC; 
  signal romo2addro0_s_1_DXMUX : STD_LOGIC; 
  signal romo2addro0_s_1_DYMUX : STD_LOGIC; 
  signal romo2addro0_s_1_SRINV : STD_LOGIC; 
  signal romo2addro0_s_1_CLKINV : STD_LOGIC; 
  signal romo2addro0_s_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_7_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_7_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_7_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_7_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_7_CEINV : STD_LOGIC; 
  signal romo2addro0_s_3_DXMUX : STD_LOGIC; 
  signal romo2addro0_s_3_DYMUX : STD_LOGIC; 
  signal romo2addro0_s_3_SRINV : STD_LOGIC; 
  signal romo2addro0_s_3_CLKINV : STD_LOGIC; 
  signal romo2addro0_s_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_1_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_1_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_1_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_1_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_1_CEINV : STD_LOGIC; 
  signal romo2addro1_s_1_DXMUX : STD_LOGIC; 
  signal romo2addro1_s_1_DYMUX : STD_LOGIC; 
  signal romo2addro1_s_1_SRINV : STD_LOGIC; 
  signal romo2addro1_s_1_CLKINV : STD_LOGIC; 
  signal romo2addro1_s_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_3_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_3_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_3_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_3_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_3_CEINV : STD_LOGIC; 
  signal romo2addro1_s_3_DXMUX : STD_LOGIC; 
  signal romo2addro1_s_3_DYMUX : STD_LOGIC; 
  signal romo2addro1_s_3_SRINV : STD_LOGIC; 
  signal romo2addro1_s_3_CLKINV : STD_LOGIC; 
  signal romo2addro1_s_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_5_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_5_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_5_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_5_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_5_CEINV : STD_LOGIC; 
  signal romo2addro2_s_1_DXMUX : STD_LOGIC; 
  signal romo2addro2_s_1_DYMUX : STD_LOGIC; 
  signal romo2addro2_s_1_SRINV : STD_LOGIC; 
  signal romo2addro2_s_1_CLKINV : STD_LOGIC; 
  signal romo2addro2_s_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_7_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_7_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_7_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_7_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_7_CEINV : STD_LOGIC; 
  signal romo2addro2_s_3_DXMUX : STD_LOGIC; 
  signal romo2addro2_s_3_DYMUX : STD_LOGIC; 
  signal romo2addro2_s_3_SRINV : STD_LOGIC; 
  signal romo2addro2_s_3_CLKINV : STD_LOGIC; 
  signal romo2addro2_s_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_1_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_1_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_1_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_1_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_1_CEINV : STD_LOGIC; 
  signal romo2addro3_s_1_DXMUX : STD_LOGIC; 
  signal romo2addro3_s_1_DYMUX : STD_LOGIC; 
  signal romo2addro3_s_1_SRINV : STD_LOGIC; 
  signal romo2addro3_s_1_CLKINV : STD_LOGIC; 
  signal romo2addro3_s_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_3_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_3_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_3_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_3_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_3_CEINV : STD_LOGIC; 
  signal romo2addro3_s_3_DXMUX : STD_LOGIC; 
  signal romo2addro3_s_3_DYMUX : STD_LOGIC; 
  signal romo2addro3_s_3_SRINV : STD_LOGIC; 
  signal romo2addro3_s_3_CLKINV : STD_LOGIC; 
  signal romo2addro3_s_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_5_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_5_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_5_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_5_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_5_CEINV : STD_LOGIC; 
  signal romo2addro4_s_1_DXMUX : STD_LOGIC; 
  signal romo2addro4_s_1_DYMUX : STD_LOGIC; 
  signal romo2addro4_s_1_SRINV : STD_LOGIC; 
  signal romo2addro4_s_1_CLKINV : STD_LOGIC; 
  signal romo2addro4_s_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_7_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_7_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_7_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_7_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_7_CEINV : STD_LOGIC; 
  signal romo2addro4_s_3_DXMUX : STD_LOGIC; 
  signal romo2addro4_s_3_DYMUX : STD_LOGIC; 
  signal romo2addro4_s_3_SRINV : STD_LOGIC; 
  signal romo2addro4_s_3_CLKINV : STD_LOGIC; 
  signal romo2addro4_s_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_1_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_1_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_1_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_1_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_1_CEINV : STD_LOGIC; 
  signal romo2addro5_s_1_DXMUX : STD_LOGIC; 
  signal romo2addro5_s_1_DYMUX : STD_LOGIC; 
  signal romo2addro5_s_1_SRINV : STD_LOGIC; 
  signal romo2addro5_s_1_CLKINV : STD_LOGIC; 
  signal romo2addro5_s_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_3_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_3_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_3_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_3_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_3_CEINV : STD_LOGIC; 
  signal romo2addro5_s_3_DXMUX : STD_LOGIC; 
  signal romo2addro5_s_3_DYMUX : STD_LOGIC; 
  signal romo2addro5_s_3_SRINV : STD_LOGIC; 
  signal romo2addro5_s_3_CLKINV : STD_LOGIC; 
  signal romo2addro5_s_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_5_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_5_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_5_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_5_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_5_CEINV : STD_LOGIC; 
  signal romo2addro6_s_1_DXMUX : STD_LOGIC; 
  signal romo2addro6_s_1_DYMUX : STD_LOGIC; 
  signal romo2addro6_s_1_SRINV : STD_LOGIC; 
  signal romo2addro6_s_1_CLKINV : STD_LOGIC; 
  signal romo2addro6_s_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_7_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_7_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_7_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_7_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_7_CEINV : STD_LOGIC; 
  signal romo2addro6_s_3_DXMUX : STD_LOGIC; 
  signal romo2addro6_s_3_DYMUX : STD_LOGIC; 
  signal romo2addro6_s_3_SRINV : STD_LOGIC; 
  signal romo2addro6_s_3_CLKINV : STD_LOGIC; 
  signal romo2addro6_s_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_1_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_1_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_1_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_1_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_1_CEINV : STD_LOGIC; 
  signal romo2addro7_s_1_DXMUX : STD_LOGIC; 
  signal romo2addro7_s_1_DYMUX : STD_LOGIC; 
  signal romo2addro7_s_1_SRINV : STD_LOGIC; 
  signal romo2addro7_s_1_CLKINV : STD_LOGIC; 
  signal romo2addro7_s_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_3_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_3_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_3_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_3_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_3_CEINV : STD_LOGIC; 
  signal romo2addro7_s_3_DXMUX : STD_LOGIC; 
  signal romo2addro7_s_3_DYMUX : STD_LOGIC; 
  signal romo2addro7_s_3_SRINV : STD_LOGIC; 
  signal romo2addro7_s_3_CLKINV : STD_LOGIC; 
  signal romo2addro7_s_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_5_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_5_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_5_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_5_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_5_CEINV : STD_LOGIC; 
  signal romo2addro8_s_1_DXMUX : STD_LOGIC; 
  signal romo2addro8_s_1_DYMUX : STD_LOGIC; 
  signal romo2addro8_s_1_SRINV : STD_LOGIC; 
  signal romo2addro8_s_1_CLKINV : STD_LOGIC; 
  signal romo2addro8_s_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_7_DXMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_7_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_7_SRINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_7_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_7_CEINV : STD_LOGIC; 
  signal romo2addro8_s_3_DXMUX : STD_LOGIC; 
  signal romo2addro8_s_3_DYMUX : STD_LOGIC; 
  signal romo2addro8_s_3_SRINV : STD_LOGIC; 
  signal romo2addro8_s_3_CLKINV : STD_LOGIC; 
  signal romo2addro8_s_3_CEINV : STD_LOGIC; 
  signal romo2addro9_s_1_DXMUX : STD_LOGIC; 
  signal romo2addro9_s_1_DYMUX : STD_LOGIC; 
  signal romo2addro9_s_1_SRINV : STD_LOGIC; 
  signal romo2addro9_s_1_CLKINV : STD_LOGIC; 
  signal romo2addro9_s_1_CEINV : STD_LOGIC; 
  signal romo2addro9_s_3_DXMUX : STD_LOGIC; 
  signal romo2addro9_s_3_DYMUX : STD_LOGIC; 
  signal romo2addro9_s_3_SRINV : STD_LOGIC; 
  signal romo2addro9_s_3_CLKINV : STD_LOGIC; 
  signal romo2addro9_s_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_7_7_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_7_7_BYINVNOT : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_7_7_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_7_7_CEINV : STD_LOGIC; 
  signal U_DCT2D_rtlc2n579_G : STD_LOGIC; 
  signal U_DCT2D_latch_done_reg_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latch_done_reg_BYINVNOT : STD_LOGIC; 
  signal U_DCT2D_latch_done_reg_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latch_done_reg_CEINV : STD_LOGIC; 
  signal U_DCT2D_nx6411z1_F : STD_LOGIC; 
  signal U_DCT2D_nx6411z1_G : STD_LOGIC; 
  signal U_DCT2D_nx41892z2_F : STD_LOGIC; 
  signal U_DCT2D_nx41892z2_G : STD_LOGIC; 
  signal U_DCT1D_row_reg_0_DXMUX : STD_LOGIC; 
  signal U_DCT1D_row_reg_0_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_row_reg_0_DYMUX : STD_LOGIC; 
  signal U_DCT1D_nx52040z1 : STD_LOGIC; 
  signal U_DCT1D_row_reg_0_SRINV : STD_LOGIC; 
  signal U_DCT1D_row_reg_0_CLKINV : STD_LOGIC; 
  signal U_DCT1D_row_reg_0_CEINV : STD_LOGIC; 
  signal U_DCT2D_state_reg_1_DXMUX : STD_LOGIC; 
  signal U_DCT2D_state_reg_1_DYMUX : STD_LOGIC; 
  signal U_DCT2D_state_reg_1_G : STD_LOGIC; 
  signal U_DCT2D_state_reg_1_BYINVNOT : STD_LOGIC; 
  signal U_DCT2D_state_reg_1_SRINV : STD_LOGIC; 
  signal U_DCT2D_state_reg_1_CLKINV : STD_LOGIC; 
  signal U_DCT2D_state_reg_1_CEINV : STD_LOGIC; 
  signal rome2addro10_s_1_DXMUX : STD_LOGIC; 
  signal rome2addro10_s_1_DYMUX : STD_LOGIC; 
  signal rome2addro10_s_1_SRINV : STD_LOGIC; 
  signal rome2addro10_s_1_CLKINV : STD_LOGIC; 
  signal rome2addro10_s_1_CEINV : STD_LOGIC; 
  signal rome2addro10_s_3_DXMUX : STD_LOGIC; 
  signal rome2addro10_s_3_DYMUX : STD_LOGIC; 
  signal rome2addro10_s_3_SRINV : STD_LOGIC; 
  signal rome2addro10_s_3_CLKINV : STD_LOGIC; 
  signal rome2addro10_s_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1684_F : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1684_G : STD_LOGIC; 
  signal romeaddro0_s_1_DXMUX : STD_LOGIC; 
  signal romeaddro0_s_1_DYMUX : STD_LOGIC; 
  signal romeaddro0_s_1_SRINV : STD_LOGIC; 
  signal romeaddro0_s_1_CLKINV : STD_LOGIC; 
  signal romeaddro0_s_1_CEINV : STD_LOGIC; 
  signal romeaddro0_s_3_DXMUX : STD_LOGIC; 
  signal romeaddro0_s_3_DYMUX : STD_LOGIC; 
  signal romeaddro0_s_3_SRINV : STD_LOGIC; 
  signal romeaddro0_s_3_CLKINV : STD_LOGIC; 
  signal romeaddro0_s_3_CEINV : STD_LOGIC; 
  signal romeaddro1_s_1_DXMUX : STD_LOGIC; 
  signal romeaddro1_s_1_DYMUX : STD_LOGIC; 
  signal romeaddro1_s_1_SRINV : STD_LOGIC; 
  signal romeaddro1_s_1_CLKINV : STD_LOGIC; 
  signal romeaddro1_s_1_CEINV : STD_LOGIC; 
  signal romeaddro1_s_3_DXMUX : STD_LOGIC; 
  signal romeaddro1_s_3_DYMUX : STD_LOGIC; 
  signal romeaddro1_s_3_SRINV : STD_LOGIC; 
  signal romeaddro1_s_3_CLKINV : STD_LOGIC; 
  signal romeaddro1_s_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_2_FFX_RST : STD_LOGIC; 
  signal romeaddro2_s_1_DXMUX : STD_LOGIC; 
  signal romeaddro2_s_1_DYMUX : STD_LOGIC; 
  signal romeaddro2_s_1_SRINV : STD_LOGIC; 
  signal romeaddro2_s_1_CLKINV : STD_LOGIC; 
  signal romeaddro2_s_1_CEINV : STD_LOGIC; 
  signal romeaddro2_s_3_DXMUX : STD_LOGIC; 
  signal romeaddro2_s_3_DYMUX : STD_LOGIC; 
  signal romeaddro2_s_3_SRINV : STD_LOGIC; 
  signal romeaddro2_s_3_CLKINV : STD_LOGIC; 
  signal romeaddro2_s_3_CEINV : STD_LOGIC; 
  signal romeaddro3_s_1_DXMUX : STD_LOGIC; 
  signal romeaddro3_s_1_DYMUX : STD_LOGIC; 
  signal romeaddro3_s_1_SRINV : STD_LOGIC; 
  signal romeaddro3_s_1_CLKINV : STD_LOGIC; 
  signal romeaddro3_s_1_CEINV : STD_LOGIC; 
  signal romeaddro3_s_3_DXMUX : STD_LOGIC; 
  signal romeaddro3_s_3_DYMUX : STD_LOGIC; 
  signal romeaddro3_s_3_SRINV : STD_LOGIC; 
  signal romeaddro3_s_3_CLKINV : STD_LOGIC; 
  signal romeaddro3_s_3_CEINV : STD_LOGIC; 
  signal romeaddro4_s_1_DXMUX : STD_LOGIC; 
  signal romeaddro4_s_1_DYMUX : STD_LOGIC; 
  signal romeaddro4_s_1_SRINV : STD_LOGIC; 
  signal romeaddro4_s_1_CLKINV : STD_LOGIC; 
  signal romeaddro4_s_1_CEINV : STD_LOGIC; 
  signal romeaddro4_s_3_DXMUX : STD_LOGIC; 
  signal romeaddro4_s_3_DYMUX : STD_LOGIC; 
  signal romeaddro4_s_3_SRINV : STD_LOGIC; 
  signal romeaddro4_s_3_CLKINV : STD_LOGIC; 
  signal romeaddro4_s_3_CEINV : STD_LOGIC; 
  signal romeaddro5_s_1_DXMUX : STD_LOGIC; 
  signal romeaddro5_s_1_DYMUX : STD_LOGIC; 
  signal romeaddro5_s_1_SRINV : STD_LOGIC; 
  signal romeaddro5_s_1_CLKINV : STD_LOGIC; 
  signal romeaddro5_s_1_CEINV : STD_LOGIC; 
  signal romeaddro5_s_3_DXMUX : STD_LOGIC; 
  signal romeaddro5_s_3_DYMUX : STD_LOGIC; 
  signal romeaddro5_s_3_SRINV : STD_LOGIC; 
  signal romeaddro5_s_3_CLKINV : STD_LOGIC; 
  signal romeaddro5_s_3_CEINV : STD_LOGIC; 
  signal romo2addro10_s_1_DXMUX : STD_LOGIC; 
  signal romo2addro10_s_1_DYMUX : STD_LOGIC; 
  signal romo2addro10_s_1_SRINV : STD_LOGIC; 
  signal romo2addro10_s_1_CLKINV : STD_LOGIC; 
  signal romo2addro10_s_1_CEINV : STD_LOGIC; 
  signal romeaddro6_s_1_DXMUX : STD_LOGIC; 
  signal romeaddro6_s_1_DYMUX : STD_LOGIC; 
  signal romeaddro6_s_1_SRINV : STD_LOGIC; 
  signal romeaddro6_s_1_CLKINV : STD_LOGIC; 
  signal romeaddro6_s_1_CEINV : STD_LOGIC; 
  signal romo2addro10_s_3_DXMUX : STD_LOGIC; 
  signal romo2addro10_s_3_DYMUX : STD_LOGIC; 
  signal romo2addro10_s_3_SRINV : STD_LOGIC; 
  signal romo2addro10_s_3_CLKINV : STD_LOGIC; 
  signal romo2addro10_s_3_CEINV : STD_LOGIC; 
  signal romeaddro6_s_3_DXMUX : STD_LOGIC; 
  signal romeaddro6_s_3_DYMUX : STD_LOGIC; 
  signal romeaddro6_s_3_SRINV : STD_LOGIC; 
  signal romeaddro6_s_3_CLKINV : STD_LOGIC; 
  signal romeaddro6_s_3_CEINV : STD_LOGIC; 
  signal romo2addro0_s_5_DXMUX : STD_LOGIC; 
  signal romo2addro0_s_5_DYMUX : STD_LOGIC; 
  signal romo2addro0_s_5_SRINV : STD_LOGIC; 
  signal romo2addro0_s_5_CLKINV : STD_LOGIC; 
  signal romo2addro0_s_5_CEINV : STD_LOGIC; 
  signal romeaddro7_s_1_DXMUX : STD_LOGIC; 
  signal romeaddro7_s_1_DYMUX : STD_LOGIC; 
  signal romeaddro7_s_1_SRINV : STD_LOGIC; 
  signal romeaddro7_s_1_CLKINV : STD_LOGIC; 
  signal romeaddro7_s_1_CEINV : STD_LOGIC; 
  signal romeaddro7_s_3_DXMUX : STD_LOGIC; 
  signal romeaddro7_s_3_DYMUX : STD_LOGIC; 
  signal romeaddro7_s_3_SRINV : STD_LOGIC; 
  signal romeaddro7_s_3_CLKINV : STD_LOGIC; 
  signal romeaddro7_s_3_CEINV : STD_LOGIC; 
  signal romeaddro8_s_1_DXMUX : STD_LOGIC; 
  signal romeaddro8_s_1_DYMUX : STD_LOGIC; 
  signal romeaddro8_s_1_SRINV : STD_LOGIC; 
  signal romeaddro8_s_1_CLKINV : STD_LOGIC; 
  signal romeaddro8_s_1_CEINV : STD_LOGIC; 
  signal romeaddro8_s_3_DXMUX : STD_LOGIC; 
  signal romeaddro8_s_3_DYMUX : STD_LOGIC; 
  signal romeaddro8_s_3_SRINV : STD_LOGIC; 
  signal romeaddro8_s_3_CLKINV : STD_LOGIC; 
  signal romeaddro8_s_3_CEINV : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1854_F : STD_LOGIC; 
  signal U_DCT2D_rtlc5n1854_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z1_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z253_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z5_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z78_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z79_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z42_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z572_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z572_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z583_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z296_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z586_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z215_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z215_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z297_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z121_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z595_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z604_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z580_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z589_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z598_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z607_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z413_G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_nx65206z592_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z224_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z601_F : STD_LOGIC; 
  signal U_DCT2D_nx65206z233_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z221_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z230_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z239_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z227_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z334_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z248_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z236_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z245_G : STD_LOGIC; 
  signal U_DCT2D_nx65206z242_G : STD_LOGIC; 
  signal requestrd_s_DYMUX : STD_LOGIC; 
  signal requestrd_s_BYINVNOT : STD_LOGIC; 
  signal requestrd_s_CLKINV : STD_LOGIC; 
  signal requestrd_s_CEINV : STD_LOGIC; 
  signal U_DCT2D_rtlc2n446_F : STD_LOGIC; 
  signal U_DCT2D_rtlc2n446_G : STD_LOGIC; 
  signal U_DCT2D_nx40895z2_F : STD_LOGIC; 
  signal U_DCT2D_nx40895z2_G : STD_LOGIC; 
  signal U_DCT1D_nx52393z1_F : STD_LOGIC; 
  signal U_DCT1D_nx52393z1_G : STD_LOGIC; 
  signal U_DCT1D_rtlc2n293_F : STD_LOGIC; 
  signal U_DCT1D_rtlc2n293_G : STD_LOGIC; 
  signal U_DCT1D_rtlc2n468_F : STD_LOGIC; 
  signal U_DCT1D_rtlc2n468_G : STD_LOGIC; 
  signal U_DCT2D_colram_reg_3_DYMUX : STD_LOGIC; 
  signal U_DCT2D_colram_reg_3_BYINVNOT : STD_LOGIC; 
  signal U_DCT2D_colram_reg_3_CLKINV : STD_LOGIC; 
  signal U_DCT2D_colram_reg_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1558_F : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1558_G : STD_LOGIC; 
  signal releasewr_s_DYMUX : STD_LOGIC; 
  signal releasewr_s_CLKINV : STD_LOGIC; 
  signal releasewr_s_CEINV : STD_LOGIC; 
  signal U_DCT1D_latch_done_reg_DYMUX : STD_LOGIC; 
  signal U_DCT1D_latch_done_reg_BYINVNOT : STD_LOGIC; 
  signal U_DCT1D_latch_done_reg_CLKINV : STD_LOGIC; 
  signal U_DCT1D_latch_done_reg_CEINV : STD_LOGIC; 
  signal U_DCT1D_NOT_rtlcs2_F : STD_LOGIC; 
  signal U_DCT1D_NOT_rtlcs2_G : STD_LOGIC; 
  signal U_DCT1D_nx62663z1_F : STD_LOGIC; 
  signal U_DCT1D_nx62663z1_G : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1612_F : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1612_G : STD_LOGIC; 
  signal U_DCT2D_completed_reg_DYMUX : STD_LOGIC; 
  signal U_DCT2D_completed_reg_BYINVNOT : STD_LOGIC; 
  signal U_DCT2D_completed_reg_CLKINV : STD_LOGIC; 
  signal U_DCT2D_completed_reg_CEINV : STD_LOGIC; 
  signal U_DCT2D_col_tmp_reg_1_DXMUX : STD_LOGIC; 
  signal U_DCT2D_col_tmp_reg_1_BXINVNOT : STD_LOGIC; 
  signal U_DCT2D_col_tmp_reg_1_DYMUX : STD_LOGIC; 
  signal U_DCT2D_col_tmp_reg_1_SRINV : STD_LOGIC; 
  signal U_DCT2D_col_tmp_reg_1_CLKINV : STD_LOGIC; 
  signal U_DCT2D_col_tmp_reg_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_nx57528z1_F : STD_LOGIC; 
  signal U_DCT1D_nx57528z1_G : STD_LOGIC; 
  signal ramwaddro_s_1_DXMUX : STD_LOGIC; 
  signal ramwaddro_s_1_DYMUX : STD_LOGIC; 
  signal ramwaddro_s_1_SRINV : STD_LOGIC; 
  signal ramwaddro_s_1_CLKINV : STD_LOGIC; 
  signal ramwaddro_s_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_4_FFX_RST : STD_LOGIC; 
  signal ramwaddro_s_3_DXMUX : STD_LOGIC; 
  signal ramwaddro_s_3_DYMUX : STD_LOGIC; 
  signal ramwaddro_s_3_SRINV : STD_LOGIC; 
  signal ramwaddro_s_3_CLKINV : STD_LOGIC; 
  signal ramwaddro_s_3_CEINV : STD_LOGIC; 
  signal ramwaddro_s_5_DXMUX : STD_LOGIC; 
  signal ramwaddro_s_5_DYMUX : STD_LOGIC; 
  signal ramwaddro_s_5_SRINV : STD_LOGIC; 
  signal ramwaddro_s_5_CLKINV : STD_LOGIC; 
  signal ramwaddro_s_5_CEINV : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_0_DXMUX : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_0_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_0_DYMUX : STD_LOGIC; 
  signal U_DCT1D_nx58996z1 : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_0_SRINV : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_0_CLKINV : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_0_CEINV : STD_LOGIC; 
  signal ramwe_s_DYMUX : STD_LOGIC; 
  signal ramwe_s_CLKINV : STD_LOGIC; 
  signal ramwe_s_CEINV : STD_LOGIC; 
  signal rome2addro0_s_1_DXMUX : STD_LOGIC; 
  signal rome2addro0_s_1_DYMUX : STD_LOGIC; 
  signal rome2addro0_s_1_SRINV : STD_LOGIC; 
  signal rome2addro0_s_1_CLKINV : STD_LOGIC; 
  signal rome2addro0_s_1_CEINV : STD_LOGIC; 
  signal rome2addro0_s_3_DXMUX : STD_LOGIC; 
  signal rome2addro0_s_3_DYMUX : STD_LOGIC; 
  signal rome2addro0_s_3_SRINV : STD_LOGIC; 
  signal rome2addro0_s_3_CLKINV : STD_LOGIC; 
  signal rome2addro0_s_3_CEINV : STD_LOGIC; 
  signal rome2addro1_s_1_DXMUX : STD_LOGIC; 
  signal rome2addro1_s_1_DYMUX : STD_LOGIC; 
  signal rome2addro1_s_1_SRINV : STD_LOGIC; 
  signal rome2addro1_s_1_CLKINV : STD_LOGIC; 
  signal rome2addro1_s_1_CEINV : STD_LOGIC; 
  signal rome2addro1_s_3_DXMUX : STD_LOGIC; 
  signal rome2addro1_s_3_DYMUX : STD_LOGIC; 
  signal rome2addro1_s_3_SRINV : STD_LOGIC; 
  signal rome2addro1_s_3_CLKINV : STD_LOGIC; 
  signal rome2addro1_s_3_CEINV : STD_LOGIC; 
  signal rome2addro2_s_1_DXMUX : STD_LOGIC; 
  signal rome2addro2_s_1_DYMUX : STD_LOGIC; 
  signal rome2addro2_s_1_SRINV : STD_LOGIC; 
  signal rome2addro2_s_1_CLKINV : STD_LOGIC; 
  signal rome2addro2_s_1_CEINV : STD_LOGIC; 
  signal rome2addro2_s_3_DXMUX : STD_LOGIC; 
  signal rome2addro2_s_3_DYMUX : STD_LOGIC; 
  signal rome2addro2_s_3_SRINV : STD_LOGIC; 
  signal rome2addro2_s_3_CLKINV : STD_LOGIC; 
  signal rome2addro2_s_3_CEINV : STD_LOGIC; 
  signal rome2addro3_s_1_DXMUX : STD_LOGIC; 
  signal rome2addro3_s_1_DYMUX : STD_LOGIC; 
  signal rome2addro3_s_1_SRINV : STD_LOGIC; 
  signal rome2addro3_s_1_CLKINV : STD_LOGIC; 
  signal rome2addro3_s_1_CEINV : STD_LOGIC; 
  signal rome2addro3_s_3_DXMUX : STD_LOGIC; 
  signal rome2addro3_s_3_DYMUX : STD_LOGIC; 
  signal rome2addro3_s_3_SRINV : STD_LOGIC; 
  signal rome2addro3_s_3_CLKINV : STD_LOGIC; 
  signal rome2addro3_s_3_CEINV : STD_LOGIC; 
  signal rome2addro4_s_1_DXMUX : STD_LOGIC; 
  signal rome2addro4_s_1_DYMUX : STD_LOGIC; 
  signal rome2addro4_s_1_SRINV : STD_LOGIC; 
  signal rome2addro4_s_1_CLKINV : STD_LOGIC; 
  signal rome2addro4_s_1_CEINV : STD_LOGIC; 
  signal rome2addro4_s_3_DXMUX : STD_LOGIC; 
  signal rome2addro4_s_3_DYMUX : STD_LOGIC; 
  signal rome2addro4_s_3_SRINV : STD_LOGIC; 
  signal rome2addro4_s_3_CLKINV : STD_LOGIC; 
  signal rome2addro4_s_3_CEINV : STD_LOGIC; 
  signal rome2addro5_s_1_DXMUX : STD_LOGIC; 
  signal rome2addro5_s_1_DYMUX : STD_LOGIC; 
  signal rome2addro5_s_1_SRINV : STD_LOGIC; 
  signal rome2addro5_s_1_CLKINV : STD_LOGIC; 
  signal rome2addro5_s_1_CEINV : STD_LOGIC; 
  signal rome2addro5_s_3_DXMUX : STD_LOGIC; 
  signal rome2addro5_s_3_DYMUX : STD_LOGIC; 
  signal rome2addro5_s_3_SRINV : STD_LOGIC; 
  signal rome2addro5_s_3_CLKINV : STD_LOGIC; 
  signal rome2addro5_s_3_CEINV : STD_LOGIC; 
  signal rome2addro6_s_1_DXMUX : STD_LOGIC; 
  signal rome2addro6_s_1_DYMUX : STD_LOGIC; 
  signal rome2addro6_s_1_SRINV : STD_LOGIC; 
  signal rome2addro6_s_1_CLKINV : STD_LOGIC; 
  signal rome2addro6_s_1_CEINV : STD_LOGIC; 
  signal rome2addro6_s_3_DXMUX : STD_LOGIC; 
  signal rome2addro6_s_3_DYMUX : STD_LOGIC; 
  signal rome2addro6_s_3_SRINV : STD_LOGIC; 
  signal rome2addro6_s_3_CLKINV : STD_LOGIC; 
  signal rome2addro6_s_3_CEINV : STD_LOGIC; 
  signal rome2addro7_s_1_DXMUX : STD_LOGIC; 
  signal rome2addro7_s_1_DYMUX : STD_LOGIC; 
  signal rome2addro7_s_1_SRINV : STD_LOGIC; 
  signal rome2addro7_s_1_CLKINV : STD_LOGIC; 
  signal rome2addro7_s_1_CEINV : STD_LOGIC; 
  signal rome2addro7_s_3_DXMUX : STD_LOGIC; 
  signal rome2addro7_s_3_DYMUX : STD_LOGIC; 
  signal rome2addro7_s_3_SRINV : STD_LOGIC; 
  signal rome2addro7_s_3_CLKINV : STD_LOGIC; 
  signal rome2addro7_s_3_CEINV : STD_LOGIC; 
  signal rome2addro8_s_1_DXMUX : STD_LOGIC; 
  signal rome2addro8_s_1_DYMUX : STD_LOGIC; 
  signal rome2addro8_s_1_SRINV : STD_LOGIC; 
  signal rome2addro8_s_1_CLKINV : STD_LOGIC; 
  signal rome2addro8_s_1_CEINV : STD_LOGIC; 
  signal rome2addro8_s_3_DXMUX : STD_LOGIC; 
  signal rome2addro8_s_3_DYMUX : STD_LOGIC; 
  signal rome2addro8_s_3_SRINV : STD_LOGIC; 
  signal rome2addro8_s_3_CLKINV : STD_LOGIC; 
  signal rome2addro8_s_3_CEINV : STD_LOGIC; 
  signal rome2addro9_s_1_DXMUX : STD_LOGIC; 
  signal rome2addro9_s_1_DYMUX : STD_LOGIC; 
  signal rome2addro9_s_1_SRINV : STD_LOGIC; 
  signal rome2addro9_s_1_CLKINV : STD_LOGIC; 
  signal rome2addro9_s_1_CEINV : STD_LOGIC; 
  signal rome2addro9_s_3_DXMUX : STD_LOGIC; 
  signal rome2addro9_s_3_DYMUX : STD_LOGIC; 
  signal rome2addro9_s_3_SRINV : STD_LOGIC; 
  signal rome2addro9_s_3_CLKINV : STD_LOGIC; 
  signal rome2addro9_s_3_CEINV : STD_LOGIC; 
  signal U_DCT1D_rtlc2n471_F : STD_LOGIC; 
  signal U_DCT1D_rtlc2n471_G : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_1_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_1_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_1_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_1_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_1_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_3_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_3_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_3_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_3_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_3_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_5_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_5_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_5_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_5_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_5_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_7_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_7_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_7_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_7_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_7_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_10_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_10_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_10_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_1_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_1_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_1_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_1_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_1_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_3_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_3_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_3_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_3_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_3_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_5_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_5_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_5_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_5_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_5_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_7_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_7_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_7_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_7_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_7_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_10_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_10_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_10_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_1_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_1_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_1_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_1_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_1_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_3_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_3_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_3_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_3_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_3_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_5_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_5_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_5_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_5_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_5_CEINV : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_7_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_7_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_7_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_7_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_7_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_10_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_10_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_10_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_1_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_1_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_1_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_1_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_1_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_3_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_3_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_3_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_3_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_3_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_5_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_5_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_5_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_5_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_5_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_7_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_7_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_7_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_7_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_7_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_10_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_10_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_10_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_1_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_1_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_1_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_1_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_1_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_3_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_3_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_3_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_3_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_3_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_5_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_5_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_5_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_5_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_5_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_7_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_7_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_7_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_7_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_7_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_10_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_10_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_10_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_1_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_1_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_1_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_1_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_1_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_3_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_3_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_3_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_3_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_3_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_5_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_5_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_5_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_5_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_5_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_7_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_7_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_7_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_7_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_7_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_10_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_10_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_10_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_1_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_1_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_1_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_1_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_1_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_3_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_3_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_3_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_3_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_3_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_5_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_5_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_5_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_5_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_5_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_7_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_7_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_7_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_7_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_7_CEINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_10_DXMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_10_DYMUX : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_10_SRINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_10_CLKINV : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_10_CEINV : STD_LOGIC; 
  signal U_DCT1D_rtlc5n1685_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z303_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z303_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z1_G : STD_LOGIC; 
  signal U_DCT1D_col_tmp_reg_1_DXMUX : STD_LOGIC; 
  signal U_DCT1D_col_tmp_reg_1_BXINVNOT : STD_LOGIC; 
  signal U_DCT1D_col_tmp_reg_1_DYMUX : STD_LOGIC; 
  signal U_DCT1D_col_tmp_reg_1_SRINV : STD_LOGIC; 
  signal U_DCT1D_col_tmp_reg_1_CLKINV : STD_LOGIC; 
  signal U_DCT1D_col_tmp_reg_1_CEINV : STD_LOGIC; 
  signal U_DCT1D_nx59700z333_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z333_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z251_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z251_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z218_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z218_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z348_F : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_6_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_nx59700z357_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z366_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z342_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z351_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z360_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z369_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z345_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z354_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z363_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z5_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z78_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z79_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z42_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z215_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z215_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z121_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z224_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z233_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z221_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z230_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z306_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z300_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z255_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z239_G : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_8_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_1_8_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT1D_nx59700z227_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z248_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z236_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z321_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z315_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z309_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z245_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z242_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z330_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z324_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z318_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z312_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z327_G : STD_LOGIC; 
  signal U_DCT1D_nx59700z334_F : STD_LOGIC; 
  signal U_DCT1D_nx59700z334_G : STD_LOGIC; 
  signal releaserd_s_DYMUX : STD_LOGIC; 
  signal releaserd_s_BYINVNOT : STD_LOGIC; 
  signal releaserd_s_CLKINV : STD_LOGIC; 
  signal releaserd_s_CEINV : STD_LOGIC; 
  signal romoaddro0_s_1_DXMUX : STD_LOGIC; 
  signal romoaddro0_s_1_DYMUX : STD_LOGIC; 
  signal romoaddro0_s_1_SRINV : STD_LOGIC; 
  signal romoaddro0_s_1_CLKINV : STD_LOGIC; 
  signal romoaddro0_s_1_CEINV : STD_LOGIC; 
  signal romoaddro0_s_3_DXMUX : STD_LOGIC; 
  signal romoaddro0_s_3_DYMUX : STD_LOGIC; 
  signal romoaddro0_s_3_SRINV : STD_LOGIC; 
  signal romoaddro0_s_3_CLKINV : STD_LOGIC; 
  signal romoaddro0_s_3_CEINV : STD_LOGIC; 
  signal romoaddro1_s_1_DXMUX : STD_LOGIC; 
  signal romoaddro1_s_1_DYMUX : STD_LOGIC; 
  signal romoaddro1_s_1_SRINV : STD_LOGIC; 
  signal romoaddro1_s_1_CLKINV : STD_LOGIC; 
  signal romoaddro1_s_1_CEINV : STD_LOGIC; 
  signal romoaddro1_s_3_DXMUX : STD_LOGIC; 
  signal romoaddro1_s_3_DYMUX : STD_LOGIC; 
  signal romoaddro1_s_3_SRINV : STD_LOGIC; 
  signal romoaddro1_s_3_CLKINV : STD_LOGIC; 
  signal romoaddro1_s_3_CEINV : STD_LOGIC; 
  signal romoaddro2_s_1_DXMUX : STD_LOGIC; 
  signal romoaddro2_s_1_DYMUX : STD_LOGIC; 
  signal romoaddro2_s_1_SRINV : STD_LOGIC; 
  signal romoaddro2_s_1_CLKINV : STD_LOGIC; 
  signal romoaddro2_s_1_CEINV : STD_LOGIC; 
  signal romoaddro2_s_3_DXMUX : STD_LOGIC; 
  signal romoaddro2_s_3_DYMUX : STD_LOGIC; 
  signal romoaddro2_s_3_SRINV : STD_LOGIC; 
  signal romoaddro2_s_3_CLKINV : STD_LOGIC; 
  signal romoaddro2_s_3_CEINV : STD_LOGIC; 
  signal romoaddro3_s_1_DXMUX : STD_LOGIC; 
  signal romoaddro3_s_1_DYMUX : STD_LOGIC; 
  signal romoaddro3_s_1_SRINV : STD_LOGIC; 
  signal romoaddro3_s_1_CLKINV : STD_LOGIC; 
  signal romoaddro3_s_1_CEINV : STD_LOGIC; 
  signal romoaddro3_s_3_DXMUX : STD_LOGIC; 
  signal romoaddro3_s_3_DYMUX : STD_LOGIC; 
  signal romoaddro3_s_3_SRINV : STD_LOGIC; 
  signal romoaddro3_s_3_CLKINV : STD_LOGIC; 
  signal romoaddro3_s_3_CEINV : STD_LOGIC; 
  signal romoaddro4_s_1_DXMUX : STD_LOGIC; 
  signal romoaddro4_s_1_DYMUX : STD_LOGIC; 
  signal romoaddro4_s_1_SRINV : STD_LOGIC; 
  signal romoaddro4_s_1_CLKINV : STD_LOGIC; 
  signal romoaddro4_s_1_CEINV : STD_LOGIC; 
  signal romoaddro4_s_3_DXMUX : STD_LOGIC; 
  signal romoaddro4_s_3_DYMUX : STD_LOGIC; 
  signal romoaddro4_s_3_SRINV : STD_LOGIC; 
  signal romoaddro4_s_3_CLKINV : STD_LOGIC; 
  signal romoaddro4_s_3_CEINV : STD_LOGIC; 
  signal romoaddro5_s_1_DXMUX : STD_LOGIC; 
  signal romoaddro5_s_1_DYMUX : STD_LOGIC; 
  signal romoaddro5_s_1_SRINV : STD_LOGIC; 
  signal romoaddro5_s_1_CLKINV : STD_LOGIC; 
  signal romoaddro5_s_1_CEINV : STD_LOGIC; 
  signal romoaddro5_s_3_DXMUX : STD_LOGIC; 
  signal romoaddro5_s_3_DYMUX : STD_LOGIC; 
  signal romoaddro5_s_3_SRINV : STD_LOGIC; 
  signal romoaddro5_s_3_CLKINV : STD_LOGIC; 
  signal romoaddro5_s_3_CEINV : STD_LOGIC; 
  signal romoaddro6_s_1_DXMUX : STD_LOGIC; 
  signal romoaddro6_s_1_DYMUX : STD_LOGIC; 
  signal romoaddro6_s_1_SRINV : STD_LOGIC; 
  signal romoaddro6_s_1_CLKINV : STD_LOGIC; 
  signal romoaddro6_s_1_CEINV : STD_LOGIC; 
  signal romoaddro6_s_3_DXMUX : STD_LOGIC; 
  signal romoaddro6_s_3_DYMUX : STD_LOGIC; 
  signal romoaddro6_s_3_SRINV : STD_LOGIC; 
  signal romoaddro6_s_3_CLKINV : STD_LOGIC; 
  signal romoaddro6_s_3_CEINV : STD_LOGIC; 
  signal romoaddro7_s_1_DXMUX : STD_LOGIC; 
  signal romoaddro7_s_1_DYMUX : STD_LOGIC; 
  signal romoaddro7_s_1_SRINV : STD_LOGIC; 
  signal romoaddro7_s_1_CLKINV : STD_LOGIC; 
  signal romoaddro7_s_1_CEINV : STD_LOGIC; 
  signal romoaddro7_s_3_DXMUX : STD_LOGIC; 
  signal romoaddro7_s_3_DYMUX : STD_LOGIC; 
  signal romoaddro7_s_3_SRINV : STD_LOGIC; 
  signal romoaddro7_s_3_CLKINV : STD_LOGIC; 
  signal romoaddro7_s_3_CEINV : STD_LOGIC; 
  signal romoaddro8_s_1_DXMUX : STD_LOGIC; 
  signal romoaddro8_s_1_DYMUX : STD_LOGIC; 
  signal romoaddro8_s_1_SRINV : STD_LOGIC; 
  signal romoaddro8_s_1_CLKINV : STD_LOGIC; 
  signal romoaddro8_s_1_CEINV : STD_LOGIC; 
  signal romoaddro8_s_3_DXMUX : STD_LOGIC; 
  signal romoaddro8_s_3_DYMUX : STD_LOGIC; 
  signal romoaddro8_s_3_SRINV : STD_LOGIC; 
  signal romoaddro8_s_3_CLKINV : STD_LOGIC; 
  signal romoaddro8_s_3_CEINV : STD_LOGIC; 
  signal romoaddro0_s_5_DXMUX : STD_LOGIC; 
  signal romoaddro0_s_5_DYMUX : STD_LOGIC; 
  signal romoaddro0_s_5_SRINV : STD_LOGIC; 
  signal romoaddro0_s_5_CLKINV : STD_LOGIC; 
  signal romoaddro0_s_5_CEINV : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_8_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_10_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_4_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_4_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_1_0_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_0_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_2_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_4_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_6_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_8_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_8_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_8_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_10_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_8_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_8_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_2_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_0_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_4_2_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_6_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_0_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_2_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_0_6_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_6_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_8_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_7_8_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_0_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_2_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_4_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_8_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_8_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_8_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_0_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_6_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_8_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_8_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_6_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_10_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_0_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_6_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_8_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_10_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_3_4_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_0_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_8_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_10_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_0_0_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_2_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_6_4_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_2_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_5_4_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_4_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_6_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_6_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_8_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_8_FFX_RSTAND : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_4_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_6_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_databuf_reg_5_2_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_3_2_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_0_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_2_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_databuf_reg_6_4_FFX_RST : STD_LOGIC; 
  signal ramdatai_s_4_FFY_RST : STD_LOGIC; 
  signal ramdatai_s_4_FFX_RST : STD_LOGIC; 
  signal ramdatai_s_0_FFY_RST : STD_LOGIC; 
  signal ramdatai_s_6_FFY_RST : STD_LOGIC; 
  signal ramdatai_s_6_FFX_RST : STD_LOGIC; 
  signal ramdatai_s_8_FFY_RST : STD_LOGIC; 
  signal ramdatai_s_8_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_5_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_7_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_7_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_1_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_3_FFY_RST : STD_LOGIC; 
  signal romo2addro5_s_1_FFY_RST : STD_LOGIC; 
  signal romo2addro5_s_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_3_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_3_FFX_RST : STD_LOGIC; 
  signal romo2addro5_s_3_FFY_RST : STD_LOGIC; 
  signal romo2addro5_s_3_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_5_FFY_RST : STD_LOGIC; 
  signal odv1_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal ramwe_repl0 : STD_LOGIC; 
  signal odv1_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal odv1_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal odv1_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal odv1_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcti_0_IFF_IFF1_RST : STD_LOGIC; 
  signal dcti_0_IFF_ISR_USED : STD_LOGIC; 
  signal dcti_0_IFF_ICLK1INV : STD_LOGIC; 
  signal dcti_0_IFF_ICEINV : STD_LOGIC; 
  signal dcti_0_IFF_IFFDMUX : STD_LOGIC; 
  signal dcti_1_IFF_ICLK1INV : STD_LOGIC; 
  signal dcti_1_IFF_ICEINV : STD_LOGIC; 
  signal dcti_1_IFF_IFFDMUX : STD_LOGIC; 
  signal dcti_1_IFF_IFF1_RST : STD_LOGIC; 
  signal dcti_1_IFF_IFF1_RSTAND : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_3_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_5_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_5_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_7_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_7_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_10_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_10_FFX_RST : STD_LOGIC; 
  signal ready_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal ready_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal ready_repl0 : STD_LOGIC; 
  signal ready_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal ready_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal ready_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto_10_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto_10_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto_10_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto_10_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto_10_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto_11_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto_11_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto_11_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto_11_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto_11_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto_4_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto_4_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto_4_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto_4_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto_4_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto_5_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto_5_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto_5_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto_5_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto_5_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto_6_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto_6_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto_6_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto_6_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto_6_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto1_10_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto1_10_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal ramdatai_9_repl1 : STD_LOGIC; 
  signal dcto1_10_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto1_10_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto1_10_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal U_DCT1D_istate_reg_1_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_istate_reg_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_2_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_2_FFY_RSTAND : STD_LOGIC; 
  signal reqrdfail_s_FFY_RST : STD_LOGIC; 
  signal reqrdfail_s_FFY_RSTAND : STD_LOGIC; 
  signal dcto_1_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto_1_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto_1_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto_1_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto_1_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto_2_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto_2_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto_2_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto_2_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto_2_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto_3_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto_3_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto_3_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto_3_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto_3_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcti_6_IFF_ICLK1INV : STD_LOGIC; 
  signal dcti_6_IFF_ICEINV : STD_LOGIC; 
  signal dcti_6_IFF_IFFDMUX : STD_LOGIC; 
  signal dcti_6_IFF_IFF1_RST : STD_LOGIC; 
  signal dcti_6_IFF_IFF1_RSTAND : STD_LOGIC; 
  signal dcto_0_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto_0_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto_0_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto_0_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto_0_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal rome2addro1_s_1_FFY_RST : STD_LOGIC; 
  signal rome2addro1_s_1_FFX_RST : STD_LOGIC; 
  signal rome2addro1_s_3_FFY_RST : STD_LOGIC; 
  signal rome2addro1_s_3_FFX_RST : STD_LOGIC; 
  signal rome2addro2_s_1_FFY_RST : STD_LOGIC; 
  signal rome2addro2_s_1_FFX_RST : STD_LOGIC; 
  signal dcto1_11_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto1_11_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal ramdatai_9_repl2 : STD_LOGIC; 
  signal dcto1_11_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto1_11_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto1_11_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal odv_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal odv_dup0 : STD_LOGIC; 
  signal odv_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal odv_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal odv_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal odv_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto1_0_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto1_0_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal ramdatai_0_repl0 : STD_LOGIC; 
  signal dcto1_0_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto1_0_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto1_0_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto1_1_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto1_1_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal ramdatai_1_repl0 : STD_LOGIC; 
  signal dcto1_1_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto1_1_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto1_1_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto1_2_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto1_2_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal ramdatai_2_repl0 : STD_LOGIC; 
  signal dcto1_2_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto1_2_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto1_2_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcti_2_IFF_ICLK1INV : STD_LOGIC; 
  signal dcti_2_IFF_ICEINV : STD_LOGIC; 
  signal dcti_2_IFF_IFFDMUX : STD_LOGIC; 
  signal dcti_2_IFF_IFF1_RST : STD_LOGIC; 
  signal dcti_2_IFF_IFF1_RSTAND : STD_LOGIC; 
  signal dcti_3_IFF_ICLK1INV : STD_LOGIC; 
  signal dcti_3_IFF_ICEINV : STD_LOGIC; 
  signal dcti_3_IFF_IFFDMUX : STD_LOGIC; 
  signal dcti_3_IFF_IFF1_RST : STD_LOGIC; 
  signal dcti_3_IFF_IFF1_RSTAND : STD_LOGIC; 
  signal dcti_5_IFF_IFF1_RST : STD_LOGIC; 
  signal dcti_5_IFF_ISR_USED : STD_LOGIC; 
  signal dcti_5_IFF_ICLK1INV : STD_LOGIC; 
  signal dcti_5_IFF_ICEINV : STD_LOGIC; 
  signal dcti_5_IFF_IFFDMUX : STD_LOGIC; 
  signal dcti_4_IFF_ICLK1INV : STD_LOGIC; 
  signal dcti_4_IFF_ICEINV : STD_LOGIC; 
  signal dcti_4_IFF_IFFDMUX : STD_LOGIC; 
  signal dcti_4_IFF_IFF1_RST : STD_LOGIC; 
  signal dcti_4_IFF_IFF1_RSTAND : STD_LOGIC; 
  signal dcto_7_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto_7_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto_7_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto_7_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto_7_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto_8_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto_8_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto_8_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto_8_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto_8_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto_9_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto_9_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto_9_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto_9_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto_9_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto1_3_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto1_3_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal ramdatai_3_repl0 : STD_LOGIC; 
  signal dcto1_3_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto1_3_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto1_3_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto1_4_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto1_4_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal ramdatai_4_repl0 : STD_LOGIC; 
  signal dcto1_4_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto1_4_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto1_4_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto1_5_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto1_5_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal ramdatai_5_repl0 : STD_LOGIC; 
  signal dcto1_5_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto1_9_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto1_9_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal ramdatai_9_repl0 : STD_LOGIC; 
  signal dcto1_9_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto1_9_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto1_9_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto1_5_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto1_5_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto1_6_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto1_6_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal ramdatai_6_repl0 : STD_LOGIC; 
  signal dcto1_6_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto1_6_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto1_6_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto1_7_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto1_7_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal ramdatai_7_repl0 : STD_LOGIC; 
  signal dcto1_7_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal dcto1_7_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto1_7_OUTPUT_OFF_OFF1_RSTAND : STD_LOGIC; 
  signal dcto1_8_OUTPUT_OFF_OFF1_RST : STD_LOGIC; 
  signal dcto1_8_OUTPUT_OFF_O1INV : STD_LOGIC; 
  signal dcto1_8_OUTPUT_OFF_OCEINV : STD_LOGIC; 
  signal dcto1_8_OUTPUT_OFF_OSR_USED : STD_LOGIC; 
  signal ramdatai_8_repl0 : STD_LOGIC; 
  signal dcto1_8_OUTPUT_OTCLK1INV : STD_LOGIC; 
  signal U_DCT2D_istate_reg_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_istate_reg_1_FFX_RST : STD_LOGIC; 
  signal memswitchrd_s_FFX_RST : STD_LOGIC; 
  signal memswitchrd_s_FFX_RSTAND : STD_LOGIC; 
  signal ramraddro_s_5_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_col_reg_0_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_col_reg_0_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_col_reg_0_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_5_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_5_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_7_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_7_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_col_reg_2_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_col_reg_2_FFY_RSTAND : STD_LOGIC; 
  signal U_DCT1D_col_reg_2_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_col_reg_2_FFY_RSTAND : STD_LOGIC; 
  signal U_DCT1D_ready_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_ready_FFY_RSTAND : STD_LOGIC; 
  signal ramraddro_s_5_FFX_RST : STD_LOGIC; 
  signal memswitchwr_s_FFY_RST : STD_LOGIC; 
  signal memswitchwr_s_FFY_RSTAND : STD_LOGIC; 
  signal U_DBUFCTL_mem1_full_reg_FFY_RST : STD_LOGIC; 
  signal U_DBUFCTL_mem1_full_reg_FFY_RSTAND : STD_LOGIC; 
  signal U_DCT1D_row_reg_2_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_row_reg_2_FFY_RSTAND : STD_LOGIC; 
  signal rome2addro0_s_5_FFY_RST : STD_LOGIC; 
  signal rome2addro0_s_5_FFX_RST : STD_LOGIC; 
  signal romeaddro0_s_5_FFY_RST : STD_LOGIC; 
  signal romeaddro0_s_5_FFX_RST : STD_LOGIC; 
  signal U_DBUFCTL_mem1_lock_reg_FFY_RST : STD_LOGIC; 
  signal U_DBUFCTL_mem1_lock_reg_FFY_RSTAND : STD_LOGIC; 
  signal U_DBUFCTL_mem2_full_reg_FFY_RST : STD_LOGIC; 
  signal U_DBUFCTL_mem2_full_reg_FFY_RSTAND : STD_LOGIC; 
  signal U_DBUFCTL_mem2_lock_reg_FFY_RST : STD_LOGIC; 
  signal U_DBUFCTL_mem2_lock_reg_FFY_RSTAND : STD_LOGIC; 
  signal ramraddro_s_0_FFY_RST : STD_LOGIC; 
  signal ramraddro_s_0_FFY_RSTAND : STD_LOGIC; 
  signal ramraddro_s_1_FFY_RST : STD_LOGIC; 
  signal ramraddro_s_1_FFY_RSTAND : STD_LOGIC; 
  signal ramraddro_s_2_FFY_RST : STD_LOGIC; 
  signal ramraddro_s_2_FFY_RSTAND : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_1_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_1_FFX_RST : STD_LOGIC; 
  signal romo2addro3_s_1_FFY_RST : STD_LOGIC; 
  signal romo2addro3_s_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_3_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_3_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_10_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_10_FFX_RST : STD_LOGIC; 
  signal ramraddro_s_3_FFY_RST : STD_LOGIC; 
  signal ramraddro_s_3_FFY_RSTAND : STD_LOGIC; 
  signal requestwr_s_FFY_RST : STD_LOGIC; 
  signal requestwr_s_FFY_RSTAND : STD_LOGIC; 
  signal reqwrfail_s_FFY_RST : STD_LOGIC; 
  signal reqwrfail_s_FFY_RSTAND : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_1_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_3_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_7_3_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_col_reg_0_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_completed_reg_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_completed_reg_FFY_RSTAND : STD_LOGIC; 
  signal U_DCT1D_state_reg_1_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_state_reg_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_1_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_3_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_3_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_5_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_5_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_7_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_0_7_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_1_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_3_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_3_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_1_5_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_7_FFX_RST : STD_LOGIC; 
  signal romo2addro0_s_3_FFY_RST : STD_LOGIC; 
  signal romo2addro0_s_3_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_1_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_1_FFX_RST : STD_LOGIC; 
  signal romo2addro1_s_1_FFY_RST : STD_LOGIC; 
  signal romo2addro1_s_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_3_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_3_FFX_RST : STD_LOGIC; 
  signal romo2addro1_s_3_FFY_RST : STD_LOGIC; 
  signal romo2addro1_s_3_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_5_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_5_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_3_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_5_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_5_FFX_RST : STD_LOGIC; 
  signal romo2addro0_s_1_FFY_RST : STD_LOGIC; 
  signal romo2addro0_s_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_7_FFY_RST : STD_LOGIC; 
  signal romo2addro8_s_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_7_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_7_FFX_RST : STD_LOGIC; 
  signal romo2addro8_s_3_FFY_RST : STD_LOGIC; 
  signal romo2addro8_s_3_FFX_RST : STD_LOGIC; 
  signal romo2addro9_s_1_FFY_RST : STD_LOGIC; 
  signal romo2addro2_s_1_FFY_RST : STD_LOGIC; 
  signal romo2addro2_s_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_7_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_3_7_FFX_RST : STD_LOGIC; 
  signal romo2addro2_s_3_FFY_RST : STD_LOGIC; 
  signal romo2addro2_s_3_FFX_RST : STD_LOGIC; 
  signal romo2addro3_s_3_FFY_RST : STD_LOGIC; 
  signal romo2addro3_s_3_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_5_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_5_FFX_RST : STD_LOGIC; 
  signal romo2addro4_s_1_FFY_RST : STD_LOGIC; 
  signal romo2addro4_s_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_5_FFX_RST : STD_LOGIC; 
  signal romo2addro6_s_1_FFY_RST : STD_LOGIC; 
  signal romo2addro6_s_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_7_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_7_FFX_RST : STD_LOGIC; 
  signal romo2addro6_s_3_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_7_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_4_7_FFX_RST : STD_LOGIC; 
  signal romo2addro4_s_3_FFY_RST : STD_LOGIC; 
  signal romo2addro4_s_3_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_1_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_5_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_3_FFX_RST : STD_LOGIC; 
  signal romo2addro7_s_3_FFY_RST : STD_LOGIC; 
  signal romo2addro7_s_3_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_5_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_5_FFX_RST : STD_LOGIC; 
  signal romo2addro8_s_1_FFY_RST : STD_LOGIC; 
  signal romo2addro9_s_1_FFX_RST : STD_LOGIC; 
  signal romo2addro9_s_3_FFY_RST : STD_LOGIC; 
  signal romo2addro9_s_3_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_7_7_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_7_7_FFY_RSTAND : STD_LOGIC; 
  signal U_DCT2D_latch_done_reg_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latch_done_reg_FFY_RSTAND : STD_LOGIC; 
  signal romeaddro6_s_3_FFX_RST : STD_LOGIC; 
  signal romo2addro0_s_5_FFY_RST : STD_LOGIC; 
  signal romo2addro0_s_5_FFX_RST : STD_LOGIC; 
  signal romeaddro7_s_1_FFY_RST : STD_LOGIC; 
  signal romeaddro7_s_1_FFX_RST : STD_LOGIC; 
  signal romeaddro7_s_3_FFY_RST : STD_LOGIC; 
  signal romeaddro7_s_3_FFX_RST : STD_LOGIC; 
  signal romoaddro1_s_3_FFX_RST : STD_LOGIC; 
  signal romoaddro2_s_1_FFY_RST : STD_LOGIC; 
  signal romoaddro2_s_1_FFX_RST : STD_LOGIC; 
  signal romoaddro2_s_3_FFY_RST : STD_LOGIC; 
  signal romoaddro2_s_3_FFX_RST : STD_LOGIC; 
  signal romoaddro3_s_1_FFY_RST : STD_LOGIC; 
  signal romoaddro3_s_1_FFX_RST : STD_LOGIC; 
  signal romo2addro6_s_3_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_1_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_1_FFX_RST : STD_LOGIC; 
  signal romo2addro7_s_1_FFY_RST : STD_LOGIC; 
  signal romo2addro7_s_1_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_6_3_FFY_RST : STD_LOGIC; 
  signal romeaddro3_s_1_FFX_RST : STD_LOGIC; 
  signal romeaddro3_s_3_FFY_RST : STD_LOGIC; 
  signal romeaddro3_s_3_FFX_RST : STD_LOGIC; 
  signal romeaddro4_s_1_FFY_RST : STD_LOGIC; 
  signal romeaddro4_s_1_FFX_RST : STD_LOGIC; 
  signal romeaddro4_s_3_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_row_reg_0_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_row_reg_0_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_state_reg_1_FFY_RST : STD_LOGIC; 
  signal rome2addro4_s_1_FFY_RST : STD_LOGIC; 
  signal rome2addro4_s_1_FFX_RST : STD_LOGIC; 
  signal rome2addro4_s_3_FFY_RST : STD_LOGIC; 
  signal rome2addro4_s_3_FFX_RST : STD_LOGIC; 
  signal rome2addro5_s_1_FFY_RST : STD_LOGIC; 
  signal rome2addro5_s_1_FFX_RST : STD_LOGIC; 
  signal romeaddro8_s_1_FFY_RST : STD_LOGIC; 
  signal romeaddro8_s_1_FFX_RST : STD_LOGIC; 
  signal romeaddro8_s_3_FFY_RST : STD_LOGIC; 
  signal romeaddro8_s_3_FFX_RST : STD_LOGIC; 
  signal romeaddro4_s_3_FFX_RST : STD_LOGIC; 
  signal romeaddro5_s_1_FFY_RST : STD_LOGIC; 
  signal romeaddro5_s_1_FFX_RST : STD_LOGIC; 
  signal romeaddro5_s_3_FFY_RST : STD_LOGIC; 
  signal romeaddro5_s_3_FFX_RST : STD_LOGIC; 
  signal romo2addro10_s_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_state_reg_1_FFX_RST : STD_LOGIC; 
  signal rome2addro10_s_1_FFY_RST : STD_LOGIC; 
  signal rome2addro10_s_1_FFX_RST : STD_LOGIC; 
  signal rome2addro10_s_3_FFY_RST : STD_LOGIC; 
  signal rome2addro10_s_3_FFX_RST : STD_LOGIC; 
  signal romeaddro1_s_3_FFX_RST : STD_LOGIC; 
  signal romeaddro2_s_1_FFY_RST : STD_LOGIC; 
  signal romeaddro2_s_1_FFX_RST : STD_LOGIC; 
  signal romeaddro2_s_3_FFY_RST : STD_LOGIC; 
  signal romeaddro2_s_3_FFX_RST : STD_LOGIC; 
  signal romeaddro3_s_1_FFY_RST : STD_LOGIC; 
  signal romeaddro0_s_1_FFY_RST : STD_LOGIC; 
  signal romeaddro0_s_1_FFX_RST : STD_LOGIC; 
  signal romeaddro0_s_3_FFY_RST : STD_LOGIC; 
  signal romeaddro0_s_3_FFX_RST : STD_LOGIC; 
  signal romeaddro1_s_1_FFY_RST : STD_LOGIC; 
  signal romeaddro1_s_1_FFX_RST : STD_LOGIC; 
  signal romeaddro1_s_3_FFY_RST : STD_LOGIC; 
  signal romo2addro10_s_1_FFX_RST : STD_LOGIC; 
  signal romeaddro6_s_1_FFY_RST : STD_LOGIC; 
  signal romeaddro6_s_1_FFX_RST : STD_LOGIC; 
  signal romo2addro10_s_3_FFY_RST : STD_LOGIC; 
  signal romo2addro10_s_3_FFX_RST : STD_LOGIC; 
  signal romeaddro6_s_3_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_0_FFX_RST : STD_LOGIC; 
  signal ramwe_s_FFY_RST : STD_LOGIC; 
  signal ramwe_s_FFY_RSTAND : STD_LOGIC; 
  signal rome2addro0_s_1_FFY_RST : STD_LOGIC; 
  signal rome2addro0_s_1_FFX_RST : STD_LOGIC; 
  signal rome2addro0_s_3_FFY_RST : STD_LOGIC; 
  signal rome2addro0_s_3_FFX_RST : STD_LOGIC; 
  signal requestrd_s_FFY_RST : STD_LOGIC; 
  signal requestrd_s_FFY_RSTAND : STD_LOGIC; 
  signal ramwaddro_s_1_FFX_RST : STD_LOGIC; 
  signal ramwaddro_s_3_FFY_RST : STD_LOGIC; 
  signal ramwaddro_s_3_FFX_RST : STD_LOGIC; 
  signal ramwaddro_s_5_FFY_RST : STD_LOGIC; 
  signal ramwaddro_s_5_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_inpcnt_reg_0_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_completed_reg_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_completed_reg_FFY_RSTAND : STD_LOGIC; 
  signal U_DCT2D_col_tmp_reg_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_col_tmp_reg_1_FFX_RST : STD_LOGIC; 
  signal ramwaddro_s_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_1_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_3_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_3_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_5_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_5_FFX_RST : STD_LOGIC; 
  signal releasewr_s_FFY_RST : STD_LOGIC; 
  signal releasewr_s_FFY_RSTAND : STD_LOGIC; 
  signal U_DCT1D_latch_done_reg_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_latch_done_reg_FFY_RSTAND : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_7_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_10_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_1_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_4_3_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_colram_reg_3_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_colram_reg_3_FFY_RSTAND : STD_LOGIC; 
  signal rome2addro5_s_3_FFY_RST : STD_LOGIC; 
  signal rome2addro5_s_3_FFX_RST : STD_LOGIC; 
  signal rome2addro6_s_1_FFY_RST : STD_LOGIC; 
  signal rome2addro6_s_1_FFX_RST : STD_LOGIC; 
  signal rome2addro6_s_3_FFY_RST : STD_LOGIC; 
  signal rome2addro6_s_3_FFX_RST : STD_LOGIC; 
  signal rome2addro7_s_1_FFY_RST : STD_LOGIC; 
  signal rome2addro2_s_3_FFY_RST : STD_LOGIC; 
  signal rome2addro2_s_3_FFX_RST : STD_LOGIC; 
  signal rome2addro3_s_1_FFY_RST : STD_LOGIC; 
  signal rome2addro3_s_1_FFX_RST : STD_LOGIC; 
  signal rome2addro3_s_3_FFY_RST : STD_LOGIC; 
  signal rome2addro3_s_3_FFX_RST : STD_LOGIC; 
  signal rome2addro7_s_1_FFX_RST : STD_LOGIC; 
  signal rome2addro7_s_3_FFY_RST : STD_LOGIC; 
  signal rome2addro7_s_3_FFX_RST : STD_LOGIC; 
  signal rome2addro8_s_1_FFY_RST : STD_LOGIC; 
  signal rome2addro8_s_1_FFX_RST : STD_LOGIC; 
  signal rome2addro8_s_3_FFY_RST : STD_LOGIC; 
  signal rome2addro8_s_3_FFX_RST : STD_LOGIC; 
  signal rome2addro9_s_1_FFY_RST : STD_LOGIC; 
  signal rome2addro9_s_1_FFX_RST : STD_LOGIC; 
  signal rome2addro9_s_3_FFY_RST : STD_LOGIC; 
  signal rome2addro9_s_3_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_3_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_3_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_5_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_5_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_7_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_7_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_10_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_1_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_3_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_3_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_5_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_5_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_7_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_7_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_10_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_0_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_1_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_5_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_7_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_7_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_10_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_1_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_1_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_3_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_3_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_2_5_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_7_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_7_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_10_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_5_10_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_1_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_1_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_3_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_3_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_5_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_5_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_3_7_FFY_RST : STD_LOGIC; 
  signal releaserd_s_FFY_RST : STD_LOGIC; 
  signal releaserd_s_FFY_RSTAND : STD_LOGIC; 
  signal romoaddro0_s_1_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_3_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_3_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_5_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_5_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_7_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_7_FFX_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_10_FFY_RST : STD_LOGIC; 
  signal U_DCT2D_latchbuf_reg_6_10_FFX_RST : STD_LOGIC; 
  signal U_DCT1D_col_tmp_reg_1_FFY_RST : STD_LOGIC; 
  signal U_DCT1D_col_tmp_reg_1_FFX_RST : STD_LOGIC; 
  signal romoaddro0_s_1_FFX_RST : STD_LOGIC; 
  signal romoaddro0_s_3_FFY_RST : STD_LOGIC; 
  signal romoaddro0_s_3_FFX_RST : STD_LOGIC; 
  signal romoaddro1_s_1_FFY_RST : STD_LOGIC; 
  signal romoaddro1_s_1_FFX_RST : STD_LOGIC; 
  signal romoaddro1_s_3_FFY_RST : STD_LOGIC; 
  signal romoaddro6_s_3_FFY_RST : STD_LOGIC; 
  signal romoaddro6_s_3_FFX_RST : STD_LOGIC; 
  signal romoaddro7_s_1_FFY_RST : STD_LOGIC; 
  signal romoaddro7_s_1_FFX_RST : STD_LOGIC; 
  signal romoaddro7_s_3_FFY_RST : STD_LOGIC; 
  signal romoaddro7_s_3_FFX_RST : STD_LOGIC; 
  signal romoaddro8_s_1_FFY_RST : STD_LOGIC; 
  signal romoaddro8_s_1_FFX_RST : STD_LOGIC; 
  signal romoaddro8_s_3_FFY_RST : STD_LOGIC; 
  signal romoaddro8_s_3_FFX_RST : STD_LOGIC; 
  signal romoaddro0_s_5_FFY_RST : STD_LOGIC; 
  signal romoaddro0_s_5_FFX_RST : STD_LOGIC; 
  signal romoaddro5_s_1_FFY_RST : STD_LOGIC; 
  signal romoaddro5_s_1_FFX_RST : STD_LOGIC; 
  signal romoaddro5_s_3_FFY_RST : STD_LOGIC; 
  signal romoaddro5_s_3_FFX_RST : STD_LOGIC; 
  signal romoaddro6_s_1_FFY_RST : STD_LOGIC; 
  signal romoaddro6_s_1_FFX_RST : STD_LOGIC; 
  signal romoaddro3_s_3_FFY_RST : STD_LOGIC; 
  signal romoaddro3_s_3_FFX_RST : STD_LOGIC; 
  signal romoaddro4_s_1_FFY_RST : STD_LOGIC; 
  signal romoaddro4_s_1_FFX_RST : STD_LOGIC; 
  signal romoaddro4_s_3_FFY_RST : STD_LOGIC; 
  signal romoaddro4_s_3_FFX_RST : STD_LOGIC; 
  signal PWR_GND_0_G : STD_LOGIC; 
  signal PWR_GND_1_G : STD_LOGIC; 
  signal PWR_GND_2_G : STD_LOGIC; 
  signal PWR_GND_3_G : STD_LOGIC; 
  signal PWR_GND_4_G : STD_LOGIC; 
  signal GND : STD_LOGIC; 
  signal VCC : STD_LOGIC; 
  signal U_DCT1D_latchbuf_reg_2_Q : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal U_DCT1D_latchbuf_reg_5_Q : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal U_DCT1D_databuf_reg_2_Q : STD_LOGIC_VECTOR ( 8 downto 0 ); 
  signal U_DCT2D_databuf_reg_2_Q : STD_LOGIC_VECTOR ( 10 downto 0 ); 
  signal U_DCT2D_databuf_reg_4_Q : STD_LOGIC_VECTOR ( 10 downto 0 ); 
  signal U_DCT2D_databuf_reg_7_Q : STD_LOGIC_VECTOR ( 10 downto 0 ); 
  signal U_DCT1D_latchbuf_reg_1_Q : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal U_DCT1D_latchbuf_reg_6_Q : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal U_DCT1D_databuf_reg_1_Q : STD_LOGIC_VECTOR ( 8 downto 0 ); 
  signal U_DCT2D_rtlc5n1484 : STD_LOGIC_VECTOR ( 23 downto 9 ); 
  signal romo2datao10_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal U_DCT2D_state_reg : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal U_DCT2D_rtlc5n1501 : STD_LOGIC_VECTOR ( 23 downto 10 ); 
  signal rome2datao10_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal romo2datao8_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal romo2datao9_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal rome2datao8_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal rome2datao9_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal U_DCT2D_databuf_reg_1_Q : STD_LOGIC_VECTOR ( 10 downto 0 ); 
  signal U_DCT1D_latchbuf_reg_0_Q : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal U_DCT1D_latchbuf_reg_7_Q : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal U_DCT1D_databuf_reg_4_Q : STD_LOGIC_VECTOR ( 8 downto 0 ); 
  signal romo2datao0_s : STD_LOGIC_VECTOR ( 13 downto 1 ); 
  signal romo2datao1_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal U_DCT2D_rtlc5n1480 : STD_LOGIC_VECTOR ( 15 downto 2 ); 
  signal U_DCT1D_latchbuf_reg_3_Q : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal U_DCT1D_latchbuf_reg_4_Q : STD_LOGIC_VECTOR ( 7 downto 0 ); 
  signal U_DCT1D_databuf_reg_7_Q : STD_LOGIC_VECTOR ( 8 downto 0 ); 
  signal U_DCT2D_databuf_reg_0_Q : STD_LOGIC_VECTOR ( 10 downto 0 ); 
  signal romo2datao2_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal U_DCT2D_rtlc5n1481 : STD_LOGIC_VECTOR ( 17 downto 3 ); 
  signal U_DCT2D_rtlc5n1485 : STD_LOGIC_VECTOR ( 18 downto 4 ); 
  signal romo2datao6_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal romo2datao7_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal U_DCT2D_rtlc5n1483 : STD_LOGIC_VECTOR ( 21 downto 7 ); 
  signal U_DCT2D_databuf_reg_3_Q : STD_LOGIC_VECTOR ( 10 downto 0 ); 
  signal rome2datao2_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal rome2datao3_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal U_DCT2D_rtlc5n1493 : STD_LOGIC_VECTOR ( 17 downto 5 ); 
  signal U_DCT1D_state_reg : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal romodatao6_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal U_DCT1D_rtlc5n1346 : STD_LOGIC_VECTOR ( 19 downto 5 ); 
  signal romedatao4_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal U_DCT1D_rtlc5n1347 : STD_LOGIC_VECTOR ( 21 downto 7 ); 
  signal U_DCT1D_rtlc5n1359 : STD_LOGIC_VECTOR ( 21 downto 6 ); 
  signal U_DCT2D_databuf_reg_6_Q : STD_LOGIC_VECTOR ( 10 downto 0 ); 
  signal U_DCT1D_databuf_reg_0_Q : STD_LOGIC_VECTOR ( 8 downto 0 ); 
  signal U_DCT1D_databuf_reg_5_Q : STD_LOGIC_VECTOR ( 8 downto 0 ); 
  signal U_DCT2D_databuf_reg_5_Q : STD_LOGIC_VECTOR ( 10 downto 0 ); 
  signal U_DCT1D_databuf_reg_3_Q : STD_LOGIC_VECTOR ( 8 downto 0 ); 
  signal rome2datao0_s : STD_LOGIC_VECTOR ( 13 downto 3 ); 
  signal rome2datao1_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal U_DCT2D_rtlc5n1492 : STD_LOGIC_VECTOR ( 15 downto 4 ); 
  signal rome2datao6_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal rome2datao7_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal U_DCT2D_rtlc5n1495 : STD_LOGIC_VECTOR ( 21 downto 9 ); 
  signal U_DCT1D_databuf_reg_6_Q : STD_LOGIC_VECTOR ( 8 downto 0 ); 
  signal romodatao2_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal romodatao3_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal U_DCT1D_rtlc5n1345 : STD_LOGIC_VECTOR ( 17 downto 3 ); 
  signal romo2datao4_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal U_DCT2D_rtlc5n1482 : STD_LOGIC_VECTOR ( 19 downto 5 ); 
  signal U_DCT2D_nx115_bus : STD_LOGIC_VECTOR ( 18 downto 2 ); 
  signal U_DCT2D_rtlc5n1499 : STD_LOGIC_VECTOR ( 23 downto 8 ); 
  signal U_DCT2D_rtlc5n1491 : STD_LOGIC_VECTOR ( 23 downto 12 ); 
  signal romodatao4_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal U_DCT1D_rtlc5n1350 : STD_LOGIC_VECTOR ( 21 downto 8 ); 
  signal romedatao2_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal romedatao3_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal U_DCT1D_rtlc5n1355 : STD_LOGIC_VECTOR ( 17 downto 5 ); 
  signal rome2datao4_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal U_DCT2D_rtlc5n1494 : STD_LOGIC_VECTOR ( 19 downto 7 ); 
  signal U_DCT2D_rtlc5n1498 : STD_LOGIC_VECTOR ( 22 downto 8 ); 
  signal romodatao5_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal romedatao5_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal rome2datao5_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal romodatao0_s : STD_LOGIC_VECTOR ( 13 downto 1 ); 
  signal romodatao1_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal U_DCT1D_rtlc5n1344 : STD_LOGIC_VECTOR ( 15 downto 2 ); 
  signal romo2datao3_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal romedatao0_s : STD_LOGIC_VECTOR ( 13 downto 3 ); 
  signal romedatao1_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal U_DCT1D_rtlc5n1354 : STD_LOGIC_VECTOR ( 15 downto 4 ); 
  signal U_DCT1D_rtlc5n1348 : STD_LOGIC_VECTOR ( 18 downto 4 ); 
  signal romodatao8_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal romedatao8_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal ramdatai_s : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal romodatao7_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal romedatao6_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal romedatao7_s : STD_LOGIC_VECTOR ( 13 downto 2 ); 
  signal romo2datao5_s : STD_LOGIC_VECTOR ( 13 downto 0 ); 
  signal rome2addro0_s : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal rome2addro9_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal rome2addro8_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal rome2addro10_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal rome2addro2_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal rome2addro1_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romo2addro0_s : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal romo2addro1_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romo2addro7_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romo2addro8_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romo2addro9_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal rome2addro4_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romo2addro2_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal rome2addro3_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romo2addro3_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal rome2addro5_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal rome2addro6_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romo2addro10_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romo2addro4_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal rome2addro7_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romo2addro6_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romo2addro5_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romeaddro0_s : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal romoaddro0_s : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal romeaddro8_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romeaddro2_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romoaddro1_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romeaddro1_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romoaddro8_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romoaddro2_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romeaddro4_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romeaddro3_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romeaddro5_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romoaddro5_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romoaddro4_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romoaddro3_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romeaddro6_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romoaddro6_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romeaddro7_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal romoaddro7_s : STD_LOGIC_VECTOR ( 3 downto 0 ); 
  signal dcti_int : STD_LOGIC_VECTOR ( 7 downto 7 ); 
  signal U_DCT1D_istate_reg : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal ramwaddro_s : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal ramraddro_s : STD_LOGIC_VECTOR ( 5 downto 0 ); 
  signal ramdatao2_s : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal ramdatao1_s : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal U_DCT2D_istate_reg : STD_LOGIC_VECTOR ( 1 downto 0 ); 
  signal U_DCT2D_col_reg : STD_LOGIC_VECTOR ( 2 downto 0 ); 
  signal U_DCT1D_col_reg : STD_LOGIC_VECTOR ( 2 downto 0 ); 
  signal U_DCT1D_row_reg : STD_LOGIC_VECTOR ( 2 downto 0 ); 
  signal U_DCT2D_col_tmp_reg : STD_LOGIC_VECTOR ( 2 downto 1 ); 
  signal U_DCT1D_col_tmp_reg : STD_LOGIC_VECTOR ( 2 downto 1 ); 
  signal U_DCT2D_colram_reg : STD_LOGIC_VECTOR ( 3 downto 3 ); 
  signal U_DCT1D_inpcnt_reg : STD_LOGIC_VECTOR ( 2 downto 0 ); 
  signal U_DCT2D_rtlc2_istate_reg_fsm_SS9_n171 : STD_LOGIC_VECTOR ( 0 downto 0 ); 
  signal U_DCT2D_rtlc5_romeaddro0_SS3_n342 : STD_LOGIC_VECTOR ( 5 downto 4 ); 
  signal U_DCT1D_rtlc5_romeaddro0_SS4_n350 : STD_LOGIC_VECTOR ( 5 downto 4 ); 
  signal ramdatao_s : STD_LOGIC_VECTOR ( 9 downto 0 ); 
  signal U_DCT1D_rtlc5_state_reg_fsm_SS4_n374 : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal U_DCT2D_rtlc5_state_reg_fsm_SS3_n367 : STD_LOGIC_VECTOR ( 1 downto 1 ); 
  signal U_DCT2D_rtlc5n942 : STD_LOGIC_VECTOR ( 2 downto 2 ); 
  signal U_DCT1D_rtlc5n875 : STD_LOGIC_VECTOR ( 2 downto 2 ); 
  signal dcto_dup0 : STD_LOGIC_VECTOR ( 11 downto 0 ); 
begin
  U_DCT1D_databuf_reg_2_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_2_0_FFY_RST
    );
  U_DCT1D_reg_databuf_reg_2_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_2_0_DYMUX,
      CE => U_DCT1D_databuf_reg_2_0_CEINV,
      CLK => U_DCT1D_databuf_reg_2_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_2_0_FFY_RST,
      O => U_DCT1D_databuf_reg_2_Q(1)
    );
  U_DCT1D_ix60819z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_2_Q(1),
      ADR1 => U_DCT1D_latchbuf_reg_5_Q(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx60819z1
    );
  U_DCT1D_databuf_reg_2_0_DXMUX_0 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_0_XORF,
      O => U_DCT1D_databuf_reg_2_0_DXMUX
    );
  U_DCT1D_databuf_reg_2_0_XORF_1 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_0_CYINIT,
      I1 => U_DCT1D_nx59822z1,
      O => U_DCT1D_databuf_reg_2_0_XORF
    );
  U_DCT1D_databuf_reg_2_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_0_CY0F,
      IB => U_DCT1D_databuf_reg_2_0_CYINIT,
      SEL => U_DCT1D_databuf_reg_2_0_CYSELF,
      O => U_DCT1D_rtlc5_1421_add_10_ix60819z63342_O
    );
  U_DCT1D_databuf_reg_2_0_CYINIT_2 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_0_BXINVNOT,
      O => U_DCT1D_databuf_reg_2_0_CYINIT
    );
  U_DCT1D_databuf_reg_2_0_CY0F_3 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(0),
      O => U_DCT1D_databuf_reg_2_0_CY0F
    );
  U_DCT1D_databuf_reg_2_0_CYSELF_4 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59822z1,
      O => U_DCT1D_databuf_reg_2_0_CYSELF
    );
  U_DCT1D_databuf_reg_2_0_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_16,
      O => U_DCT1D_databuf_reg_2_0_BXINVNOT
    );
  U_DCT1D_databuf_reg_2_0_DYMUX_5 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_0_XORG,
      O => U_DCT1D_databuf_reg_2_0_DYMUX
    );
  U_DCT1D_databuf_reg_2_0_XORG_6 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1421_add_10_ix60819z63342_O,
      I1 => U_DCT1D_nx60819z1,
      O => U_DCT1D_databuf_reg_2_0_XORG
    );
  U_DCT1D_databuf_reg_2_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_0_CYMUXG,
      O => U_DCT1D_rtlc5_1421_add_10_ix61816z63342_O
    );
  U_DCT1D_databuf_reg_2_0_CYMUXG_7 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_0_CY0G,
      IB => U_DCT1D_rtlc5_1421_add_10_ix60819z63342_O,
      SEL => U_DCT1D_databuf_reg_2_0_CYSELG,
      O => U_DCT1D_databuf_reg_2_0_CYMUXG
    );
  U_DCT1D_databuf_reg_2_0_CY0G_8 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(1),
      O => U_DCT1D_databuf_reg_2_0_CY0G
    );
  U_DCT1D_databuf_reg_2_0_CYSELG_9 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx60819z1,
      O => U_DCT1D_databuf_reg_2_0_CYSELG
    );
  U_DCT1D_databuf_reg_2_0_SRINV_10 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_2_0_SRINV
    );
  U_DCT1D_databuf_reg_2_0_CLKINV_11 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_2_0_CLKINV
    );
  U_DCT1D_databuf_reg_2_0_CEINV_12 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_2_0_CEINV
    );
  U_DCT1D_databuf_reg_2_2_DXMUX_13 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_2_XORF,
      O => U_DCT1D_databuf_reg_2_2_DXMUX
    );
  U_DCT1D_databuf_reg_2_2_XORF_14 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_2_CYINIT,
      I1 => U_DCT1D_nx61816z1,
      O => U_DCT1D_databuf_reg_2_2_XORF
    );
  U_DCT1D_databuf_reg_2_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_2_CY0F,
      IB => U_DCT1D_databuf_reg_2_2_CYINIT,
      SEL => U_DCT1D_databuf_reg_2_2_CYSELF,
      O => U_DCT1D_rtlc5_1421_add_10_ix62813z63342_O
    );
  U_DCT1D_databuf_reg_2_2_CYMUXF2_15 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_2_CY0F,
      IB => U_DCT1D_databuf_reg_2_2_CY0F,
      SEL => U_DCT1D_databuf_reg_2_2_CYSELF,
      O => U_DCT1D_databuf_reg_2_2_CYMUXF2
    );
  U_DCT1D_databuf_reg_2_2_CYINIT_16 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1421_add_10_ix61816z63342_O,
      O => U_DCT1D_databuf_reg_2_2_CYINIT
    );
  U_DCT1D_databuf_reg_2_2_CY0F_17 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(2),
      O => U_DCT1D_databuf_reg_2_2_CY0F
    );
  U_DCT1D_databuf_reg_2_2_CYSELF_18 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx61816z1,
      O => U_DCT1D_databuf_reg_2_2_CYSELF
    );
  U_DCT1D_databuf_reg_2_2_DYMUX_19 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_2_XORG,
      O => U_DCT1D_databuf_reg_2_2_DYMUX
    );
  U_DCT1D_databuf_reg_2_2_XORG_20 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1421_add_10_ix62813z63342_O,
      I1 => U_DCT1D_nx62813z1,
      O => U_DCT1D_databuf_reg_2_2_XORG
    );
  U_DCT1D_databuf_reg_2_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_2_CYMUXFAST,
      O => U_DCT1D_rtlc5_1421_add_10_ix63810z63342_O
    );
  U_DCT1D_databuf_reg_2_2_FASTCARRY_21 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1421_add_10_ix61816z63342_O,
      O => U_DCT1D_databuf_reg_2_2_FASTCARRY
    );
  U_DCT1D_databuf_reg_2_2_CYAND_22 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_2_2_CYSELG,
      I1 => U_DCT1D_databuf_reg_2_2_CYSELF,
      O => U_DCT1D_databuf_reg_2_2_CYAND
    );
  U_DCT1D_databuf_reg_2_2_CYMUXFAST_23 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_2_CYMUXG2,
      IB => U_DCT1D_databuf_reg_2_2_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_2_2_CYAND,
      O => U_DCT1D_databuf_reg_2_2_CYMUXFAST
    );
  U_DCT1D_databuf_reg_2_2_CYMUXG2_24 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_2_CY0G,
      IB => U_DCT1D_databuf_reg_2_2_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_2_2_CYSELG,
      O => U_DCT1D_databuf_reg_2_2_CYMUXG2
    );
  U_DCT1D_databuf_reg_2_2_CY0G_25 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(3),
      O => U_DCT1D_databuf_reg_2_2_CY0G
    );
  U_DCT1D_databuf_reg_2_2_CYSELG_26 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx62813z1,
      O => U_DCT1D_databuf_reg_2_2_CYSELG
    );
  U_DCT1D_databuf_reg_2_2_SRINV_27 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_2_2_SRINV
    );
  U_DCT1D_databuf_reg_2_2_CLKINV_28 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_2_2_CLKINV
    );
  U_DCT1D_databuf_reg_2_2_CEINV_29 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_2_2_CEINV
    );
  U_DCT1D_databuf_reg_2_4_DXMUX_30 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_4_XORF,
      O => U_DCT1D_databuf_reg_2_4_DXMUX
    );
  U_DCT1D_databuf_reg_2_4_XORF_31 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_4_CYINIT,
      I1 => U_DCT1D_nx63810z1,
      O => U_DCT1D_databuf_reg_2_4_XORF
    );
  U_DCT1D_databuf_reg_2_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_4_CY0F,
      IB => U_DCT1D_databuf_reg_2_4_CYINIT,
      SEL => U_DCT1D_databuf_reg_2_4_CYSELF,
      O => U_DCT1D_rtlc5_1421_add_10_ix64807z63342_O
    );
  U_DCT1D_databuf_reg_2_4_CYMUXF2_32 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_4_CY0F,
      IB => U_DCT1D_databuf_reg_2_4_CY0F,
      SEL => U_DCT1D_databuf_reg_2_4_CYSELF,
      O => U_DCT1D_databuf_reg_2_4_CYMUXF2
    );
  U_DCT1D_databuf_reg_2_4_CYINIT_33 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1421_add_10_ix63810z63342_O,
      O => U_DCT1D_databuf_reg_2_4_CYINIT
    );
  U_DCT1D_databuf_reg_2_4_CY0F_34 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(4),
      O => U_DCT1D_databuf_reg_2_4_CY0F
    );
  U_DCT1D_databuf_reg_2_4_CYSELF_35 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx63810z1,
      O => U_DCT1D_databuf_reg_2_4_CYSELF
    );
  U_DCT1D_databuf_reg_2_4_DYMUX_36 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_4_XORG,
      O => U_DCT1D_databuf_reg_2_4_DYMUX
    );
  U_DCT1D_databuf_reg_2_4_XORG_37 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1421_add_10_ix64807z63342_O,
      I1 => U_DCT1D_nx64807z1,
      O => U_DCT1D_databuf_reg_2_4_XORG
    );
  U_DCT1D_databuf_reg_2_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_4_CYMUXFAST,
      O => U_DCT1D_rtlc5_1421_add_10_ix268z63342_O
    );
  U_DCT1D_databuf_reg_2_4_FASTCARRY_38 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1421_add_10_ix63810z63342_O,
      O => U_DCT1D_databuf_reg_2_4_FASTCARRY
    );
  U_DCT1D_databuf_reg_2_4_CYAND_39 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_2_4_CYSELG,
      I1 => U_DCT1D_databuf_reg_2_4_CYSELF,
      O => U_DCT1D_databuf_reg_2_4_CYAND
    );
  U_DCT1D_databuf_reg_2_4_CYMUXFAST_40 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_4_CYMUXG2,
      IB => U_DCT1D_databuf_reg_2_4_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_2_4_CYAND,
      O => U_DCT1D_databuf_reg_2_4_CYMUXFAST
    );
  U_DCT1D_databuf_reg_2_4_CYMUXG2_41 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_4_CY0G,
      IB => U_DCT1D_databuf_reg_2_4_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_2_4_CYSELG,
      O => U_DCT1D_databuf_reg_2_4_CYMUXG2
    );
  U_DCT1D_databuf_reg_2_4_CY0G_42 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(5),
      O => U_DCT1D_databuf_reg_2_4_CY0G
    );
  U_DCT1D_databuf_reg_2_4_CYSELG_43 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx64807z1,
      O => U_DCT1D_databuf_reg_2_4_CYSELG
    );
  U_DCT1D_databuf_reg_2_4_SRINV_44 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_2_4_SRINV
    );
  U_DCT1D_databuf_reg_2_4_CLKINV_45 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_2_4_CLKINV
    );
  U_DCT1D_databuf_reg_2_4_CEINV_46 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_2_4_CEINV
    );
  U_DCT1D_databuf_reg_2_6_DXMUX_47 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_6_XORF,
      O => U_DCT1D_databuf_reg_2_6_DXMUX
    );
  U_DCT1D_databuf_reg_2_6_XORF_48 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_6_CYINIT,
      I1 => U_DCT1D_nx268z1,
      O => U_DCT1D_databuf_reg_2_6_XORF
    );
  U_DCT1D_databuf_reg_2_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_6_CY0F,
      IB => U_DCT1D_databuf_reg_2_6_CYINIT,
      SEL => U_DCT1D_databuf_reg_2_6_CYSELF,
      O => U_DCT1D_rtlc5_1421_add_10_ix1265z63342_O
    );
  U_DCT1D_databuf_reg_2_6_CYMUXF2_49 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_6_CY0F,
      IB => U_DCT1D_databuf_reg_2_6_CY0F,
      SEL => U_DCT1D_databuf_reg_2_6_CYSELF,
      O => U_DCT1D_databuf_reg_2_6_CYMUXF2
    );
  U_DCT1D_databuf_reg_2_6_CYINIT_50 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1421_add_10_ix268z63342_O,
      O => U_DCT1D_databuf_reg_2_6_CYINIT
    );
  U_DCT1D_databuf_reg_2_6_CY0F_51 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(6),
      O => U_DCT1D_databuf_reg_2_6_CY0F
    );
  U_DCT1D_databuf_reg_2_6_CYSELF_52 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx268z1,
      O => U_DCT1D_databuf_reg_2_6_CYSELF
    );
  U_DCT1D_databuf_reg_2_6_DYMUX_53 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_6_XORG,
      O => U_DCT1D_databuf_reg_2_6_DYMUX
    );
  U_DCT1D_databuf_reg_2_6_XORG_54 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1421_add_10_ix1265z63342_O,
      I1 => U_DCT1D_nx1265z1,
      O => U_DCT1D_databuf_reg_2_6_XORG
    );
  U_DCT1D_databuf_reg_2_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_6_CYMUXFAST,
      O => U_DCT1D_rtlc5_1421_add_10_ix2262z63342_O
    );
  U_DCT1D_databuf_reg_2_6_FASTCARRY_55 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1421_add_10_ix268z63342_O,
      O => U_DCT1D_databuf_reg_2_6_FASTCARRY
    );
  U_DCT1D_databuf_reg_2_6_CYAND_56 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_2_6_CYSELG,
      I1 => U_DCT1D_databuf_reg_2_6_CYSELF,
      O => U_DCT1D_databuf_reg_2_6_CYAND
    );
  U_DCT1D_databuf_reg_2_6_CYMUXFAST_57 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_6_CYMUXG2,
      IB => U_DCT1D_databuf_reg_2_6_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_2_6_CYAND,
      O => U_DCT1D_databuf_reg_2_6_CYMUXFAST
    );
  U_DCT1D_databuf_reg_2_6_CYMUXG2_58 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_2_6_CY0G,
      IB => U_DCT1D_databuf_reg_2_6_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_2_6_CYSELG,
      O => U_DCT1D_databuf_reg_2_6_CYMUXG2
    );
  U_DCT1D_databuf_reg_2_6_CY0G_59 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(7),
      O => U_DCT1D_databuf_reg_2_6_CY0G
    );
  U_DCT1D_databuf_reg_2_6_CYSELG_60 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx1265z1,
      O => U_DCT1D_databuf_reg_2_6_CYSELG
    );
  U_DCT1D_databuf_reg_2_6_SRINV_61 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_2_6_SRINV
    );
  U_DCT1D_databuf_reg_2_6_CLKINV_62 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_2_6_CLKINV
    );
  U_DCT1D_databuf_reg_2_6_CEINV_63 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_2_6_CEINV
    );
  U_DCT1D_databuf_reg_2_8_DXMUX_64 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_8_XORF,
      O => U_DCT1D_databuf_reg_2_8_DXMUX
    );
  U_DCT1D_databuf_reg_2_8_XORF_65 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_8_CYINIT,
      I1 => U_DCT1D_nx2262z1_rt,
      O => U_DCT1D_databuf_reg_2_8_XORF
    );
  U_DCT1D_databuf_reg_2_8_CYINIT_66 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1421_add_10_ix2262z63342_O,
      O => U_DCT1D_databuf_reg_2_8_CYINIT
    );
  U_DCT1D_databuf_reg_2_8_CLKINV_67 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_2_8_CLKINV
    );
  U_DCT1D_databuf_reg_2_8_CEINV_68 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_2_8_CEINV
    );
  U_DCT2D_databuf_reg_2_0_DXMUX_69 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_0_XORF,
      O => U_DCT2D_databuf_reg_2_0_DXMUX
    );
  U_DCT2D_databuf_reg_2_0_XORF_70 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_0_CYINIT,
      I1 => U_DCT2D_nx59822z1,
      O => U_DCT2D_databuf_reg_2_0_XORF
    );
  U_DCT2D_databuf_reg_2_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_0_CY0F,
      IB => U_DCT2D_databuf_reg_2_0_CYINIT,
      SEL => U_DCT2D_databuf_reg_2_0_CYSELF,
      O => U_DCT2D_rtlc5_1580_add_47_ix60819z63342_O
    );
  U_DCT2D_databuf_reg_2_0_CYINIT_71 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_0_BXINVNOT,
      O => U_DCT2D_databuf_reg_2_0_CYINIT
    );
  U_DCT2D_databuf_reg_2_0_CY0F_72 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_0_Q,
      O => U_DCT2D_databuf_reg_2_0_CY0F
    );
  U_DCT2D_databuf_reg_2_0_CYSELF_73 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx59822z1,
      O => U_DCT2D_databuf_reg_2_0_CYSELF
    );
  U_DCT2D_databuf_reg_2_0_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_26,
      O => U_DCT2D_databuf_reg_2_0_BXINVNOT
    );
  U_DCT2D_databuf_reg_2_0_DYMUX_74 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_0_XORG,
      O => U_DCT2D_databuf_reg_2_0_DYMUX
    );
  U_DCT2D_databuf_reg_2_0_XORG_75 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1580_add_47_ix60819z63342_O,
      I1 => U_DCT2D_nx60819z1,
      O => U_DCT2D_databuf_reg_2_0_XORG
    );
  U_DCT2D_databuf_reg_2_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_0_CYMUXG,
      O => U_DCT2D_rtlc5_1580_add_47_ix61816z63342_O
    );
  U_DCT2D_databuf_reg_2_0_CYMUXG_76 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_0_CY0G,
      IB => U_DCT2D_rtlc5_1580_add_47_ix60819z63342_O,
      SEL => U_DCT2D_databuf_reg_2_0_CYSELG,
      O => U_DCT2D_databuf_reg_2_0_CYMUXG
    );
  U_DCT2D_databuf_reg_2_0_CY0G_77 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_1_Q,
      O => U_DCT2D_databuf_reg_2_0_CY0G
    );
  U_DCT2D_databuf_reg_2_0_CYSELG_78 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx60819z1,
      O => U_DCT2D_databuf_reg_2_0_CYSELG
    );
  U_DCT2D_databuf_reg_2_0_SRINV_79 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_2_0_SRINV
    );
  U_DCT2D_databuf_reg_2_0_CLKINV_80 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_2_0_CLKINV
    );
  U_DCT2D_databuf_reg_2_0_CEINV_81 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_2_0_CEINV
    );
  U_DCT2D_databuf_reg_2_2_DXMUX_82 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_2_XORF,
      O => U_DCT2D_databuf_reg_2_2_DXMUX
    );
  U_DCT2D_databuf_reg_2_2_XORF_83 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_2_CYINIT,
      I1 => U_DCT2D_nx61816z1,
      O => U_DCT2D_databuf_reg_2_2_XORF
    );
  U_DCT2D_databuf_reg_2_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_2_CY0F,
      IB => U_DCT2D_databuf_reg_2_2_CYINIT,
      SEL => U_DCT2D_databuf_reg_2_2_CYSELF,
      O => U_DCT2D_rtlc5_1580_add_47_ix62813z63342_O
    );
  U_DCT2D_databuf_reg_2_2_CYMUXF2_84 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_2_CY0F,
      IB => U_DCT2D_databuf_reg_2_2_CY0F,
      SEL => U_DCT2D_databuf_reg_2_2_CYSELF,
      O => U_DCT2D_databuf_reg_2_2_CYMUXF2
    );
  U_DCT2D_databuf_reg_2_2_CYINIT_85 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1580_add_47_ix61816z63342_O,
      O => U_DCT2D_databuf_reg_2_2_CYINIT
    );
  U_DCT2D_databuf_reg_2_2_CY0F_86 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_2_Q,
      O => U_DCT2D_databuf_reg_2_2_CY0F
    );
  U_DCT2D_databuf_reg_2_2_CYSELF_87 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx61816z1,
      O => U_DCT2D_databuf_reg_2_2_CYSELF
    );
  U_DCT2D_databuf_reg_2_2_DYMUX_88 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_2_XORG,
      O => U_DCT2D_databuf_reg_2_2_DYMUX
    );
  U_DCT2D_databuf_reg_2_2_XORG_89 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1580_add_47_ix62813z63342_O,
      I1 => U_DCT2D_nx62813z1,
      O => U_DCT2D_databuf_reg_2_2_XORG
    );
  U_DCT2D_databuf_reg_2_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_2_CYMUXFAST,
      O => U_DCT2D_rtlc5_1580_add_47_ix63810z63342_O
    );
  U_DCT2D_databuf_reg_2_2_FASTCARRY_90 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1580_add_47_ix61816z63342_O,
      O => U_DCT2D_databuf_reg_2_2_FASTCARRY
    );
  U_DCT2D_databuf_reg_2_2_CYAND_91 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_2_2_CYSELG,
      I1 => U_DCT2D_databuf_reg_2_2_CYSELF,
      O => U_DCT2D_databuf_reg_2_2_CYAND
    );
  U_DCT2D_databuf_reg_2_2_CYMUXFAST_92 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_2_CYMUXG2,
      IB => U_DCT2D_databuf_reg_2_2_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_2_2_CYAND,
      O => U_DCT2D_databuf_reg_2_2_CYMUXFAST
    );
  U_DCT2D_databuf_reg_2_2_CYMUXG2_93 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_2_CY0G,
      IB => U_DCT2D_databuf_reg_2_2_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_2_2_CYSELG,
      O => U_DCT2D_databuf_reg_2_2_CYMUXG2
    );
  U_DCT2D_databuf_reg_2_2_CY0G_94 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_3_Q,
      O => U_DCT2D_databuf_reg_2_2_CY0G
    );
  U_DCT2D_databuf_reg_2_2_CYSELG_95 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx62813z1,
      O => U_DCT2D_databuf_reg_2_2_CYSELG
    );
  U_DCT2D_databuf_reg_2_2_SRINV_96 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_2_2_SRINV
    );
  U_DCT2D_databuf_reg_2_2_CLKINV_97 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_2_2_CLKINV
    );
  U_DCT2D_databuf_reg_2_2_CEINV_98 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_2_2_CEINV
    );
  U_DCT2D_databuf_reg_2_4_DXMUX_99 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_4_XORF,
      O => U_DCT2D_databuf_reg_2_4_DXMUX
    );
  U_DCT2D_databuf_reg_2_4_XORF_100 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_4_CYINIT,
      I1 => U_DCT2D_nx63810z1,
      O => U_DCT2D_databuf_reg_2_4_XORF
    );
  U_DCT2D_databuf_reg_2_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_4_CY0F,
      IB => U_DCT2D_databuf_reg_2_4_CYINIT,
      SEL => U_DCT2D_databuf_reg_2_4_CYSELF,
      O => U_DCT2D_rtlc5_1580_add_47_ix64807z63342_O
    );
  U_DCT2D_databuf_reg_2_4_CYMUXF2_101 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_4_CY0F,
      IB => U_DCT2D_databuf_reg_2_4_CY0F,
      SEL => U_DCT2D_databuf_reg_2_4_CYSELF,
      O => U_DCT2D_databuf_reg_2_4_CYMUXF2
    );
  U_DCT2D_databuf_reg_2_4_CYINIT_102 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1580_add_47_ix63810z63342_O,
      O => U_DCT2D_databuf_reg_2_4_CYINIT
    );
  U_DCT2D_databuf_reg_2_4_CY0F_103 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_4_Q,
      O => U_DCT2D_databuf_reg_2_4_CY0F
    );
  U_DCT2D_databuf_reg_2_4_CYSELF_104 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx63810z1,
      O => U_DCT2D_databuf_reg_2_4_CYSELF
    );
  U_DCT2D_databuf_reg_2_4_DYMUX_105 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_4_XORG,
      O => U_DCT2D_databuf_reg_2_4_DYMUX
    );
  U_DCT2D_databuf_reg_2_4_XORG_106 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1580_add_47_ix64807z63342_O,
      I1 => U_DCT2D_nx64807z1,
      O => U_DCT2D_databuf_reg_2_4_XORG
    );
  U_DCT2D_databuf_reg_2_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_4_CYMUXFAST,
      O => U_DCT2D_rtlc5_1580_add_47_ix268z63342_O
    );
  U_DCT2D_databuf_reg_2_4_FASTCARRY_107 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1580_add_47_ix63810z63342_O,
      O => U_DCT2D_databuf_reg_2_4_FASTCARRY
    );
  U_DCT2D_databuf_reg_2_4_CYAND_108 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_2_4_CYSELG,
      I1 => U_DCT2D_databuf_reg_2_4_CYSELF,
      O => U_DCT2D_databuf_reg_2_4_CYAND
    );
  U_DCT2D_databuf_reg_2_4_CYMUXFAST_109 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_4_CYMUXG2,
      IB => U_DCT2D_databuf_reg_2_4_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_2_4_CYAND,
      O => U_DCT2D_databuf_reg_2_4_CYMUXFAST
    );
  U_DCT2D_databuf_reg_2_4_CYMUXG2_110 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_4_CY0G,
      IB => U_DCT2D_databuf_reg_2_4_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_2_4_CYSELG,
      O => U_DCT2D_databuf_reg_2_4_CYMUXG2
    );
  U_DCT2D_databuf_reg_2_4_CY0G_111 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_5_Q,
      O => U_DCT2D_databuf_reg_2_4_CY0G
    );
  U_DCT2D_databuf_reg_2_4_CYSELG_112 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx64807z1,
      O => U_DCT2D_databuf_reg_2_4_CYSELG
    );
  U_DCT2D_databuf_reg_2_4_SRINV_113 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_2_4_SRINV
    );
  U_DCT2D_databuf_reg_2_4_CLKINV_114 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_2_4_CLKINV
    );
  U_DCT2D_databuf_reg_2_4_CEINV_115 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_2_4_CEINV
    );
  U_DCT2D_databuf_reg_2_6_DXMUX_116 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_6_XORF,
      O => U_DCT2D_databuf_reg_2_6_DXMUX
    );
  U_DCT2D_databuf_reg_2_6_XORF_117 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_6_CYINIT,
      I1 => U_DCT2D_nx268z1,
      O => U_DCT2D_databuf_reg_2_6_XORF
    );
  U_DCT2D_databuf_reg_2_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_6_CY0F,
      IB => U_DCT2D_databuf_reg_2_6_CYINIT,
      SEL => U_DCT2D_databuf_reg_2_6_CYSELF,
      O => U_DCT2D_rtlc5_1580_add_47_ix1265z63342_O
    );
  U_DCT2D_databuf_reg_2_6_CYMUXF2_118 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_6_CY0F,
      IB => U_DCT2D_databuf_reg_2_6_CY0F,
      SEL => U_DCT2D_databuf_reg_2_6_CYSELF,
      O => U_DCT2D_databuf_reg_2_6_CYMUXF2
    );
  U_DCT2D_databuf_reg_2_6_CYINIT_119 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1580_add_47_ix268z63342_O,
      O => U_DCT2D_databuf_reg_2_6_CYINIT
    );
  U_DCT2D_databuf_reg_2_6_CY0F_120 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_6_Q,
      O => U_DCT2D_databuf_reg_2_6_CY0F
    );
  U_DCT2D_databuf_reg_2_6_CYSELF_121 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx268z1,
      O => U_DCT2D_databuf_reg_2_6_CYSELF
    );
  U_DCT2D_databuf_reg_2_6_DYMUX_122 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_6_XORG,
      O => U_DCT2D_databuf_reg_2_6_DYMUX
    );
  U_DCT2D_databuf_reg_2_6_XORG_123 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1580_add_47_ix1265z63342_O,
      I1 => U_DCT2D_nx1265z1,
      O => U_DCT2D_databuf_reg_2_6_XORG
    );
  U_DCT2D_databuf_reg_2_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_6_CYMUXFAST,
      O => U_DCT2D_rtlc5_1580_add_47_ix2262z63342_O
    );
  U_DCT2D_databuf_reg_2_6_FASTCARRY_124 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1580_add_47_ix268z63342_O,
      O => U_DCT2D_databuf_reg_2_6_FASTCARRY
    );
  U_DCT2D_databuf_reg_2_6_CYAND_125 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_2_6_CYSELG,
      I1 => U_DCT2D_databuf_reg_2_6_CYSELF,
      O => U_DCT2D_databuf_reg_2_6_CYAND
    );
  U_DCT2D_databuf_reg_2_6_CYMUXFAST_126 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_6_CYMUXG2,
      IB => U_DCT2D_databuf_reg_2_6_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_2_6_CYAND,
      O => U_DCT2D_databuf_reg_2_6_CYMUXFAST
    );
  U_DCT2D_databuf_reg_2_6_CYMUXG2_127 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_6_CY0G,
      IB => U_DCT2D_databuf_reg_2_6_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_2_6_CYSELG,
      O => U_DCT2D_databuf_reg_2_6_CYMUXG2
    );
  U_DCT2D_databuf_reg_2_6_CY0G_128 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_7_Q,
      O => U_DCT2D_databuf_reg_2_6_CY0G
    );
  U_DCT2D_databuf_reg_2_6_CYSELG_129 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx1265z1,
      O => U_DCT2D_databuf_reg_2_6_CYSELG
    );
  U_DCT2D_databuf_reg_2_6_SRINV_130 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_2_6_SRINV
    );
  U_DCT2D_databuf_reg_2_6_CLKINV_131 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_2_6_CLKINV
    );
  U_DCT2D_databuf_reg_2_6_CEINV_132 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_2_6_CEINV
    );
  U_DCT2D_databuf_reg_2_8_DXMUX_133 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_8_XORF,
      O => U_DCT2D_databuf_reg_2_8_DXMUX
    );
  U_DCT2D_databuf_reg_2_8_XORF_134 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_8_CYINIT,
      I1 => U_DCT2D_nx2262z1,
      O => U_DCT2D_databuf_reg_2_8_XORF
    );
  U_DCT2D_databuf_reg_2_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_8_CY0F,
      IB => U_DCT2D_databuf_reg_2_8_CYINIT,
      SEL => U_DCT2D_databuf_reg_2_8_CYSELF,
      O => U_DCT2D_rtlc5_1580_add_47_ix3259z63342_O
    );
  U_DCT2D_databuf_reg_2_8_CYMUXF2_135 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_8_CY0F,
      IB => U_DCT2D_databuf_reg_2_8_CY0F,
      SEL => U_DCT2D_databuf_reg_2_8_CYSELF,
      O => U_DCT2D_databuf_reg_2_8_CYMUXF2
    );
  U_DCT2D_databuf_reg_2_8_CYINIT_136 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1580_add_47_ix2262z63342_O,
      O => U_DCT2D_databuf_reg_2_8_CYINIT
    );
  U_DCT2D_databuf_reg_2_8_CY0F_137 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_8_Q,
      O => U_DCT2D_databuf_reg_2_8_CY0F
    );
  U_DCT2D_databuf_reg_2_8_CYSELF_138 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx2262z1,
      O => U_DCT2D_databuf_reg_2_8_CYSELF
    );
  U_DCT2D_databuf_reg_2_8_DYMUX_139 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_8_XORG,
      O => U_DCT2D_databuf_reg_2_8_DYMUX
    );
  U_DCT2D_databuf_reg_2_8_XORG_140 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1580_add_47_ix3259z63342_O,
      I1 => U_DCT2D_nx3259z1,
      O => U_DCT2D_databuf_reg_2_8_XORG
    );
  U_DCT2D_databuf_reg_2_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_8_CYMUXFAST,
      O => U_DCT2D_rtlc5_1580_add_47_ix22763z63342_O
    );
  U_DCT2D_databuf_reg_2_8_FASTCARRY_141 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1580_add_47_ix2262z63342_O,
      O => U_DCT2D_databuf_reg_2_8_FASTCARRY
    );
  U_DCT2D_databuf_reg_2_8_CYAND_142 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_2_8_CYSELG,
      I1 => U_DCT2D_databuf_reg_2_8_CYSELF,
      O => U_DCT2D_databuf_reg_2_8_CYAND
    );
  U_DCT2D_databuf_reg_2_8_CYMUXFAST_143 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_8_CYMUXG2,
      IB => U_DCT2D_databuf_reg_2_8_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_2_8_CYAND,
      O => U_DCT2D_databuf_reg_2_8_CYMUXFAST
    );
  U_DCT2D_databuf_reg_2_8_CYMUXG2_144 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_2_8_CY0G,
      IB => U_DCT2D_databuf_reg_2_8_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_2_8_CYSELG,
      O => U_DCT2D_databuf_reg_2_8_CYMUXG2
    );
  U_DCT2D_databuf_reg_2_8_CY0G_145 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_10_Q,
      O => U_DCT2D_databuf_reg_2_8_CY0G
    );
  U_DCT2D_databuf_reg_2_8_CYSELG_146 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx3259z1,
      O => U_DCT2D_databuf_reg_2_8_CYSELG
    );
  U_DCT2D_databuf_reg_2_8_SRINV_147 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_2_8_SRINV
    );
  U_DCT2D_databuf_reg_2_8_CLKINV_148 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_2_8_CLKINV
    );
  U_DCT2D_databuf_reg_2_8_CEINV_149 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_2_8_CEINV
    );
  U_DCT2D_nx22763z1_rt_150 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_nx22763z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx22763z1_rt
    );
  U_DCT2D_databuf_reg_2_10_DXMUX_151 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_10_XORF,
      O => U_DCT2D_databuf_reg_2_10_DXMUX
    );
  U_DCT2D_databuf_reg_2_10_XORF_152 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_10_CYINIT,
      I1 => U_DCT2D_nx22763z1_rt,
      O => U_DCT2D_databuf_reg_2_10_XORF
    );
  U_DCT2D_databuf_reg_2_10_CYINIT_153 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1580_add_47_ix22763z63342_O,
      O => U_DCT2D_databuf_reg_2_10_CYINIT
    );
  U_DCT2D_databuf_reg_2_10_CLKINV_154 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_2_10_CLKINV
    );
  U_DCT2D_databuf_reg_2_10_CEINV_155 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_2_10_CEINV
    );
  U_DCT2D_databuf_reg_4_0_DXMUX_156 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_0_XORF,
      O => U_DCT2D_databuf_reg_4_0_DXMUX
    );
  U_DCT2D_databuf_reg_4_0_XORF_157 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_0_CYINIT,
      I1 => U_DCT2D_nx49552z1,
      O => U_DCT2D_databuf_reg_4_0_XORF
    );
  U_DCT2D_databuf_reg_4_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_0_CY0F,
      IB => U_DCT2D_databuf_reg_4_0_CYINIT,
      SEL => U_DCT2D_databuf_reg_4_0_CYSELF,
      O => U_DCT2D_rtlc5_97_sub_41_ix50549z63342_O
    );
  U_DCT2D_databuf_reg_4_0_CYINIT_158 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GLOBAL_LOGIC1_23,
      O => U_DCT2D_databuf_reg_4_0_CYINIT
    );
  U_DCT2D_databuf_reg_4_0_CY0F_159 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_0_Q,
      O => U_DCT2D_databuf_reg_4_0_CY0F
    );
  U_DCT2D_databuf_reg_4_0_CYSELF_160 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx49552z1,
      O => U_DCT2D_databuf_reg_4_0_CYSELF
    );
  U_DCT2D_databuf_reg_4_0_DYMUX_161 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_0_XORG,
      O => U_DCT2D_databuf_reg_4_0_DYMUX
    );
  U_DCT2D_databuf_reg_4_0_XORG_162 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_97_sub_41_ix50549z63342_O,
      I1 => U_DCT2D_nx50549z1,
      O => U_DCT2D_databuf_reg_4_0_XORG
    );
  U_DCT2D_databuf_reg_4_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_0_CYMUXG,
      O => U_DCT2D_rtlc5_97_sub_41_ix51546z63342_O
    );
  U_DCT2D_databuf_reg_4_0_CYMUXG_163 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_0_CY0G,
      IB => U_DCT2D_rtlc5_97_sub_41_ix50549z63342_O,
      SEL => U_DCT2D_databuf_reg_4_0_CYSELG,
      O => U_DCT2D_databuf_reg_4_0_CYMUXG
    );
  U_DCT2D_databuf_reg_4_0_CY0G_164 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_1_Q,
      O => U_DCT2D_databuf_reg_4_0_CY0G
    );
  U_DCT2D_databuf_reg_4_0_CYSELG_165 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx50549z1,
      O => U_DCT2D_databuf_reg_4_0_CYSELG
    );
  U_DCT2D_databuf_reg_4_0_SRINV_166 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_4_0_SRINV
    );
  U_DCT2D_databuf_reg_4_0_CLKINV_167 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_4_0_CLKINV
    );
  U_DCT2D_databuf_reg_4_0_CEINV_168 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_4_0_CEINV
    );
  U_DCT2D_databuf_reg_4_2_DXMUX_169 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_2_XORF,
      O => U_DCT2D_databuf_reg_4_2_DXMUX
    );
  U_DCT2D_databuf_reg_4_2_XORF_170 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_2_CYINIT,
      I1 => U_DCT2D_nx51546z1,
      O => U_DCT2D_databuf_reg_4_2_XORF
    );
  U_DCT2D_databuf_reg_4_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_2_CY0F,
      IB => U_DCT2D_databuf_reg_4_2_CYINIT,
      SEL => U_DCT2D_databuf_reg_4_2_CYSELF,
      O => U_DCT2D_rtlc5_97_sub_41_ix52543z63342_O
    );
  U_DCT2D_databuf_reg_4_2_CYMUXF2_171 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_2_CY0F,
      IB => U_DCT2D_databuf_reg_4_2_CY0F,
      SEL => U_DCT2D_databuf_reg_4_2_CYSELF,
      O => U_DCT2D_databuf_reg_4_2_CYMUXF2
    );
  U_DCT2D_databuf_reg_4_2_CYINIT_172 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_97_sub_41_ix51546z63342_O,
      O => U_DCT2D_databuf_reg_4_2_CYINIT
    );
  U_DCT2D_databuf_reg_4_2_CY0F_173 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_2_Q,
      O => U_DCT2D_databuf_reg_4_2_CY0F
    );
  U_DCT2D_databuf_reg_4_2_CYSELF_174 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx51546z1,
      O => U_DCT2D_databuf_reg_4_2_CYSELF
    );
  U_DCT2D_databuf_reg_4_2_DYMUX_175 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_2_XORG,
      O => U_DCT2D_databuf_reg_4_2_DYMUX
    );
  U_DCT2D_databuf_reg_4_2_XORG_176 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_97_sub_41_ix52543z63342_O,
      I1 => U_DCT2D_nx52543z1,
      O => U_DCT2D_databuf_reg_4_2_XORG
    );
  U_DCT2D_databuf_reg_4_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_2_CYMUXFAST,
      O => U_DCT2D_rtlc5_97_sub_41_ix53540z63342_O
    );
  U_DCT2D_databuf_reg_4_2_FASTCARRY_177 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_97_sub_41_ix51546z63342_O,
      O => U_DCT2D_databuf_reg_4_2_FASTCARRY
    );
  U_DCT2D_databuf_reg_4_2_CYAND_178 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_4_2_CYSELG,
      I1 => U_DCT2D_databuf_reg_4_2_CYSELF,
      O => U_DCT2D_databuf_reg_4_2_CYAND
    );
  U_DCT2D_databuf_reg_4_2_CYMUXFAST_179 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_2_CYMUXG2,
      IB => U_DCT2D_databuf_reg_4_2_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_4_2_CYAND,
      O => U_DCT2D_databuf_reg_4_2_CYMUXFAST
    );
  U_DCT2D_databuf_reg_4_2_CYMUXG2_180 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_2_CY0G,
      IB => U_DCT2D_databuf_reg_4_2_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_4_2_CYSELG,
      O => U_DCT2D_databuf_reg_4_2_CYMUXG2
    );
  U_DCT2D_databuf_reg_4_2_CY0G_181 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_3_Q,
      O => U_DCT2D_databuf_reg_4_2_CY0G
    );
  U_DCT2D_databuf_reg_4_2_CYSELG_182 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx52543z1,
      O => U_DCT2D_databuf_reg_4_2_CYSELG
    );
  U_DCT2D_databuf_reg_4_2_SRINV_183 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_4_2_SRINV
    );
  U_DCT2D_databuf_reg_4_2_CLKINV_184 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_4_2_CLKINV
    );
  U_DCT2D_databuf_reg_4_2_CEINV_185 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_4_2_CEINV
    );
  U_DCT2D_databuf_reg_4_4_DXMUX_186 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_4_XORF,
      O => U_DCT2D_databuf_reg_4_4_DXMUX
    );
  U_DCT2D_databuf_reg_4_4_XORF_187 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_4_CYINIT,
      I1 => U_DCT2D_nx53540z1,
      O => U_DCT2D_databuf_reg_4_4_XORF
    );
  U_DCT2D_databuf_reg_4_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_4_CY0F,
      IB => U_DCT2D_databuf_reg_4_4_CYINIT,
      SEL => U_DCT2D_databuf_reg_4_4_CYSELF,
      O => U_DCT2D_rtlc5_97_sub_41_ix54537z63342_O
    );
  U_DCT2D_databuf_reg_4_4_CYMUXF2_188 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_4_CY0F,
      IB => U_DCT2D_databuf_reg_4_4_CY0F,
      SEL => U_DCT2D_databuf_reg_4_4_CYSELF,
      O => U_DCT2D_databuf_reg_4_4_CYMUXF2
    );
  U_DCT2D_databuf_reg_4_4_CYINIT_189 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_97_sub_41_ix53540z63342_O,
      O => U_DCT2D_databuf_reg_4_4_CYINIT
    );
  U_DCT2D_databuf_reg_4_4_CY0F_190 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_4_Q,
      O => U_DCT2D_databuf_reg_4_4_CY0F
    );
  U_DCT2D_databuf_reg_4_4_CYSELF_191 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx53540z1,
      O => U_DCT2D_databuf_reg_4_4_CYSELF
    );
  U_DCT2D_databuf_reg_4_4_DYMUX_192 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_4_XORG,
      O => U_DCT2D_databuf_reg_4_4_DYMUX
    );
  U_DCT2D_databuf_reg_4_4_XORG_193 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_97_sub_41_ix54537z63342_O,
      I1 => U_DCT2D_nx54537z1,
      O => U_DCT2D_databuf_reg_4_4_XORG
    );
  U_DCT2D_databuf_reg_4_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_4_CYMUXFAST,
      O => U_DCT2D_rtlc5_97_sub_41_ix55534z63342_O
    );
  U_DCT2D_databuf_reg_4_4_FASTCARRY_194 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_97_sub_41_ix53540z63342_O,
      O => U_DCT2D_databuf_reg_4_4_FASTCARRY
    );
  U_DCT2D_databuf_reg_4_4_CYAND_195 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_4_4_CYSELG,
      I1 => U_DCT2D_databuf_reg_4_4_CYSELF,
      O => U_DCT2D_databuf_reg_4_4_CYAND
    );
  U_DCT2D_databuf_reg_4_4_CYMUXFAST_196 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_4_CYMUXG2,
      IB => U_DCT2D_databuf_reg_4_4_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_4_4_CYAND,
      O => U_DCT2D_databuf_reg_4_4_CYMUXFAST
    );
  U_DCT2D_databuf_reg_4_4_CYMUXG2_197 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_4_CY0G,
      IB => U_DCT2D_databuf_reg_4_4_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_4_4_CYSELG,
      O => U_DCT2D_databuf_reg_4_4_CYMUXG2
    );
  U_DCT2D_databuf_reg_4_4_CY0G_198 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_5_Q,
      O => U_DCT2D_databuf_reg_4_4_CY0G
    );
  U_DCT2D_databuf_reg_4_4_CYSELG_199 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx54537z1,
      O => U_DCT2D_databuf_reg_4_4_CYSELG
    );
  U_DCT2D_databuf_reg_4_4_SRINV_200 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_4_4_SRINV
    );
  U_DCT2D_databuf_reg_4_4_CLKINV_201 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_4_4_CLKINV
    );
  U_DCT2D_databuf_reg_4_4_CEINV_202 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_4_4_CEINV
    );
  U_DCT2D_databuf_reg_4_6_DXMUX_203 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_6_XORF,
      O => U_DCT2D_databuf_reg_4_6_DXMUX
    );
  U_DCT2D_databuf_reg_4_6_XORF_204 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_6_CYINIT,
      I1 => U_DCT2D_nx55534z1,
      O => U_DCT2D_databuf_reg_4_6_XORF
    );
  U_DCT2D_databuf_reg_4_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_6_CY0F,
      IB => U_DCT2D_databuf_reg_4_6_CYINIT,
      SEL => U_DCT2D_databuf_reg_4_6_CYSELF,
      O => U_DCT2D_rtlc5_97_sub_41_ix56531z63342_O
    );
  U_DCT2D_databuf_reg_4_6_CYMUXF2_205 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_6_CY0F,
      IB => U_DCT2D_databuf_reg_4_6_CY0F,
      SEL => U_DCT2D_databuf_reg_4_6_CYSELF,
      O => U_DCT2D_databuf_reg_4_6_CYMUXF2
    );
  U_DCT2D_databuf_reg_4_6_CYINIT_206 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_97_sub_41_ix55534z63342_O,
      O => U_DCT2D_databuf_reg_4_6_CYINIT
    );
  U_DCT2D_databuf_reg_4_6_CY0F_207 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_6_Q,
      O => U_DCT2D_databuf_reg_4_6_CY0F
    );
  U_DCT2D_databuf_reg_4_6_CYSELF_208 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx55534z1,
      O => U_DCT2D_databuf_reg_4_6_CYSELF
    );
  U_DCT2D_databuf_reg_4_6_DYMUX_209 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_6_XORG,
      O => U_DCT2D_databuf_reg_4_6_DYMUX
    );
  U_DCT2D_databuf_reg_4_6_XORG_210 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_97_sub_41_ix56531z63342_O,
      I1 => U_DCT2D_nx56531z1,
      O => U_DCT2D_databuf_reg_4_6_XORG
    );
  U_DCT2D_databuf_reg_4_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_6_CYMUXFAST,
      O => U_DCT2D_rtlc5_97_sub_41_ix57528z63342_O
    );
  U_DCT2D_databuf_reg_4_6_FASTCARRY_211 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_97_sub_41_ix55534z63342_O,
      O => U_DCT2D_databuf_reg_4_6_FASTCARRY
    );
  U_DCT2D_databuf_reg_4_6_CYAND_212 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_4_6_CYSELG,
      I1 => U_DCT2D_databuf_reg_4_6_CYSELF,
      O => U_DCT2D_databuf_reg_4_6_CYAND
    );
  U_DCT2D_databuf_reg_4_6_CYMUXFAST_213 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_6_CYMUXG2,
      IB => U_DCT2D_databuf_reg_4_6_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_4_6_CYAND,
      O => U_DCT2D_databuf_reg_4_6_CYMUXFAST
    );
  U_DCT2D_databuf_reg_4_6_CYMUXG2_214 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_6_CY0G,
      IB => U_DCT2D_databuf_reg_4_6_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_4_6_CYSELG,
      O => U_DCT2D_databuf_reg_4_6_CYMUXG2
    );
  U_DCT2D_databuf_reg_4_6_CY0G_215 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_7_Q,
      O => U_DCT2D_databuf_reg_4_6_CY0G
    );
  U_DCT2D_databuf_reg_4_6_CYSELG_216 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx56531z1,
      O => U_DCT2D_databuf_reg_4_6_CYSELG
    );
  U_DCT2D_databuf_reg_4_6_SRINV_217 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_4_6_SRINV
    );
  U_DCT2D_databuf_reg_4_6_CLKINV_218 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_4_6_CLKINV
    );
  U_DCT2D_databuf_reg_4_6_CEINV_219 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_4_6_CEINV
    );
  U_DCT2D_databuf_reg_4_8_DXMUX_220 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_8_XORF,
      O => U_DCT2D_databuf_reg_4_8_DXMUX
    );
  U_DCT2D_databuf_reg_4_8_XORF_221 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_8_CYINIT,
      I1 => U_DCT2D_nx57528z1,
      O => U_DCT2D_databuf_reg_4_8_XORF
    );
  U_DCT2D_databuf_reg_4_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_8_CY0F,
      IB => U_DCT2D_databuf_reg_4_8_CYINIT,
      SEL => U_DCT2D_databuf_reg_4_8_CYSELF,
      O => U_DCT2D_rtlc5_97_sub_41_ix58525z63342_O
    );
  U_DCT2D_databuf_reg_4_8_CYMUXF2_222 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_8_CY0F,
      IB => U_DCT2D_databuf_reg_4_8_CY0F,
      SEL => U_DCT2D_databuf_reg_4_8_CYSELF,
      O => U_DCT2D_databuf_reg_4_8_CYMUXF2
    );
  U_DCT2D_databuf_reg_4_8_CYINIT_223 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_97_sub_41_ix57528z63342_O,
      O => U_DCT2D_databuf_reg_4_8_CYINIT
    );
  U_DCT2D_databuf_reg_4_8_CY0F_224 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_8_Q,
      O => U_DCT2D_databuf_reg_4_8_CY0F
    );
  U_DCT2D_databuf_reg_4_8_CYSELF_225 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx57528z1,
      O => U_DCT2D_databuf_reg_4_8_CYSELF
    );
  U_DCT2D_databuf_reg_4_8_DYMUX_226 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_8_XORG,
      O => U_DCT2D_databuf_reg_4_8_DYMUX
    );
  U_DCT2D_databuf_reg_4_8_XORG_227 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_97_sub_41_ix58525z63342_O,
      I1 => U_DCT2D_nx58525z1,
      O => U_DCT2D_databuf_reg_4_8_XORG
    );
  U_DCT2D_databuf_reg_4_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_8_CYMUXFAST,
      O => U_DCT2D_rtlc5_97_sub_41_ix7189z63342_O
    );
  U_DCT2D_databuf_reg_4_8_FASTCARRY_228 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_97_sub_41_ix57528z63342_O,
      O => U_DCT2D_databuf_reg_4_8_FASTCARRY
    );
  U_DCT2D_databuf_reg_4_8_CYAND_229 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_4_8_CYSELG,
      I1 => U_DCT2D_databuf_reg_4_8_CYSELF,
      O => U_DCT2D_databuf_reg_4_8_CYAND
    );
  U_DCT2D_databuf_reg_4_8_CYMUXFAST_230 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_8_CYMUXG2,
      IB => U_DCT2D_databuf_reg_4_8_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_4_8_CYAND,
      O => U_DCT2D_databuf_reg_4_8_CYMUXFAST
    );
  U_DCT2D_databuf_reg_4_8_CYMUXG2_231 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_4_8_CY0G,
      IB => U_DCT2D_databuf_reg_4_8_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_4_8_CYSELG,
      O => U_DCT2D_databuf_reg_4_8_CYMUXG2
    );
  U_DCT2D_databuf_reg_4_8_CY0G_232 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_10_Q,
      O => U_DCT2D_databuf_reg_4_8_CY0G
    );
  U_DCT2D_databuf_reg_4_8_CYSELG_233 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx58525z1,
      O => U_DCT2D_databuf_reg_4_8_CYSELG
    );
  U_DCT2D_databuf_reg_4_8_SRINV_234 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_4_8_SRINV
    );
  U_DCT2D_databuf_reg_4_8_CLKINV_235 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_4_8_CLKINV
    );
  U_DCT2D_databuf_reg_4_8_CEINV_236 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_4_8_CEINV
    );
  U_DCT2D_nx7189z1_rt_237 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT2D_nx7189z1,
      ADR3 => VCC,
      O => U_DCT2D_nx7189z1_rt
    );
  U_DCT2D_databuf_reg_4_10_DXMUX_238 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_10_XORF,
      O => U_DCT2D_databuf_reg_4_10_DXMUX
    );
  U_DCT2D_databuf_reg_4_10_XORF_239 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_10_CYINIT,
      I1 => U_DCT2D_nx7189z1_rt,
      O => U_DCT2D_databuf_reg_4_10_XORF
    );
  U_DCT2D_databuf_reg_4_10_CYINIT_240 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_97_sub_41_ix7189z63342_O,
      O => U_DCT2D_databuf_reg_4_10_CYINIT
    );
  U_DCT2D_databuf_reg_4_10_CLKINV_241 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_4_10_CLKINV
    );
  U_DCT2D_databuf_reg_4_10_CEINV_242 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_4_10_CEINV
    );
  U_DCT2D_databuf_reg_7_0_DXMUX_243 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_0_XORF,
      O => U_DCT2D_databuf_reg_7_0_DXMUX
    );
  U_DCT2D_databuf_reg_7_0_XORF_244 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_0_CYINIT,
      I1 => U_DCT2D_nx34147z1,
      O => U_DCT2D_databuf_reg_7_0_XORF
    );
  U_DCT2D_databuf_reg_7_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_0_CY0F,
      IB => U_DCT2D_databuf_reg_7_0_CYINIT,
      SEL => U_DCT2D_databuf_reg_7_0_CYSELF,
      O => U_DCT2D_rtlc5_100_sub_44_ix35144z63342_O
    );
  U_DCT2D_databuf_reg_7_0_CYINIT_245 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GLOBAL_LOGIC1_28,
      O => U_DCT2D_databuf_reg_7_0_CYINIT
    );
  U_DCT2D_databuf_reg_7_0_CY0F_246 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_0_Q,
      O => U_DCT2D_databuf_reg_7_0_CY0F
    );
  U_DCT2D_databuf_reg_7_0_CYSELF_247 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx34147z1,
      O => U_DCT2D_databuf_reg_7_0_CYSELF
    );
  U_DCT2D_databuf_reg_7_0_DYMUX_248 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_0_XORG,
      O => U_DCT2D_databuf_reg_7_0_DYMUX
    );
  U_DCT2D_databuf_reg_7_0_XORG_249 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_100_sub_44_ix35144z63342_O,
      I1 => U_DCT2D_nx35144z1,
      O => U_DCT2D_databuf_reg_7_0_XORG
    );
  U_DCT2D_databuf_reg_7_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_0_CYMUXG,
      O => U_DCT2D_rtlc5_100_sub_44_ix36141z63342_O
    );
  U_DCT2D_databuf_reg_7_0_CYMUXG_250 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_0_CY0G,
      IB => U_DCT2D_rtlc5_100_sub_44_ix35144z63342_O,
      SEL => U_DCT2D_databuf_reg_7_0_CYSELG,
      O => U_DCT2D_databuf_reg_7_0_CYMUXG
    );
  U_DCT2D_databuf_reg_7_0_CY0G_251 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_1_Q,
      O => U_DCT2D_databuf_reg_7_0_CY0G
    );
  U_DCT2D_databuf_reg_7_0_CYSELG_252 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx35144z1,
      O => U_DCT2D_databuf_reg_7_0_CYSELG
    );
  U_DCT2D_databuf_reg_7_0_SRINV_253 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_7_0_SRINV
    );
  U_DCT2D_databuf_reg_7_0_CLKINV_254 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_7_0_CLKINV
    );
  U_DCT2D_databuf_reg_7_0_CEINV_255 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_7_0_CEINV
    );
  U_DCT2D_databuf_reg_7_2_DXMUX_256 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_2_XORF,
      O => U_DCT2D_databuf_reg_7_2_DXMUX
    );
  U_DCT2D_databuf_reg_7_2_XORF_257 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_2_CYINIT,
      I1 => U_DCT2D_nx36141z1,
      O => U_DCT2D_databuf_reg_7_2_XORF
    );
  U_DCT2D_databuf_reg_7_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_2_CY0F,
      IB => U_DCT2D_databuf_reg_7_2_CYINIT,
      SEL => U_DCT2D_databuf_reg_7_2_CYSELF,
      O => U_DCT2D_rtlc5_100_sub_44_ix37138z63342_O
    );
  U_DCT2D_databuf_reg_7_2_CYMUXF2_258 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_2_CY0F,
      IB => U_DCT2D_databuf_reg_7_2_CY0F,
      SEL => U_DCT2D_databuf_reg_7_2_CYSELF,
      O => U_DCT2D_databuf_reg_7_2_CYMUXF2
    );
  U_DCT2D_databuf_reg_7_2_CYINIT_259 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_100_sub_44_ix36141z63342_O,
      O => U_DCT2D_databuf_reg_7_2_CYINIT
    );
  U_DCT2D_databuf_reg_7_2_CY0F_260 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_2_Q,
      O => U_DCT2D_databuf_reg_7_2_CY0F
    );
  U_DCT2D_databuf_reg_7_2_CYSELF_261 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx36141z1,
      O => U_DCT2D_databuf_reg_7_2_CYSELF
    );
  U_DCT2D_databuf_reg_7_2_DYMUX_262 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_2_XORG,
      O => U_DCT2D_databuf_reg_7_2_DYMUX
    );
  U_DCT2D_databuf_reg_7_2_XORG_263 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_100_sub_44_ix37138z63342_O,
      I1 => U_DCT2D_nx37138z1,
      O => U_DCT2D_databuf_reg_7_2_XORG
    );
  U_DCT2D_databuf_reg_7_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_2_CYMUXFAST,
      O => U_DCT2D_rtlc5_100_sub_44_ix38135z63342_O
    );
  U_DCT2D_databuf_reg_7_2_FASTCARRY_264 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_100_sub_44_ix36141z63342_O,
      O => U_DCT2D_databuf_reg_7_2_FASTCARRY
    );
  U_DCT2D_databuf_reg_7_2_CYAND_265 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_7_2_CYSELG,
      I1 => U_DCT2D_databuf_reg_7_2_CYSELF,
      O => U_DCT2D_databuf_reg_7_2_CYAND
    );
  U_DCT2D_databuf_reg_7_2_CYMUXFAST_266 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_2_CYMUXG2,
      IB => U_DCT2D_databuf_reg_7_2_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_7_2_CYAND,
      O => U_DCT2D_databuf_reg_7_2_CYMUXFAST
    );
  U_DCT2D_databuf_reg_7_2_CYMUXG2_267 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_2_CY0G,
      IB => U_DCT2D_databuf_reg_7_2_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_7_2_CYSELG,
      O => U_DCT2D_databuf_reg_7_2_CYMUXG2
    );
  U_DCT2D_databuf_reg_7_2_CY0G_268 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_3_Q,
      O => U_DCT2D_databuf_reg_7_2_CY0G
    );
  U_DCT2D_databuf_reg_7_2_CYSELG_269 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx37138z1,
      O => U_DCT2D_databuf_reg_7_2_CYSELG
    );
  U_DCT2D_databuf_reg_7_2_SRINV_270 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_7_2_SRINV
    );
  U_DCT2D_databuf_reg_7_2_CLKINV_271 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_7_2_CLKINV
    );
  U_DCT2D_databuf_reg_7_2_CEINV_272 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_7_2_CEINV
    );
  U_DCT1D_ix59822z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_2_Q(0),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_5_Q(0),
      O => U_DCT1D_nx59822z1
    );
  U_DCT2D_databuf_reg_7_4_DXMUX_273 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_4_XORF,
      O => U_DCT2D_databuf_reg_7_4_DXMUX
    );
  U_DCT2D_databuf_reg_7_4_XORF_274 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_4_CYINIT,
      I1 => U_DCT2D_nx38135z1,
      O => U_DCT2D_databuf_reg_7_4_XORF
    );
  U_DCT2D_databuf_reg_7_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_4_CY0F,
      IB => U_DCT2D_databuf_reg_7_4_CYINIT,
      SEL => U_DCT2D_databuf_reg_7_4_CYSELF,
      O => U_DCT2D_rtlc5_100_sub_44_ix39132z63342_O
    );
  U_DCT2D_databuf_reg_7_4_CYMUXF2_275 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_4_CY0F,
      IB => U_DCT2D_databuf_reg_7_4_CY0F,
      SEL => U_DCT2D_databuf_reg_7_4_CYSELF,
      O => U_DCT2D_databuf_reg_7_4_CYMUXF2
    );
  U_DCT2D_databuf_reg_7_4_CYINIT_276 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_100_sub_44_ix38135z63342_O,
      O => U_DCT2D_databuf_reg_7_4_CYINIT
    );
  U_DCT2D_databuf_reg_7_4_CY0F_277 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_4_Q,
      O => U_DCT2D_databuf_reg_7_4_CY0F
    );
  U_DCT2D_databuf_reg_7_4_CYSELF_278 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx38135z1,
      O => U_DCT2D_databuf_reg_7_4_CYSELF
    );
  U_DCT2D_databuf_reg_7_4_DYMUX_279 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_4_XORG,
      O => U_DCT2D_databuf_reg_7_4_DYMUX
    );
  U_DCT2D_databuf_reg_7_4_XORG_280 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_100_sub_44_ix39132z63342_O,
      I1 => U_DCT2D_nx39132z1,
      O => U_DCT2D_databuf_reg_7_4_XORG
    );
  U_DCT2D_databuf_reg_7_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_4_CYMUXFAST,
      O => U_DCT2D_rtlc5_100_sub_44_ix40129z63342_O
    );
  U_DCT2D_databuf_reg_7_4_FASTCARRY_281 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_100_sub_44_ix38135z63342_O,
      O => U_DCT2D_databuf_reg_7_4_FASTCARRY
    );
  U_DCT2D_databuf_reg_7_4_CYAND_282 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_7_4_CYSELG,
      I1 => U_DCT2D_databuf_reg_7_4_CYSELF,
      O => U_DCT2D_databuf_reg_7_4_CYAND
    );
  U_DCT2D_databuf_reg_7_4_CYMUXFAST_283 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_4_CYMUXG2,
      IB => U_DCT2D_databuf_reg_7_4_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_7_4_CYAND,
      O => U_DCT2D_databuf_reg_7_4_CYMUXFAST
    );
  U_DCT2D_databuf_reg_7_4_CYMUXG2_284 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_4_CY0G,
      IB => U_DCT2D_databuf_reg_7_4_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_7_4_CYSELG,
      O => U_DCT2D_databuf_reg_7_4_CYMUXG2
    );
  U_DCT2D_databuf_reg_7_4_CY0G_285 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_5_Q,
      O => U_DCT2D_databuf_reg_7_4_CY0G
    );
  U_DCT2D_databuf_reg_7_4_CYSELG_286 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx39132z1,
      O => U_DCT2D_databuf_reg_7_4_CYSELG
    );
  U_DCT2D_databuf_reg_7_4_SRINV_287 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_7_4_SRINV
    );
  U_DCT2D_databuf_reg_7_4_CLKINV_288 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_7_4_CLKINV
    );
  U_DCT2D_databuf_reg_7_4_CEINV_289 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_7_4_CEINV
    );
  U_DCT2D_databuf_reg_7_6_DXMUX_290 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_6_XORF,
      O => U_DCT2D_databuf_reg_7_6_DXMUX
    );
  U_DCT2D_databuf_reg_7_6_XORF_291 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_6_CYINIT,
      I1 => U_DCT2D_nx40129z1,
      O => U_DCT2D_databuf_reg_7_6_XORF
    );
  U_DCT2D_databuf_reg_7_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_6_CY0F,
      IB => U_DCT2D_databuf_reg_7_6_CYINIT,
      SEL => U_DCT2D_databuf_reg_7_6_CYSELF,
      O => U_DCT2D_rtlc5_100_sub_44_ix41126z63342_O
    );
  U_DCT2D_databuf_reg_7_6_CYMUXF2_292 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_6_CY0F,
      IB => U_DCT2D_databuf_reg_7_6_CY0F,
      SEL => U_DCT2D_databuf_reg_7_6_CYSELF,
      O => U_DCT2D_databuf_reg_7_6_CYMUXF2
    );
  U_DCT2D_databuf_reg_7_6_CYINIT_293 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_100_sub_44_ix40129z63342_O,
      O => U_DCT2D_databuf_reg_7_6_CYINIT
    );
  U_DCT2D_databuf_reg_7_6_CY0F_294 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_6_Q,
      O => U_DCT2D_databuf_reg_7_6_CY0F
    );
  U_DCT2D_databuf_reg_7_6_CYSELF_295 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx40129z1,
      O => U_DCT2D_databuf_reg_7_6_CYSELF
    );
  U_DCT2D_databuf_reg_7_6_DYMUX_296 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_6_XORG,
      O => U_DCT2D_databuf_reg_7_6_DYMUX
    );
  U_DCT2D_databuf_reg_7_6_XORG_297 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_100_sub_44_ix41126z63342_O,
      I1 => U_DCT2D_nx41126z1,
      O => U_DCT2D_databuf_reg_7_6_XORG
    );
  U_DCT2D_databuf_reg_7_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_6_CYMUXFAST,
      O => U_DCT2D_rtlc5_100_sub_44_ix42123z63342_O
    );
  U_DCT2D_databuf_reg_7_6_FASTCARRY_298 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_100_sub_44_ix40129z63342_O,
      O => U_DCT2D_databuf_reg_7_6_FASTCARRY
    );
  U_DCT2D_databuf_reg_7_6_CYAND_299 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_7_6_CYSELG,
      I1 => U_DCT2D_databuf_reg_7_6_CYSELF,
      O => U_DCT2D_databuf_reg_7_6_CYAND
    );
  U_DCT2D_databuf_reg_7_6_CYMUXFAST_300 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_6_CYMUXG2,
      IB => U_DCT2D_databuf_reg_7_6_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_7_6_CYAND,
      O => U_DCT2D_databuf_reg_7_6_CYMUXFAST
    );
  U_DCT2D_databuf_reg_7_6_CYMUXG2_301 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_6_CY0G,
      IB => U_DCT2D_databuf_reg_7_6_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_7_6_CYSELG,
      O => U_DCT2D_databuf_reg_7_6_CYMUXG2
    );
  U_DCT2D_databuf_reg_7_6_CY0G_302 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_7_Q,
      O => U_DCT2D_databuf_reg_7_6_CY0G
    );
  U_DCT2D_databuf_reg_7_6_CYSELG_303 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx41126z1,
      O => U_DCT2D_databuf_reg_7_6_CYSELG
    );
  U_DCT2D_databuf_reg_7_6_SRINV_304 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_7_6_SRINV
    );
  U_DCT2D_databuf_reg_7_6_CLKINV_305 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_7_6_CLKINV
    );
  U_DCT2D_databuf_reg_7_6_CEINV_306 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_7_6_CEINV
    );
  U_DCT2D_databuf_reg_7_8_DXMUX_307 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_8_XORF,
      O => U_DCT2D_databuf_reg_7_8_DXMUX
    );
  U_DCT2D_databuf_reg_7_8_XORF_308 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_8_CYINIT,
      I1 => U_DCT2D_nx42123z1,
      O => U_DCT2D_databuf_reg_7_8_XORF
    );
  U_DCT2D_databuf_reg_7_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_8_CY0F,
      IB => U_DCT2D_databuf_reg_7_8_CYINIT,
      SEL => U_DCT2D_databuf_reg_7_8_CYSELF,
      O => U_DCT2D_rtlc5_100_sub_44_ix43120z63342_O
    );
  U_DCT2D_databuf_reg_7_8_CYMUXF2_309 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_8_CY0F,
      IB => U_DCT2D_databuf_reg_7_8_CY0F,
      SEL => U_DCT2D_databuf_reg_7_8_CYSELF,
      O => U_DCT2D_databuf_reg_7_8_CYMUXF2
    );
  U_DCT2D_databuf_reg_7_8_CYINIT_310 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_100_sub_44_ix42123z63342_O,
      O => U_DCT2D_databuf_reg_7_8_CYINIT
    );
  U_DCT2D_databuf_reg_7_8_CY0F_311 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_8_Q,
      O => U_DCT2D_databuf_reg_7_8_CY0F
    );
  U_DCT2D_databuf_reg_7_8_CYSELF_312 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx42123z1,
      O => U_DCT2D_databuf_reg_7_8_CYSELF
    );
  U_DCT2D_databuf_reg_7_8_DYMUX_313 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_8_XORG,
      O => U_DCT2D_databuf_reg_7_8_DYMUX
    );
  U_DCT2D_databuf_reg_7_8_XORG_314 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_100_sub_44_ix43120z63342_O,
      I1 => U_DCT2D_nx43120z1,
      O => U_DCT2D_databuf_reg_7_8_XORG
    );
  U_DCT2D_databuf_reg_7_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_8_CYMUXFAST,
      O => U_DCT2D_rtlc5_100_sub_44_ix16172z63342_O
    );
  U_DCT2D_databuf_reg_7_8_FASTCARRY_315 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_100_sub_44_ix42123z63342_O,
      O => U_DCT2D_databuf_reg_7_8_FASTCARRY
    );
  U_DCT2D_databuf_reg_7_8_CYAND_316 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_7_8_CYSELG,
      I1 => U_DCT2D_databuf_reg_7_8_CYSELF,
      O => U_DCT2D_databuf_reg_7_8_CYAND
    );
  U_DCT2D_databuf_reg_7_8_CYMUXFAST_317 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_8_CYMUXG2,
      IB => U_DCT2D_databuf_reg_7_8_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_7_8_CYAND,
      O => U_DCT2D_databuf_reg_7_8_CYMUXFAST
    );
  U_DCT2D_databuf_reg_7_8_CYMUXG2_318 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_7_8_CY0G,
      IB => U_DCT2D_databuf_reg_7_8_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_7_8_CYSELG,
      O => U_DCT2D_databuf_reg_7_8_CYMUXG2
    );
  U_DCT2D_databuf_reg_7_8_CY0G_319 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_10_Q,
      O => U_DCT2D_databuf_reg_7_8_CY0G
    );
  U_DCT2D_databuf_reg_7_8_CYSELG_320 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx43120z1,
      O => U_DCT2D_databuf_reg_7_8_CYSELG
    );
  U_DCT2D_databuf_reg_7_8_SRINV_321 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_7_8_SRINV
    );
  U_DCT2D_databuf_reg_7_8_CLKINV_322 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_7_8_CLKINV
    );
  U_DCT2D_databuf_reg_7_8_CEINV_323 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_7_8_CEINV
    );
  U_DCT2D_nx16172z1_rt_324 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT2D_nx16172z1,
      ADR3 => VCC,
      O => U_DCT2D_nx16172z1_rt
    );
  U_DCT2D_databuf_reg_7_10_DXMUX_325 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_10_XORF,
      O => U_DCT2D_databuf_reg_7_10_DXMUX
    );
  U_DCT2D_databuf_reg_7_10_XORF_326 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_10_CYINIT,
      I1 => U_DCT2D_nx16172z1_rt,
      O => U_DCT2D_databuf_reg_7_10_XORF
    );
  U_DCT2D_databuf_reg_7_10_CYINIT_327 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_100_sub_44_ix16172z63342_O,
      O => U_DCT2D_databuf_reg_7_10_CYINIT
    );
  U_DCT2D_databuf_reg_7_10_CLKINV_328 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_7_10_CLKINV
    );
  U_DCT2D_databuf_reg_7_10_CEINV_329 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_7_10_CEINV
    );
  U_DCT1D_databuf_reg_1_0_DXMUX_330 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_0_XORF,
      O => U_DCT1D_databuf_reg_1_0_DXMUX
    );
  U_DCT1D_databuf_reg_1_0_XORF_331 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_0_CYINIT,
      I1 => U_DCT1D_nx64957z1,
      O => U_DCT1D_databuf_reg_1_0_XORF
    );
  U_DCT1D_databuf_reg_1_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_0_CY0F,
      IB => U_DCT1D_databuf_reg_1_0_CYINIT,
      SEL => U_DCT1D_databuf_reg_1_0_CYSELF,
      O => U_DCT1D_rtlc5_1420_add_9_ix418z63342_O
    );
  U_DCT1D_databuf_reg_1_0_CYINIT_332 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_0_BXINVNOT,
      O => U_DCT1D_databuf_reg_1_0_CYINIT
    );
  U_DCT1D_databuf_reg_1_0_CY0F_333 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(0),
      O => U_DCT1D_databuf_reg_1_0_CY0F
    );
  U_DCT1D_databuf_reg_1_0_CYSELF_334 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx64957z1,
      O => U_DCT1D_databuf_reg_1_0_CYSELF
    );
  U_DCT1D_databuf_reg_1_0_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_12,
      O => U_DCT1D_databuf_reg_1_0_BXINVNOT
    );
  U_DCT1D_databuf_reg_1_0_DYMUX_335 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_0_XORG,
      O => U_DCT1D_databuf_reg_1_0_DYMUX
    );
  U_DCT1D_databuf_reg_1_0_XORG_336 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1420_add_9_ix418z63342_O,
      I1 => U_DCT1D_nx418z1,
      O => U_DCT1D_databuf_reg_1_0_XORG
    );
  U_DCT1D_databuf_reg_1_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_0_CYMUXG,
      O => U_DCT1D_rtlc5_1420_add_9_ix1415z63342_O
    );
  U_DCT1D_databuf_reg_1_0_CYMUXG_337 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_0_CY0G,
      IB => U_DCT1D_rtlc5_1420_add_9_ix418z63342_O,
      SEL => U_DCT1D_databuf_reg_1_0_CYSELG,
      O => U_DCT1D_databuf_reg_1_0_CYMUXG
    );
  U_DCT1D_databuf_reg_1_0_CY0G_338 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(1),
      O => U_DCT1D_databuf_reg_1_0_CY0G
    );
  U_DCT1D_databuf_reg_1_0_CYSELG_339 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx418z1,
      O => U_DCT1D_databuf_reg_1_0_CYSELG
    );
  U_DCT1D_databuf_reg_1_0_SRINV_340 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_1_0_SRINV
    );
  U_DCT1D_databuf_reg_1_0_CLKINV_341 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_1_0_CLKINV
    );
  U_DCT1D_databuf_reg_1_0_CEINV_342 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_1_0_CEINV
    );
  U_DCT1D_databuf_reg_1_2_DXMUX_343 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_2_XORF,
      O => U_DCT1D_databuf_reg_1_2_DXMUX
    );
  U_DCT1D_databuf_reg_1_2_XORF_344 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_2_CYINIT,
      I1 => U_DCT1D_nx1415z1,
      O => U_DCT1D_databuf_reg_1_2_XORF
    );
  U_DCT1D_databuf_reg_1_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_2_CY0F,
      IB => U_DCT1D_databuf_reg_1_2_CYINIT,
      SEL => U_DCT1D_databuf_reg_1_2_CYSELF,
      O => U_DCT1D_rtlc5_1420_add_9_ix2412z63342_O
    );
  U_DCT1D_databuf_reg_1_2_CYMUXF2_345 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_2_CY0F,
      IB => U_DCT1D_databuf_reg_1_2_CY0F,
      SEL => U_DCT1D_databuf_reg_1_2_CYSELF,
      O => U_DCT1D_databuf_reg_1_2_CYMUXF2
    );
  U_DCT1D_databuf_reg_1_2_CYINIT_346 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1420_add_9_ix1415z63342_O,
      O => U_DCT1D_databuf_reg_1_2_CYINIT
    );
  U_DCT1D_databuf_reg_1_2_CY0F_347 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(2),
      O => U_DCT1D_databuf_reg_1_2_CY0F
    );
  U_DCT1D_databuf_reg_1_2_CYSELF_348 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx1415z1,
      O => U_DCT1D_databuf_reg_1_2_CYSELF
    );
  U_DCT1D_databuf_reg_1_2_DYMUX_349 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_2_XORG,
      O => U_DCT1D_databuf_reg_1_2_DYMUX
    );
  U_DCT1D_databuf_reg_1_2_XORG_350 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1420_add_9_ix2412z63342_O,
      I1 => U_DCT1D_nx2412z1,
      O => U_DCT1D_databuf_reg_1_2_XORG
    );
  U_DCT1D_databuf_reg_1_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_2_CYMUXFAST,
      O => U_DCT1D_rtlc5_1420_add_9_ix3409z63342_O
    );
  U_DCT1D_databuf_reg_1_2_FASTCARRY_351 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1420_add_9_ix1415z63342_O,
      O => U_DCT1D_databuf_reg_1_2_FASTCARRY
    );
  U_DCT1D_databuf_reg_1_2_CYAND_352 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_1_2_CYSELG,
      I1 => U_DCT1D_databuf_reg_1_2_CYSELF,
      O => U_DCT1D_databuf_reg_1_2_CYAND
    );
  U_DCT1D_databuf_reg_1_2_CYMUXFAST_353 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_2_CYMUXG2,
      IB => U_DCT1D_databuf_reg_1_2_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_1_2_CYAND,
      O => U_DCT1D_databuf_reg_1_2_CYMUXFAST
    );
  U_DCT1D_databuf_reg_1_2_CYMUXG2_354 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_2_CY0G,
      IB => U_DCT1D_databuf_reg_1_2_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_1_2_CYSELG,
      O => U_DCT1D_databuf_reg_1_2_CYMUXG2
    );
  U_DCT1D_databuf_reg_1_2_CY0G_355 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(3),
      O => U_DCT1D_databuf_reg_1_2_CY0G
    );
  U_DCT1D_databuf_reg_1_2_CYSELG_356 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx2412z1,
      O => U_DCT1D_databuf_reg_1_2_CYSELG
    );
  U_DCT1D_databuf_reg_1_2_SRINV_357 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_1_2_SRINV
    );
  U_DCT1D_databuf_reg_1_2_CLKINV_358 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_1_2_CLKINV
    );
  U_DCT1D_databuf_reg_1_2_CEINV_359 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_1_2_CEINV
    );
  U_DCT1D_databuf_reg_1_4_DXMUX_360 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_4_XORF,
      O => U_DCT1D_databuf_reg_1_4_DXMUX
    );
  U_DCT1D_databuf_reg_1_4_XORF_361 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_4_CYINIT,
      I1 => U_DCT1D_nx3409z1,
      O => U_DCT1D_databuf_reg_1_4_XORF
    );
  U_DCT1D_databuf_reg_1_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_4_CY0F,
      IB => U_DCT1D_databuf_reg_1_4_CYINIT,
      SEL => U_DCT1D_databuf_reg_1_4_CYSELF,
      O => U_DCT1D_rtlc5_1420_add_9_ix4406z63342_O
    );
  U_DCT1D_databuf_reg_1_4_CYMUXF2_362 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_4_CY0F,
      IB => U_DCT1D_databuf_reg_1_4_CY0F,
      SEL => U_DCT1D_databuf_reg_1_4_CYSELF,
      O => U_DCT1D_databuf_reg_1_4_CYMUXF2
    );
  U_DCT1D_databuf_reg_1_4_CYINIT_363 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1420_add_9_ix3409z63342_O,
      O => U_DCT1D_databuf_reg_1_4_CYINIT
    );
  U_DCT1D_databuf_reg_1_4_CY0F_364 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(4),
      O => U_DCT1D_databuf_reg_1_4_CY0F
    );
  U_DCT1D_databuf_reg_1_4_CYSELF_365 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx3409z1,
      O => U_DCT1D_databuf_reg_1_4_CYSELF
    );
  U_DCT1D_databuf_reg_1_4_DYMUX_366 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_4_XORG,
      O => U_DCT1D_databuf_reg_1_4_DYMUX
    );
  U_DCT1D_databuf_reg_1_4_XORG_367 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1420_add_9_ix4406z63342_O,
      I1 => U_DCT1D_nx4406z1,
      O => U_DCT1D_databuf_reg_1_4_XORG
    );
  U_DCT1D_databuf_reg_1_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_4_CYMUXFAST,
      O => U_DCT1D_rtlc5_1420_add_9_ix5403z63342_O
    );
  U_DCT1D_databuf_reg_1_4_FASTCARRY_368 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1420_add_9_ix3409z63342_O,
      O => U_DCT1D_databuf_reg_1_4_FASTCARRY
    );
  U_DCT1D_databuf_reg_1_4_CYAND_369 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_1_4_CYSELG,
      I1 => U_DCT1D_databuf_reg_1_4_CYSELF,
      O => U_DCT1D_databuf_reg_1_4_CYAND
    );
  U_DCT1D_databuf_reg_1_4_CYMUXFAST_370 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_4_CYMUXG2,
      IB => U_DCT1D_databuf_reg_1_4_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_1_4_CYAND,
      O => U_DCT1D_databuf_reg_1_4_CYMUXFAST
    );
  U_DCT1D_databuf_reg_1_4_CYMUXG2_371 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_4_CY0G,
      IB => U_DCT1D_databuf_reg_1_4_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_1_4_CYSELG,
      O => U_DCT1D_databuf_reg_1_4_CYMUXG2
    );
  U_DCT1D_databuf_reg_1_4_CY0G_372 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(5),
      O => U_DCT1D_databuf_reg_1_4_CY0G
    );
  U_DCT1D_databuf_reg_1_4_CYSELG_373 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx4406z1,
      O => U_DCT1D_databuf_reg_1_4_CYSELG
    );
  U_DCT1D_databuf_reg_1_4_SRINV_374 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_1_4_SRINV
    );
  U_DCT1D_databuf_reg_1_4_CLKINV_375 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_1_4_CLKINV
    );
  U_DCT1D_databuf_reg_1_4_CEINV_376 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_1_4_CEINV
    );
  U_DCT1D_databuf_reg_1_6_DXMUX_377 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_6_XORF,
      O => U_DCT1D_databuf_reg_1_6_DXMUX
    );
  U_DCT1D_databuf_reg_1_6_XORF_378 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_6_CYINIT,
      I1 => U_DCT1D_nx5403z1,
      O => U_DCT1D_databuf_reg_1_6_XORF
    );
  U_DCT1D_databuf_reg_1_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_6_CY0F,
      IB => U_DCT1D_databuf_reg_1_6_CYINIT,
      SEL => U_DCT1D_databuf_reg_1_6_CYSELF,
      O => U_DCT1D_rtlc5_1420_add_9_ix6400z63342_O
    );
  U_DCT1D_databuf_reg_1_6_CYMUXF2_379 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_6_CY0F,
      IB => U_DCT1D_databuf_reg_1_6_CY0F,
      SEL => U_DCT1D_databuf_reg_1_6_CYSELF,
      O => U_DCT1D_databuf_reg_1_6_CYMUXF2
    );
  U_DCT1D_databuf_reg_1_6_CYINIT_380 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1420_add_9_ix5403z63342_O,
      O => U_DCT1D_databuf_reg_1_6_CYINIT
    );
  U_DCT1D_databuf_reg_1_6_CY0F_381 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(6),
      O => U_DCT1D_databuf_reg_1_6_CY0F
    );
  U_DCT1D_databuf_reg_1_6_CYSELF_382 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx5403z1,
      O => U_DCT1D_databuf_reg_1_6_CYSELF
    );
  U_DCT1D_databuf_reg_1_6_DYMUX_383 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_6_XORG,
      O => U_DCT1D_databuf_reg_1_6_DYMUX
    );
  U_DCT1D_databuf_reg_1_6_XORG_384 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1420_add_9_ix6400z63342_O,
      I1 => U_DCT1D_nx6400z1,
      O => U_DCT1D_databuf_reg_1_6_XORG
    );
  U_DCT1D_databuf_reg_1_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_6_CYMUXFAST,
      O => U_DCT1D_rtlc5_1420_add_9_ix7397z63342_O
    );
  U_DCT1D_databuf_reg_1_6_FASTCARRY_385 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1420_add_9_ix5403z63342_O,
      O => U_DCT1D_databuf_reg_1_6_FASTCARRY
    );
  U_DCT1D_databuf_reg_1_6_CYAND_386 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_1_6_CYSELG,
      I1 => U_DCT1D_databuf_reg_1_6_CYSELF,
      O => U_DCT1D_databuf_reg_1_6_CYAND
    );
  U_DCT1D_databuf_reg_1_6_CYMUXFAST_387 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_6_CYMUXG2,
      IB => U_DCT1D_databuf_reg_1_6_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_1_6_CYAND,
      O => U_DCT1D_databuf_reg_1_6_CYMUXFAST
    );
  U_DCT1D_databuf_reg_1_6_CYMUXG2_388 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_1_6_CY0G,
      IB => U_DCT1D_databuf_reg_1_6_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_1_6_CYSELG,
      O => U_DCT1D_databuf_reg_1_6_CYMUXG2
    );
  U_DCT1D_databuf_reg_1_6_CY0G_389 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(7),
      O => U_DCT1D_databuf_reg_1_6_CY0G
    );
  U_DCT1D_databuf_reg_1_6_CYSELG_390 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx6400z1,
      O => U_DCT1D_databuf_reg_1_6_CYSELG
    );
  U_DCT1D_databuf_reg_1_6_SRINV_391 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_1_6_SRINV
    );
  U_DCT1D_databuf_reg_1_6_CLKINV_392 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_1_6_CLKINV
    );
  U_DCT1D_databuf_reg_1_6_CEINV_393 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_1_6_CEINV
    );
  U_DCT1D_databuf_reg_1_8_DXMUX_394 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_8_XORF,
      O => U_DCT1D_databuf_reg_1_8_DXMUX
    );
  U_DCT1D_databuf_reg_1_8_XORF_395 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_8_CYINIT,
      I1 => U_DCT1D_nx7397z1_rt,
      O => U_DCT1D_databuf_reg_1_8_XORF
    );
  U_DCT1D_databuf_reg_1_8_CYINIT_396 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1420_add_9_ix7397z63342_O,
      O => U_DCT1D_databuf_reg_1_8_CYINIT
    );
  U_DCT1D_databuf_reg_1_8_CLKINV_397 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_1_8_CLKINV
    );
  U_DCT1D_databuf_reg_1_8_CEINV_398 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_1_8_CEINV
    );
  U_DCT2D_ix65206z2345 : X_LUT4
    generic map(
      INIT => X"9595"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1484(11),
      ADR1 => romo2datao10_s(1),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z648
    );
  U_DCT2D_rtlc5n1501_10_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_10_XORF,
      O => U_DCT2D_rtlc5n1501(10)
    );
  U_DCT2D_rtlc5n1501_10_XORF_399 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1501_10_CYINIT,
      I1 => U_DCT2D_nx65206z651,
      O => U_DCT2D_rtlc5n1501_10_XORF
    );
  U_DCT2D_rtlc5n1501_10_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_10_CY0F,
      IB => U_DCT2D_rtlc5n1501_10_CYINIT,
      SEL => U_DCT2D_rtlc5n1501_10_CYSELF,
      O => U_DCT2D_ix65206z64239_O
    );
  U_DCT2D_rtlc5n1501_10_CYINIT_400 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GLOBAL_LOGIC1_39,
      O => U_DCT2D_rtlc5n1501_10_CYINIT
    );
  U_DCT2D_rtlc5n1501_10_CY0F_401 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(10),
      O => U_DCT2D_rtlc5n1501_10_CY0F
    );
  U_DCT2D_rtlc5n1501_10_CYSELF_402 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z651,
      O => U_DCT2D_rtlc5n1501_10_CYSELF
    );
  U_DCT2D_rtlc5n1501_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_10_XORG,
      O => U_DCT2D_rtlc5n1501(11)
    );
  U_DCT2D_rtlc5n1501_10_XORG_403 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64239_O,
      I1 => U_DCT2D_nx65206z648,
      O => U_DCT2D_rtlc5n1501_10_XORG
    );
  U_DCT2D_rtlc5n1501_10_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_10_CYMUXG,
      O => U_DCT2D_ix65206z64235_O
    );
  U_DCT2D_rtlc5n1501_10_CYMUXG_404 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_10_CY0G,
      IB => U_DCT2D_ix65206z64239_O,
      SEL => U_DCT2D_rtlc5n1501_10_CYSELG,
      O => U_DCT2D_rtlc5n1501_10_CYMUXG
    );
  U_DCT2D_rtlc5n1501_10_CY0G_405 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(11),
      O => U_DCT2D_rtlc5n1501_10_CY0G
    );
  U_DCT2D_rtlc5n1501_10_CYSELG_406 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z648,
      O => U_DCT2D_rtlc5n1501_10_CYSELG
    );
  U_DCT2D_ix65206z45555 : X_LUT4
    generic map(
      INIT => X"A959"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1484(13),
      ADR1 => rome2datao10_s(3),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao10_s(3),
      O => U_DCT2D_nx65206z642
    );
  U_DCT2D_rtlc5n1501_12_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_12_XORF,
      O => U_DCT2D_rtlc5n1501(12)
    );
  U_DCT2D_rtlc5n1501_12_XORF_407 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1501_12_CYINIT,
      I1 => U_DCT2D_nx65206z645,
      O => U_DCT2D_rtlc5n1501_12_XORF
    );
  U_DCT2D_rtlc5n1501_12_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_12_CY0F,
      IB => U_DCT2D_rtlc5n1501_12_CYINIT,
      SEL => U_DCT2D_rtlc5n1501_12_CYSELF,
      O => U_DCT2D_ix65206z64231_O
    );
  U_DCT2D_rtlc5n1501_12_CYMUXF2_408 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_12_CY0F,
      IB => U_DCT2D_rtlc5n1501_12_CY0F,
      SEL => U_DCT2D_rtlc5n1501_12_CYSELF,
      O => U_DCT2D_rtlc5n1501_12_CYMUXF2
    );
  U_DCT2D_rtlc5n1501_12_CYINIT_409 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64235_O,
      O => U_DCT2D_rtlc5n1501_12_CYINIT
    );
  U_DCT2D_rtlc5n1501_12_CY0F_410 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(12),
      O => U_DCT2D_rtlc5n1501_12_CY0F
    );
  U_DCT2D_rtlc5n1501_12_CYSELF_411 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z645,
      O => U_DCT2D_rtlc5n1501_12_CYSELF
    );
  U_DCT2D_rtlc5n1501_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_12_XORG,
      O => U_DCT2D_rtlc5n1501(13)
    );
  U_DCT2D_rtlc5n1501_12_XORG_412 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64231_O,
      I1 => U_DCT2D_nx65206z642,
      O => U_DCT2D_rtlc5n1501_12_XORG
    );
  U_DCT2D_rtlc5n1501_12_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_12_CYMUXFAST,
      O => U_DCT2D_ix65206z64227_O
    );
  U_DCT2D_rtlc5n1501_12_FASTCARRY_413 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64235_O,
      O => U_DCT2D_rtlc5n1501_12_FASTCARRY
    );
  U_DCT2D_rtlc5n1501_12_CYAND_414 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1501_12_CYSELG,
      I1 => U_DCT2D_rtlc5n1501_12_CYSELF,
      O => U_DCT2D_rtlc5n1501_12_CYAND
    );
  U_DCT2D_rtlc5n1501_12_CYMUXFAST_415 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_12_CYMUXG2,
      IB => U_DCT2D_rtlc5n1501_12_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1501_12_CYAND,
      O => U_DCT2D_rtlc5n1501_12_CYMUXFAST
    );
  U_DCT2D_rtlc5n1501_12_CYMUXG2_416 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_12_CY0G,
      IB => U_DCT2D_rtlc5n1501_12_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1501_12_CYSELG,
      O => U_DCT2D_rtlc5n1501_12_CYMUXG2
    );
  U_DCT2D_rtlc5n1501_12_CY0G_417 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(13),
      O => U_DCT2D_rtlc5n1501_12_CY0G
    );
  U_DCT2D_rtlc5n1501_12_CYSELG_418 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z642,
      O => U_DCT2D_rtlc5n1501_12_CYSELG
    );
  U_DCT2D_ix65206z45547 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => rome2datao10_s(5),
      ADR1 => U_DCT2D_rtlc5n1484(15),
      ADR2 => romo2datao10_s(5),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z636
    );
  U_DCT2D_rtlc5n1501_14_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_14_XORF,
      O => U_DCT2D_rtlc5n1501(14)
    );
  U_DCT2D_rtlc5n1501_14_XORF_419 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1501_14_CYINIT,
      I1 => U_DCT2D_nx65206z639,
      O => U_DCT2D_rtlc5n1501_14_XORF
    );
  U_DCT2D_rtlc5n1501_14_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_14_CY0F,
      IB => U_DCT2D_rtlc5n1501_14_CYINIT,
      SEL => U_DCT2D_rtlc5n1501_14_CYSELF,
      O => U_DCT2D_ix65206z64223_O
    );
  U_DCT2D_rtlc5n1501_14_CYMUXF2_420 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_14_CY0F,
      IB => U_DCT2D_rtlc5n1501_14_CY0F,
      SEL => U_DCT2D_rtlc5n1501_14_CYSELF,
      O => U_DCT2D_rtlc5n1501_14_CYMUXF2
    );
  U_DCT2D_rtlc5n1501_14_CYINIT_421 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64227_O,
      O => U_DCT2D_rtlc5n1501_14_CYINIT
    );
  U_DCT2D_rtlc5n1501_14_CY0F_422 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(14),
      O => U_DCT2D_rtlc5n1501_14_CY0F
    );
  U_DCT2D_rtlc5n1501_14_CYSELF_423 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z639,
      O => U_DCT2D_rtlc5n1501_14_CYSELF
    );
  U_DCT2D_rtlc5n1501_14_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_14_XORG,
      O => U_DCT2D_rtlc5n1501(15)
    );
  U_DCT2D_rtlc5n1501_14_XORG_424 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64223_O,
      I1 => U_DCT2D_nx65206z636,
      O => U_DCT2D_rtlc5n1501_14_XORG
    );
  U_DCT2D_rtlc5n1501_14_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_14_CYMUXFAST,
      O => U_DCT2D_ix65206z64219_O
    );
  U_DCT2D_rtlc5n1501_14_FASTCARRY_425 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64227_O,
      O => U_DCT2D_rtlc5n1501_14_FASTCARRY
    );
  U_DCT2D_rtlc5n1501_14_CYAND_426 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1501_14_CYSELG,
      I1 => U_DCT2D_rtlc5n1501_14_CYSELF,
      O => U_DCT2D_rtlc5n1501_14_CYAND
    );
  U_DCT2D_rtlc5n1501_14_CYMUXFAST_427 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_14_CYMUXG2,
      IB => U_DCT2D_rtlc5n1501_14_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1501_14_CYAND,
      O => U_DCT2D_rtlc5n1501_14_CYMUXFAST
    );
  U_DCT2D_rtlc5n1501_14_CYMUXG2_428 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_14_CY0G,
      IB => U_DCT2D_rtlc5n1501_14_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1501_14_CYSELG,
      O => U_DCT2D_rtlc5n1501_14_CYMUXG2
    );
  U_DCT2D_rtlc5n1501_14_CY0G_429 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(15),
      O => U_DCT2D_rtlc5n1501_14_CY0G
    );
  U_DCT2D_rtlc5n1501_14_CYSELG_430 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z636,
      O => U_DCT2D_rtlc5n1501_14_CYSELG
    );
  U_DCT2D_ix65206z45539 : X_LUT4
    generic map(
      INIT => X"A959"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1484(17),
      ADR1 => rome2datao10_s(7),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao10_s(7),
      O => U_DCT2D_nx65206z630
    );
  U_DCT2D_rtlc5n1501_16_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_16_XORF,
      O => U_DCT2D_rtlc5n1501(16)
    );
  U_DCT2D_rtlc5n1501_16_XORF_431 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1501_16_CYINIT,
      I1 => U_DCT2D_nx65206z633,
      O => U_DCT2D_rtlc5n1501_16_XORF
    );
  U_DCT2D_rtlc5n1501_16_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_16_CY0F,
      IB => U_DCT2D_rtlc5n1501_16_CYINIT,
      SEL => U_DCT2D_rtlc5n1501_16_CYSELF,
      O => U_DCT2D_ix65206z64215_O
    );
  U_DCT2D_rtlc5n1501_16_CYMUXF2_432 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_16_CY0F,
      IB => U_DCT2D_rtlc5n1501_16_CY0F,
      SEL => U_DCT2D_rtlc5n1501_16_CYSELF,
      O => U_DCT2D_rtlc5n1501_16_CYMUXF2
    );
  U_DCT2D_rtlc5n1501_16_CYINIT_433 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64219_O,
      O => U_DCT2D_rtlc5n1501_16_CYINIT
    );
  U_DCT2D_rtlc5n1501_16_CY0F_434 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(16),
      O => U_DCT2D_rtlc5n1501_16_CY0F
    );
  U_DCT2D_rtlc5n1501_16_CYSELF_435 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z633,
      O => U_DCT2D_rtlc5n1501_16_CYSELF
    );
  U_DCT2D_rtlc5n1501_16_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_16_XORG,
      O => U_DCT2D_rtlc5n1501(17)
    );
  U_DCT2D_rtlc5n1501_16_XORG_436 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64215_O,
      I1 => U_DCT2D_nx65206z630,
      O => U_DCT2D_rtlc5n1501_16_XORG
    );
  U_DCT2D_rtlc5n1501_16_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_16_CYMUXFAST,
      O => U_DCT2D_ix65206z64211_O
    );
  U_DCT2D_rtlc5n1501_16_FASTCARRY_437 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64219_O,
      O => U_DCT2D_rtlc5n1501_16_FASTCARRY
    );
  U_DCT2D_rtlc5n1501_16_CYAND_438 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1501_16_CYSELG,
      I1 => U_DCT2D_rtlc5n1501_16_CYSELF,
      O => U_DCT2D_rtlc5n1501_16_CYAND
    );
  U_DCT2D_rtlc5n1501_16_CYMUXFAST_439 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_16_CYMUXG2,
      IB => U_DCT2D_rtlc5n1501_16_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1501_16_CYAND,
      O => U_DCT2D_rtlc5n1501_16_CYMUXFAST
    );
  U_DCT2D_rtlc5n1501_16_CYMUXG2_440 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_16_CY0G,
      IB => U_DCT2D_rtlc5n1501_16_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1501_16_CYSELG,
      O => U_DCT2D_rtlc5n1501_16_CYMUXG2
    );
  U_DCT2D_rtlc5n1501_16_CY0G_441 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(17),
      O => U_DCT2D_rtlc5n1501_16_CY0G
    );
  U_DCT2D_rtlc5n1501_16_CYSELG_442 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z630,
      O => U_DCT2D_rtlc5n1501_16_CYSELG
    );
  U_DCT2D_ix65206z45531 : X_LUT4
    generic map(
      INIT => X"A959"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1484(19),
      ADR1 => rome2datao10_s(9),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao10_s(9),
      O => U_DCT2D_nx65206z624
    );
  U_DCT2D_rtlc5n1501_18_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_18_XORF,
      O => U_DCT2D_rtlc5n1501(18)
    );
  U_DCT2D_rtlc5n1501_18_XORF_443 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1501_18_CYINIT,
      I1 => U_DCT2D_nx65206z627,
      O => U_DCT2D_rtlc5n1501_18_XORF
    );
  U_DCT2D_rtlc5n1501_18_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_18_CY0F,
      IB => U_DCT2D_rtlc5n1501_18_CYINIT,
      SEL => U_DCT2D_rtlc5n1501_18_CYSELF,
      O => U_DCT2D_ix65206z64207_O
    );
  U_DCT2D_rtlc5n1501_18_CYMUXF2_444 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_18_CY0F,
      IB => U_DCT2D_rtlc5n1501_18_CY0F,
      SEL => U_DCT2D_rtlc5n1501_18_CYSELF,
      O => U_DCT2D_rtlc5n1501_18_CYMUXF2
    );
  U_DCT2D_rtlc5n1501_18_CYINIT_445 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64211_O,
      O => U_DCT2D_rtlc5n1501_18_CYINIT
    );
  U_DCT2D_rtlc5n1501_18_CY0F_446 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(18),
      O => U_DCT2D_rtlc5n1501_18_CY0F
    );
  U_DCT2D_rtlc5n1501_18_CYSELF_447 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z627,
      O => U_DCT2D_rtlc5n1501_18_CYSELF
    );
  U_DCT2D_rtlc5n1501_18_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_18_XORG,
      O => U_DCT2D_rtlc5n1501(19)
    );
  U_DCT2D_rtlc5n1501_18_XORG_448 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64207_O,
      I1 => U_DCT2D_nx65206z624,
      O => U_DCT2D_rtlc5n1501_18_XORG
    );
  U_DCT2D_rtlc5n1501_18_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_18_CYMUXFAST,
      O => U_DCT2D_ix65206z64203_O
    );
  U_DCT2D_rtlc5n1501_18_FASTCARRY_449 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64211_O,
      O => U_DCT2D_rtlc5n1501_18_FASTCARRY
    );
  U_DCT2D_rtlc5n1501_18_CYAND_450 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1501_18_CYSELG,
      I1 => U_DCT2D_rtlc5n1501_18_CYSELF,
      O => U_DCT2D_rtlc5n1501_18_CYAND
    );
  U_DCT2D_rtlc5n1501_18_CYMUXFAST_451 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_18_CYMUXG2,
      IB => U_DCT2D_rtlc5n1501_18_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1501_18_CYAND,
      O => U_DCT2D_rtlc5n1501_18_CYMUXFAST
    );
  U_DCT2D_rtlc5n1501_18_CYMUXG2_452 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_18_CY0G,
      IB => U_DCT2D_rtlc5n1501_18_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1501_18_CYSELG,
      O => U_DCT2D_rtlc5n1501_18_CYMUXG2
    );
  U_DCT2D_rtlc5n1501_18_CY0G_453 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(19),
      O => U_DCT2D_rtlc5n1501_18_CY0G
    );
  U_DCT2D_rtlc5n1501_18_CYSELG_454 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z624,
      O => U_DCT2D_rtlc5n1501_18_CYSELG
    );
  U_DCT2D_ix65206z45523 : X_LUT4
    generic map(
      INIT => X"A959"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1484(21),
      ADR1 => rome2datao10_s(11),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao10_s(11),
      O => U_DCT2D_nx65206z618
    );
  U_DCT2D_rtlc5n1501_20_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_20_XORF,
      O => U_DCT2D_rtlc5n1501(20)
    );
  U_DCT2D_rtlc5n1501_20_XORF_455 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1501_20_CYINIT,
      I1 => U_DCT2D_nx65206z621,
      O => U_DCT2D_rtlc5n1501_20_XORF
    );
  U_DCT2D_rtlc5n1501_20_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_20_CY0F,
      IB => U_DCT2D_rtlc5n1501_20_CYINIT,
      SEL => U_DCT2D_rtlc5n1501_20_CYSELF,
      O => U_DCT2D_ix65206z64199_O
    );
  U_DCT2D_rtlc5n1501_20_CYMUXF2_456 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_20_CY0F,
      IB => U_DCT2D_rtlc5n1501_20_CY0F,
      SEL => U_DCT2D_rtlc5n1501_20_CYSELF,
      O => U_DCT2D_rtlc5n1501_20_CYMUXF2
    );
  U_DCT2D_rtlc5n1501_20_CYINIT_457 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64203_O,
      O => U_DCT2D_rtlc5n1501_20_CYINIT
    );
  U_DCT2D_rtlc5n1501_20_CY0F_458 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(20),
      O => U_DCT2D_rtlc5n1501_20_CY0F
    );
  U_DCT2D_rtlc5n1501_20_CYSELF_459 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z621,
      O => U_DCT2D_rtlc5n1501_20_CYSELF
    );
  U_DCT2D_rtlc5n1501_20_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_20_XORG,
      O => U_DCT2D_rtlc5n1501(21)
    );
  U_DCT2D_rtlc5n1501_20_XORG_460 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64199_O,
      I1 => U_DCT2D_nx65206z618,
      O => U_DCT2D_rtlc5n1501_20_XORG
    );
  U_DCT2D_rtlc5n1501_20_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_20_CYMUXFAST,
      O => U_DCT2D_ix65206z64195_O
    );
  U_DCT2D_rtlc5n1501_20_FASTCARRY_461 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64203_O,
      O => U_DCT2D_rtlc5n1501_20_FASTCARRY
    );
  U_DCT2D_rtlc5n1501_20_CYAND_462 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1501_20_CYSELG,
      I1 => U_DCT2D_rtlc5n1501_20_CYSELF,
      O => U_DCT2D_rtlc5n1501_20_CYAND
    );
  U_DCT2D_rtlc5n1501_20_CYMUXFAST_463 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_20_CYMUXG2,
      IB => U_DCT2D_rtlc5n1501_20_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1501_20_CYAND,
      O => U_DCT2D_rtlc5n1501_20_CYMUXFAST
    );
  U_DCT2D_rtlc5n1501_20_CYMUXG2_464 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_20_CY0G,
      IB => U_DCT2D_rtlc5n1501_20_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1501_20_CYSELG,
      O => U_DCT2D_rtlc5n1501_20_CYMUXG2
    );
  U_DCT2D_rtlc5n1501_20_CY0G_465 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(21),
      O => U_DCT2D_rtlc5n1501_20_CY0G
    );
  U_DCT2D_rtlc5n1501_20_CYSELG_466 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z618,
      O => U_DCT2D_rtlc5n1501_20_CYSELG
    );
  U_DCT2D_nx65206z571_rt_467 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_nx65206z571,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z571_rt
    );
  U_DCT2D_rtlc5n1501_22_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_22_XORF,
      O => U_DCT2D_rtlc5n1501(22)
    );
  U_DCT2D_rtlc5n1501_22_XORF_468 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1501_22_CYINIT,
      I1 => U_DCT2D_nx65206z615,
      O => U_DCT2D_rtlc5n1501_22_XORF
    );
  U_DCT2D_rtlc5n1501_22_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1501_22_CY0F,
      IB => U_DCT2D_rtlc5n1501_22_CYINIT,
      SEL => U_DCT2D_rtlc5n1501_22_CYSELF,
      O => U_DCT2D_ix65206z64191_O
    );
  U_DCT2D_rtlc5n1501_22_CYINIT_469 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64195_O,
      O => U_DCT2D_rtlc5n1501_22_CYINIT
    );
  U_DCT2D_rtlc5n1501_22_CY0F_470 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484(22),
      O => U_DCT2D_rtlc5n1501_22_CY0F
    );
  U_DCT2D_rtlc5n1501_22_CYSELF_471 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z615,
      O => U_DCT2D_rtlc5n1501_22_CYSELF
    );
  U_DCT2D_rtlc5n1501_22_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1501_22_XORG,
      O => U_DCT2D_rtlc5n1501(23)
    );
  U_DCT2D_rtlc5n1501_22_XORG_472 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64191_O,
      I1 => U_DCT2D_nx65206z571_rt,
      O => U_DCT2D_rtlc5n1501_22_XORG
    );
  U_DCT2D_ix65206z32040 : X_LUT4
    generic map(
      INIT => X"74B8"
    )
    port map (
      ADR0 => romo2datao9_s(1),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => rome2datao8_s(2),
      ADR3 => romo2datao8_s(2),
      O => U_DCT2D_nx65206z609
    );
  U_DCT2D_ix65206z2235 : X_LUT4
    generic map(
      INIT => X"4848"
    )
    port map (
      ADR0 => romo2datao8_s(1),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => romo2datao9_s(0),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z612
    );
  U_DCT2D_rtlc5n1484_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_9_XORF,
      O => U_DCT2D_rtlc5n1484(9)
    );
  U_DCT2D_rtlc5n1484_9_XORF_473 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1484_9_CYINIT,
      I1 => U_DCT2D_nx65206z612,
      O => U_DCT2D_rtlc5n1484_9_XORF
    );
  U_DCT2D_rtlc5n1484_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_9_CY0F,
      IB => U_DCT2D_rtlc5n1484_9_CYINIT,
      SEL => U_DCT2D_rtlc5n1484_9_CYSELF,
      O => U_DCT2D_ix65206z64188_O
    );
  U_DCT2D_rtlc5n1484_9_CYINIT_474 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_9_BXINVNOT,
      O => U_DCT2D_rtlc5n1484_9_CYINIT
    );
  U_DCT2D_rtlc5n1484_9_CY0F_475 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z613,
      O => U_DCT2D_rtlc5n1484_9_CY0F
    );
  U_DCT2D_rtlc5n1484_9_FAND : X_AND2
    port map (
      I0 => U_DCT2D_state_reg(0),
      I1 => romo2datao8_s(1),
      O => U_DCT2D_nx65206z613
    );
  U_DCT2D_rtlc5n1484_9_CYSELF_476 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z612,
      O => U_DCT2D_rtlc5n1484_9_CYSELF
    );
  U_DCT2D_rtlc5n1484_9_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_33,
      O => U_DCT2D_rtlc5n1484_9_BXINVNOT
    );
  U_DCT2D_rtlc5n1484_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_9_XORG,
      O => U_DCT2D_rtlc5n1484(10)
    );
  U_DCT2D_rtlc5n1484_9_XORG_477 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64188_O,
      I1 => U_DCT2D_nx65206z609,
      O => U_DCT2D_rtlc5n1484_9_XORG
    );
  U_DCT2D_rtlc5n1484_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_9_CYMUXG,
      O => U_DCT2D_ix65206z64185_O
    );
  U_DCT2D_rtlc5n1484_9_CYMUXG_478 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_9_CY0G,
      IB => U_DCT2D_ix65206z64188_O,
      SEL => U_DCT2D_rtlc5n1484_9_CYSELG,
      O => U_DCT2D_rtlc5n1484_9_CYMUXG
    );
  U_DCT2D_rtlc5n1484_9_CY0G_479 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z610,
      O => U_DCT2D_rtlc5n1484_9_CY0G
    );
  U_DCT2D_rtlc5n1484_9_GAND : X_AND2
    port map (
      I0 => U_DCT2D_state_reg(0),
      I1 => romo2datao9_s(1),
      O => U_DCT2D_nx65206z610
    );
  U_DCT2D_rtlc5n1484_9_CYSELG_480 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z609,
      O => U_DCT2D_rtlc5n1484_9_CYSELG
    );
  U_DCT2D_ix65206z24336 : X_LUT4
    generic map(
      INIT => X"36C6"
    )
    port map (
      ADR0 => rome2datao9_s(3),
      ADR1 => U_DCT2D_nx65206z604,
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao9_s(3),
      O => U_DCT2D_nx65206z603
    );
  U_DCT2D_ix65206z24339 : X_LUT4
    generic map(
      INIT => X"56A6"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z607,
      ADR1 => rome2datao9_s(2),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao9_s(2),
      O => U_DCT2D_nx65206z606
    );
  U_DCT2D_rtlc5n1484_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_11_XORF,
      O => U_DCT2D_rtlc5n1484(11)
    );
  U_DCT2D_rtlc5n1484_11_XORF_481 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1484_11_CYINIT,
      I1 => U_DCT2D_nx65206z606,
      O => U_DCT2D_rtlc5n1484_11_XORF
    );
  U_DCT2D_rtlc5n1484_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_11_CY0F,
      IB => U_DCT2D_rtlc5n1484_11_CYINIT,
      SEL => U_DCT2D_rtlc5n1484_11_CYSELF,
      O => U_DCT2D_ix65206z64182_O
    );
  U_DCT2D_rtlc5n1484_11_CYMUXF2_482 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_11_CY0F,
      IB => U_DCT2D_rtlc5n1484_11_CY0F,
      SEL => U_DCT2D_rtlc5n1484_11_CYSELF,
      O => U_DCT2D_rtlc5n1484_11_CYMUXF2
    );
  U_DCT2D_rtlc5n1484_11_CYINIT_483 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64185_O,
      O => U_DCT2D_rtlc5n1484_11_CYINIT
    );
  U_DCT2D_rtlc5n1484_11_CY0F_484 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z607,
      O => U_DCT2D_rtlc5n1484_11_CY0F
    );
  U_DCT2D_rtlc5n1484_11_CYSELF_485 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z606,
      O => U_DCT2D_rtlc5n1484_11_CYSELF
    );
  U_DCT2D_rtlc5n1484_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_11_XORG,
      O => U_DCT2D_rtlc5n1484(12)
    );
  U_DCT2D_rtlc5n1484_11_XORG_486 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64182_O,
      I1 => U_DCT2D_nx65206z603,
      O => U_DCT2D_rtlc5n1484_11_XORG
    );
  U_DCT2D_rtlc5n1484_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_11_CYMUXFAST,
      O => U_DCT2D_ix65206z64179_O
    );
  U_DCT2D_rtlc5n1484_11_FASTCARRY_487 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64185_O,
      O => U_DCT2D_rtlc5n1484_11_FASTCARRY
    );
  U_DCT2D_rtlc5n1484_11_CYAND_488 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1484_11_CYSELG,
      I1 => U_DCT2D_rtlc5n1484_11_CYSELF,
      O => U_DCT2D_rtlc5n1484_11_CYAND
    );
  U_DCT2D_rtlc5n1484_11_CYMUXFAST_489 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_11_CYMUXG2,
      IB => U_DCT2D_rtlc5n1484_11_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1484_11_CYAND,
      O => U_DCT2D_rtlc5n1484_11_CYMUXFAST
    );
  U_DCT2D_rtlc5n1484_11_CYMUXG2_490 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_11_CY0G,
      IB => U_DCT2D_rtlc5n1484_11_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1484_11_CYSELG,
      O => U_DCT2D_rtlc5n1484_11_CYMUXG2
    );
  U_DCT2D_rtlc5n1484_11_CY0G_491 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z604,
      O => U_DCT2D_rtlc5n1484_11_CY0G
    );
  U_DCT2D_rtlc5n1484_11_CYSELG_492 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z603,
      O => U_DCT2D_rtlc5n1484_11_CYSELG
    );
  U_DCT1D_reg_databuf_reg_2_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_2_0_DXMUX,
      CE => U_DCT1D_databuf_reg_2_0_CEINV,
      CLK => U_DCT1D_databuf_reg_2_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_2_0_FFX_RST,
      O => U_DCT1D_databuf_reg_2_Q(0)
    );
  U_DCT1D_databuf_reg_2_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_2_0_FFX_RST
    );
  U_DCT2D_ix65206z24330 : X_LUT4
    generic map(
      INIT => X"5A66"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z598,
      ADR1 => rome2datao9_s(5),
      ADR2 => romo2datao9_s(5),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z597
    );
  U_DCT2D_rtlc5n1484_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_13_XORF,
      O => U_DCT2D_rtlc5n1484(13)
    );
  U_DCT2D_rtlc5n1484_13_XORF_493 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1484_13_CYINIT,
      I1 => U_DCT2D_nx65206z600,
      O => U_DCT2D_rtlc5n1484_13_XORF
    );
  U_DCT2D_rtlc5n1484_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_13_CY0F,
      IB => U_DCT2D_rtlc5n1484_13_CYINIT,
      SEL => U_DCT2D_rtlc5n1484_13_CYSELF,
      O => U_DCT2D_ix65206z64176_O
    );
  U_DCT2D_rtlc5n1484_13_CYMUXF2_494 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_13_CY0F,
      IB => U_DCT2D_rtlc5n1484_13_CY0F,
      SEL => U_DCT2D_rtlc5n1484_13_CYSELF,
      O => U_DCT2D_rtlc5n1484_13_CYMUXF2
    );
  U_DCT2D_rtlc5n1484_13_CYINIT_495 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64179_O,
      O => U_DCT2D_rtlc5n1484_13_CYINIT
    );
  U_DCT2D_rtlc5n1484_13_CY0F_496 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z601,
      O => U_DCT2D_rtlc5n1484_13_CY0F
    );
  U_DCT2D_rtlc5n1484_13_CYSELF_497 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z600,
      O => U_DCT2D_rtlc5n1484_13_CYSELF
    );
  U_DCT2D_rtlc5n1484_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_13_XORG,
      O => U_DCT2D_rtlc5n1484(14)
    );
  U_DCT2D_rtlc5n1484_13_XORG_498 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64176_O,
      I1 => U_DCT2D_nx65206z597,
      O => U_DCT2D_rtlc5n1484_13_XORG
    );
  U_DCT2D_rtlc5n1484_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_13_CYMUXFAST,
      O => U_DCT2D_ix65206z64173_O
    );
  U_DCT2D_rtlc5n1484_13_FASTCARRY_499 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64179_O,
      O => U_DCT2D_rtlc5n1484_13_FASTCARRY
    );
  U_DCT2D_rtlc5n1484_13_CYAND_500 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1484_13_CYSELG,
      I1 => U_DCT2D_rtlc5n1484_13_CYSELF,
      O => U_DCT2D_rtlc5n1484_13_CYAND
    );
  U_DCT2D_rtlc5n1484_13_CYMUXFAST_501 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_13_CYMUXG2,
      IB => U_DCT2D_rtlc5n1484_13_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1484_13_CYAND,
      O => U_DCT2D_rtlc5n1484_13_CYMUXFAST
    );
  U_DCT2D_rtlc5n1484_13_CYMUXG2_502 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_13_CY0G,
      IB => U_DCT2D_rtlc5n1484_13_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1484_13_CYSELG,
      O => U_DCT2D_rtlc5n1484_13_CYMUXG2
    );
  U_DCT2D_rtlc5n1484_13_CY0G_503 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z598,
      O => U_DCT2D_rtlc5n1484_13_CY0G
    );
  U_DCT2D_rtlc5n1484_13_CYSELG_504 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z597,
      O => U_DCT2D_rtlc5n1484_13_CYSELG
    );
  U_DCT2D_ix65206z24324 : X_LUT4
    generic map(
      INIT => X"5A66"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z592,
      ADR1 => rome2datao9_s(7),
      ADR2 => romo2datao9_s(7),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z591
    );
  U_DCT2D_rtlc5n1484_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_15_XORF,
      O => U_DCT2D_rtlc5n1484(15)
    );
  U_DCT2D_rtlc5n1484_15_XORF_505 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1484_15_CYINIT,
      I1 => U_DCT2D_nx65206z594,
      O => U_DCT2D_rtlc5n1484_15_XORF
    );
  U_DCT2D_rtlc5n1484_15_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_15_CY0F,
      IB => U_DCT2D_rtlc5n1484_15_CYINIT,
      SEL => U_DCT2D_rtlc5n1484_15_CYSELF,
      O => U_DCT2D_ix65206z64170_O
    );
  U_DCT2D_rtlc5n1484_15_CYMUXF2_506 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_15_CY0F,
      IB => U_DCT2D_rtlc5n1484_15_CY0F,
      SEL => U_DCT2D_rtlc5n1484_15_CYSELF,
      O => U_DCT2D_rtlc5n1484_15_CYMUXF2
    );
  U_DCT2D_rtlc5n1484_15_CYINIT_507 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64173_O,
      O => U_DCT2D_rtlc5n1484_15_CYINIT
    );
  U_DCT2D_rtlc5n1484_15_CY0F_508 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z595,
      O => U_DCT2D_rtlc5n1484_15_CY0F
    );
  U_DCT2D_rtlc5n1484_15_CYSELF_509 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z594,
      O => U_DCT2D_rtlc5n1484_15_CYSELF
    );
  U_DCT2D_rtlc5n1484_15_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_15_XORG,
      O => U_DCT2D_rtlc5n1484(16)
    );
  U_DCT2D_rtlc5n1484_15_XORG_510 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64170_O,
      I1 => U_DCT2D_nx65206z591,
      O => U_DCT2D_rtlc5n1484_15_XORG
    );
  U_DCT2D_rtlc5n1484_15_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_15_CYMUXFAST,
      O => U_DCT2D_ix65206z64167_O
    );
  U_DCT2D_rtlc5n1484_15_FASTCARRY_511 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64173_O,
      O => U_DCT2D_rtlc5n1484_15_FASTCARRY
    );
  U_DCT2D_rtlc5n1484_15_CYAND_512 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1484_15_CYSELG,
      I1 => U_DCT2D_rtlc5n1484_15_CYSELF,
      O => U_DCT2D_rtlc5n1484_15_CYAND
    );
  U_DCT2D_rtlc5n1484_15_CYMUXFAST_513 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_15_CYMUXG2,
      IB => U_DCT2D_rtlc5n1484_15_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1484_15_CYAND,
      O => U_DCT2D_rtlc5n1484_15_CYMUXFAST
    );
  U_DCT2D_rtlc5n1484_15_CYMUXG2_514 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_15_CY0G,
      IB => U_DCT2D_rtlc5n1484_15_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1484_15_CYSELG,
      O => U_DCT2D_rtlc5n1484_15_CYMUXG2
    );
  U_DCT2D_rtlc5n1484_15_CY0G_515 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z592,
      O => U_DCT2D_rtlc5n1484_15_CY0G
    );
  U_DCT2D_rtlc5n1484_15_CYSELG_516 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z591,
      O => U_DCT2D_rtlc5n1484_15_CYSELG
    );
  U_DCT2D_ix65206z24318 : X_LUT4
    generic map(
      INIT => X"5A66"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z586,
      ADR1 => rome2datao9_s(9),
      ADR2 => romo2datao9_s(9),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z585
    );
  U_DCT2D_rtlc5n1484_17_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_17_XORF,
      O => U_DCT2D_rtlc5n1484(17)
    );
  U_DCT2D_rtlc5n1484_17_XORF_517 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1484_17_CYINIT,
      I1 => U_DCT2D_nx65206z588,
      O => U_DCT2D_rtlc5n1484_17_XORF
    );
  U_DCT2D_rtlc5n1484_17_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_17_CY0F,
      IB => U_DCT2D_rtlc5n1484_17_CYINIT,
      SEL => U_DCT2D_rtlc5n1484_17_CYSELF,
      O => U_DCT2D_ix65206z64164_O
    );
  U_DCT2D_rtlc5n1484_17_CYMUXF2_518 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_17_CY0F,
      IB => U_DCT2D_rtlc5n1484_17_CY0F,
      SEL => U_DCT2D_rtlc5n1484_17_CYSELF,
      O => U_DCT2D_rtlc5n1484_17_CYMUXF2
    );
  U_DCT2D_rtlc5n1484_17_CYINIT_519 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64167_O,
      O => U_DCT2D_rtlc5n1484_17_CYINIT
    );
  U_DCT2D_rtlc5n1484_17_CY0F_520 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z589,
      O => U_DCT2D_rtlc5n1484_17_CY0F
    );
  U_DCT2D_rtlc5n1484_17_CYSELF_521 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z588,
      O => U_DCT2D_rtlc5n1484_17_CYSELF
    );
  U_DCT2D_rtlc5n1484_17_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_17_XORG,
      O => U_DCT2D_rtlc5n1484(18)
    );
  U_DCT2D_rtlc5n1484_17_XORG_522 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64164_O,
      I1 => U_DCT2D_nx65206z585,
      O => U_DCT2D_rtlc5n1484_17_XORG
    );
  U_DCT2D_rtlc5n1484_17_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_17_CYMUXFAST,
      O => U_DCT2D_ix65206z64161_O
    );
  U_DCT2D_rtlc5n1484_17_FASTCARRY_523 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64167_O,
      O => U_DCT2D_rtlc5n1484_17_FASTCARRY
    );
  U_DCT2D_rtlc5n1484_17_CYAND_524 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1484_17_CYSELG,
      I1 => U_DCT2D_rtlc5n1484_17_CYSELF,
      O => U_DCT2D_rtlc5n1484_17_CYAND
    );
  U_DCT2D_rtlc5n1484_17_CYMUXFAST_525 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_17_CYMUXG2,
      IB => U_DCT2D_rtlc5n1484_17_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1484_17_CYAND,
      O => U_DCT2D_rtlc5n1484_17_CYMUXFAST
    );
  U_DCT2D_rtlc5n1484_17_CYMUXG2_526 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_17_CY0G,
      IB => U_DCT2D_rtlc5n1484_17_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1484_17_CYSELG,
      O => U_DCT2D_rtlc5n1484_17_CYMUXG2
    );
  U_DCT2D_rtlc5n1484_17_CY0G_527 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z586,
      O => U_DCT2D_rtlc5n1484_17_CY0G
    );
  U_DCT2D_rtlc5n1484_17_CYSELG_528 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z585,
      O => U_DCT2D_rtlc5n1484_17_CYSELG
    );
  U_DCT2D_ix65206z24312 : X_LUT4
    generic map(
      INIT => X"56A6"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z580,
      ADR1 => rome2datao9_s(11),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao9_s(11),
      O => U_DCT2D_nx65206z579
    );
  U_DCT2D_rtlc5n1484_19_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_19_XORF,
      O => U_DCT2D_rtlc5n1484(19)
    );
  U_DCT2D_rtlc5n1484_19_XORF_529 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1484_19_CYINIT,
      I1 => U_DCT2D_nx65206z582,
      O => U_DCT2D_rtlc5n1484_19_XORF
    );
  U_DCT2D_rtlc5n1484_19_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_19_CY0F,
      IB => U_DCT2D_rtlc5n1484_19_CYINIT,
      SEL => U_DCT2D_rtlc5n1484_19_CYSELF,
      O => U_DCT2D_ix65206z64158_O
    );
  U_DCT2D_rtlc5n1484_19_CYMUXF2_530 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_19_CY0F,
      IB => U_DCT2D_rtlc5n1484_19_CY0F,
      SEL => U_DCT2D_rtlc5n1484_19_CYSELF,
      O => U_DCT2D_rtlc5n1484_19_CYMUXF2
    );
  U_DCT2D_rtlc5n1484_19_CYINIT_531 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64161_O,
      O => U_DCT2D_rtlc5n1484_19_CYINIT
    );
  U_DCT2D_rtlc5n1484_19_CY0F_532 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z583,
      O => U_DCT2D_rtlc5n1484_19_CY0F
    );
  U_DCT2D_rtlc5n1484_19_CYSELF_533 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z582,
      O => U_DCT2D_rtlc5n1484_19_CYSELF
    );
  U_DCT2D_rtlc5n1484_19_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_19_XORG,
      O => U_DCT2D_rtlc5n1484(20)
    );
  U_DCT2D_rtlc5n1484_19_XORG_534 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64158_O,
      I1 => U_DCT2D_nx65206z579,
      O => U_DCT2D_rtlc5n1484_19_XORG
    );
  U_DCT2D_rtlc5n1484_19_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_19_CYMUXFAST,
      O => U_DCT2D_ix65206z64155_O
    );
  U_DCT2D_rtlc5n1484_19_FASTCARRY_535 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64161_O,
      O => U_DCT2D_rtlc5n1484_19_FASTCARRY
    );
  U_DCT2D_rtlc5n1484_19_CYAND_536 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1484_19_CYSELG,
      I1 => U_DCT2D_rtlc5n1484_19_CYSELF,
      O => U_DCT2D_rtlc5n1484_19_CYAND
    );
  U_DCT2D_rtlc5n1484_19_CYMUXFAST_537 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_19_CYMUXG2,
      IB => U_DCT2D_rtlc5n1484_19_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1484_19_CYAND,
      O => U_DCT2D_rtlc5n1484_19_CYMUXFAST
    );
  U_DCT2D_rtlc5n1484_19_CYMUXG2_538 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_19_CY0G,
      IB => U_DCT2D_rtlc5n1484_19_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1484_19_CYSELG,
      O => U_DCT2D_rtlc5n1484_19_CYMUXG2
    );
  U_DCT2D_rtlc5n1484_19_CY0G_539 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z580,
      O => U_DCT2D_rtlc5n1484_19_CY0G
    );
  U_DCT2D_rtlc5n1484_19_CYSELG_540 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z579,
      O => U_DCT2D_rtlc5n1484_19_CYSELG
    );
  U_DCT2D_ix65206z24308 : X_LUT4
    generic map(
      INIT => X"5A66"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z573,
      ADR1 => rome2datao9_s(13),
      ADR2 => romo2datao9_s(13),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z575
    );
  U_DCT2D_rtlc5n1484_21_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_21_XORF,
      O => U_DCT2D_rtlc5n1484(21)
    );
  U_DCT2D_rtlc5n1484_21_XORF_541 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1484_21_CYINIT,
      I1 => U_DCT2D_nx65206z577,
      O => U_DCT2D_rtlc5n1484_21_XORF
    );
  U_DCT2D_rtlc5n1484_21_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_21_CY0F,
      IB => U_DCT2D_rtlc5n1484_21_CYINIT,
      SEL => U_DCT2D_rtlc5n1484_21_CYSELF,
      O => U_DCT2D_ix65206z64153_O
    );
  U_DCT2D_rtlc5n1484_21_CYMUXF2_542 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_21_CY0F,
      IB => U_DCT2D_rtlc5n1484_21_CY0F,
      SEL => U_DCT2D_rtlc5n1484_21_CYSELF,
      O => U_DCT2D_rtlc5n1484_21_CYMUXF2
    );
  U_DCT2D_rtlc5n1484_21_CYINIT_543 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64155_O,
      O => U_DCT2D_rtlc5n1484_21_CYINIT
    );
  U_DCT2D_rtlc5n1484_21_CY0F_544 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z573,
      O => U_DCT2D_rtlc5n1484_21_CY0F
    );
  U_DCT2D_rtlc5n1484_21_CYSELF_545 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z577,
      O => U_DCT2D_rtlc5n1484_21_CYSELF
    );
  U_DCT2D_rtlc5n1484_21_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_21_XORG,
      O => U_DCT2D_rtlc5n1484(22)
    );
  U_DCT2D_rtlc5n1484_21_XORG_546 : X_XOR2
    port map (
      I0 => U_DCT2D_ix65206z64153_O,
      I1 => U_DCT2D_nx65206z575,
      O => U_DCT2D_rtlc5n1484_21_XORG
    );
  U_DCT2D_rtlc5n1484_21_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_21_CYMUXFAST,
      O => U_DCT2D_ix65206z64151_O
    );
  U_DCT2D_rtlc5n1484_21_FASTCARRY_547 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64155_O,
      O => U_DCT2D_rtlc5n1484_21_FASTCARRY
    );
  U_DCT2D_rtlc5n1484_21_CYAND_548 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1484_21_CYSELG,
      I1 => U_DCT2D_rtlc5n1484_21_CYSELF,
      O => U_DCT2D_rtlc5n1484_21_CYAND
    );
  U_DCT2D_rtlc5n1484_21_CYMUXFAST_549 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_21_CYMUXG2,
      IB => U_DCT2D_rtlc5n1484_21_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1484_21_CYAND,
      O => U_DCT2D_rtlc5n1484_21_CYMUXFAST
    );
  U_DCT2D_rtlc5n1484_21_CYMUXG2_550 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1484_21_CY0G,
      IB => U_DCT2D_rtlc5n1484_21_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1484_21_CYSELG,
      O => U_DCT2D_rtlc5n1484_21_CYMUXG2
    );
  U_DCT2D_rtlc5n1484_21_CY0G_551 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z573,
      O => U_DCT2D_rtlc5n1484_21_CY0G
    );
  U_DCT2D_rtlc5n1484_21_CYSELG_552 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z575,
      O => U_DCT2D_rtlc5n1484_21_CYSELG
    );
  U_DCT2D_rtlc5n1484_23_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1484_23_XORF,
      O => U_DCT2D_rtlc5n1484(23)
    );
  U_DCT2D_rtlc5n1484_23_XORF_553 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1484_23_CYINIT,
      I1 => U_DCT2D_nx65206z572_rt,
      O => U_DCT2D_rtlc5n1484_23_XORF
    );
  U_DCT2D_rtlc5n1484_23_CYINIT_554 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix65206z64151_O,
      O => U_DCT2D_rtlc5n1484_23_CYINIT
    );
  U_DCT2D_databuf_reg_1_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_1_0_FFX_RST
    );
  U_DCT2D_reg_databuf_reg_1_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_1_0_DXMUX,
      CE => U_DCT2D_databuf_reg_1_0_CEINV,
      CLK => U_DCT2D_databuf_reg_1_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_1_0_FFX_RST,
      O => U_DCT2D_databuf_reg_1_Q(0)
    );
  U_DCT2D_databuf_reg_1_0_DXMUX_555 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_0_XORF,
      O => U_DCT2D_databuf_reg_1_0_DXMUX
    );
  U_DCT2D_databuf_reg_1_0_XORF_556 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_0_CYINIT,
      I1 => U_DCT2D_nx64957z1,
      O => U_DCT2D_databuf_reg_1_0_XORF
    );
  U_DCT2D_databuf_reg_1_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_0_CY0F,
      IB => U_DCT2D_databuf_reg_1_0_CYINIT,
      SEL => U_DCT2D_databuf_reg_1_0_CYSELF,
      O => U_DCT2D_rtlc5_1579_add_46_ix418z63342_O
    );
  U_DCT2D_databuf_reg_1_0_CYINIT_557 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_0_BXINVNOT,
      O => U_DCT2D_databuf_reg_1_0_CYINIT
    );
  U_DCT2D_databuf_reg_1_0_CY0F_558 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_0_Q,
      O => U_DCT2D_databuf_reg_1_0_CY0F
    );
  U_DCT2D_databuf_reg_1_0_CYSELF_559 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx64957z1,
      O => U_DCT2D_databuf_reg_1_0_CYSELF
    );
  U_DCT2D_databuf_reg_1_0_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_25,
      O => U_DCT2D_databuf_reg_1_0_BXINVNOT
    );
  U_DCT2D_databuf_reg_1_0_DYMUX_560 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_0_XORG,
      O => U_DCT2D_databuf_reg_1_0_DYMUX
    );
  U_DCT2D_databuf_reg_1_0_XORG_561 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1579_add_46_ix418z63342_O,
      I1 => U_DCT2D_nx418z1,
      O => U_DCT2D_databuf_reg_1_0_XORG
    );
  U_DCT2D_databuf_reg_1_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_0_CYMUXG,
      O => U_DCT2D_rtlc5_1579_add_46_ix1415z63342_O
    );
  U_DCT2D_databuf_reg_1_0_CYMUXG_562 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_0_CY0G,
      IB => U_DCT2D_rtlc5_1579_add_46_ix418z63342_O,
      SEL => U_DCT2D_databuf_reg_1_0_CYSELG,
      O => U_DCT2D_databuf_reg_1_0_CYMUXG
    );
  U_DCT2D_databuf_reg_1_0_CY0G_563 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_1_Q,
      O => U_DCT2D_databuf_reg_1_0_CY0G
    );
  U_DCT2D_databuf_reg_1_0_CYSELG_564 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx418z1,
      O => U_DCT2D_databuf_reg_1_0_CYSELG
    );
  U_DCT2D_databuf_reg_1_0_SRINV_565 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_1_0_SRINV
    );
  U_DCT2D_databuf_reg_1_0_CLKINV_566 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_1_0_CLKINV
    );
  U_DCT2D_databuf_reg_1_0_CEINV_567 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_1_0_CEINV
    );
  U_DCT2D_databuf_reg_1_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_1_2_FFX_RST
    );
  U_DCT2D_reg_databuf_reg_1_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_1_2_DXMUX,
      CE => U_DCT2D_databuf_reg_1_2_CEINV,
      CLK => U_DCT2D_databuf_reg_1_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_1_2_FFX_RST,
      O => U_DCT2D_databuf_reg_1_Q(2)
    );
  U_DCT2D_ix1415z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_6_2_Q,
      ADR1 => U_DCT2D_latchbuf_reg_1_2_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx1415z1
    );
  U_DCT2D_databuf_reg_1_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_1_2_FFY_RST
    );
  U_DCT2D_reg_databuf_reg_1_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_1_2_DYMUX,
      CE => U_DCT2D_databuf_reg_1_2_CEINV,
      CLK => U_DCT2D_databuf_reg_1_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_1_2_FFY_RST,
      O => U_DCT2D_databuf_reg_1_Q(3)
    );
  U_DCT2D_ix2412z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_1_3_Q,
      ADR1 => U_DCT2D_latchbuf_reg_6_3_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx2412z1
    );
  U_DCT2D_databuf_reg_1_2_DXMUX_568 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_2_XORF,
      O => U_DCT2D_databuf_reg_1_2_DXMUX
    );
  U_DCT2D_databuf_reg_1_2_XORF_569 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_2_CYINIT,
      I1 => U_DCT2D_nx1415z1,
      O => U_DCT2D_databuf_reg_1_2_XORF
    );
  U_DCT2D_databuf_reg_1_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_2_CY0F,
      IB => U_DCT2D_databuf_reg_1_2_CYINIT,
      SEL => U_DCT2D_databuf_reg_1_2_CYSELF,
      O => U_DCT2D_rtlc5_1579_add_46_ix2412z63342_O
    );
  U_DCT2D_databuf_reg_1_2_CYMUXF2_570 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_2_CY0F,
      IB => U_DCT2D_databuf_reg_1_2_CY0F,
      SEL => U_DCT2D_databuf_reg_1_2_CYSELF,
      O => U_DCT2D_databuf_reg_1_2_CYMUXF2
    );
  U_DCT2D_databuf_reg_1_2_CYINIT_571 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1579_add_46_ix1415z63342_O,
      O => U_DCT2D_databuf_reg_1_2_CYINIT
    );
  U_DCT2D_databuf_reg_1_2_CY0F_572 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_2_Q,
      O => U_DCT2D_databuf_reg_1_2_CY0F
    );
  U_DCT2D_databuf_reg_1_2_CYSELF_573 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx1415z1,
      O => U_DCT2D_databuf_reg_1_2_CYSELF
    );
  U_DCT2D_databuf_reg_1_2_DYMUX_574 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_2_XORG,
      O => U_DCT2D_databuf_reg_1_2_DYMUX
    );
  U_DCT2D_databuf_reg_1_2_XORG_575 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1579_add_46_ix2412z63342_O,
      I1 => U_DCT2D_nx2412z1,
      O => U_DCT2D_databuf_reg_1_2_XORG
    );
  U_DCT2D_databuf_reg_1_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_2_CYMUXFAST,
      O => U_DCT2D_rtlc5_1579_add_46_ix3409z63342_O
    );
  U_DCT2D_databuf_reg_1_2_FASTCARRY_576 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1579_add_46_ix1415z63342_O,
      O => U_DCT2D_databuf_reg_1_2_FASTCARRY
    );
  U_DCT2D_databuf_reg_1_2_CYAND_577 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_1_2_CYSELG,
      I1 => U_DCT2D_databuf_reg_1_2_CYSELF,
      O => U_DCT2D_databuf_reg_1_2_CYAND
    );
  U_DCT2D_databuf_reg_1_2_CYMUXFAST_578 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_2_CYMUXG2,
      IB => U_DCT2D_databuf_reg_1_2_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_1_2_CYAND,
      O => U_DCT2D_databuf_reg_1_2_CYMUXFAST
    );
  U_DCT2D_databuf_reg_1_2_CYMUXG2_579 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_2_CY0G,
      IB => U_DCT2D_databuf_reg_1_2_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_1_2_CYSELG,
      O => U_DCT2D_databuf_reg_1_2_CYMUXG2
    );
  U_DCT2D_databuf_reg_1_2_CY0G_580 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_3_Q,
      O => U_DCT2D_databuf_reg_1_2_CY0G
    );
  U_DCT2D_databuf_reg_1_2_CYSELG_581 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx2412z1,
      O => U_DCT2D_databuf_reg_1_2_CYSELG
    );
  U_DCT2D_databuf_reg_1_2_SRINV_582 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_1_2_SRINV
    );
  U_DCT2D_databuf_reg_1_2_CLKINV_583 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_1_2_CLKINV
    );
  U_DCT2D_databuf_reg_1_2_CEINV_584 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_1_2_CEINV
    );
  U_DCT2D_databuf_reg_1_4_DXMUX_585 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_4_XORF,
      O => U_DCT2D_databuf_reg_1_4_DXMUX
    );
  U_DCT2D_databuf_reg_1_4_XORF_586 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_4_CYINIT,
      I1 => U_DCT2D_nx3409z1,
      O => U_DCT2D_databuf_reg_1_4_XORF
    );
  U_DCT2D_databuf_reg_1_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_4_CY0F,
      IB => U_DCT2D_databuf_reg_1_4_CYINIT,
      SEL => U_DCT2D_databuf_reg_1_4_CYSELF,
      O => U_DCT2D_rtlc5_1579_add_46_ix4406z63342_O
    );
  U_DCT2D_databuf_reg_1_4_CYMUXF2_587 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_4_CY0F,
      IB => U_DCT2D_databuf_reg_1_4_CY0F,
      SEL => U_DCT2D_databuf_reg_1_4_CYSELF,
      O => U_DCT2D_databuf_reg_1_4_CYMUXF2
    );
  U_DCT2D_databuf_reg_1_4_CYINIT_588 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1579_add_46_ix3409z63342_O,
      O => U_DCT2D_databuf_reg_1_4_CYINIT
    );
  U_DCT2D_databuf_reg_1_4_CY0F_589 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_4_Q,
      O => U_DCT2D_databuf_reg_1_4_CY0F
    );
  U_DCT2D_databuf_reg_1_4_CYSELF_590 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx3409z1,
      O => U_DCT2D_databuf_reg_1_4_CYSELF
    );
  U_DCT2D_databuf_reg_1_4_DYMUX_591 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_4_XORG,
      O => U_DCT2D_databuf_reg_1_4_DYMUX
    );
  U_DCT2D_databuf_reg_1_4_XORG_592 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1579_add_46_ix4406z63342_O,
      I1 => U_DCT2D_nx4406z1,
      O => U_DCT2D_databuf_reg_1_4_XORG
    );
  U_DCT2D_databuf_reg_1_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_4_CYMUXFAST,
      O => U_DCT2D_rtlc5_1579_add_46_ix5403z63342_O
    );
  U_DCT2D_databuf_reg_1_4_FASTCARRY_593 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1579_add_46_ix3409z63342_O,
      O => U_DCT2D_databuf_reg_1_4_FASTCARRY
    );
  U_DCT2D_databuf_reg_1_4_CYAND_594 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_1_4_CYSELG,
      I1 => U_DCT2D_databuf_reg_1_4_CYSELF,
      O => U_DCT2D_databuf_reg_1_4_CYAND
    );
  U_DCT2D_databuf_reg_1_4_CYMUXFAST_595 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_4_CYMUXG2,
      IB => U_DCT2D_databuf_reg_1_4_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_1_4_CYAND,
      O => U_DCT2D_databuf_reg_1_4_CYMUXFAST
    );
  U_DCT2D_databuf_reg_1_4_CYMUXG2_596 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_4_CY0G,
      IB => U_DCT2D_databuf_reg_1_4_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_1_4_CYSELG,
      O => U_DCT2D_databuf_reg_1_4_CYMUXG2
    );
  U_DCT2D_databuf_reg_1_4_CY0G_597 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_5_Q,
      O => U_DCT2D_databuf_reg_1_4_CY0G
    );
  U_DCT2D_databuf_reg_1_4_CYSELG_598 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx4406z1,
      O => U_DCT2D_databuf_reg_1_4_CYSELG
    );
  U_DCT2D_databuf_reg_1_4_SRINV_599 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_1_4_SRINV
    );
  U_DCT2D_databuf_reg_1_4_CLKINV_600 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_1_4_CLKINV
    );
  U_DCT2D_databuf_reg_1_4_CEINV_601 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_1_4_CEINV
    );
  U_DCT1D_ix62813z1321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_2_Q(3),
      ADR2 => U_DCT1D_latchbuf_reg_5_Q(3),
      ADR3 => VCC,
      O => U_DCT1D_nx62813z1
    );
  U_DCT2D_databuf_reg_1_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_1_6_FFX_RST
    );
  U_DCT2D_reg_databuf_reg_1_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_1_6_DXMUX,
      CE => U_DCT2D_databuf_reg_1_6_CEINV,
      CLK => U_DCT2D_databuf_reg_1_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_1_6_FFX_RST,
      O => U_DCT2D_databuf_reg_1_Q(6)
    );
  U_DCT2D_ix5403z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_1_6_Q,
      ADR1 => U_DCT2D_latchbuf_reg_6_6_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx5403z1
    );
  U_DCT2D_databuf_reg_1_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_1_6_FFY_RST
    );
  U_DCT2D_reg_databuf_reg_1_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_1_6_DYMUX,
      CE => U_DCT2D_databuf_reg_1_6_CEINV,
      CLK => U_DCT2D_databuf_reg_1_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_1_6_FFY_RST,
      O => U_DCT2D_databuf_reg_1_Q(7)
    );
  U_DCT2D_databuf_reg_1_6_DXMUX_602 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_6_XORF,
      O => U_DCT2D_databuf_reg_1_6_DXMUX
    );
  U_DCT2D_databuf_reg_1_6_XORF_603 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_6_CYINIT,
      I1 => U_DCT2D_nx5403z1,
      O => U_DCT2D_databuf_reg_1_6_XORF
    );
  U_DCT2D_databuf_reg_1_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_6_CY0F,
      IB => U_DCT2D_databuf_reg_1_6_CYINIT,
      SEL => U_DCT2D_databuf_reg_1_6_CYSELF,
      O => U_DCT2D_rtlc5_1579_add_46_ix6400z63342_O
    );
  U_DCT2D_databuf_reg_1_6_CYMUXF2_604 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_6_CY0F,
      IB => U_DCT2D_databuf_reg_1_6_CY0F,
      SEL => U_DCT2D_databuf_reg_1_6_CYSELF,
      O => U_DCT2D_databuf_reg_1_6_CYMUXF2
    );
  U_DCT2D_databuf_reg_1_6_CYINIT_605 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1579_add_46_ix5403z63342_O,
      O => U_DCT2D_databuf_reg_1_6_CYINIT
    );
  U_DCT2D_databuf_reg_1_6_CY0F_606 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_6_Q,
      O => U_DCT2D_databuf_reg_1_6_CY0F
    );
  U_DCT2D_databuf_reg_1_6_CYSELF_607 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx5403z1,
      O => U_DCT2D_databuf_reg_1_6_CYSELF
    );
  U_DCT2D_databuf_reg_1_6_DYMUX_608 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_6_XORG,
      O => U_DCT2D_databuf_reg_1_6_DYMUX
    );
  U_DCT2D_databuf_reg_1_6_XORG_609 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1579_add_46_ix6400z63342_O,
      I1 => U_DCT2D_nx6400z1,
      O => U_DCT2D_databuf_reg_1_6_XORG
    );
  U_DCT2D_databuf_reg_1_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_6_CYMUXFAST,
      O => U_DCT2D_rtlc5_1579_add_46_ix7397z63342_O
    );
  U_DCT2D_databuf_reg_1_6_FASTCARRY_610 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1579_add_46_ix5403z63342_O,
      O => U_DCT2D_databuf_reg_1_6_FASTCARRY
    );
  U_DCT2D_databuf_reg_1_6_CYAND_611 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_1_6_CYSELG,
      I1 => U_DCT2D_databuf_reg_1_6_CYSELF,
      O => U_DCT2D_databuf_reg_1_6_CYAND
    );
  U_DCT2D_databuf_reg_1_6_CYMUXFAST_612 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_6_CYMUXG2,
      IB => U_DCT2D_databuf_reg_1_6_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_1_6_CYAND,
      O => U_DCT2D_databuf_reg_1_6_CYMUXFAST
    );
  U_DCT2D_databuf_reg_1_6_CYMUXG2_613 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_6_CY0G,
      IB => U_DCT2D_databuf_reg_1_6_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_1_6_CYSELG,
      O => U_DCT2D_databuf_reg_1_6_CYMUXG2
    );
  U_DCT2D_databuf_reg_1_6_CY0G_614 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_7_Q,
      O => U_DCT2D_databuf_reg_1_6_CY0G
    );
  U_DCT2D_databuf_reg_1_6_CYSELG_615 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx6400z1,
      O => U_DCT2D_databuf_reg_1_6_CYSELG
    );
  U_DCT2D_databuf_reg_1_6_SRINV_616 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_1_6_SRINV
    );
  U_DCT2D_databuf_reg_1_6_CLKINV_617 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_1_6_CLKINV
    );
  U_DCT2D_databuf_reg_1_6_CEINV_618 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_1_6_CEINV
    );
  U_DCT2D_databuf_reg_1_8_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_1_8_FFY_RST
    );
  U_DCT2D_reg_databuf_reg_1_9_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_1_8_DYMUX,
      CE => U_DCT2D_databuf_reg_1_8_CEINV,
      CLK => U_DCT2D_databuf_reg_1_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_1_8_FFY_RST,
      O => U_DCT2D_databuf_reg_1_Q(9)
    );
  U_DCT2D_ix8394z1321 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_1_10_Q,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_6_10_Q,
      O => U_DCT2D_nx8394z1
    );
  U_DCT2D_databuf_reg_1_8_DXMUX_619 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_8_XORF,
      O => U_DCT2D_databuf_reg_1_8_DXMUX
    );
  U_DCT2D_databuf_reg_1_8_XORF_620 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_8_CYINIT,
      I1 => U_DCT2D_nx7397z1,
      O => U_DCT2D_databuf_reg_1_8_XORF
    );
  U_DCT2D_databuf_reg_1_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_8_CY0F,
      IB => U_DCT2D_databuf_reg_1_8_CYINIT,
      SEL => U_DCT2D_databuf_reg_1_8_CYSELF,
      O => U_DCT2D_rtlc5_1579_add_46_ix8394z63342_O
    );
  U_DCT2D_databuf_reg_1_8_CYMUXF2_621 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_8_CY0F,
      IB => U_DCT2D_databuf_reg_1_8_CY0F,
      SEL => U_DCT2D_databuf_reg_1_8_CYSELF,
      O => U_DCT2D_databuf_reg_1_8_CYMUXF2
    );
  U_DCT2D_databuf_reg_1_8_CYINIT_622 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1579_add_46_ix7397z63342_O,
      O => U_DCT2D_databuf_reg_1_8_CYINIT
    );
  U_DCT2D_databuf_reg_1_8_CY0F_623 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_8_Q,
      O => U_DCT2D_databuf_reg_1_8_CY0F
    );
  U_DCT2D_databuf_reg_1_8_CYSELF_624 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx7397z1,
      O => U_DCT2D_databuf_reg_1_8_CYSELF
    );
  U_DCT2D_databuf_reg_1_8_DYMUX_625 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_8_XORG,
      O => U_DCT2D_databuf_reg_1_8_DYMUX
    );
  U_DCT2D_databuf_reg_1_8_XORG_626 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1579_add_46_ix8394z63342_O,
      I1 => U_DCT2D_nx8394z1,
      O => U_DCT2D_databuf_reg_1_8_XORG
    );
  U_DCT2D_databuf_reg_1_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_8_CYMUXFAST,
      O => U_DCT2D_rtlc5_1579_add_46_ix30550z63342_O
    );
  U_DCT2D_databuf_reg_1_8_FASTCARRY_627 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1579_add_46_ix7397z63342_O,
      O => U_DCT2D_databuf_reg_1_8_FASTCARRY
    );
  U_DCT2D_databuf_reg_1_8_CYAND_628 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_1_8_CYSELG,
      I1 => U_DCT2D_databuf_reg_1_8_CYSELF,
      O => U_DCT2D_databuf_reg_1_8_CYAND
    );
  U_DCT2D_databuf_reg_1_8_CYMUXFAST_629 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_8_CYMUXG2,
      IB => U_DCT2D_databuf_reg_1_8_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_1_8_CYAND,
      O => U_DCT2D_databuf_reg_1_8_CYMUXFAST
    );
  U_DCT2D_databuf_reg_1_8_CYMUXG2_630 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_1_8_CY0G,
      IB => U_DCT2D_databuf_reg_1_8_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_1_8_CYSELG,
      O => U_DCT2D_databuf_reg_1_8_CYMUXG2
    );
  U_DCT2D_databuf_reg_1_8_CY0G_631 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_10_Q,
      O => U_DCT2D_databuf_reg_1_8_CY0G
    );
  U_DCT2D_databuf_reg_1_8_CYSELG_632 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx8394z1,
      O => U_DCT2D_databuf_reg_1_8_CYSELG
    );
  U_DCT2D_databuf_reg_1_8_SRINV_633 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_1_8_SRINV
    );
  U_DCT2D_databuf_reg_1_8_CLKINV_634 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_1_8_CLKINV
    );
  U_DCT2D_databuf_reg_1_8_CEINV_635 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_1_8_CEINV
    );
  U_DCT2D_nx30550z1_rt_636 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_nx30550z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx30550z1_rt
    );
  U_DCT2D_databuf_reg_1_10_DXMUX_637 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_10_XORF,
      O => U_DCT2D_databuf_reg_1_10_DXMUX
    );
  U_DCT2D_databuf_reg_1_10_XORF_638 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_10_CYINIT,
      I1 => U_DCT2D_nx30550z1_rt,
      O => U_DCT2D_databuf_reg_1_10_XORF
    );
  U_DCT2D_databuf_reg_1_10_CYINIT_639 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1579_add_46_ix30550z63342_O,
      O => U_DCT2D_databuf_reg_1_10_CYINIT
    );
  U_DCT2D_databuf_reg_1_10_CLKINV_640 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_1_10_CLKINV
    );
  U_DCT2D_databuf_reg_1_10_CEINV_641 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_1_10_CEINV
    );
  U_DCT1D_databuf_reg_4_0_DXMUX_642 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_0_XORF,
      O => U_DCT1D_databuf_reg_4_0_DXMUX
    );
  U_DCT1D_databuf_reg_4_0_XORF_643 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_0_CYINIT,
      I1 => U_DCT1D_nx49552z1,
      O => U_DCT1D_databuf_reg_4_0_XORF
    );
  U_DCT1D_databuf_reg_4_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_0_CY0F,
      IB => U_DCT1D_databuf_reg_4_0_CYINIT,
      SEL => U_DCT1D_databuf_reg_4_0_CYSELF,
      O => U_DCT1D_rtlc5_83_sub_4_ix50549z63342_O
    );
  U_DCT1D_databuf_reg_4_0_CYINIT_644 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GLOBAL_LOGIC1_5,
      O => U_DCT1D_databuf_reg_4_0_CYINIT
    );
  U_DCT1D_databuf_reg_4_0_CY0F_645 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(0),
      O => U_DCT1D_databuf_reg_4_0_CY0F
    );
  U_DCT1D_databuf_reg_4_0_CYSELF_646 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx49552z1,
      O => U_DCT1D_databuf_reg_4_0_CYSELF
    );
  U_DCT1D_databuf_reg_4_0_DYMUX_647 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_0_XORG,
      O => U_DCT1D_databuf_reg_4_0_DYMUX
    );
  U_DCT1D_databuf_reg_4_0_XORG_648 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_83_sub_4_ix50549z63342_O,
      I1 => U_DCT1D_nx50549z1,
      O => U_DCT1D_databuf_reg_4_0_XORG
    );
  U_DCT1D_databuf_reg_4_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_0_CYMUXG,
      O => U_DCT1D_rtlc5_83_sub_4_ix51546z63342_O
    );
  U_DCT1D_databuf_reg_4_0_CYMUXG_649 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_0_CY0G,
      IB => U_DCT1D_rtlc5_83_sub_4_ix50549z63342_O,
      SEL => U_DCT1D_databuf_reg_4_0_CYSELG,
      O => U_DCT1D_databuf_reg_4_0_CYMUXG
    );
  U_DCT1D_databuf_reg_4_0_CY0G_650 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(1),
      O => U_DCT1D_databuf_reg_4_0_CY0G
    );
  U_DCT1D_databuf_reg_4_0_CYSELG_651 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx50549z1,
      O => U_DCT1D_databuf_reg_4_0_CYSELG
    );
  U_DCT1D_databuf_reg_4_0_SRINV_652 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_4_0_SRINV
    );
  U_DCT1D_databuf_reg_4_0_CLKINV_653 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_4_0_CLKINV
    );
  U_DCT1D_databuf_reg_4_0_CEINV_654 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_4_0_CEINV
    );
  U_DCT1D_databuf_reg_4_2_DXMUX_655 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_2_XORF,
      O => U_DCT1D_databuf_reg_4_2_DXMUX
    );
  U_DCT1D_databuf_reg_4_2_XORF_656 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_2_CYINIT,
      I1 => U_DCT1D_nx51546z1,
      O => U_DCT1D_databuf_reg_4_2_XORF
    );
  U_DCT1D_databuf_reg_4_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_2_CY0F,
      IB => U_DCT1D_databuf_reg_4_2_CYINIT,
      SEL => U_DCT1D_databuf_reg_4_2_CYSELF,
      O => U_DCT1D_rtlc5_83_sub_4_ix52543z63342_O
    );
  U_DCT1D_databuf_reg_4_2_CYMUXF2_657 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_2_CY0F,
      IB => U_DCT1D_databuf_reg_4_2_CY0F,
      SEL => U_DCT1D_databuf_reg_4_2_CYSELF,
      O => U_DCT1D_databuf_reg_4_2_CYMUXF2
    );
  U_DCT1D_databuf_reg_4_2_CYINIT_658 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_83_sub_4_ix51546z63342_O,
      O => U_DCT1D_databuf_reg_4_2_CYINIT
    );
  U_DCT1D_databuf_reg_4_2_CY0F_659 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(2),
      O => U_DCT1D_databuf_reg_4_2_CY0F
    );
  U_DCT1D_databuf_reg_4_2_CYSELF_660 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx51546z1,
      O => U_DCT1D_databuf_reg_4_2_CYSELF
    );
  U_DCT1D_databuf_reg_4_2_DYMUX_661 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_2_XORG,
      O => U_DCT1D_databuf_reg_4_2_DYMUX
    );
  U_DCT1D_databuf_reg_4_2_XORG_662 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_83_sub_4_ix52543z63342_O,
      I1 => U_DCT1D_nx52543z1,
      O => U_DCT1D_databuf_reg_4_2_XORG
    );
  U_DCT1D_databuf_reg_4_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_2_CYMUXFAST,
      O => U_DCT1D_rtlc5_83_sub_4_ix53540z63342_O
    );
  U_DCT1D_databuf_reg_4_2_FASTCARRY_663 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_83_sub_4_ix51546z63342_O,
      O => U_DCT1D_databuf_reg_4_2_FASTCARRY
    );
  U_DCT1D_databuf_reg_4_2_CYAND_664 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_4_2_CYSELG,
      I1 => U_DCT1D_databuf_reg_4_2_CYSELF,
      O => U_DCT1D_databuf_reg_4_2_CYAND
    );
  U_DCT1D_databuf_reg_4_2_CYMUXFAST_665 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_2_CYMUXG2,
      IB => U_DCT1D_databuf_reg_4_2_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_4_2_CYAND,
      O => U_DCT1D_databuf_reg_4_2_CYMUXFAST
    );
  U_DCT1D_databuf_reg_4_2_CYMUXG2_666 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_2_CY0G,
      IB => U_DCT1D_databuf_reg_4_2_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_4_2_CYSELG,
      O => U_DCT1D_databuf_reg_4_2_CYMUXG2
    );
  U_DCT1D_databuf_reg_4_2_CY0G_667 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(3),
      O => U_DCT1D_databuf_reg_4_2_CY0G
    );
  U_DCT1D_databuf_reg_4_2_CYSELG_668 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx52543z1,
      O => U_DCT1D_databuf_reg_4_2_CYSELG
    );
  U_DCT1D_databuf_reg_4_2_SRINV_669 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_4_2_SRINV
    );
  U_DCT1D_databuf_reg_4_2_CLKINV_670 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_4_2_CLKINV
    );
  U_DCT1D_databuf_reg_4_2_CEINV_671 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_4_2_CEINV
    );
  U_DCT1D_databuf_reg_4_4_DXMUX_672 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_4_XORF,
      O => U_DCT1D_databuf_reg_4_4_DXMUX
    );
  U_DCT1D_databuf_reg_4_4_XORF_673 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_4_CYINIT,
      I1 => U_DCT1D_nx53540z1,
      O => U_DCT1D_databuf_reg_4_4_XORF
    );
  U_DCT1D_databuf_reg_4_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_4_CY0F,
      IB => U_DCT1D_databuf_reg_4_4_CYINIT,
      SEL => U_DCT1D_databuf_reg_4_4_CYSELF,
      O => U_DCT1D_rtlc5_83_sub_4_ix54537z63342_O
    );
  U_DCT1D_databuf_reg_4_4_CYMUXF2_674 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_4_CY0F,
      IB => U_DCT1D_databuf_reg_4_4_CY0F,
      SEL => U_DCT1D_databuf_reg_4_4_CYSELF,
      O => U_DCT1D_databuf_reg_4_4_CYMUXF2
    );
  U_DCT1D_databuf_reg_4_4_CYINIT_675 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_83_sub_4_ix53540z63342_O,
      O => U_DCT1D_databuf_reg_4_4_CYINIT
    );
  U_DCT1D_databuf_reg_4_4_CY0F_676 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(4),
      O => U_DCT1D_databuf_reg_4_4_CY0F
    );
  U_DCT1D_databuf_reg_4_4_CYSELF_677 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx53540z1,
      O => U_DCT1D_databuf_reg_4_4_CYSELF
    );
  U_DCT1D_databuf_reg_4_4_DYMUX_678 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_4_XORG,
      O => U_DCT1D_databuf_reg_4_4_DYMUX
    );
  U_DCT1D_databuf_reg_4_4_XORG_679 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_83_sub_4_ix54537z63342_O,
      I1 => U_DCT1D_nx54537z1,
      O => U_DCT1D_databuf_reg_4_4_XORG
    );
  U_DCT1D_databuf_reg_4_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_4_CYMUXFAST,
      O => U_DCT1D_rtlc5_83_sub_4_ix55534z63342_O
    );
  U_DCT1D_databuf_reg_4_4_FASTCARRY_680 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_83_sub_4_ix53540z63342_O,
      O => U_DCT1D_databuf_reg_4_4_FASTCARRY
    );
  U_DCT1D_databuf_reg_4_4_CYAND_681 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_4_4_CYSELG,
      I1 => U_DCT1D_databuf_reg_4_4_CYSELF,
      O => U_DCT1D_databuf_reg_4_4_CYAND
    );
  U_DCT1D_databuf_reg_4_4_CYMUXFAST_682 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_4_CYMUXG2,
      IB => U_DCT1D_databuf_reg_4_4_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_4_4_CYAND,
      O => U_DCT1D_databuf_reg_4_4_CYMUXFAST
    );
  U_DCT1D_databuf_reg_4_4_CYMUXG2_683 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_4_CY0G,
      IB => U_DCT1D_databuf_reg_4_4_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_4_4_CYSELG,
      O => U_DCT1D_databuf_reg_4_4_CYMUXG2
    );
  U_DCT1D_databuf_reg_4_4_CY0G_684 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(5),
      O => U_DCT1D_databuf_reg_4_4_CY0G
    );
  U_DCT1D_databuf_reg_4_4_CYSELG_685 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx54537z1,
      O => U_DCT1D_databuf_reg_4_4_CYSELG
    );
  U_DCT1D_databuf_reg_4_4_SRINV_686 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_4_4_SRINV
    );
  U_DCT1D_databuf_reg_4_4_CLKINV_687 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_4_4_CLKINV
    );
  U_DCT1D_databuf_reg_4_4_CEINV_688 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_4_4_CEINV
    );
  U_DCT1D_databuf_reg_4_6_DXMUX_689 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_6_XORF,
      O => U_DCT1D_databuf_reg_4_6_DXMUX
    );
  U_DCT1D_databuf_reg_4_6_XORF_690 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_6_CYINIT,
      I1 => U_DCT1D_nx55534z1,
      O => U_DCT1D_databuf_reg_4_6_XORF
    );
  U_DCT1D_databuf_reg_4_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_6_CY0F,
      IB => U_DCT1D_databuf_reg_4_6_CYINIT,
      SEL => U_DCT1D_databuf_reg_4_6_CYSELF,
      O => U_DCT1D_rtlc5_83_sub_4_ix56531z63342_O
    );
  U_DCT1D_databuf_reg_4_6_CYMUXF2_691 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_6_CY0F,
      IB => U_DCT1D_databuf_reg_4_6_CY0F,
      SEL => U_DCT1D_databuf_reg_4_6_CYSELF,
      O => U_DCT1D_databuf_reg_4_6_CYMUXF2
    );
  U_DCT1D_databuf_reg_4_6_CYINIT_692 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_83_sub_4_ix55534z63342_O,
      O => U_DCT1D_databuf_reg_4_6_CYINIT
    );
  U_DCT1D_databuf_reg_4_6_CY0F_693 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(6),
      O => U_DCT1D_databuf_reg_4_6_CY0F
    );
  U_DCT1D_databuf_reg_4_6_CYSELF_694 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx55534z1,
      O => U_DCT1D_databuf_reg_4_6_CYSELF
    );
  U_DCT1D_databuf_reg_4_6_DYMUX_695 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_6_XORG,
      O => U_DCT1D_databuf_reg_4_6_DYMUX
    );
  U_DCT1D_databuf_reg_4_6_XORG_696 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_83_sub_4_ix56531z63342_O,
      I1 => U_DCT1D_nx56531z1,
      O => U_DCT1D_databuf_reg_4_6_XORG
    );
  U_DCT1D_databuf_reg_4_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_6_CYMUXFAST,
      O => U_DCT1D_rtlc5_83_sub_4_ix57528z63342_O
    );
  U_DCT1D_databuf_reg_4_6_FASTCARRY_697 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_83_sub_4_ix55534z63342_O,
      O => U_DCT1D_databuf_reg_4_6_FASTCARRY
    );
  U_DCT1D_databuf_reg_4_6_CYAND_698 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_4_6_CYSELG,
      I1 => U_DCT1D_databuf_reg_4_6_CYSELF,
      O => U_DCT1D_databuf_reg_4_6_CYAND
    );
  U_DCT1D_databuf_reg_4_6_CYMUXFAST_699 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_6_CYMUXG2,
      IB => U_DCT1D_databuf_reg_4_6_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_4_6_CYAND,
      O => U_DCT1D_databuf_reg_4_6_CYMUXFAST
    );
  U_DCT1D_databuf_reg_4_6_CYMUXG2_700 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_4_6_CY0G,
      IB => U_DCT1D_databuf_reg_4_6_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_4_6_CYSELG,
      O => U_DCT1D_databuf_reg_4_6_CYMUXG2
    );
  U_DCT1D_databuf_reg_4_6_CY0G_701 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(7),
      O => U_DCT1D_databuf_reg_4_6_CY0G
    );
  U_DCT1D_databuf_reg_4_6_CYSELG_702 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx56531z1,
      O => U_DCT1D_databuf_reg_4_6_CYSELG
    );
  U_DCT1D_databuf_reg_4_6_SRINV_703 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_4_6_SRINV
    );
  U_DCT1D_databuf_reg_4_6_CLKINV_704 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_4_6_CLKINV
    );
  U_DCT1D_databuf_reg_4_6_CEINV_705 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_4_6_CEINV
    );
  U_DCT1D_databuf_reg_4_8_DXMUX_706 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_8_XORF,
      O => U_DCT1D_databuf_reg_4_8_DXMUX
    );
  U_DCT1D_databuf_reg_4_8_XORF_707 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_8_CYINIT,
      I1 => U_DCT1D_nx57528z1_rt,
      O => U_DCT1D_databuf_reg_4_8_XORF
    );
  U_DCT1D_databuf_reg_4_8_CYINIT_708 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_83_sub_4_ix57528z63342_O,
      O => U_DCT1D_databuf_reg_4_8_CYINIT
    );
  U_DCT1D_databuf_reg_4_8_CLKINV_709 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_4_8_CLKINV
    );
  U_DCT1D_databuf_reg_4_8_CEINV_710 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_4_8_CEINV
    );
  U_DCT2D_ix65206z1463 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao0_s(2),
      ADR2 => romo2datao1_s(1),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z117
    );
  U_DCT2D_ix65206z1466 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao0_s(1),
      ADR2 => romo2datao1_s(0),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z120
    );
  U_DCT2D_rtlc5n1480_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_2_CY0F,
      IB => U_DCT2D_rtlc5n1480_2_CYINIT,
      SEL => U_DCT2D_rtlc5n1480_2_CYSELF,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63485_O
    );
  U_DCT2D_rtlc5n1480_2_CYINIT_711 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_2_BXINVNOT,
      O => U_DCT2D_rtlc5n1480_2_CYINIT
    );
  U_DCT2D_rtlc5n1480_2_CY0F_712 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(1),
      O => U_DCT2D_rtlc5n1480_2_CY0F
    );
  U_DCT2D_rtlc5n1480_2_CYSELF_713 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z120,
      O => U_DCT2D_rtlc5n1480_2_CYSELF
    );
  U_DCT2D_rtlc5n1480_2_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_31,
      O => U_DCT2D_rtlc5n1480_2_BXINVNOT
    );
  U_DCT2D_rtlc5n1480_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_2_XORG,
      O => U_DCT2D_rtlc5n1480(2)
    );
  U_DCT2D_rtlc5n1480_2_XORG_714 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_331_add_54_ix65206z63485_O,
      I1 => U_DCT2D_nx65206z117,
      O => U_DCT2D_rtlc5n1480_2_XORG
    );
  U_DCT2D_rtlc5n1480_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_2_CYMUXG,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63482_O
    );
  U_DCT2D_rtlc5n1480_2_CYMUXG_715 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_2_CY0G,
      IB => U_DCT2D_rtlc_331_add_54_ix65206z63485_O,
      SEL => U_DCT2D_rtlc5n1480_2_CYSELG,
      O => U_DCT2D_rtlc5n1480_2_CYMUXG
    );
  U_DCT2D_rtlc5n1480_2_CY0G_716 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(2),
      O => U_DCT2D_rtlc5n1480_2_CY0G
    );
  U_DCT2D_rtlc5n1480_2_CYSELG_717 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z117,
      O => U_DCT2D_rtlc5n1480_2_CYSELG
    );
  U_DCT2D_ix65206z1455 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao1_s(3),
      ADR1 => romo2datao0_s(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z111
    );
  U_DCT2D_ix65206z1601 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao0_s(3),
      ADR1 => romo2datao1_s(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z114
    );
  U_DCT2D_rtlc5n1480_3_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_3_XORF,
      O => U_DCT2D_rtlc5n1480(3)
    );
  U_DCT2D_rtlc5n1480_3_XORF_718 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1480_3_CYINIT,
      I1 => U_DCT2D_nx65206z114,
      O => U_DCT2D_rtlc5n1480_3_XORF
    );
  U_DCT2D_rtlc5n1480_3_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_3_CY0F,
      IB => U_DCT2D_rtlc5n1480_3_CYINIT,
      SEL => U_DCT2D_rtlc5n1480_3_CYSELF,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63478_O
    );
  U_DCT2D_rtlc5n1480_3_CYMUXF2_719 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_3_CY0F,
      IB => U_DCT2D_rtlc5n1480_3_CY0F,
      SEL => U_DCT2D_rtlc5n1480_3_CYSELF,
      O => U_DCT2D_rtlc5n1480_3_CYMUXF2
    );
  U_DCT2D_rtlc5n1480_3_CYINIT_720 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63482_O,
      O => U_DCT2D_rtlc5n1480_3_CYINIT
    );
  U_DCT2D_rtlc5n1480_3_CY0F_721 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(3),
      O => U_DCT2D_rtlc5n1480_3_CY0F
    );
  U_DCT2D_rtlc5n1480_3_CYSELF_722 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z114,
      O => U_DCT2D_rtlc5n1480_3_CYSELF
    );
  U_DCT2D_rtlc5n1480_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_3_XORG,
      O => U_DCT2D_rtlc5n1480(4)
    );
  U_DCT2D_rtlc5n1480_3_XORG_723 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_331_add_54_ix65206z63478_O,
      I1 => U_DCT2D_nx65206z111,
      O => U_DCT2D_rtlc5n1480_3_XORG
    );
  U_DCT2D_rtlc5n1480_3_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_3_CYMUXFAST,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63474_O
    );
  U_DCT2D_rtlc5n1480_3_FASTCARRY_724 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63482_O,
      O => U_DCT2D_rtlc5n1480_3_FASTCARRY
    );
  U_DCT2D_rtlc5n1480_3_CYAND_725 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1480_3_CYSELG,
      I1 => U_DCT2D_rtlc5n1480_3_CYSELF,
      O => U_DCT2D_rtlc5n1480_3_CYAND
    );
  U_DCT2D_rtlc5n1480_3_CYMUXFAST_726 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_3_CYMUXG2,
      IB => U_DCT2D_rtlc5n1480_3_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1480_3_CYAND,
      O => U_DCT2D_rtlc5n1480_3_CYMUXFAST
    );
  U_DCT2D_rtlc5n1480_3_CYMUXG2_727 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_3_CY0G,
      IB => U_DCT2D_rtlc5n1480_3_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1480_3_CYSELG,
      O => U_DCT2D_rtlc5n1480_3_CYMUXG2
    );
  U_DCT2D_rtlc5n1480_3_CY0G_728 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(4),
      O => U_DCT2D_rtlc5n1480_3_CY0G
    );
  U_DCT2D_rtlc5n1480_3_CYSELG_729 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z111,
      O => U_DCT2D_rtlc5n1480_3_CYSELG
    );
  U_DCT2D_ix65206z1452 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao0_s(5),
      ADR2 => romo2datao1_s(4),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z108
    );
  U_DCT2D_ix65206z1448 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao0_s(6),
      ADR1 => romo2datao1_s(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z105
    );
  U_DCT2D_rtlc5n1480_5_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_5_XORF,
      O => U_DCT2D_rtlc5n1480(5)
    );
  U_DCT2D_rtlc5n1480_5_XORF_730 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1480_5_CYINIT,
      I1 => U_DCT2D_nx65206z108,
      O => U_DCT2D_rtlc5n1480_5_XORF
    );
  U_DCT2D_rtlc5n1480_5_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_5_CY0F,
      IB => U_DCT2D_rtlc5n1480_5_CYINIT,
      SEL => U_DCT2D_rtlc5n1480_5_CYSELF,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63471_O
    );
  U_DCT2D_rtlc5n1480_5_CYMUXF2_731 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_5_CY0F,
      IB => U_DCT2D_rtlc5n1480_5_CY0F,
      SEL => U_DCT2D_rtlc5n1480_5_CYSELF,
      O => U_DCT2D_rtlc5n1480_5_CYMUXF2
    );
  U_DCT2D_rtlc5n1480_5_CYINIT_732 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63474_O,
      O => U_DCT2D_rtlc5n1480_5_CYINIT
    );
  U_DCT2D_rtlc5n1480_5_CY0F_733 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(5),
      O => U_DCT2D_rtlc5n1480_5_CY0F
    );
  U_DCT2D_rtlc5n1480_5_CYSELF_734 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z108,
      O => U_DCT2D_rtlc5n1480_5_CYSELF
    );
  U_DCT2D_rtlc5n1480_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_5_XORG,
      O => U_DCT2D_rtlc5n1480(6)
    );
  U_DCT2D_rtlc5n1480_5_XORG_735 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_331_add_54_ix65206z63471_O,
      I1 => U_DCT2D_nx65206z105,
      O => U_DCT2D_rtlc5n1480_5_XORG
    );
  U_DCT2D_rtlc5n1480_5_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_5_CYMUXFAST,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63467_O
    );
  U_DCT2D_rtlc5n1480_5_FASTCARRY_736 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63474_O,
      O => U_DCT2D_rtlc5n1480_5_FASTCARRY
    );
  U_DCT2D_rtlc5n1480_5_CYAND_737 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1480_5_CYSELG,
      I1 => U_DCT2D_rtlc5n1480_5_CYSELF,
      O => U_DCT2D_rtlc5n1480_5_CYAND
    );
  U_DCT2D_rtlc5n1480_5_CYMUXFAST_738 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_5_CYMUXG2,
      IB => U_DCT2D_rtlc5n1480_5_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1480_5_CYAND,
      O => U_DCT2D_rtlc5n1480_5_CYMUXFAST
    );
  U_DCT2D_rtlc5n1480_5_CYMUXG2_739 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_5_CY0G,
      IB => U_DCT2D_rtlc5n1480_5_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1480_5_CYSELG,
      O => U_DCT2D_rtlc5n1480_5_CYMUXG2
    );
  U_DCT2D_rtlc5n1480_5_CY0G_740 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(6),
      O => U_DCT2D_rtlc5n1480_5_CY0G
    );
  U_DCT2D_rtlc5n1480_5_CYSELG_741 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z105,
      O => U_DCT2D_rtlc5n1480_5_CYSELG
    );
  U_DCT2D_ix65206z1444 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2datao0_s(7),
      ADR1 => VCC,
      ADR2 => romo2datao1_s(6),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z102
    );
  U_DCT2D_ix65206z1441 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao0_s(8),
      ADR2 => VCC,
      ADR3 => romo2datao1_s(7),
      O => U_DCT2D_nx65206z99
    );
  U_DCT2D_rtlc5n1480_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_7_XORF,
      O => U_DCT2D_rtlc5n1480(7)
    );
  U_DCT2D_rtlc5n1480_7_XORF_742 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1480_7_CYINIT,
      I1 => U_DCT2D_nx65206z102,
      O => U_DCT2D_rtlc5n1480_7_XORF
    );
  U_DCT2D_rtlc5n1480_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_7_CY0F,
      IB => U_DCT2D_rtlc5n1480_7_CYINIT,
      SEL => U_DCT2D_rtlc5n1480_7_CYSELF,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63463_O
    );
  U_DCT2D_rtlc5n1480_7_CYMUXF2_743 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_7_CY0F,
      IB => U_DCT2D_rtlc5n1480_7_CY0F,
      SEL => U_DCT2D_rtlc5n1480_7_CYSELF,
      O => U_DCT2D_rtlc5n1480_7_CYMUXF2
    );
  U_DCT2D_rtlc5n1480_7_CYINIT_744 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63467_O,
      O => U_DCT2D_rtlc5n1480_7_CYINIT
    );
  U_DCT2D_rtlc5n1480_7_CY0F_745 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(7),
      O => U_DCT2D_rtlc5n1480_7_CY0F
    );
  U_DCT2D_rtlc5n1480_7_CYSELF_746 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z102,
      O => U_DCT2D_rtlc5n1480_7_CYSELF
    );
  U_DCT2D_rtlc5n1480_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_7_XORG,
      O => U_DCT2D_rtlc5n1480(8)
    );
  U_DCT2D_rtlc5n1480_7_XORG_747 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_331_add_54_ix65206z63463_O,
      I1 => U_DCT2D_nx65206z99,
      O => U_DCT2D_rtlc5n1480_7_XORG
    );
  U_DCT2D_rtlc5n1480_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_7_CYMUXFAST,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63460_O
    );
  U_DCT2D_rtlc5n1480_7_FASTCARRY_748 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63467_O,
      O => U_DCT2D_rtlc5n1480_7_FASTCARRY
    );
  U_DCT2D_rtlc5n1480_7_CYAND_749 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1480_7_CYSELG,
      I1 => U_DCT2D_rtlc5n1480_7_CYSELF,
      O => U_DCT2D_rtlc5n1480_7_CYAND
    );
  U_DCT2D_rtlc5n1480_7_CYMUXFAST_750 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_7_CYMUXG2,
      IB => U_DCT2D_rtlc5n1480_7_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1480_7_CYAND,
      O => U_DCT2D_rtlc5n1480_7_CYMUXFAST
    );
  U_DCT2D_rtlc5n1480_7_CYMUXG2_751 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_7_CY0G,
      IB => U_DCT2D_rtlc5n1480_7_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1480_7_CYSELG,
      O => U_DCT2D_rtlc5n1480_7_CYMUXG2
    );
  U_DCT2D_rtlc5n1480_7_CY0G_752 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(8),
      O => U_DCT2D_rtlc5n1480_7_CY0G
    );
  U_DCT2D_rtlc5n1480_7_CYSELG_753 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z99,
      O => U_DCT2D_rtlc5n1480_7_CYSELG
    );
  U_DCT2D_ix65206z1434 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao1_s(9),
      ADR1 => romo2datao0_s(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z93
    );
  U_DCT2D_rtlc5n1480_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_9_XORF,
      O => U_DCT2D_rtlc5n1480(9)
    );
  U_DCT2D_rtlc5n1480_9_XORF_754 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1480_9_CYINIT,
      I1 => U_DCT2D_nx65206z96,
      O => U_DCT2D_rtlc5n1480_9_XORF
    );
  U_DCT2D_rtlc5n1480_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_9_CY0F,
      IB => U_DCT2D_rtlc5n1480_9_CYINIT,
      SEL => U_DCT2D_rtlc5n1480_9_CYSELF,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63456_O
    );
  U_DCT2D_rtlc5n1480_9_CYMUXF2_755 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_9_CY0F,
      IB => U_DCT2D_rtlc5n1480_9_CY0F,
      SEL => U_DCT2D_rtlc5n1480_9_CYSELF,
      O => U_DCT2D_rtlc5n1480_9_CYMUXF2
    );
  U_DCT2D_rtlc5n1480_9_CYINIT_756 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63460_O,
      O => U_DCT2D_rtlc5n1480_9_CYINIT
    );
  U_DCT2D_rtlc5n1480_9_CY0F_757 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(9),
      O => U_DCT2D_rtlc5n1480_9_CY0F
    );
  U_DCT2D_rtlc5n1480_9_CYSELF_758 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z96,
      O => U_DCT2D_rtlc5n1480_9_CYSELF
    );
  U_DCT2D_rtlc5n1480_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_9_XORG,
      O => U_DCT2D_rtlc5n1480(10)
    );
  U_DCT2D_rtlc5n1480_9_XORG_759 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_331_add_54_ix65206z63456_O,
      I1 => U_DCT2D_nx65206z93,
      O => U_DCT2D_rtlc5n1480_9_XORG
    );
  U_DCT2D_rtlc5n1480_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_9_CYMUXFAST,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63453_O
    );
  U_DCT2D_rtlc5n1480_9_FASTCARRY_760 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63460_O,
      O => U_DCT2D_rtlc5n1480_9_FASTCARRY
    );
  U_DCT2D_rtlc5n1480_9_CYAND_761 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1480_9_CYSELG,
      I1 => U_DCT2D_rtlc5n1480_9_CYSELF,
      O => U_DCT2D_rtlc5n1480_9_CYAND
    );
  U_DCT2D_rtlc5n1480_9_CYMUXFAST_762 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_9_CYMUXG2,
      IB => U_DCT2D_rtlc5n1480_9_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1480_9_CYAND,
      O => U_DCT2D_rtlc5n1480_9_CYMUXFAST
    );
  U_DCT2D_rtlc5n1480_9_CYMUXG2_763 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_9_CY0G,
      IB => U_DCT2D_rtlc5n1480_9_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1480_9_CYSELG,
      O => U_DCT2D_rtlc5n1480_9_CYMUXG2
    );
  U_DCT2D_rtlc5n1480_9_CY0G_764 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(10),
      O => U_DCT2D_rtlc5n1480_9_CY0G
    );
  U_DCT2D_rtlc5n1480_9_CYSELG_765 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z93,
      O => U_DCT2D_rtlc5n1480_9_CYSELG
    );
  U_DCT2D_ix65206z1427 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao0_s(12),
      ADR2 => VCC,
      ADR3 => romo2datao1_s(11),
      O => U_DCT2D_nx65206z87
    );
  U_DCT2D_rtlc5n1480_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_11_XORF,
      O => U_DCT2D_rtlc5n1480(11)
    );
  U_DCT2D_rtlc5n1480_11_XORF_766 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1480_11_CYINIT,
      I1 => U_DCT2D_nx65206z90,
      O => U_DCT2D_rtlc5n1480_11_XORF
    );
  U_DCT2D_rtlc5n1480_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_11_CY0F,
      IB => U_DCT2D_rtlc5n1480_11_CYINIT,
      SEL => U_DCT2D_rtlc5n1480_11_CYSELF,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63449_O
    );
  U_DCT2D_rtlc5n1480_11_CYMUXF2_767 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_11_CY0F,
      IB => U_DCT2D_rtlc5n1480_11_CY0F,
      SEL => U_DCT2D_rtlc5n1480_11_CYSELF,
      O => U_DCT2D_rtlc5n1480_11_CYMUXF2
    );
  U_DCT2D_rtlc5n1480_11_CYINIT_768 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63453_O,
      O => U_DCT2D_rtlc5n1480_11_CYINIT
    );
  U_DCT2D_rtlc5n1480_11_CY0F_769 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(11),
      O => U_DCT2D_rtlc5n1480_11_CY0F
    );
  U_DCT2D_rtlc5n1480_11_CYSELF_770 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z90,
      O => U_DCT2D_rtlc5n1480_11_CYSELF
    );
  U_DCT2D_rtlc5n1480_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_11_XORG,
      O => U_DCT2D_rtlc5n1480(12)
    );
  U_DCT2D_rtlc5n1480_11_XORG_771 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_331_add_54_ix65206z63449_O,
      I1 => U_DCT2D_nx65206z87,
      O => U_DCT2D_rtlc5n1480_11_XORG
    );
  U_DCT2D_rtlc5n1480_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_11_CYMUXFAST,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63446_O
    );
  U_DCT2D_rtlc5n1480_11_FASTCARRY_772 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63453_O,
      O => U_DCT2D_rtlc5n1480_11_FASTCARRY
    );
  U_DCT2D_rtlc5n1480_11_CYAND_773 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1480_11_CYSELG,
      I1 => U_DCT2D_rtlc5n1480_11_CYSELF,
      O => U_DCT2D_rtlc5n1480_11_CYAND
    );
  U_DCT2D_rtlc5n1480_11_CYMUXFAST_774 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_11_CYMUXG2,
      IB => U_DCT2D_rtlc5n1480_11_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1480_11_CYAND,
      O => U_DCT2D_rtlc5n1480_11_CYMUXFAST
    );
  U_DCT2D_rtlc5n1480_11_CYMUXG2_775 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_11_CY0G,
      IB => U_DCT2D_rtlc5n1480_11_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1480_11_CYSELG,
      O => U_DCT2D_rtlc5n1480_11_CYMUXG2
    );
  U_DCT2D_rtlc5n1480_11_CY0G_776 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(12),
      O => U_DCT2D_rtlc5n1480_11_CY0G
    );
  U_DCT2D_rtlc5n1480_11_CYSELG_777 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z87,
      O => U_DCT2D_rtlc5n1480_11_CYSELG
    );
  U_DCT2D_rtlc5n1480_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_13_XORF,
      O => U_DCT2D_rtlc5n1480(13)
    );
  U_DCT2D_rtlc5n1480_13_XORF_778 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1480_13_CYINIT,
      I1 => U_DCT2D_nx65206z84,
      O => U_DCT2D_rtlc5n1480_13_XORF
    );
  U_DCT2D_rtlc5n1480_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_13_CY0F,
      IB => U_DCT2D_rtlc5n1480_13_CYINIT,
      SEL => U_DCT2D_rtlc5n1480_13_CYSELF,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63442_O
    );
  U_DCT2D_rtlc5n1480_13_CYMUXF2_779 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_13_CY0F,
      IB => U_DCT2D_rtlc5n1480_13_CY0F,
      SEL => U_DCT2D_rtlc5n1480_13_CYSELF,
      O => U_DCT2D_rtlc5n1480_13_CYMUXF2
    );
  U_DCT2D_rtlc5n1480_13_CYINIT_780 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63446_O,
      O => U_DCT2D_rtlc5n1480_13_CYINIT
    );
  U_DCT2D_rtlc5n1480_13_CY0F_781 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(13),
      O => U_DCT2D_rtlc5n1480_13_CY0F
    );
  U_DCT2D_rtlc5n1480_13_CYSELF_782 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z84,
      O => U_DCT2D_rtlc5n1480_13_CYSELF
    );
  U_DCT2D_rtlc5n1480_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_13_XORG,
      O => U_DCT2D_rtlc5n1480(14)
    );
  U_DCT2D_rtlc5n1480_13_XORG_783 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_331_add_54_ix65206z63442_O,
      I1 => U_DCT2D_nx65206z81,
      O => U_DCT2D_rtlc5n1480_13_XORG
    );
  U_DCT2D_rtlc5n1480_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_13_CYMUXFAST,
      O => U_DCT2D_rtlc_331_add_54_ix65206z63439_O
    );
  U_DCT2D_rtlc5n1480_13_FASTCARRY_784 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63446_O,
      O => U_DCT2D_rtlc5n1480_13_FASTCARRY
    );
  U_DCT2D_rtlc5n1480_13_CYAND_785 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1480_13_CYSELG,
      I1 => U_DCT2D_rtlc5n1480_13_CYSELF,
      O => U_DCT2D_rtlc5n1480_13_CYAND
    );
  U_DCT2D_rtlc5n1480_13_CYMUXFAST_786 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_13_CYMUXG2,
      IB => U_DCT2D_rtlc5n1480_13_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1480_13_CYAND,
      O => U_DCT2D_rtlc5n1480_13_CYMUXFAST
    );
  U_DCT2D_rtlc5n1480_13_CYMUXG2_787 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1480_13_CY0G,
      IB => U_DCT2D_rtlc5n1480_13_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1480_13_CYSELG,
      O => U_DCT2D_rtlc5n1480_13_CYMUXG2
    );
  U_DCT2D_rtlc5n1480_13_CY0G_788 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s(13),
      O => U_DCT2D_rtlc5n1480_13_CY0G
    );
  U_DCT2D_rtlc5n1480_13_CYSELG_789 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z81,
      O => U_DCT2D_rtlc5n1480_13_CYSELG
    );
  U_DCT2D_nx65206z79_rt_790 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z79,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z79_rt
    );
  U_DCT2D_rtlc5n1480_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480_15_XORF,
      O => U_DCT2D_rtlc5n1480(15)
    );
  U_DCT2D_rtlc5n1480_15_XORF_791 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1480_15_CYINIT,
      I1 => U_DCT2D_nx65206z79_rt,
      O => U_DCT2D_rtlc5n1480_15_XORF
    );
  U_DCT2D_rtlc5n1480_15_CYINIT_792 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_331_add_54_ix65206z63439_O,
      O => U_DCT2D_rtlc5n1480_15_CYINIT
    );
  U_DCT1D_databuf_reg_7_0_DXMUX_793 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_0_XORF,
      O => U_DCT1D_databuf_reg_7_0_DXMUX
    );
  U_DCT1D_databuf_reg_7_0_XORF_794 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_0_CYINIT,
      I1 => U_DCT1D_nx34147z1,
      O => U_DCT1D_databuf_reg_7_0_XORF
    );
  U_DCT1D_databuf_reg_7_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_0_CY0F,
      IB => U_DCT1D_databuf_reg_7_0_CYINIT,
      SEL => U_DCT1D_databuf_reg_7_0_CYSELF,
      O => U_DCT1D_rtlc5_86_sub_7_ix35144z63342_O
    );
  U_DCT1D_databuf_reg_7_0_CYINIT_795 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GLOBAL_LOGIC1_11,
      O => U_DCT1D_databuf_reg_7_0_CYINIT
    );
  U_DCT1D_databuf_reg_7_0_CY0F_796 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(0),
      O => U_DCT1D_databuf_reg_7_0_CY0F
    );
  U_DCT1D_databuf_reg_7_0_CYSELF_797 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx34147z1,
      O => U_DCT1D_databuf_reg_7_0_CYSELF
    );
  U_DCT1D_databuf_reg_7_0_DYMUX_798 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_0_XORG,
      O => U_DCT1D_databuf_reg_7_0_DYMUX
    );
  U_DCT1D_databuf_reg_7_0_XORG_799 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_86_sub_7_ix35144z63342_O,
      I1 => U_DCT1D_nx35144z1,
      O => U_DCT1D_databuf_reg_7_0_XORG
    );
  U_DCT1D_databuf_reg_7_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_0_CYMUXG,
      O => U_DCT1D_rtlc5_86_sub_7_ix36141z63342_O
    );
  U_DCT1D_databuf_reg_7_0_CYMUXG_800 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_0_CY0G,
      IB => U_DCT1D_rtlc5_86_sub_7_ix35144z63342_O,
      SEL => U_DCT1D_databuf_reg_7_0_CYSELG,
      O => U_DCT1D_databuf_reg_7_0_CYMUXG
    );
  U_DCT1D_databuf_reg_7_0_CY0G_801 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(1),
      O => U_DCT1D_databuf_reg_7_0_CY0G
    );
  U_DCT1D_databuf_reg_7_0_CYSELG_802 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx35144z1,
      O => U_DCT1D_databuf_reg_7_0_CYSELG
    );
  U_DCT1D_databuf_reg_7_0_SRINV_803 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_7_0_SRINV
    );
  U_DCT1D_databuf_reg_7_0_CLKINV_804 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_7_0_CLKINV
    );
  U_DCT1D_databuf_reg_7_0_CEINV_805 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_7_0_CEINV
    );
  U_DCT1D_databuf_reg_7_2_DXMUX_806 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_2_XORF,
      O => U_DCT1D_databuf_reg_7_2_DXMUX
    );
  U_DCT1D_databuf_reg_7_2_XORF_807 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_2_CYINIT,
      I1 => U_DCT1D_nx36141z1,
      O => U_DCT1D_databuf_reg_7_2_XORF
    );
  U_DCT1D_databuf_reg_7_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_2_CY0F,
      IB => U_DCT1D_databuf_reg_7_2_CYINIT,
      SEL => U_DCT1D_databuf_reg_7_2_CYSELF,
      O => U_DCT1D_rtlc5_86_sub_7_ix37138z63342_O
    );
  U_DCT1D_databuf_reg_7_2_CYMUXF2_808 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_2_CY0F,
      IB => U_DCT1D_databuf_reg_7_2_CY0F,
      SEL => U_DCT1D_databuf_reg_7_2_CYSELF,
      O => U_DCT1D_databuf_reg_7_2_CYMUXF2
    );
  U_DCT1D_databuf_reg_7_2_CYINIT_809 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_86_sub_7_ix36141z63342_O,
      O => U_DCT1D_databuf_reg_7_2_CYINIT
    );
  U_DCT1D_databuf_reg_7_2_CY0F_810 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(2),
      O => U_DCT1D_databuf_reg_7_2_CY0F
    );
  U_DCT1D_databuf_reg_7_2_CYSELF_811 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx36141z1,
      O => U_DCT1D_databuf_reg_7_2_CYSELF
    );
  U_DCT1D_databuf_reg_7_2_DYMUX_812 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_2_XORG,
      O => U_DCT1D_databuf_reg_7_2_DYMUX
    );
  U_DCT1D_databuf_reg_7_2_XORG_813 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_86_sub_7_ix37138z63342_O,
      I1 => U_DCT1D_nx37138z1,
      O => U_DCT1D_databuf_reg_7_2_XORG
    );
  U_DCT1D_databuf_reg_7_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_2_CYMUXFAST,
      O => U_DCT1D_rtlc5_86_sub_7_ix38135z63342_O
    );
  U_DCT1D_databuf_reg_7_2_FASTCARRY_814 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_86_sub_7_ix36141z63342_O,
      O => U_DCT1D_databuf_reg_7_2_FASTCARRY
    );
  U_DCT1D_databuf_reg_7_2_CYAND_815 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_7_2_CYSELG,
      I1 => U_DCT1D_databuf_reg_7_2_CYSELF,
      O => U_DCT1D_databuf_reg_7_2_CYAND
    );
  U_DCT1D_databuf_reg_7_2_CYMUXFAST_816 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_2_CYMUXG2,
      IB => U_DCT1D_databuf_reg_7_2_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_7_2_CYAND,
      O => U_DCT1D_databuf_reg_7_2_CYMUXFAST
    );
  U_DCT1D_databuf_reg_7_2_CYMUXG2_817 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_2_CY0G,
      IB => U_DCT1D_databuf_reg_7_2_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_7_2_CYSELG,
      O => U_DCT1D_databuf_reg_7_2_CYMUXG2
    );
  U_DCT1D_databuf_reg_7_2_CY0G_818 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(3),
      O => U_DCT1D_databuf_reg_7_2_CY0G
    );
  U_DCT1D_databuf_reg_7_2_CYSELG_819 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx37138z1,
      O => U_DCT1D_databuf_reg_7_2_CYSELG
    );
  U_DCT1D_databuf_reg_7_2_SRINV_820 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_7_2_SRINV
    );
  U_DCT1D_databuf_reg_7_2_CLKINV_821 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_7_2_CLKINV
    );
  U_DCT1D_databuf_reg_7_2_CEINV_822 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_7_2_CEINV
    );
  U_DCT1D_databuf_reg_7_4_DXMUX_823 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_4_XORF,
      O => U_DCT1D_databuf_reg_7_4_DXMUX
    );
  U_DCT1D_databuf_reg_7_4_XORF_824 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_4_CYINIT,
      I1 => U_DCT1D_nx38135z1,
      O => U_DCT1D_databuf_reg_7_4_XORF
    );
  U_DCT1D_databuf_reg_7_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_4_CY0F,
      IB => U_DCT1D_databuf_reg_7_4_CYINIT,
      SEL => U_DCT1D_databuf_reg_7_4_CYSELF,
      O => U_DCT1D_rtlc5_86_sub_7_ix39132z63342_O
    );
  U_DCT1D_databuf_reg_7_4_CYMUXF2_825 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_4_CY0F,
      IB => U_DCT1D_databuf_reg_7_4_CY0F,
      SEL => U_DCT1D_databuf_reg_7_4_CYSELF,
      O => U_DCT1D_databuf_reg_7_4_CYMUXF2
    );
  U_DCT1D_databuf_reg_7_4_CYINIT_826 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_86_sub_7_ix38135z63342_O,
      O => U_DCT1D_databuf_reg_7_4_CYINIT
    );
  U_DCT1D_databuf_reg_7_4_CY0F_827 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(4),
      O => U_DCT1D_databuf_reg_7_4_CY0F
    );
  U_DCT1D_databuf_reg_7_4_CYSELF_828 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx38135z1,
      O => U_DCT1D_databuf_reg_7_4_CYSELF
    );
  U_DCT1D_databuf_reg_7_4_DYMUX_829 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_4_XORG,
      O => U_DCT1D_databuf_reg_7_4_DYMUX
    );
  U_DCT1D_databuf_reg_7_4_XORG_830 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_86_sub_7_ix39132z63342_O,
      I1 => U_DCT1D_nx39132z1,
      O => U_DCT1D_databuf_reg_7_4_XORG
    );
  U_DCT1D_databuf_reg_7_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_4_CYMUXFAST,
      O => U_DCT1D_rtlc5_86_sub_7_ix40129z63342_O
    );
  U_DCT1D_databuf_reg_7_4_FASTCARRY_831 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_86_sub_7_ix38135z63342_O,
      O => U_DCT1D_databuf_reg_7_4_FASTCARRY
    );
  U_DCT1D_databuf_reg_7_4_CYAND_832 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_7_4_CYSELG,
      I1 => U_DCT1D_databuf_reg_7_4_CYSELF,
      O => U_DCT1D_databuf_reg_7_4_CYAND
    );
  U_DCT1D_databuf_reg_7_4_CYMUXFAST_833 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_4_CYMUXG2,
      IB => U_DCT1D_databuf_reg_7_4_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_7_4_CYAND,
      O => U_DCT1D_databuf_reg_7_4_CYMUXFAST
    );
  U_DCT1D_databuf_reg_7_4_CYMUXG2_834 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_4_CY0G,
      IB => U_DCT1D_databuf_reg_7_4_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_7_4_CYSELG,
      O => U_DCT1D_databuf_reg_7_4_CYMUXG2
    );
  U_DCT1D_databuf_reg_7_4_CY0G_835 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(5),
      O => U_DCT1D_databuf_reg_7_4_CY0G
    );
  U_DCT1D_databuf_reg_7_4_CYSELG_836 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx39132z1,
      O => U_DCT1D_databuf_reg_7_4_CYSELG
    );
  U_DCT1D_databuf_reg_7_4_SRINV_837 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_7_4_SRINV
    );
  U_DCT1D_databuf_reg_7_4_CLKINV_838 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_7_4_CLKINV
    );
  U_DCT1D_databuf_reg_7_4_CEINV_839 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_7_4_CEINV
    );
  U_DCT1D_databuf_reg_7_6_DXMUX_840 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_6_XORF,
      O => U_DCT1D_databuf_reg_7_6_DXMUX
    );
  U_DCT1D_databuf_reg_7_6_XORF_841 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_6_CYINIT,
      I1 => U_DCT1D_nx40129z1,
      O => U_DCT1D_databuf_reg_7_6_XORF
    );
  U_DCT1D_databuf_reg_7_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_6_CY0F,
      IB => U_DCT1D_databuf_reg_7_6_CYINIT,
      SEL => U_DCT1D_databuf_reg_7_6_CYSELF,
      O => U_DCT1D_rtlc5_86_sub_7_ix41126z63342_O
    );
  U_DCT1D_databuf_reg_7_6_CYMUXF2_842 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_6_CY0F,
      IB => U_DCT1D_databuf_reg_7_6_CY0F,
      SEL => U_DCT1D_databuf_reg_7_6_CYSELF,
      O => U_DCT1D_databuf_reg_7_6_CYMUXF2
    );
  U_DCT1D_databuf_reg_7_6_CYINIT_843 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_86_sub_7_ix40129z63342_O,
      O => U_DCT1D_databuf_reg_7_6_CYINIT
    );
  U_DCT1D_databuf_reg_7_6_CY0F_844 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(6),
      O => U_DCT1D_databuf_reg_7_6_CY0F
    );
  U_DCT1D_databuf_reg_7_6_CYSELF_845 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx40129z1,
      O => U_DCT1D_databuf_reg_7_6_CYSELF
    );
  U_DCT1D_databuf_reg_7_6_DYMUX_846 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_6_XORG,
      O => U_DCT1D_databuf_reg_7_6_DYMUX
    );
  U_DCT1D_databuf_reg_7_6_XORG_847 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_86_sub_7_ix41126z63342_O,
      I1 => U_DCT1D_nx41126z1,
      O => U_DCT1D_databuf_reg_7_6_XORG
    );
  U_DCT1D_databuf_reg_7_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_6_CYMUXFAST,
      O => U_DCT1D_rtlc5_86_sub_7_ix42123z63342_O
    );
  U_DCT1D_databuf_reg_7_6_FASTCARRY_848 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_86_sub_7_ix40129z63342_O,
      O => U_DCT1D_databuf_reg_7_6_FASTCARRY
    );
  U_DCT1D_databuf_reg_7_6_CYAND_849 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_7_6_CYSELG,
      I1 => U_DCT1D_databuf_reg_7_6_CYSELF,
      O => U_DCT1D_databuf_reg_7_6_CYAND
    );
  U_DCT1D_databuf_reg_7_6_CYMUXFAST_850 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_6_CYMUXG2,
      IB => U_DCT1D_databuf_reg_7_6_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_7_6_CYAND,
      O => U_DCT1D_databuf_reg_7_6_CYMUXFAST
    );
  U_DCT1D_databuf_reg_7_6_CYMUXG2_851 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_7_6_CY0G,
      IB => U_DCT1D_databuf_reg_7_6_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_7_6_CYSELG,
      O => U_DCT1D_databuf_reg_7_6_CYMUXG2
    );
  U_DCT1D_databuf_reg_7_6_CY0G_852 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(7),
      O => U_DCT1D_databuf_reg_7_6_CY0G
    );
  U_DCT1D_databuf_reg_7_6_CYSELG_853 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx41126z1,
      O => U_DCT1D_databuf_reg_7_6_CYSELG
    );
  U_DCT1D_databuf_reg_7_6_SRINV_854 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_7_6_SRINV
    );
  U_DCT1D_databuf_reg_7_6_CLKINV_855 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_7_6_CLKINV
    );
  U_DCT1D_databuf_reg_7_6_CEINV_856 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_7_6_CEINV
    );
  U_DCT1D_nx42123z1_rt_857 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx42123z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx42123z1_rt
    );
  U_DCT1D_databuf_reg_7_8_DXMUX_858 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_8_XORF,
      O => U_DCT1D_databuf_reg_7_8_DXMUX
    );
  U_DCT1D_databuf_reg_7_8_XORF_859 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_8_CYINIT,
      I1 => U_DCT1D_nx42123z1_rt,
      O => U_DCT1D_databuf_reg_7_8_XORF
    );
  U_DCT1D_databuf_reg_7_8_CYINIT_860 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_86_sub_7_ix42123z63342_O,
      O => U_DCT1D_databuf_reg_7_8_CYINIT
    );
  U_DCT1D_databuf_reg_7_8_CLKINV_861 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_7_8_CLKINV
    );
  U_DCT1D_databuf_reg_7_8_CEINV_862 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_7_8_CEINV
    );
  U_DCT2D_databuf_reg_0_0_DXMUX_863 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_0_XORF,
      O => U_DCT2D_databuf_reg_0_0_DXMUX
    );
  U_DCT2D_databuf_reg_0_0_XORF_864 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_0_CYINIT,
      I1 => U_DCT2D_nx60980z1,
      O => U_DCT2D_databuf_reg_0_0_XORF
    );
  U_DCT2D_databuf_reg_0_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_0_CY0F,
      IB => U_DCT2D_databuf_reg_0_0_CYINIT,
      SEL => U_DCT2D_databuf_reg_0_0_CYSELF,
      O => U_DCT2D_rtlc5_1578_add_45_ix59983z63342_O
    );
  U_DCT2D_databuf_reg_0_0_CYINIT_865 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_0_BXINVNOT,
      O => U_DCT2D_databuf_reg_0_0_CYINIT
    );
  U_DCT2D_databuf_reg_0_0_CY0F_866 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_0_Q,
      O => U_DCT2D_databuf_reg_0_0_CY0F
    );
  U_DCT2D_databuf_reg_0_0_CYSELF_867 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx60980z1,
      O => U_DCT2D_databuf_reg_0_0_CYSELF
    );
  U_DCT2D_databuf_reg_0_0_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_22,
      O => U_DCT2D_databuf_reg_0_0_BXINVNOT
    );
  U_DCT2D_databuf_reg_0_0_DYMUX_868 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_0_XORG,
      O => U_DCT2D_databuf_reg_0_0_DYMUX
    );
  U_DCT2D_databuf_reg_0_0_XORG_869 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1578_add_45_ix59983z63342_O,
      I1 => U_DCT2D_nx59983z1,
      O => U_DCT2D_databuf_reg_0_0_XORG
    );
  U_DCT2D_databuf_reg_0_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_0_CYMUXG,
      O => U_DCT2D_rtlc5_1578_add_45_ix58986z63342_O
    );
  U_DCT2D_databuf_reg_0_0_CYMUXG_870 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_0_CY0G,
      IB => U_DCT2D_rtlc5_1578_add_45_ix59983z63342_O,
      SEL => U_DCT2D_databuf_reg_0_0_CYSELG,
      O => U_DCT2D_databuf_reg_0_0_CYMUXG
    );
  U_DCT2D_databuf_reg_0_0_CY0G_871 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_1_Q,
      O => U_DCT2D_databuf_reg_0_0_CY0G
    );
  U_DCT2D_databuf_reg_0_0_CYSELG_872 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx59983z1,
      O => U_DCT2D_databuf_reg_0_0_CYSELG
    );
  U_DCT2D_databuf_reg_0_0_SRINV_873 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_0_0_SRINV
    );
  U_DCT2D_databuf_reg_0_0_CLKINV_874 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_0_0_CLKINV
    );
  U_DCT2D_databuf_reg_0_0_CEINV_875 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_0_0_CEINV
    );
  U_DCT2D_databuf_reg_0_2_DXMUX_876 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_2_XORF,
      O => U_DCT2D_databuf_reg_0_2_DXMUX
    );
  U_DCT2D_databuf_reg_0_2_XORF_877 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_2_CYINIT,
      I1 => U_DCT2D_nx58986z1,
      O => U_DCT2D_databuf_reg_0_2_XORF
    );
  U_DCT2D_databuf_reg_0_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_2_CY0F,
      IB => U_DCT2D_databuf_reg_0_2_CYINIT,
      SEL => U_DCT2D_databuf_reg_0_2_CYSELF,
      O => U_DCT2D_rtlc5_1578_add_45_ix57989z63342_O
    );
  U_DCT2D_databuf_reg_0_2_CYMUXF2_878 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_2_CY0F,
      IB => U_DCT2D_databuf_reg_0_2_CY0F,
      SEL => U_DCT2D_databuf_reg_0_2_CYSELF,
      O => U_DCT2D_databuf_reg_0_2_CYMUXF2
    );
  U_DCT2D_databuf_reg_0_2_CYINIT_879 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1578_add_45_ix58986z63342_O,
      O => U_DCT2D_databuf_reg_0_2_CYINIT
    );
  U_DCT2D_databuf_reg_0_2_CY0F_880 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_2_Q,
      O => U_DCT2D_databuf_reg_0_2_CY0F
    );
  U_DCT2D_databuf_reg_0_2_CYSELF_881 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx58986z1,
      O => U_DCT2D_databuf_reg_0_2_CYSELF
    );
  U_DCT2D_databuf_reg_0_2_DYMUX_882 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_2_XORG,
      O => U_DCT2D_databuf_reg_0_2_DYMUX
    );
  U_DCT2D_databuf_reg_0_2_XORG_883 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1578_add_45_ix57989z63342_O,
      I1 => U_DCT2D_nx57989z1,
      O => U_DCT2D_databuf_reg_0_2_XORG
    );
  U_DCT2D_databuf_reg_0_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_2_CYMUXFAST,
      O => U_DCT2D_rtlc5_1578_add_45_ix56992z63342_O
    );
  U_DCT2D_databuf_reg_0_2_FASTCARRY_884 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1578_add_45_ix58986z63342_O,
      O => U_DCT2D_databuf_reg_0_2_FASTCARRY
    );
  U_DCT2D_databuf_reg_0_2_CYAND_885 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_0_2_CYSELG,
      I1 => U_DCT2D_databuf_reg_0_2_CYSELF,
      O => U_DCT2D_databuf_reg_0_2_CYAND
    );
  U_DCT2D_databuf_reg_0_2_CYMUXFAST_886 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_2_CYMUXG2,
      IB => U_DCT2D_databuf_reg_0_2_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_0_2_CYAND,
      O => U_DCT2D_databuf_reg_0_2_CYMUXFAST
    );
  U_DCT2D_databuf_reg_0_2_CYMUXG2_887 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_2_CY0G,
      IB => U_DCT2D_databuf_reg_0_2_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_0_2_CYSELG,
      O => U_DCT2D_databuf_reg_0_2_CYMUXG2
    );
  U_DCT2D_databuf_reg_0_2_CY0G_888 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_3_Q,
      O => U_DCT2D_databuf_reg_0_2_CY0G
    );
  U_DCT2D_databuf_reg_0_2_CYSELG_889 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx57989z1,
      O => U_DCT2D_databuf_reg_0_2_CYSELG
    );
  U_DCT2D_databuf_reg_0_2_SRINV_890 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_0_2_SRINV
    );
  U_DCT2D_databuf_reg_0_2_CLKINV_891 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_0_2_CLKINV
    );
  U_DCT2D_databuf_reg_0_2_CEINV_892 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_0_2_CEINV
    );
  U_DCT2D_databuf_reg_0_4_DXMUX_893 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_4_XORF,
      O => U_DCT2D_databuf_reg_0_4_DXMUX
    );
  U_DCT2D_databuf_reg_0_4_XORF_894 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_4_CYINIT,
      I1 => U_DCT2D_nx56992z1,
      O => U_DCT2D_databuf_reg_0_4_XORF
    );
  U_DCT2D_databuf_reg_0_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_4_CY0F,
      IB => U_DCT2D_databuf_reg_0_4_CYINIT,
      SEL => U_DCT2D_databuf_reg_0_4_CYSELF,
      O => U_DCT2D_rtlc5_1578_add_45_ix55995z63342_O
    );
  U_DCT2D_databuf_reg_0_4_CYMUXF2_895 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_4_CY0F,
      IB => U_DCT2D_databuf_reg_0_4_CY0F,
      SEL => U_DCT2D_databuf_reg_0_4_CYSELF,
      O => U_DCT2D_databuf_reg_0_4_CYMUXF2
    );
  U_DCT2D_databuf_reg_0_4_CYINIT_896 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1578_add_45_ix56992z63342_O,
      O => U_DCT2D_databuf_reg_0_4_CYINIT
    );
  U_DCT2D_databuf_reg_0_4_CY0F_897 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_4_Q,
      O => U_DCT2D_databuf_reg_0_4_CY0F
    );
  U_DCT2D_databuf_reg_0_4_CYSELF_898 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx56992z1,
      O => U_DCT2D_databuf_reg_0_4_CYSELF
    );
  U_DCT2D_databuf_reg_0_4_DYMUX_899 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_4_XORG,
      O => U_DCT2D_databuf_reg_0_4_DYMUX
    );
  U_DCT2D_databuf_reg_0_4_XORG_900 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1578_add_45_ix55995z63342_O,
      I1 => U_DCT2D_nx55995z1,
      O => U_DCT2D_databuf_reg_0_4_XORG
    );
  U_DCT2D_databuf_reg_0_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_4_CYMUXFAST,
      O => U_DCT2D_rtlc5_1578_add_45_ix54998z63342_O
    );
  U_DCT2D_databuf_reg_0_4_FASTCARRY_901 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1578_add_45_ix56992z63342_O,
      O => U_DCT2D_databuf_reg_0_4_FASTCARRY
    );
  U_DCT2D_databuf_reg_0_4_CYAND_902 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_0_4_CYSELG,
      I1 => U_DCT2D_databuf_reg_0_4_CYSELF,
      O => U_DCT2D_databuf_reg_0_4_CYAND
    );
  U_DCT2D_databuf_reg_0_4_CYMUXFAST_903 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_4_CYMUXG2,
      IB => U_DCT2D_databuf_reg_0_4_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_0_4_CYAND,
      O => U_DCT2D_databuf_reg_0_4_CYMUXFAST
    );
  U_DCT2D_databuf_reg_0_4_CYMUXG2_904 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_4_CY0G,
      IB => U_DCT2D_databuf_reg_0_4_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_0_4_CYSELG,
      O => U_DCT2D_databuf_reg_0_4_CYMUXG2
    );
  U_DCT2D_databuf_reg_0_4_CY0G_905 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_5_Q,
      O => U_DCT2D_databuf_reg_0_4_CY0G
    );
  U_DCT2D_databuf_reg_0_4_CYSELG_906 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx55995z1,
      O => U_DCT2D_databuf_reg_0_4_CYSELG
    );
  U_DCT2D_databuf_reg_0_4_SRINV_907 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_0_4_SRINV
    );
  U_DCT2D_databuf_reg_0_4_CLKINV_908 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_0_4_CLKINV
    );
  U_DCT2D_databuf_reg_0_4_CEINV_909 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_0_4_CEINV
    );
  U_DCT2D_databuf_reg_0_6_DXMUX_910 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_6_XORF,
      O => U_DCT2D_databuf_reg_0_6_DXMUX
    );
  U_DCT2D_databuf_reg_0_6_XORF_911 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_6_CYINIT,
      I1 => U_DCT2D_nx54998z1,
      O => U_DCT2D_databuf_reg_0_6_XORF
    );
  U_DCT2D_databuf_reg_0_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_6_CY0F,
      IB => U_DCT2D_databuf_reg_0_6_CYINIT,
      SEL => U_DCT2D_databuf_reg_0_6_CYSELF,
      O => U_DCT2D_rtlc5_1578_add_45_ix54001z63342_O
    );
  U_DCT2D_databuf_reg_0_6_CYMUXF2_912 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_6_CY0F,
      IB => U_DCT2D_databuf_reg_0_6_CY0F,
      SEL => U_DCT2D_databuf_reg_0_6_CYSELF,
      O => U_DCT2D_databuf_reg_0_6_CYMUXF2
    );
  U_DCT2D_databuf_reg_0_6_CYINIT_913 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1578_add_45_ix54998z63342_O,
      O => U_DCT2D_databuf_reg_0_6_CYINIT
    );
  U_DCT2D_databuf_reg_0_6_CY0F_914 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_6_Q,
      O => U_DCT2D_databuf_reg_0_6_CY0F
    );
  U_DCT2D_databuf_reg_0_6_CYSELF_915 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx54998z1,
      O => U_DCT2D_databuf_reg_0_6_CYSELF
    );
  U_DCT2D_databuf_reg_0_6_DYMUX_916 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_6_XORG,
      O => U_DCT2D_databuf_reg_0_6_DYMUX
    );
  U_DCT2D_databuf_reg_0_6_XORG_917 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1578_add_45_ix54001z63342_O,
      I1 => U_DCT2D_nx54001z1,
      O => U_DCT2D_databuf_reg_0_6_XORG
    );
  U_DCT2D_databuf_reg_0_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_6_CYMUXFAST,
      O => U_DCT2D_rtlc5_1578_add_45_ix53004z63342_O
    );
  U_DCT2D_databuf_reg_0_6_FASTCARRY_918 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1578_add_45_ix54998z63342_O,
      O => U_DCT2D_databuf_reg_0_6_FASTCARRY
    );
  U_DCT2D_databuf_reg_0_6_CYAND_919 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_0_6_CYSELG,
      I1 => U_DCT2D_databuf_reg_0_6_CYSELF,
      O => U_DCT2D_databuf_reg_0_6_CYAND
    );
  U_DCT2D_databuf_reg_0_6_CYMUXFAST_920 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_6_CYMUXG2,
      IB => U_DCT2D_databuf_reg_0_6_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_0_6_CYAND,
      O => U_DCT2D_databuf_reg_0_6_CYMUXFAST
    );
  U_DCT2D_databuf_reg_0_6_CYMUXG2_921 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_6_CY0G,
      IB => U_DCT2D_databuf_reg_0_6_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_0_6_CYSELG,
      O => U_DCT2D_databuf_reg_0_6_CYMUXG2
    );
  U_DCT2D_databuf_reg_0_6_CY0G_922 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_7_Q,
      O => U_DCT2D_databuf_reg_0_6_CY0G
    );
  U_DCT2D_databuf_reg_0_6_CYSELG_923 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx54001z1,
      O => U_DCT2D_databuf_reg_0_6_CYSELG
    );
  U_DCT2D_databuf_reg_0_6_SRINV_924 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_0_6_SRINV
    );
  U_DCT2D_databuf_reg_0_6_CLKINV_925 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_0_6_CLKINV
    );
  U_DCT2D_databuf_reg_0_6_CEINV_926 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_0_6_CEINV
    );
  U_DCT2D_databuf_reg_0_8_DXMUX_927 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_8_XORF,
      O => U_DCT2D_databuf_reg_0_8_DXMUX
    );
  U_DCT2D_databuf_reg_0_8_XORF_928 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_8_CYINIT,
      I1 => U_DCT2D_nx53004z1,
      O => U_DCT2D_databuf_reg_0_8_XORF
    );
  U_DCT2D_databuf_reg_0_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_8_CY0F,
      IB => U_DCT2D_databuf_reg_0_8_CYINIT,
      SEL => U_DCT2D_databuf_reg_0_8_CYSELF,
      O => U_DCT2D_rtlc5_1578_add_45_ix52007z63342_O
    );
  U_DCT2D_databuf_reg_0_8_CYMUXF2_929 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_8_CY0F,
      IB => U_DCT2D_databuf_reg_0_8_CY0F,
      SEL => U_DCT2D_databuf_reg_0_8_CYSELF,
      O => U_DCT2D_databuf_reg_0_8_CYMUXF2
    );
  U_DCT2D_databuf_reg_0_8_CYINIT_930 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1578_add_45_ix53004z63342_O,
      O => U_DCT2D_databuf_reg_0_8_CYINIT
    );
  U_DCT2D_databuf_reg_0_8_CY0F_931 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_8_Q,
      O => U_DCT2D_databuf_reg_0_8_CY0F
    );
  U_DCT2D_databuf_reg_0_8_CYSELF_932 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx53004z1,
      O => U_DCT2D_databuf_reg_0_8_CYSELF
    );
  U_DCT2D_databuf_reg_0_8_DYMUX_933 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_8_XORG,
      O => U_DCT2D_databuf_reg_0_8_DYMUX
    );
  U_DCT2D_databuf_reg_0_8_XORG_934 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1578_add_45_ix52007z63342_O,
      I1 => U_DCT2D_nx52007z1,
      O => U_DCT2D_databuf_reg_0_8_XORG
    );
  U_DCT2D_databuf_reg_0_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_8_CYMUXFAST,
      O => U_DCT2D_rtlc5_1578_add_45_ix38337z63342_O
    );
  U_DCT2D_databuf_reg_0_8_FASTCARRY_935 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1578_add_45_ix53004z63342_O,
      O => U_DCT2D_databuf_reg_0_8_FASTCARRY
    );
  U_DCT2D_databuf_reg_0_8_CYAND_936 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_0_8_CYSELG,
      I1 => U_DCT2D_databuf_reg_0_8_CYSELF,
      O => U_DCT2D_databuf_reg_0_8_CYAND
    );
  U_DCT2D_databuf_reg_0_8_CYMUXFAST_937 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_8_CYMUXG2,
      IB => U_DCT2D_databuf_reg_0_8_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_0_8_CYAND,
      O => U_DCT2D_databuf_reg_0_8_CYMUXFAST
    );
  U_DCT2D_databuf_reg_0_8_CYMUXG2_938 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_0_8_CY0G,
      IB => U_DCT2D_databuf_reg_0_8_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_0_8_CYSELG,
      O => U_DCT2D_databuf_reg_0_8_CYMUXG2
    );
  U_DCT2D_databuf_reg_0_8_CY0G_939 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_10_Q,
      O => U_DCT2D_databuf_reg_0_8_CY0G
    );
  U_DCT2D_databuf_reg_0_8_CYSELG_940 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx52007z1,
      O => U_DCT2D_databuf_reg_0_8_CYSELG
    );
  U_DCT2D_databuf_reg_0_8_SRINV_941 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_0_8_SRINV
    );
  U_DCT2D_databuf_reg_0_8_CLKINV_942 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_0_8_CLKINV
    );
  U_DCT2D_databuf_reg_0_8_CEINV_943 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_0_8_CEINV
    );
  U_DCT2D_databuf_reg_0_10_DXMUX_944 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_10_XORF,
      O => U_DCT2D_databuf_reg_0_10_DXMUX
    );
  U_DCT2D_databuf_reg_0_10_XORF_945 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_10_CYINIT,
      I1 => U_DCT2D_nx38337z1_rt,
      O => U_DCT2D_databuf_reg_0_10_XORF
    );
  U_DCT2D_databuf_reg_0_10_CYINIT_946 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1578_add_45_ix38337z63342_O,
      O => U_DCT2D_databuf_reg_0_10_CYINIT
    );
  U_DCT2D_databuf_reg_0_10_CLKINV_947 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_0_10_CLKINV
    );
  U_DCT2D_databuf_reg_0_10_CEINV_948 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_0_10_CEINV
    );
  U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CY0F,
      IB => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYINIT,
      SEL => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYSELF,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63612_O
    );
  U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYINIT_949 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_BXINVNOT,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYINIT
    );
  U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CY0F_950 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(2),
      O => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CY0F
    );
  U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYSELF_951 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z209,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYSELF
    );
  U_DCT2D_rtlc_336_add_56_ix65206z63608_O_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_32,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_BXINVNOT
    );
  U_DCT2D_rtlc_336_add_56_ix65206z63608_O_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYMUXG,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63608_O
    );
  U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYMUXG_952 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CY0G,
      IB => U_DCT2D_rtlc_336_add_56_ix65206z63612_O,
      SEL => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYSELG,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYMUXG
    );
  U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CY0G_953 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(3),
      O => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CY0G
    );
  U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYSELG_954 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z207,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63608_O_CYSELG
    );
  U_DCT2D_rtlc5n1485_4_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_4_XORF,
      O => U_DCT2D_rtlc5n1485(4)
    );
  U_DCT2D_rtlc5n1485_4_XORF_955 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1485_4_CYINIT,
      I1 => U_DCT2D_nx65206z204,
      O => U_DCT2D_rtlc5n1485_4_XORF
    );
  U_DCT2D_rtlc5n1485_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_4_CY0F,
      IB => U_DCT2D_rtlc5n1485_4_CYINIT,
      SEL => U_DCT2D_rtlc5n1485_4_CYSELF,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63603_O
    );
  U_DCT2D_rtlc5n1485_4_CYMUXF2_956 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_4_CY0F,
      IB => U_DCT2D_rtlc5n1485_4_CY0F,
      SEL => U_DCT2D_rtlc5n1485_4_CYSELF,
      O => U_DCT2D_rtlc5n1485_4_CYMUXF2
    );
  U_DCT2D_rtlc5n1485_4_CYINIT_957 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63608_O,
      O => U_DCT2D_rtlc5n1485_4_CYINIT
    );
  U_DCT2D_rtlc5n1485_4_CY0F_958 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(4),
      O => U_DCT2D_rtlc5n1485_4_CY0F
    );
  U_DCT2D_rtlc5n1485_4_CYSELF_959 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z204,
      O => U_DCT2D_rtlc5n1485_4_CYSELF
    );
  U_DCT2D_rtlc5n1485_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_4_XORG,
      O => U_DCT2D_rtlc5n1485(5)
    );
  U_DCT2D_rtlc5n1485_4_XORG_960 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_336_add_56_ix65206z63603_O,
      I1 => U_DCT2D_nx65206z201,
      O => U_DCT2D_rtlc5n1485_4_XORG
    );
  U_DCT2D_rtlc5n1485_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_4_CYMUXFAST,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63597_O
    );
  U_DCT2D_rtlc5n1485_4_FASTCARRY_961 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63608_O,
      O => U_DCT2D_rtlc5n1485_4_FASTCARRY
    );
  U_DCT2D_rtlc5n1485_4_CYAND_962 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1485_4_CYSELG,
      I1 => U_DCT2D_rtlc5n1485_4_CYSELF,
      O => U_DCT2D_rtlc5n1485_4_CYAND
    );
  U_DCT2D_rtlc5n1485_4_CYMUXFAST_963 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_4_CYMUXG2,
      IB => U_DCT2D_rtlc5n1485_4_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1485_4_CYAND,
      O => U_DCT2D_rtlc5n1485_4_CYMUXFAST
    );
  U_DCT2D_rtlc5n1485_4_CYMUXG2_964 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_4_CY0G,
      IB => U_DCT2D_rtlc5n1485_4_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1485_4_CYSELG,
      O => U_DCT2D_rtlc5n1485_4_CYMUXG2
    );
  U_DCT2D_rtlc5n1485_4_CY0G_965 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(5),
      O => U_DCT2D_rtlc5n1485_4_CY0G
    );
  U_DCT2D_rtlc5n1485_4_CYSELG_966 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z201,
      O => U_DCT2D_rtlc5n1485_4_CYSELG
    );
  U_DCT2D_rtlc5n1485_6_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_6_XORF,
      O => U_DCT2D_rtlc5n1485(6)
    );
  U_DCT2D_rtlc5n1485_6_XORF_967 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1485_6_CYINIT,
      I1 => U_DCT2D_nx65206z198,
      O => U_DCT2D_rtlc5n1485_6_XORF
    );
  U_DCT2D_rtlc5n1485_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_6_CY0F,
      IB => U_DCT2D_rtlc5n1485_6_CYINIT,
      SEL => U_DCT2D_rtlc5n1485_6_CYSELF,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63592_O
    );
  U_DCT2D_rtlc5n1485_6_CYMUXF2_968 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_6_CY0F,
      IB => U_DCT2D_rtlc5n1485_6_CY0F,
      SEL => U_DCT2D_rtlc5n1485_6_CYSELF,
      O => U_DCT2D_rtlc5n1485_6_CYMUXF2
    );
  U_DCT2D_rtlc5n1485_6_CYINIT_969 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63597_O,
      O => U_DCT2D_rtlc5n1485_6_CYINIT
    );
  U_DCT2D_rtlc5n1485_6_CY0F_970 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(6),
      O => U_DCT2D_rtlc5n1485_6_CY0F
    );
  U_DCT2D_rtlc5n1485_6_CYSELF_971 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z198,
      O => U_DCT2D_rtlc5n1485_6_CYSELF
    );
  U_DCT2D_rtlc5n1485_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_6_XORG,
      O => U_DCT2D_rtlc5n1485(7)
    );
  U_DCT2D_rtlc5n1485_6_XORG_972 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_336_add_56_ix65206z63592_O,
      I1 => U_DCT2D_nx65206z195,
      O => U_DCT2D_rtlc5n1485_6_XORG
    );
  U_DCT2D_rtlc5n1485_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_6_CYMUXFAST,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63587_O
    );
  U_DCT2D_rtlc5n1485_6_FASTCARRY_973 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63597_O,
      O => U_DCT2D_rtlc5n1485_6_FASTCARRY
    );
  U_DCT2D_rtlc5n1485_6_CYAND_974 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1485_6_CYSELG,
      I1 => U_DCT2D_rtlc5n1485_6_CYSELF,
      O => U_DCT2D_rtlc5n1485_6_CYAND
    );
  U_DCT2D_rtlc5n1485_6_CYMUXFAST_975 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_6_CYMUXG2,
      IB => U_DCT2D_rtlc5n1485_6_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1485_6_CYAND,
      O => U_DCT2D_rtlc5n1485_6_CYMUXFAST
    );
  U_DCT2D_rtlc5n1485_6_CYMUXG2_976 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_6_CY0G,
      IB => U_DCT2D_rtlc5n1485_6_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1485_6_CYSELG,
      O => U_DCT2D_rtlc5n1485_6_CYMUXG2
    );
  U_DCT2D_rtlc5n1485_6_CY0G_977 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(7),
      O => U_DCT2D_rtlc5n1485_6_CY0G
    );
  U_DCT2D_rtlc5n1485_6_CYSELG_978 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z195,
      O => U_DCT2D_rtlc5n1485_6_CYSELG
    );
  U_DCT2D_rtlc5n1485_8_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_8_XORF,
      O => U_DCT2D_rtlc5n1485(8)
    );
  U_DCT2D_rtlc5n1485_8_XORF_979 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1485_8_CYINIT,
      I1 => U_DCT2D_nx65206z192,
      O => U_DCT2D_rtlc5n1485_8_XORF
    );
  U_DCT2D_rtlc5n1485_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_8_CY0F,
      IB => U_DCT2D_rtlc5n1485_8_CYINIT,
      SEL => U_DCT2D_rtlc5n1485_8_CYSELF,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63582_O
    );
  U_DCT2D_rtlc5n1485_8_CYMUXF2_980 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_8_CY0F,
      IB => U_DCT2D_rtlc5n1485_8_CY0F,
      SEL => U_DCT2D_rtlc5n1485_8_CYSELF,
      O => U_DCT2D_rtlc5n1485_8_CYMUXF2
    );
  U_DCT2D_rtlc5n1485_8_CYINIT_981 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63587_O,
      O => U_DCT2D_rtlc5n1485_8_CYINIT
    );
  U_DCT2D_rtlc5n1485_8_CY0F_982 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(8),
      O => U_DCT2D_rtlc5n1485_8_CY0F
    );
  U_DCT2D_rtlc5n1485_8_CYSELF_983 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z192,
      O => U_DCT2D_rtlc5n1485_8_CYSELF
    );
  U_DCT2D_rtlc5n1485_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_8_XORG,
      O => U_DCT2D_rtlc5n1485(9)
    );
  U_DCT2D_rtlc5n1485_8_XORG_984 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_336_add_56_ix65206z63582_O,
      I1 => U_DCT2D_nx65206z189,
      O => U_DCT2D_rtlc5n1485_8_XORG
    );
  U_DCT2D_rtlc5n1485_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_8_CYMUXFAST,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63577_O
    );
  U_DCT2D_rtlc5n1485_8_FASTCARRY_985 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63587_O,
      O => U_DCT2D_rtlc5n1485_8_FASTCARRY
    );
  U_DCT2D_rtlc5n1485_8_CYAND_986 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1485_8_CYSELG,
      I1 => U_DCT2D_rtlc5n1485_8_CYSELF,
      O => U_DCT2D_rtlc5n1485_8_CYAND
    );
  U_DCT2D_rtlc5n1485_8_CYMUXFAST_987 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_8_CYMUXG2,
      IB => U_DCT2D_rtlc5n1485_8_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1485_8_CYAND,
      O => U_DCT2D_rtlc5n1485_8_CYMUXFAST
    );
  U_DCT2D_rtlc5n1485_8_CYMUXG2_988 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_8_CY0G,
      IB => U_DCT2D_rtlc5n1485_8_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1485_8_CYSELG,
      O => U_DCT2D_rtlc5n1485_8_CYMUXG2
    );
  U_DCT2D_rtlc5n1485_8_CY0G_989 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(9),
      O => U_DCT2D_rtlc5n1485_8_CY0G
    );
  U_DCT2D_rtlc5n1485_8_CYSELG_990 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z189,
      O => U_DCT2D_rtlc5n1485_8_CYSELG
    );
  U_DCT2D_rtlc5n1485_10_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_10_XORF,
      O => U_DCT2D_rtlc5n1485(10)
    );
  U_DCT2D_rtlc5n1485_10_XORF_991 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1485_10_CYINIT,
      I1 => U_DCT2D_nx65206z186,
      O => U_DCT2D_rtlc5n1485_10_XORF
    );
  U_DCT2D_rtlc5n1485_10_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_10_CY0F,
      IB => U_DCT2D_rtlc5n1485_10_CYINIT,
      SEL => U_DCT2D_rtlc5n1485_10_CYSELF,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63572_O
    );
  U_DCT2D_rtlc5n1485_10_CYMUXF2_992 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_10_CY0F,
      IB => U_DCT2D_rtlc5n1485_10_CY0F,
      SEL => U_DCT2D_rtlc5n1485_10_CYSELF,
      O => U_DCT2D_rtlc5n1485_10_CYMUXF2
    );
  U_DCT2D_rtlc5n1485_10_CYINIT_993 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63577_O,
      O => U_DCT2D_rtlc5n1485_10_CYINIT
    );
  U_DCT2D_rtlc5n1485_10_CY0F_994 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(10),
      O => U_DCT2D_rtlc5n1485_10_CY0F
    );
  U_DCT2D_rtlc5n1485_10_CYSELF_995 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z186,
      O => U_DCT2D_rtlc5n1485_10_CYSELF
    );
  U_DCT2D_rtlc5n1485_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_10_XORG,
      O => U_DCT2D_rtlc5n1485(11)
    );
  U_DCT2D_rtlc5n1485_10_XORG_996 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_336_add_56_ix65206z63572_O,
      I1 => U_DCT2D_nx65206z183,
      O => U_DCT2D_rtlc5n1485_10_XORG
    );
  U_DCT2D_rtlc5n1485_10_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_10_CYMUXFAST,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63567_O
    );
  U_DCT2D_rtlc5n1485_10_FASTCARRY_997 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63577_O,
      O => U_DCT2D_rtlc5n1485_10_FASTCARRY
    );
  U_DCT2D_rtlc5n1485_10_CYAND_998 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1485_10_CYSELG,
      I1 => U_DCT2D_rtlc5n1485_10_CYSELF,
      O => U_DCT2D_rtlc5n1485_10_CYAND
    );
  U_DCT2D_rtlc5n1485_10_CYMUXFAST_999 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_10_CYMUXG2,
      IB => U_DCT2D_rtlc5n1485_10_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1485_10_CYAND,
      O => U_DCT2D_rtlc5n1485_10_CYMUXFAST
    );
  U_DCT2D_rtlc5n1485_10_CYMUXG2_1000 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_10_CY0G,
      IB => U_DCT2D_rtlc5n1485_10_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1485_10_CYSELG,
      O => U_DCT2D_rtlc5n1485_10_CYMUXG2
    );
  U_DCT2D_rtlc5n1485_10_CY0G_1001 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(11),
      O => U_DCT2D_rtlc5n1485_10_CY0G
    );
  U_DCT2D_rtlc5n1485_10_CYSELG_1002 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z183,
      O => U_DCT2D_rtlc5n1485_10_CYSELG
    );
  U_DCT2D_rtlc5n1485_12_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_12_XORF,
      O => U_DCT2D_rtlc5n1485(12)
    );
  U_DCT2D_rtlc5n1485_12_XORF_1003 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1485_12_CYINIT,
      I1 => U_DCT2D_nx65206z180,
      O => U_DCT2D_rtlc5n1485_12_XORF
    );
  U_DCT2D_rtlc5n1485_12_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_12_CY0F,
      IB => U_DCT2D_rtlc5n1485_12_CYINIT,
      SEL => U_DCT2D_rtlc5n1485_12_CYSELF,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63561_O
    );
  U_DCT2D_rtlc5n1485_12_CYMUXF2_1004 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_12_CY0F,
      IB => U_DCT2D_rtlc5n1485_12_CY0F,
      SEL => U_DCT2D_rtlc5n1485_12_CYSELF,
      O => U_DCT2D_rtlc5n1485_12_CYMUXF2
    );
  U_DCT2D_rtlc5n1485_12_CYINIT_1005 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63567_O,
      O => U_DCT2D_rtlc5n1485_12_CYINIT
    );
  U_DCT2D_rtlc5n1485_12_CY0F_1006 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(12),
      O => U_DCT2D_rtlc5n1485_12_CY0F
    );
  U_DCT2D_rtlc5n1485_12_CYSELF_1007 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z180,
      O => U_DCT2D_rtlc5n1485_12_CYSELF
    );
  U_DCT2D_rtlc5n1485_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_12_XORG,
      O => U_DCT2D_rtlc5n1485(13)
    );
  U_DCT2D_rtlc5n1485_12_XORG_1008 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_336_add_56_ix65206z63561_O,
      I1 => U_DCT2D_nx65206z177,
      O => U_DCT2D_rtlc5n1485_12_XORG
    );
  U_DCT2D_rtlc5n1485_12_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_12_CYMUXFAST,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63556_O
    );
  U_DCT2D_rtlc5n1485_12_FASTCARRY_1009 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63567_O,
      O => U_DCT2D_rtlc5n1485_12_FASTCARRY
    );
  U_DCT2D_rtlc5n1485_12_CYAND_1010 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1485_12_CYSELG,
      I1 => U_DCT2D_rtlc5n1485_12_CYSELF,
      O => U_DCT2D_rtlc5n1485_12_CYAND
    );
  U_DCT2D_rtlc5n1485_12_CYMUXFAST_1011 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_12_CYMUXG2,
      IB => U_DCT2D_rtlc5n1485_12_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1485_12_CYAND,
      O => U_DCT2D_rtlc5n1485_12_CYMUXFAST
    );
  U_DCT2D_rtlc5n1485_12_CYMUXG2_1012 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_12_CY0G,
      IB => U_DCT2D_rtlc5n1485_12_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1485_12_CYSELG,
      O => U_DCT2D_rtlc5n1485_12_CYMUXG2
    );
  U_DCT2D_rtlc5n1485_12_CY0G_1013 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(13),
      O => U_DCT2D_rtlc5n1485_12_CY0G
    );
  U_DCT2D_rtlc5n1485_12_CYSELG_1014 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z177,
      O => U_DCT2D_rtlc5n1485_12_CYSELG
    );
  U_DCT2D_rtlc5n1485_14_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_14_XORF,
      O => U_DCT2D_rtlc5n1485(14)
    );
  U_DCT2D_rtlc5n1485_14_XORF_1015 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1485_14_CYINIT,
      I1 => U_DCT2D_nx65206z174,
      O => U_DCT2D_rtlc5n1485_14_XORF
    );
  U_DCT2D_rtlc5n1485_14_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_14_CY0F,
      IB => U_DCT2D_rtlc5n1485_14_CYINIT,
      SEL => U_DCT2D_rtlc5n1485_14_CYSELF,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63551_O
    );
  U_DCT2D_rtlc5n1485_14_CYMUXF2_1016 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_14_CY0F,
      IB => U_DCT2D_rtlc5n1485_14_CY0F,
      SEL => U_DCT2D_rtlc5n1485_14_CYSELF,
      O => U_DCT2D_rtlc5n1485_14_CYMUXF2
    );
  U_DCT2D_rtlc5n1485_14_CYINIT_1017 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63556_O,
      O => U_DCT2D_rtlc5n1485_14_CYINIT
    );
  U_DCT2D_rtlc5n1485_14_CY0F_1018 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(14),
      O => U_DCT2D_rtlc5n1485_14_CY0F
    );
  U_DCT2D_rtlc5n1485_14_CYSELF_1019 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z174,
      O => U_DCT2D_rtlc5n1485_14_CYSELF
    );
  U_DCT2D_rtlc5n1485_14_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_14_XORG,
      O => U_DCT2D_rtlc5n1485(15)
    );
  U_DCT2D_rtlc5n1485_14_XORG_1020 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_336_add_56_ix65206z63551_O,
      I1 => U_DCT2D_nx65206z171,
      O => U_DCT2D_rtlc5n1485_14_XORG
    );
  U_DCT2D_rtlc5n1485_14_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_14_CYMUXFAST,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63546_O
    );
  U_DCT2D_rtlc5n1485_14_FASTCARRY_1021 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63556_O,
      O => U_DCT2D_rtlc5n1485_14_FASTCARRY
    );
  U_DCT2D_rtlc5n1485_14_CYAND_1022 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1485_14_CYSELG,
      I1 => U_DCT2D_rtlc5n1485_14_CYSELF,
      O => U_DCT2D_rtlc5n1485_14_CYAND
    );
  U_DCT2D_rtlc5n1485_14_CYMUXFAST_1023 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_14_CYMUXG2,
      IB => U_DCT2D_rtlc5n1485_14_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1485_14_CYAND,
      O => U_DCT2D_rtlc5n1485_14_CYMUXFAST
    );
  U_DCT2D_rtlc5n1485_14_CYMUXG2_1024 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_14_CY0G,
      IB => U_DCT2D_rtlc5n1485_14_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1485_14_CYSELG,
      O => U_DCT2D_rtlc5n1485_14_CYMUXG2
    );
  U_DCT2D_rtlc5n1485_14_CY0G_1025 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(15),
      O => U_DCT2D_rtlc5n1485_14_CY0G
    );
  U_DCT2D_rtlc5n1485_14_CYSELG_1026 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z171,
      O => U_DCT2D_rtlc5n1485_14_CYSELG
    );
  U_DCT2D_rtlc5n1485_16_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_16_XORF,
      O => U_DCT2D_rtlc5n1485(16)
    );
  U_DCT2D_rtlc5n1485_16_XORF_1027 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1485_16_CYINIT,
      I1 => U_DCT2D_nx65206z168,
      O => U_DCT2D_rtlc5n1485_16_XORF
    );
  U_DCT2D_rtlc5n1485_16_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_16_CY0F,
      IB => U_DCT2D_rtlc5n1485_16_CYINIT,
      SEL => U_DCT2D_rtlc5n1485_16_CYSELF,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63542_O
    );
  U_DCT2D_rtlc5n1485_16_CYMUXF2_1028 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_16_CY0F,
      IB => U_DCT2D_rtlc5n1485_16_CY0F,
      SEL => U_DCT2D_rtlc5n1485_16_CYSELF,
      O => U_DCT2D_rtlc5n1485_16_CYMUXF2
    );
  U_DCT2D_rtlc5n1485_16_CYINIT_1029 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63546_O,
      O => U_DCT2D_rtlc5n1485_16_CYINIT
    );
  U_DCT2D_rtlc5n1485_16_CY0F_1030 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(15),
      O => U_DCT2D_rtlc5n1485_16_CY0F
    );
  U_DCT2D_rtlc5n1485_16_CYSELF_1031 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z168,
      O => U_DCT2D_rtlc5n1485_16_CYSELF
    );
  U_DCT2D_rtlc5n1485_16_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_16_XORG,
      O => U_DCT2D_rtlc5n1485(17)
    );
  U_DCT2D_rtlc5n1485_16_XORG_1032 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_336_add_56_ix65206z63542_O,
      I1 => U_DCT2D_nx65206z165,
      O => U_DCT2D_rtlc5n1485_16_XORG
    );
  U_DCT2D_rtlc5n1485_16_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_16_CYMUXFAST,
      O => U_DCT2D_rtlc_336_add_56_ix65206z63538_O
    );
  U_DCT2D_rtlc5n1485_16_FASTCARRY_1033 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63546_O,
      O => U_DCT2D_rtlc5n1485_16_FASTCARRY
    );
  U_DCT2D_rtlc5n1485_16_CYAND_1034 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1485_16_CYSELG,
      I1 => U_DCT2D_rtlc5n1485_16_CYSELF,
      O => U_DCT2D_rtlc5n1485_16_CYAND
    );
  U_DCT2D_rtlc5n1485_16_CYMUXFAST_1035 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_16_CYMUXG2,
      IB => U_DCT2D_rtlc5n1485_16_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1485_16_CYAND,
      O => U_DCT2D_rtlc5n1485_16_CYMUXFAST
    );
  U_DCT2D_rtlc5n1485_16_CYMUXG2_1036 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1485_16_CY0G,
      IB => U_DCT2D_rtlc5n1485_16_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1485_16_CYSELG,
      O => U_DCT2D_rtlc5n1485_16_CYMUXG2
    );
  U_DCT2D_rtlc5n1485_16_CY0G_1037 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1480(15),
      O => U_DCT2D_rtlc5n1485_16_CY0G
    );
  U_DCT2D_rtlc5n1485_16_CYSELG_1038 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z165,
      O => U_DCT2D_rtlc5n1485_16_CYSELG
    );
  U_DCT1D_reg_databuf_reg_2_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_2_2_DYMUX,
      CE => U_DCT1D_databuf_reg_2_2_CEINV,
      CLK => U_DCT1D_databuf_reg_2_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_2_2_FFY_RST,
      O => U_DCT1D_databuf_reg_2_Q(3)
    );
  U_DCT1D_databuf_reg_2_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_2_2_FFY_RST
    );
  U_DCT2D_nx65206z78_rt_1039 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z78,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z78_rt
    );
  U_DCT2D_rtlc5n1485_18_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1485_18_XORF,
      O => U_DCT2D_rtlc5n1485(18)
    );
  U_DCT2D_rtlc5n1485_18_XORF_1040 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1485_18_CYINIT,
      I1 => U_DCT2D_nx65206z78_rt,
      O => U_DCT2D_rtlc5n1485_18_XORF
    );
  U_DCT2D_rtlc5n1485_18_CYINIT_1041 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_336_add_56_ix65206z63538_O,
      O => U_DCT2D_rtlc5n1485_18_CYINIT
    );
  U_DCT2D_rtlc5n1483_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_7_XORF,
      O => U_DCT2D_rtlc5n1483(7)
    );
  U_DCT2D_rtlc5n1483_7_XORF_1042 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1483_7_CYINIT,
      I1 => U_DCT2D_nx65206z294,
      O => U_DCT2D_rtlc5n1483_7_XORF
    );
  U_DCT2D_rtlc5n1483_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_7_CY0F,
      IB => U_DCT2D_rtlc5n1483_7_CYINIT,
      SEL => U_DCT2D_rtlc5n1483_7_CYSELF,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63745_O
    );
  U_DCT2D_rtlc5n1483_7_CYINIT_1043 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_7_BXINVNOT,
      O => U_DCT2D_rtlc5n1483_7_CYINIT
    );
  U_DCT2D_rtlc5n1483_7_CY0F_1044 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(1),
      O => U_DCT2D_rtlc5n1483_7_CY0F
    );
  U_DCT2D_rtlc5n1483_7_CYSELF_1045 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z294,
      O => U_DCT2D_rtlc5n1483_7_CYSELF
    );
  U_DCT2D_rtlc5n1483_7_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_17,
      O => U_DCT2D_rtlc5n1483_7_BXINVNOT
    );
  U_DCT2D_rtlc5n1483_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_7_XORG,
      O => U_DCT2D_rtlc5n1483(8)
    );
  U_DCT2D_rtlc5n1483_7_XORG_1046 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_340_add_58_ix65206z63745_O,
      I1 => U_DCT2D_nx65206z291,
      O => U_DCT2D_rtlc5n1483_7_XORG
    );
  U_DCT2D_rtlc5n1483_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_7_CYMUXG,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63742_O
    );
  U_DCT2D_rtlc5n1483_7_CYMUXG_1047 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_7_CY0G,
      IB => U_DCT2D_rtlc_340_add_58_ix65206z63745_O,
      SEL => U_DCT2D_rtlc5n1483_7_CYSELG,
      O => U_DCT2D_rtlc5n1483_7_CYMUXG
    );
  U_DCT2D_rtlc5n1483_7_CY0G_1048 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(2),
      O => U_DCT2D_rtlc5n1483_7_CY0G
    );
  U_DCT2D_rtlc5n1483_7_CYSELG_1049 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z291,
      O => U_DCT2D_rtlc5n1483_7_CYSELG
    );
  U_DCT2D_ix65206z1716 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao6_s(4),
      ADR2 => VCC,
      ADR3 => romo2datao7_s(3),
      O => U_DCT2D_nx65206z285
    );
  U_DCT2D_rtlc5n1483_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_9_XORF,
      O => U_DCT2D_rtlc5n1483(9)
    );
  U_DCT2D_rtlc5n1483_9_XORF_1050 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1483_9_CYINIT,
      I1 => U_DCT2D_nx65206z288,
      O => U_DCT2D_rtlc5n1483_9_XORF
    );
  U_DCT2D_rtlc5n1483_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_9_CY0F,
      IB => U_DCT2D_rtlc5n1483_9_CYINIT,
      SEL => U_DCT2D_rtlc5n1483_9_CYSELF,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63738_O
    );
  U_DCT2D_rtlc5n1483_9_CYMUXF2_1051 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_9_CY0F,
      IB => U_DCT2D_rtlc5n1483_9_CY0F,
      SEL => U_DCT2D_rtlc5n1483_9_CYSELF,
      O => U_DCT2D_rtlc5n1483_9_CYMUXF2
    );
  U_DCT2D_rtlc5n1483_9_CYINIT_1052 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63742_O,
      O => U_DCT2D_rtlc5n1483_9_CYINIT
    );
  U_DCT2D_rtlc5n1483_9_CY0F_1053 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(3),
      O => U_DCT2D_rtlc5n1483_9_CY0F
    );
  U_DCT2D_rtlc5n1483_9_CYSELF_1054 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z288,
      O => U_DCT2D_rtlc5n1483_9_CYSELF
    );
  U_DCT2D_rtlc5n1483_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_9_XORG,
      O => U_DCT2D_rtlc5n1483(10)
    );
  U_DCT2D_rtlc5n1483_9_XORG_1055 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_340_add_58_ix65206z63738_O,
      I1 => U_DCT2D_nx65206z285,
      O => U_DCT2D_rtlc5n1483_9_XORG
    );
  U_DCT2D_rtlc5n1483_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_9_CYMUXFAST,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63735_O
    );
  U_DCT2D_rtlc5n1483_9_FASTCARRY_1056 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63742_O,
      O => U_DCT2D_rtlc5n1483_9_FASTCARRY
    );
  U_DCT2D_rtlc5n1483_9_CYAND_1057 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483_9_CYSELG,
      I1 => U_DCT2D_rtlc5n1483_9_CYSELF,
      O => U_DCT2D_rtlc5n1483_9_CYAND
    );
  U_DCT2D_rtlc5n1483_9_CYMUXFAST_1058 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_9_CYMUXG2,
      IB => U_DCT2D_rtlc5n1483_9_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1483_9_CYAND,
      O => U_DCT2D_rtlc5n1483_9_CYMUXFAST
    );
  U_DCT2D_rtlc5n1483_9_CYMUXG2_1059 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_9_CY0G,
      IB => U_DCT2D_rtlc5n1483_9_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1483_9_CYSELG,
      O => U_DCT2D_rtlc5n1483_9_CYMUXG2
    );
  U_DCT2D_rtlc5n1483_9_CY0G_1060 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(4),
      O => U_DCT2D_rtlc5n1483_9_CY0G
    );
  U_DCT2D_rtlc5n1483_9_CYSELG_1061 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z285,
      O => U_DCT2D_rtlc5n1483_9_CYSELG
    );
  U_DCT2D_rtlc5n1483_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_11_XORF,
      O => U_DCT2D_rtlc5n1483(11)
    );
  U_DCT2D_rtlc5n1483_11_XORF_1062 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1483_11_CYINIT,
      I1 => U_DCT2D_nx65206z282,
      O => U_DCT2D_rtlc5n1483_11_XORF
    );
  U_DCT2D_rtlc5n1483_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_11_CY0F,
      IB => U_DCT2D_rtlc5n1483_11_CYINIT,
      SEL => U_DCT2D_rtlc5n1483_11_CYSELF,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63731_O
    );
  U_DCT2D_rtlc5n1483_11_CYMUXF2_1063 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_11_CY0F,
      IB => U_DCT2D_rtlc5n1483_11_CY0F,
      SEL => U_DCT2D_rtlc5n1483_11_CYSELF,
      O => U_DCT2D_rtlc5n1483_11_CYMUXF2
    );
  U_DCT2D_rtlc5n1483_11_CYINIT_1064 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63735_O,
      O => U_DCT2D_rtlc5n1483_11_CYINIT
    );
  U_DCT2D_rtlc5n1483_11_CY0F_1065 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(5),
      O => U_DCT2D_rtlc5n1483_11_CY0F
    );
  U_DCT2D_rtlc5n1483_11_CYSELF_1066 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z282,
      O => U_DCT2D_rtlc5n1483_11_CYSELF
    );
  U_DCT2D_rtlc5n1483_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_11_XORG,
      O => U_DCT2D_rtlc5n1483(12)
    );
  U_DCT2D_rtlc5n1483_11_XORG_1067 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_340_add_58_ix65206z63731_O,
      I1 => U_DCT2D_nx65206z279,
      O => U_DCT2D_rtlc5n1483_11_XORG
    );
  U_DCT2D_rtlc5n1483_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_11_CYMUXFAST,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63728_O
    );
  U_DCT2D_rtlc5n1483_11_FASTCARRY_1068 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63735_O,
      O => U_DCT2D_rtlc5n1483_11_FASTCARRY
    );
  U_DCT2D_rtlc5n1483_11_CYAND_1069 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483_11_CYSELG,
      I1 => U_DCT2D_rtlc5n1483_11_CYSELF,
      O => U_DCT2D_rtlc5n1483_11_CYAND
    );
  U_DCT2D_rtlc5n1483_11_CYMUXFAST_1070 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_11_CYMUXG2,
      IB => U_DCT2D_rtlc5n1483_11_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1483_11_CYAND,
      O => U_DCT2D_rtlc5n1483_11_CYMUXFAST
    );
  U_DCT2D_rtlc5n1483_11_CYMUXG2_1071 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_11_CY0G,
      IB => U_DCT2D_rtlc5n1483_11_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1483_11_CYSELG,
      O => U_DCT2D_rtlc5n1483_11_CYMUXG2
    );
  U_DCT2D_rtlc5n1483_11_CY0G_1072 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(6),
      O => U_DCT2D_rtlc5n1483_11_CY0G
    );
  U_DCT2D_rtlc5n1483_11_CYSELG_1073 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z279,
      O => U_DCT2D_rtlc5n1483_11_CYSELG
    );
  U_DCT2D_rtlc5n1483_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_13_XORF,
      O => U_DCT2D_rtlc5n1483(13)
    );
  U_DCT2D_rtlc5n1483_13_XORF_1074 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1483_13_CYINIT,
      I1 => U_DCT2D_nx65206z276,
      O => U_DCT2D_rtlc5n1483_13_XORF
    );
  U_DCT2D_rtlc5n1483_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_13_CY0F,
      IB => U_DCT2D_rtlc5n1483_13_CYINIT,
      SEL => U_DCT2D_rtlc5n1483_13_CYSELF,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63724_O
    );
  U_DCT2D_rtlc5n1483_13_CYMUXF2_1075 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_13_CY0F,
      IB => U_DCT2D_rtlc5n1483_13_CY0F,
      SEL => U_DCT2D_rtlc5n1483_13_CYSELF,
      O => U_DCT2D_rtlc5n1483_13_CYMUXF2
    );
  U_DCT2D_rtlc5n1483_13_CYINIT_1076 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63728_O,
      O => U_DCT2D_rtlc5n1483_13_CYINIT
    );
  U_DCT2D_rtlc5n1483_13_CY0F_1077 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(7),
      O => U_DCT2D_rtlc5n1483_13_CY0F
    );
  U_DCT2D_rtlc5n1483_13_CYSELF_1078 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z276,
      O => U_DCT2D_rtlc5n1483_13_CYSELF
    );
  U_DCT2D_rtlc5n1483_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_13_XORG,
      O => U_DCT2D_rtlc5n1483(14)
    );
  U_DCT2D_rtlc5n1483_13_XORG_1079 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_340_add_58_ix65206z63724_O,
      I1 => U_DCT2D_nx65206z273,
      O => U_DCT2D_rtlc5n1483_13_XORG
    );
  U_DCT2D_rtlc5n1483_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_13_CYMUXFAST,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63721_O
    );
  U_DCT2D_rtlc5n1483_13_FASTCARRY_1080 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63728_O,
      O => U_DCT2D_rtlc5n1483_13_FASTCARRY
    );
  U_DCT2D_rtlc5n1483_13_CYAND_1081 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483_13_CYSELG,
      I1 => U_DCT2D_rtlc5n1483_13_CYSELF,
      O => U_DCT2D_rtlc5n1483_13_CYAND
    );
  U_DCT2D_rtlc5n1483_13_CYMUXFAST_1082 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_13_CYMUXG2,
      IB => U_DCT2D_rtlc5n1483_13_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1483_13_CYAND,
      O => U_DCT2D_rtlc5n1483_13_CYMUXFAST
    );
  U_DCT2D_rtlc5n1483_13_CYMUXG2_1083 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_13_CY0G,
      IB => U_DCT2D_rtlc5n1483_13_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1483_13_CYSELG,
      O => U_DCT2D_rtlc5n1483_13_CYMUXG2
    );
  U_DCT2D_rtlc5n1483_13_CY0G_1084 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(8),
      O => U_DCT2D_rtlc5n1483_13_CY0G
    );
  U_DCT2D_rtlc5n1483_13_CYSELG_1085 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z273,
      O => U_DCT2D_rtlc5n1483_13_CYSELG
    );
  U_DCT2D_rtlc5n1483_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_15_XORF,
      O => U_DCT2D_rtlc5n1483(15)
    );
  U_DCT2D_rtlc5n1483_15_XORF_1086 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1483_15_CYINIT,
      I1 => U_DCT2D_nx65206z270,
      O => U_DCT2D_rtlc5n1483_15_XORF
    );
  U_DCT2D_rtlc5n1483_15_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_15_CY0F,
      IB => U_DCT2D_rtlc5n1483_15_CYINIT,
      SEL => U_DCT2D_rtlc5n1483_15_CYSELF,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63717_O
    );
  U_DCT2D_rtlc5n1483_15_CYMUXF2_1087 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_15_CY0F,
      IB => U_DCT2D_rtlc5n1483_15_CY0F,
      SEL => U_DCT2D_rtlc5n1483_15_CYSELF,
      O => U_DCT2D_rtlc5n1483_15_CYMUXF2
    );
  U_DCT2D_rtlc5n1483_15_CYINIT_1088 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63721_O,
      O => U_DCT2D_rtlc5n1483_15_CYINIT
    );
  U_DCT2D_rtlc5n1483_15_CY0F_1089 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(9),
      O => U_DCT2D_rtlc5n1483_15_CY0F
    );
  U_DCT2D_rtlc5n1483_15_CYSELF_1090 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z270,
      O => U_DCT2D_rtlc5n1483_15_CYSELF
    );
  U_DCT2D_rtlc5n1483_15_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_15_XORG,
      O => U_DCT2D_rtlc5n1483(16)
    );
  U_DCT2D_rtlc5n1483_15_XORG_1091 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_340_add_58_ix65206z63717_O,
      I1 => U_DCT2D_nx65206z267,
      O => U_DCT2D_rtlc5n1483_15_XORG
    );
  U_DCT2D_rtlc5n1483_15_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_15_CYMUXFAST,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63714_O
    );
  U_DCT2D_rtlc5n1483_15_FASTCARRY_1092 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63721_O,
      O => U_DCT2D_rtlc5n1483_15_FASTCARRY
    );
  U_DCT2D_rtlc5n1483_15_CYAND_1093 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483_15_CYSELG,
      I1 => U_DCT2D_rtlc5n1483_15_CYSELF,
      O => U_DCT2D_rtlc5n1483_15_CYAND
    );
  U_DCT2D_rtlc5n1483_15_CYMUXFAST_1094 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_15_CYMUXG2,
      IB => U_DCT2D_rtlc5n1483_15_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1483_15_CYAND,
      O => U_DCT2D_rtlc5n1483_15_CYMUXFAST
    );
  U_DCT2D_rtlc5n1483_15_CYMUXG2_1095 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_15_CY0G,
      IB => U_DCT2D_rtlc5n1483_15_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1483_15_CYSELG,
      O => U_DCT2D_rtlc5n1483_15_CYMUXG2
    );
  U_DCT2D_rtlc5n1483_15_CY0G_1096 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(10),
      O => U_DCT2D_rtlc5n1483_15_CY0G
    );
  U_DCT2D_rtlc5n1483_15_CYSELG_1097 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z267,
      O => U_DCT2D_rtlc5n1483_15_CYSELG
    );
  U_DCT2D_rtlc5n1483_17_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_17_XORF,
      O => U_DCT2D_rtlc5n1483(17)
    );
  U_DCT2D_rtlc5n1483_17_XORF_1098 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1483_17_CYINIT,
      I1 => U_DCT2D_nx65206z264,
      O => U_DCT2D_rtlc5n1483_17_XORF
    );
  U_DCT2D_rtlc5n1483_17_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_17_CY0F,
      IB => U_DCT2D_rtlc5n1483_17_CYINIT,
      SEL => U_DCT2D_rtlc5n1483_17_CYSELF,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63710_O
    );
  U_DCT2D_rtlc5n1483_17_CYMUXF2_1099 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_17_CY0F,
      IB => U_DCT2D_rtlc5n1483_17_CY0F,
      SEL => U_DCT2D_rtlc5n1483_17_CYSELF,
      O => U_DCT2D_rtlc5n1483_17_CYMUXF2
    );
  U_DCT2D_rtlc5n1483_17_CYINIT_1100 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63714_O,
      O => U_DCT2D_rtlc5n1483_17_CYINIT
    );
  U_DCT2D_rtlc5n1483_17_CY0F_1101 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(11),
      O => U_DCT2D_rtlc5n1483_17_CY0F
    );
  U_DCT2D_rtlc5n1483_17_CYSELF_1102 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z264,
      O => U_DCT2D_rtlc5n1483_17_CYSELF
    );
  U_DCT2D_rtlc5n1483_17_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_17_XORG,
      O => U_DCT2D_rtlc5n1483(18)
    );
  U_DCT2D_rtlc5n1483_17_XORG_1103 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_340_add_58_ix65206z63710_O,
      I1 => U_DCT2D_nx65206z261,
      O => U_DCT2D_rtlc5n1483_17_XORG
    );
  U_DCT2D_rtlc5n1483_17_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_17_CYMUXFAST,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63706_O
    );
  U_DCT2D_rtlc5n1483_17_FASTCARRY_1104 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63714_O,
      O => U_DCT2D_rtlc5n1483_17_FASTCARRY
    );
  U_DCT2D_rtlc5n1483_17_CYAND_1105 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483_17_CYSELG,
      I1 => U_DCT2D_rtlc5n1483_17_CYSELF,
      O => U_DCT2D_rtlc5n1483_17_CYAND
    );
  U_DCT2D_rtlc5n1483_17_CYMUXFAST_1106 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_17_CYMUXG2,
      IB => U_DCT2D_rtlc5n1483_17_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1483_17_CYAND,
      O => U_DCT2D_rtlc5n1483_17_CYMUXFAST
    );
  U_DCT2D_rtlc5n1483_17_CYMUXG2_1107 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_17_CY0G,
      IB => U_DCT2D_rtlc5n1483_17_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1483_17_CYSELG,
      O => U_DCT2D_rtlc5n1483_17_CYMUXG2
    );
  U_DCT2D_rtlc5n1483_17_CY0G_1108 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(12),
      O => U_DCT2D_rtlc5n1483_17_CY0G
    );
  U_DCT2D_rtlc5n1483_17_CYSELG_1109 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z261,
      O => U_DCT2D_rtlc5n1483_17_CYSELG
    );
  U_DCT2D_rtlc5n1483_19_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_19_XORF,
      O => U_DCT2D_rtlc5n1483(19)
    );
  U_DCT2D_rtlc5n1483_19_XORF_1110 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1483_19_CYINIT,
      I1 => U_DCT2D_nx65206z258,
      O => U_DCT2D_rtlc5n1483_19_XORF
    );
  U_DCT2D_rtlc5n1483_19_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_19_CY0F,
      IB => U_DCT2D_rtlc5n1483_19_CYINIT,
      SEL => U_DCT2D_rtlc5n1483_19_CYSELF,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63703_O
    );
  U_DCT2D_rtlc5n1483_19_CYMUXF2_1111 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_19_CY0F,
      IB => U_DCT2D_rtlc5n1483_19_CY0F,
      SEL => U_DCT2D_rtlc5n1483_19_CYSELF,
      O => U_DCT2D_rtlc5n1483_19_CYMUXF2
    );
  U_DCT2D_rtlc5n1483_19_CYINIT_1112 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63706_O,
      O => U_DCT2D_rtlc5n1483_19_CYINIT
    );
  U_DCT2D_rtlc5n1483_19_CY0F_1113 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(13),
      O => U_DCT2D_rtlc5n1483_19_CY0F
    );
  U_DCT2D_rtlc5n1483_19_CYSELF_1114 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z258,
      O => U_DCT2D_rtlc5n1483_19_CYSELF
    );
  U_DCT2D_rtlc5n1483_19_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_19_XORG,
      O => U_DCT2D_rtlc5n1483(20)
    );
  U_DCT2D_rtlc5n1483_19_XORG_1115 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_340_add_58_ix65206z63703_O,
      I1 => U_DCT2D_nx65206z255,
      O => U_DCT2D_rtlc5n1483_19_XORG
    );
  U_DCT2D_rtlc5n1483_19_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_19_CYMUXFAST,
      O => U_DCT2D_rtlc_340_add_58_ix65206z63699_O
    );
  U_DCT2D_rtlc5n1483_19_FASTCARRY_1116 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63706_O,
      O => U_DCT2D_rtlc5n1483_19_FASTCARRY
    );
  U_DCT2D_rtlc5n1483_19_CYAND_1117 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483_19_CYSELG,
      I1 => U_DCT2D_rtlc5n1483_19_CYSELF,
      O => U_DCT2D_rtlc5n1483_19_CYAND
    );
  U_DCT2D_rtlc5n1483_19_CYMUXFAST_1118 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_19_CYMUXG2,
      IB => U_DCT2D_rtlc5n1483_19_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1483_19_CYAND,
      O => U_DCT2D_rtlc5n1483_19_CYMUXFAST
    );
  U_DCT2D_rtlc5n1483_19_CYMUXG2_1119 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1483_19_CY0G,
      IB => U_DCT2D_rtlc5n1483_19_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1483_19_CYSELG,
      O => U_DCT2D_rtlc5n1483_19_CYMUXG2
    );
  U_DCT2D_rtlc5n1483_19_CY0G_1120 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s(13),
      O => U_DCT2D_rtlc5n1483_19_CY0G
    );
  U_DCT2D_rtlc5n1483_19_CYSELG_1121 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z255,
      O => U_DCT2D_rtlc5n1483_19_CYSELG
    );
  U_DCT2D_nx65206z253_rt_1122 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_nx65206z253,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z253_rt
    );
  U_DCT2D_rtlc5n1483_21_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1483_21_XORF,
      O => U_DCT2D_rtlc5n1483(21)
    );
  U_DCT2D_rtlc5n1483_21_XORF_1123 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1483_21_CYINIT,
      I1 => U_DCT2D_nx65206z253_rt,
      O => U_DCT2D_rtlc5n1483_21_XORF
    );
  U_DCT2D_rtlc5n1483_21_CYINIT_1124 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_340_add_58_ix65206z63699_O,
      O => U_DCT2D_rtlc5n1483_21_CYINIT
    );
  U_DCT2D_databuf_reg_3_0_DXMUX_1125 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_0_XORF,
      O => U_DCT2D_databuf_reg_3_0_DXMUX
    );
  U_DCT2D_databuf_reg_3_0_XORF_1126 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_0_CYINIT,
      I1 => U_DCT2D_nx54687z1,
      O => U_DCT2D_databuf_reg_3_0_XORF
    );
  U_DCT2D_databuf_reg_3_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_0_CY0F,
      IB => U_DCT2D_databuf_reg_3_0_CYINIT,
      SEL => U_DCT2D_databuf_reg_3_0_CYSELF,
      O => U_DCT2D_rtlc5_1581_add_48_ix55684z63342_O
    );
  U_DCT2D_databuf_reg_3_0_CYINIT_1127 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_0_BXINVNOT,
      O => U_DCT2D_databuf_reg_3_0_CYINIT
    );
  U_DCT2D_databuf_reg_3_0_CY0F_1128 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_0_Q,
      O => U_DCT2D_databuf_reg_3_0_CY0F
    );
  U_DCT2D_databuf_reg_3_0_CYSELF_1129 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx54687z1,
      O => U_DCT2D_databuf_reg_3_0_CYSELF
    );
  U_DCT2D_databuf_reg_3_0_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_29,
      O => U_DCT2D_databuf_reg_3_0_BXINVNOT
    );
  U_DCT2D_databuf_reg_3_0_DYMUX_1130 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_0_XORG,
      O => U_DCT2D_databuf_reg_3_0_DYMUX
    );
  U_DCT2D_databuf_reg_3_0_XORG_1131 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1581_add_48_ix55684z63342_O,
      I1 => U_DCT2D_nx55684z1,
      O => U_DCT2D_databuf_reg_3_0_XORG
    );
  U_DCT2D_databuf_reg_3_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_0_CYMUXG,
      O => U_DCT2D_rtlc5_1581_add_48_ix56681z63342_O
    );
  U_DCT2D_databuf_reg_3_0_CYMUXG_1132 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_0_CY0G,
      IB => U_DCT2D_rtlc5_1581_add_48_ix55684z63342_O,
      SEL => U_DCT2D_databuf_reg_3_0_CYSELG,
      O => U_DCT2D_databuf_reg_3_0_CYMUXG
    );
  U_DCT2D_databuf_reg_3_0_CY0G_1133 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_1_Q,
      O => U_DCT2D_databuf_reg_3_0_CY0G
    );
  U_DCT2D_databuf_reg_3_0_CYSELG_1134 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx55684z1,
      O => U_DCT2D_databuf_reg_3_0_CYSELG
    );
  U_DCT2D_databuf_reg_3_0_SRINV_1135 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_3_0_SRINV
    );
  U_DCT2D_databuf_reg_3_0_CLKINV_1136 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_3_0_CLKINV
    );
  U_DCT2D_databuf_reg_3_0_CEINV_1137 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_3_0_CEINV
    );
  U_DCT1D_ix61816z1321 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_2_Q(2),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_5_Q(2),
      ADR3 => VCC,
      O => U_DCT1D_nx61816z1
    );
  U_DCT2D_databuf_reg_3_2_DXMUX_1138 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_2_XORF,
      O => U_DCT2D_databuf_reg_3_2_DXMUX
    );
  U_DCT2D_databuf_reg_3_2_XORF_1139 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_2_CYINIT,
      I1 => U_DCT2D_nx56681z1,
      O => U_DCT2D_databuf_reg_3_2_XORF
    );
  U_DCT2D_databuf_reg_3_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_2_CY0F,
      IB => U_DCT2D_databuf_reg_3_2_CYINIT,
      SEL => U_DCT2D_databuf_reg_3_2_CYSELF,
      O => U_DCT2D_rtlc5_1581_add_48_ix57678z63342_O
    );
  U_DCT2D_databuf_reg_3_2_CYMUXF2_1140 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_2_CY0F,
      IB => U_DCT2D_databuf_reg_3_2_CY0F,
      SEL => U_DCT2D_databuf_reg_3_2_CYSELF,
      O => U_DCT2D_databuf_reg_3_2_CYMUXF2
    );
  U_DCT2D_databuf_reg_3_2_CYINIT_1141 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1581_add_48_ix56681z63342_O,
      O => U_DCT2D_databuf_reg_3_2_CYINIT
    );
  U_DCT2D_databuf_reg_3_2_CY0F_1142 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_2_Q,
      O => U_DCT2D_databuf_reg_3_2_CY0F
    );
  U_DCT2D_databuf_reg_3_2_CYSELF_1143 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx56681z1,
      O => U_DCT2D_databuf_reg_3_2_CYSELF
    );
  U_DCT2D_databuf_reg_3_2_DYMUX_1144 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_2_XORG,
      O => U_DCT2D_databuf_reg_3_2_DYMUX
    );
  U_DCT2D_databuf_reg_3_2_XORG_1145 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1581_add_48_ix57678z63342_O,
      I1 => U_DCT2D_nx57678z1,
      O => U_DCT2D_databuf_reg_3_2_XORG
    );
  U_DCT2D_databuf_reg_3_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_2_CYMUXFAST,
      O => U_DCT2D_rtlc5_1581_add_48_ix58675z63342_O
    );
  U_DCT2D_databuf_reg_3_2_FASTCARRY_1146 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1581_add_48_ix56681z63342_O,
      O => U_DCT2D_databuf_reg_3_2_FASTCARRY
    );
  U_DCT2D_databuf_reg_3_2_CYAND_1147 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_3_2_CYSELG,
      I1 => U_DCT2D_databuf_reg_3_2_CYSELF,
      O => U_DCT2D_databuf_reg_3_2_CYAND
    );
  U_DCT2D_databuf_reg_3_2_CYMUXFAST_1148 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_2_CYMUXG2,
      IB => U_DCT2D_databuf_reg_3_2_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_3_2_CYAND,
      O => U_DCT2D_databuf_reg_3_2_CYMUXFAST
    );
  U_DCT2D_databuf_reg_3_2_CYMUXG2_1149 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_2_CY0G,
      IB => U_DCT2D_databuf_reg_3_2_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_3_2_CYSELG,
      O => U_DCT2D_databuf_reg_3_2_CYMUXG2
    );
  U_DCT2D_databuf_reg_3_2_CY0G_1150 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_3_Q,
      O => U_DCT2D_databuf_reg_3_2_CY0G
    );
  U_DCT2D_databuf_reg_3_2_CYSELG_1151 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx57678z1,
      O => U_DCT2D_databuf_reg_3_2_CYSELG
    );
  U_DCT2D_databuf_reg_3_2_SRINV_1152 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_3_2_SRINV
    );
  U_DCT2D_databuf_reg_3_2_CLKINV_1153 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_3_2_CLKINV
    );
  U_DCT2D_databuf_reg_3_2_CEINV_1154 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_3_2_CEINV
    );
  U_DCT2D_databuf_reg_3_4_DXMUX_1155 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_4_XORF,
      O => U_DCT2D_databuf_reg_3_4_DXMUX
    );
  U_DCT2D_databuf_reg_3_4_XORF_1156 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_4_CYINIT,
      I1 => U_DCT2D_nx58675z1,
      O => U_DCT2D_databuf_reg_3_4_XORF
    );
  U_DCT2D_databuf_reg_3_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_4_CY0F,
      IB => U_DCT2D_databuf_reg_3_4_CYINIT,
      SEL => U_DCT2D_databuf_reg_3_4_CYSELF,
      O => U_DCT2D_rtlc5_1581_add_48_ix59672z63342_O
    );
  U_DCT2D_databuf_reg_3_4_CYMUXF2_1157 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_4_CY0F,
      IB => U_DCT2D_databuf_reg_3_4_CY0F,
      SEL => U_DCT2D_databuf_reg_3_4_CYSELF,
      O => U_DCT2D_databuf_reg_3_4_CYMUXF2
    );
  U_DCT2D_databuf_reg_3_4_CYINIT_1158 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1581_add_48_ix58675z63342_O,
      O => U_DCT2D_databuf_reg_3_4_CYINIT
    );
  U_DCT2D_databuf_reg_3_4_CY0F_1159 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_4_Q,
      O => U_DCT2D_databuf_reg_3_4_CY0F
    );
  U_DCT2D_databuf_reg_3_4_CYSELF_1160 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx58675z1,
      O => U_DCT2D_databuf_reg_3_4_CYSELF
    );
  U_DCT2D_databuf_reg_3_4_DYMUX_1161 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_4_XORG,
      O => U_DCT2D_databuf_reg_3_4_DYMUX
    );
  U_DCT2D_databuf_reg_3_4_XORG_1162 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1581_add_48_ix59672z63342_O,
      I1 => U_DCT2D_nx59672z1,
      O => U_DCT2D_databuf_reg_3_4_XORG
    );
  U_DCT2D_databuf_reg_3_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_4_CYMUXFAST,
      O => U_DCT2D_rtlc5_1581_add_48_ix60669z63342_O
    );
  U_DCT2D_databuf_reg_3_4_FASTCARRY_1163 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1581_add_48_ix58675z63342_O,
      O => U_DCT2D_databuf_reg_3_4_FASTCARRY
    );
  U_DCT2D_databuf_reg_3_4_CYAND_1164 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_3_4_CYSELG,
      I1 => U_DCT2D_databuf_reg_3_4_CYSELF,
      O => U_DCT2D_databuf_reg_3_4_CYAND
    );
  U_DCT2D_databuf_reg_3_4_CYMUXFAST_1165 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_4_CYMUXG2,
      IB => U_DCT2D_databuf_reg_3_4_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_3_4_CYAND,
      O => U_DCT2D_databuf_reg_3_4_CYMUXFAST
    );
  U_DCT2D_databuf_reg_3_4_CYMUXG2_1166 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_4_CY0G,
      IB => U_DCT2D_databuf_reg_3_4_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_3_4_CYSELG,
      O => U_DCT2D_databuf_reg_3_4_CYMUXG2
    );
  U_DCT2D_databuf_reg_3_4_CY0G_1167 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_5_Q,
      O => U_DCT2D_databuf_reg_3_4_CY0G
    );
  U_DCT2D_databuf_reg_3_4_CYSELG_1168 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx59672z1,
      O => U_DCT2D_databuf_reg_3_4_CYSELG
    );
  U_DCT2D_databuf_reg_3_4_SRINV_1169 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_3_4_SRINV
    );
  U_DCT2D_databuf_reg_3_4_CLKINV_1170 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_3_4_CLKINV
    );
  U_DCT2D_databuf_reg_3_4_CEINV_1171 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_3_4_CEINV
    );
  U_DCT2D_databuf_reg_3_6_DXMUX_1172 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_6_XORF,
      O => U_DCT2D_databuf_reg_3_6_DXMUX
    );
  U_DCT2D_databuf_reg_3_6_XORF_1173 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_6_CYINIT,
      I1 => U_DCT2D_nx60669z1,
      O => U_DCT2D_databuf_reg_3_6_XORF
    );
  U_DCT2D_databuf_reg_3_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_6_CY0F,
      IB => U_DCT2D_databuf_reg_3_6_CYINIT,
      SEL => U_DCT2D_databuf_reg_3_6_CYSELF,
      O => U_DCT2D_rtlc5_1581_add_48_ix61666z63342_O
    );
  U_DCT2D_databuf_reg_3_6_CYMUXF2_1174 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_6_CY0F,
      IB => U_DCT2D_databuf_reg_3_6_CY0F,
      SEL => U_DCT2D_databuf_reg_3_6_CYSELF,
      O => U_DCT2D_databuf_reg_3_6_CYMUXF2
    );
  U_DCT2D_databuf_reg_3_6_CYINIT_1175 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1581_add_48_ix60669z63342_O,
      O => U_DCT2D_databuf_reg_3_6_CYINIT
    );
  U_DCT2D_databuf_reg_3_6_CY0F_1176 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_6_Q,
      O => U_DCT2D_databuf_reg_3_6_CY0F
    );
  U_DCT2D_databuf_reg_3_6_CYSELF_1177 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx60669z1,
      O => U_DCT2D_databuf_reg_3_6_CYSELF
    );
  U_DCT2D_databuf_reg_3_6_DYMUX_1178 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_6_XORG,
      O => U_DCT2D_databuf_reg_3_6_DYMUX
    );
  U_DCT2D_databuf_reg_3_6_XORG_1179 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1581_add_48_ix61666z63342_O,
      I1 => U_DCT2D_nx61666z1,
      O => U_DCT2D_databuf_reg_3_6_XORG
    );
  U_DCT2D_databuf_reg_3_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_6_CYMUXFAST,
      O => U_DCT2D_rtlc5_1581_add_48_ix62663z63342_O
    );
  U_DCT2D_databuf_reg_3_6_FASTCARRY_1180 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1581_add_48_ix60669z63342_O,
      O => U_DCT2D_databuf_reg_3_6_FASTCARRY
    );
  U_DCT2D_databuf_reg_3_6_CYAND_1181 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_3_6_CYSELG,
      I1 => U_DCT2D_databuf_reg_3_6_CYSELF,
      O => U_DCT2D_databuf_reg_3_6_CYAND
    );
  U_DCT2D_databuf_reg_3_6_CYMUXFAST_1182 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_6_CYMUXG2,
      IB => U_DCT2D_databuf_reg_3_6_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_3_6_CYAND,
      O => U_DCT2D_databuf_reg_3_6_CYMUXFAST
    );
  U_DCT2D_databuf_reg_3_6_CYMUXG2_1183 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_6_CY0G,
      IB => U_DCT2D_databuf_reg_3_6_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_3_6_CYSELG,
      O => U_DCT2D_databuf_reg_3_6_CYMUXG2
    );
  U_DCT2D_databuf_reg_3_6_CY0G_1184 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_7_Q,
      O => U_DCT2D_databuf_reg_3_6_CY0G
    );
  U_DCT2D_databuf_reg_3_6_CYSELG_1185 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx61666z1,
      O => U_DCT2D_databuf_reg_3_6_CYSELG
    );
  U_DCT2D_databuf_reg_3_6_SRINV_1186 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_3_6_SRINV
    );
  U_DCT2D_databuf_reg_3_6_CLKINV_1187 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_3_6_CLKINV
    );
  U_DCT2D_databuf_reg_3_6_CEINV_1188 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_3_6_CEINV
    );
  U_DCT2D_databuf_reg_3_8_DXMUX_1189 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_8_XORF,
      O => U_DCT2D_databuf_reg_3_8_DXMUX
    );
  U_DCT2D_databuf_reg_3_8_XORF_1190 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_8_CYINIT,
      I1 => U_DCT2D_nx62663z1,
      O => U_DCT2D_databuf_reg_3_8_XORF
    );
  U_DCT2D_databuf_reg_3_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_8_CY0F,
      IB => U_DCT2D_databuf_reg_3_8_CYINIT,
      SEL => U_DCT2D_databuf_reg_3_8_CYSELF,
      O => U_DCT2D_rtlc5_1581_add_48_ix63660z63342_O
    );
  U_DCT2D_databuf_reg_3_8_CYMUXF2_1191 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_8_CY0F,
      IB => U_DCT2D_databuf_reg_3_8_CY0F,
      SEL => U_DCT2D_databuf_reg_3_8_CYSELF,
      O => U_DCT2D_databuf_reg_3_8_CYMUXF2
    );
  U_DCT2D_databuf_reg_3_8_CYINIT_1192 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1581_add_48_ix62663z63342_O,
      O => U_DCT2D_databuf_reg_3_8_CYINIT
    );
  U_DCT2D_databuf_reg_3_8_CY0F_1193 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_8_Q,
      O => U_DCT2D_databuf_reg_3_8_CY0F
    );
  U_DCT2D_databuf_reg_3_8_CYSELF_1194 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx62663z1,
      O => U_DCT2D_databuf_reg_3_8_CYSELF
    );
  U_DCT2D_databuf_reg_3_8_DYMUX_1195 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_8_XORG,
      O => U_DCT2D_databuf_reg_3_8_DYMUX
    );
  U_DCT2D_databuf_reg_3_8_XORG_1196 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_1581_add_48_ix63660z63342_O,
      I1 => U_DCT2D_nx63660z1,
      O => U_DCT2D_databuf_reg_3_8_XORG
    );
  U_DCT2D_databuf_reg_3_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_8_CYMUXFAST,
      O => U_DCT2D_rtlc5_1581_add_48_ix14976z63342_O
    );
  U_DCT2D_databuf_reg_3_8_FASTCARRY_1197 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1581_add_48_ix62663z63342_O,
      O => U_DCT2D_databuf_reg_3_8_FASTCARRY
    );
  U_DCT2D_databuf_reg_3_8_CYAND_1198 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_3_8_CYSELG,
      I1 => U_DCT2D_databuf_reg_3_8_CYSELF,
      O => U_DCT2D_databuf_reg_3_8_CYAND
    );
  U_DCT2D_databuf_reg_3_8_CYMUXFAST_1199 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_8_CYMUXG2,
      IB => U_DCT2D_databuf_reg_3_8_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_3_8_CYAND,
      O => U_DCT2D_databuf_reg_3_8_CYMUXFAST
    );
  U_DCT2D_databuf_reg_3_8_CYMUXG2_1200 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_3_8_CY0G,
      IB => U_DCT2D_databuf_reg_3_8_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_3_8_CYSELG,
      O => U_DCT2D_databuf_reg_3_8_CYMUXG2
    );
  U_DCT2D_databuf_reg_3_8_CY0G_1201 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_10_Q,
      O => U_DCT2D_databuf_reg_3_8_CY0G
    );
  U_DCT2D_databuf_reg_3_8_CYSELG_1202 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx63660z1,
      O => U_DCT2D_databuf_reg_3_8_CYSELG
    );
  U_DCT2D_databuf_reg_3_8_SRINV_1203 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_3_8_SRINV
    );
  U_DCT2D_databuf_reg_3_8_CLKINV_1204 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_3_8_CLKINV
    );
  U_DCT2D_databuf_reg_3_8_CEINV_1205 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_3_8_CEINV
    );
  U_DCT2D_databuf_reg_3_10_DXMUX_1206 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_10_XORF,
      O => U_DCT2D_databuf_reg_3_10_DXMUX
    );
  U_DCT2D_databuf_reg_3_10_XORF_1207 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_10_CYINIT,
      I1 => U_DCT2D_nx14976z1_rt,
      O => U_DCT2D_databuf_reg_3_10_XORF
    );
  U_DCT2D_databuf_reg_3_10_CYINIT_1208 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_1581_add_48_ix14976z63342_O,
      O => U_DCT2D_databuf_reg_3_10_CYINIT
    );
  U_DCT2D_databuf_reg_3_10_CLKINV_1209 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_3_10_CLKINV
    );
  U_DCT2D_databuf_reg_3_10_CEINV_1210 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_3_10_CEINV
    );
  U_DCT2D_rtlc5n1493_5_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_5_XORF,
      O => U_DCT2D_rtlc5n1493(5)
    );
  U_DCT2D_rtlc5n1493_5_XORF_1211 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1493_5_CYINIT,
      I1 => U_DCT2D_nx65206z40,
      O => U_DCT2D_rtlc5n1493_5_XORF
    );
  U_DCT2D_rtlc5n1493_5_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_5_CY0F,
      IB => U_DCT2D_rtlc5n1493_5_CYINIT,
      SEL => U_DCT2D_rtlc5n1493_5_CYSELF,
      O => U_DCT2D_rtlc_389_add_65_ix65206z63386_O
    );
  U_DCT2D_rtlc5n1493_5_CYINIT_1212 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_5_BXINVNOT,
      O => U_DCT2D_rtlc5n1493_5_CYINIT
    );
  U_DCT2D_rtlc5n1493_5_CY0F_1213 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s(3),
      O => U_DCT2D_rtlc5n1493_5_CY0F
    );
  U_DCT2D_rtlc5n1493_5_CYSELF_1214 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z40,
      O => U_DCT2D_rtlc5n1493_5_CYSELF
    );
  U_DCT2D_rtlc5n1493_5_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_36,
      O => U_DCT2D_rtlc5n1493_5_BXINVNOT
    );
  U_DCT2D_rtlc5n1493_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_5_XORG,
      O => U_DCT2D_rtlc5n1493(6)
    );
  U_DCT2D_rtlc5n1493_5_XORG_1215 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_389_add_65_ix65206z63386_O,
      I1 => U_DCT2D_nx65206z37,
      O => U_DCT2D_rtlc5n1493_5_XORG
    );
  U_DCT2D_rtlc5n1493_5_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_5_CYMUXG,
      O => U_DCT2D_rtlc_389_add_65_ix65206z63383_O
    );
  U_DCT2D_rtlc5n1493_5_CYMUXG_1216 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_5_CY0G,
      IB => U_DCT2D_rtlc_389_add_65_ix65206z63386_O,
      SEL => U_DCT2D_rtlc5n1493_5_CYSELG,
      O => U_DCT2D_rtlc5n1493_5_CYMUXG
    );
  U_DCT2D_rtlc5n1493_5_CY0G_1217 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s(4),
      O => U_DCT2D_rtlc5n1493_5_CY0G
    );
  U_DCT2D_rtlc5n1493_5_CYSELG_1218 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z37,
      O => U_DCT2D_rtlc5n1493_5_CYSELG
    );
  U_DCT2D_rtlc5n1493_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_7_XORF,
      O => U_DCT2D_rtlc5n1493(7)
    );
  U_DCT2D_rtlc5n1493_7_XORF_1219 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1493_7_CYINIT,
      I1 => U_DCT2D_nx65206z34,
      O => U_DCT2D_rtlc5n1493_7_XORF
    );
  U_DCT2D_rtlc5n1493_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_7_CY0F,
      IB => U_DCT2D_rtlc5n1493_7_CYINIT,
      SEL => U_DCT2D_rtlc5n1493_7_CYSELF,
      O => U_DCT2D_rtlc_389_add_65_ix65206z63379_O
    );
  U_DCT2D_rtlc5n1493_7_CYMUXF2_1220 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_7_CY0F,
      IB => U_DCT2D_rtlc5n1493_7_CY0F,
      SEL => U_DCT2D_rtlc5n1493_7_CYSELF,
      O => U_DCT2D_rtlc5n1493_7_CYMUXF2
    );
  U_DCT2D_rtlc5n1493_7_CYINIT_1221 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_389_add_65_ix65206z63383_O,
      O => U_DCT2D_rtlc5n1493_7_CYINIT
    );
  U_DCT2D_rtlc5n1493_7_CY0F_1222 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s(5),
      O => U_DCT2D_rtlc5n1493_7_CY0F
    );
  U_DCT2D_rtlc5n1493_7_CYSELF_1223 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z34,
      O => U_DCT2D_rtlc5n1493_7_CYSELF
    );
  U_DCT2D_rtlc5n1493_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_7_XORG,
      O => U_DCT2D_rtlc5n1493(8)
    );
  U_DCT2D_rtlc5n1493_7_XORG_1224 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_389_add_65_ix65206z63379_O,
      I1 => U_DCT2D_nx65206z31,
      O => U_DCT2D_rtlc5n1493_7_XORG
    );
  U_DCT2D_rtlc5n1493_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_7_CYMUXFAST,
      O => U_DCT2D_rtlc_389_add_65_ix65206z63376_O
    );
  U_DCT2D_rtlc5n1493_7_FASTCARRY_1225 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_389_add_65_ix65206z63383_O,
      O => U_DCT2D_rtlc5n1493_7_FASTCARRY
    );
  U_DCT2D_rtlc5n1493_7_CYAND_1226 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1493_7_CYSELG,
      I1 => U_DCT2D_rtlc5n1493_7_CYSELF,
      O => U_DCT2D_rtlc5n1493_7_CYAND
    );
  U_DCT2D_rtlc5n1493_7_CYMUXFAST_1227 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_7_CYMUXG2,
      IB => U_DCT2D_rtlc5n1493_7_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1493_7_CYAND,
      O => U_DCT2D_rtlc5n1493_7_CYMUXFAST
    );
  U_DCT2D_rtlc5n1493_7_CYMUXG2_1228 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_7_CY0G,
      IB => U_DCT2D_rtlc5n1493_7_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1493_7_CYSELG,
      O => U_DCT2D_rtlc5n1493_7_CYMUXG2
    );
  U_DCT2D_rtlc5n1493_7_CY0G_1229 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s(6),
      O => U_DCT2D_rtlc5n1493_7_CY0G
    );
  U_DCT2D_rtlc5n1493_7_CYSELG_1230 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z31,
      O => U_DCT2D_rtlc5n1493_7_CYSELG
    );
  U_DCT2D_rtlc5n1493_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_9_XORF,
      O => U_DCT2D_rtlc5n1493(9)
    );
  U_DCT2D_rtlc5n1493_9_XORF_1231 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1493_9_CYINIT,
      I1 => U_DCT2D_nx65206z28,
      O => U_DCT2D_rtlc5n1493_9_XORF
    );
  U_DCT2D_rtlc5n1493_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_9_CY0F,
      IB => U_DCT2D_rtlc5n1493_9_CYINIT,
      SEL => U_DCT2D_rtlc5n1493_9_CYSELF,
      O => U_DCT2D_rtlc_389_add_65_ix65206z63372_O
    );
  U_DCT2D_rtlc5n1493_9_CYMUXF2_1232 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_9_CY0F,
      IB => U_DCT2D_rtlc5n1493_9_CY0F,
      SEL => U_DCT2D_rtlc5n1493_9_CYSELF,
      O => U_DCT2D_rtlc5n1493_9_CYMUXF2
    );
  U_DCT2D_rtlc5n1493_9_CYINIT_1233 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_389_add_65_ix65206z63376_O,
      O => U_DCT2D_rtlc5n1493_9_CYINIT
    );
  U_DCT2D_rtlc5n1493_9_CY0F_1234 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s(7),
      O => U_DCT2D_rtlc5n1493_9_CY0F
    );
  U_DCT2D_rtlc5n1493_9_CYSELF_1235 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z28,
      O => U_DCT2D_rtlc5n1493_9_CYSELF
    );
  U_DCT2D_rtlc5n1493_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_9_XORG,
      O => U_DCT2D_rtlc5n1493(10)
    );
  U_DCT2D_rtlc5n1493_9_XORG_1236 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_389_add_65_ix65206z63372_O,
      I1 => U_DCT2D_nx65206z25,
      O => U_DCT2D_rtlc5n1493_9_XORG
    );
  U_DCT2D_rtlc5n1493_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_9_CYMUXFAST,
      O => U_DCT2D_rtlc_389_add_65_ix65206z63369_O
    );
  U_DCT2D_rtlc5n1493_9_FASTCARRY_1237 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_389_add_65_ix65206z63376_O,
      O => U_DCT2D_rtlc5n1493_9_FASTCARRY
    );
  U_DCT2D_rtlc5n1493_9_CYAND_1238 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1493_9_CYSELG,
      I1 => U_DCT2D_rtlc5n1493_9_CYSELF,
      O => U_DCT2D_rtlc5n1493_9_CYAND
    );
  U_DCT2D_rtlc5n1493_9_CYMUXFAST_1239 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_9_CYMUXG2,
      IB => U_DCT2D_rtlc5n1493_9_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1493_9_CYAND,
      O => U_DCT2D_rtlc5n1493_9_CYMUXFAST
    );
  U_DCT2D_rtlc5n1493_9_CYMUXG2_1240 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_9_CY0G,
      IB => U_DCT2D_rtlc5n1493_9_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1493_9_CYSELG,
      O => U_DCT2D_rtlc5n1493_9_CYMUXG2
    );
  U_DCT2D_rtlc5n1493_9_CY0G_1241 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s(8),
      O => U_DCT2D_rtlc5n1493_9_CY0G
    );
  U_DCT2D_rtlc5n1493_9_CYSELG_1242 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z25,
      O => U_DCT2D_rtlc5n1493_9_CYSELG
    );
  U_DCT2D_rtlc5n1493_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_11_XORF,
      O => U_DCT2D_rtlc5n1493(11)
    );
  U_DCT2D_rtlc5n1493_11_XORF_1243 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1493_11_CYINIT,
      I1 => U_DCT2D_nx65206z22,
      O => U_DCT2D_rtlc5n1493_11_XORF
    );
  U_DCT2D_rtlc5n1493_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_11_CY0F,
      IB => U_DCT2D_rtlc5n1493_11_CYINIT,
      SEL => U_DCT2D_rtlc5n1493_11_CYSELF,
      O => U_DCT2D_rtlc_389_add_65_ix65206z63365_O
    );
  U_DCT2D_rtlc5n1493_11_CYMUXF2_1244 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_11_CY0F,
      IB => U_DCT2D_rtlc5n1493_11_CY0F,
      SEL => U_DCT2D_rtlc5n1493_11_CYSELF,
      O => U_DCT2D_rtlc5n1493_11_CYMUXF2
    );
  U_DCT2D_rtlc5n1493_11_CYINIT_1245 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_389_add_65_ix65206z63369_O,
      O => U_DCT2D_rtlc5n1493_11_CYINIT
    );
  U_DCT2D_rtlc5n1493_11_CY0F_1246 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s(9),
      O => U_DCT2D_rtlc5n1493_11_CY0F
    );
  U_DCT2D_rtlc5n1493_11_CYSELF_1247 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z22,
      O => U_DCT2D_rtlc5n1493_11_CYSELF
    );
  U_DCT2D_rtlc5n1493_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_11_XORG,
      O => U_DCT2D_rtlc5n1493(12)
    );
  U_DCT2D_rtlc5n1493_11_XORG_1248 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_389_add_65_ix65206z63365_O,
      I1 => U_DCT2D_nx65206z19,
      O => U_DCT2D_rtlc5n1493_11_XORG
    );
  U_DCT2D_rtlc5n1493_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_11_CYMUXFAST,
      O => U_DCT2D_rtlc_389_add_65_ix65206z63362_O
    );
  U_DCT2D_rtlc5n1493_11_FASTCARRY_1249 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_389_add_65_ix65206z63369_O,
      O => U_DCT2D_rtlc5n1493_11_FASTCARRY
    );
  U_DCT2D_rtlc5n1493_11_CYAND_1250 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1493_11_CYSELG,
      I1 => U_DCT2D_rtlc5n1493_11_CYSELF,
      O => U_DCT2D_rtlc5n1493_11_CYAND
    );
  U_DCT2D_rtlc5n1493_11_CYMUXFAST_1251 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_11_CYMUXG2,
      IB => U_DCT2D_rtlc5n1493_11_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1493_11_CYAND,
      O => U_DCT2D_rtlc5n1493_11_CYMUXFAST
    );
  U_DCT2D_rtlc5n1493_11_CYMUXG2_1252 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_11_CY0G,
      IB => U_DCT2D_rtlc5n1493_11_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1493_11_CYSELG,
      O => U_DCT2D_rtlc5n1493_11_CYMUXG2
    );
  U_DCT2D_rtlc5n1493_11_CY0G_1253 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s(10),
      O => U_DCT2D_rtlc5n1493_11_CY0G
    );
  U_DCT2D_rtlc5n1493_11_CYSELG_1254 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z19,
      O => U_DCT2D_rtlc5n1493_11_CYSELG
    );
  U_DCT2D_rtlc5n1493_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_13_XORF,
      O => U_DCT2D_rtlc5n1493(13)
    );
  U_DCT2D_rtlc5n1493_13_XORF_1255 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1493_13_CYINIT,
      I1 => U_DCT2D_nx65206z16,
      O => U_DCT2D_rtlc5n1493_13_XORF
    );
  U_DCT2D_rtlc5n1493_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_13_CY0F,
      IB => U_DCT2D_rtlc5n1493_13_CYINIT,
      SEL => U_DCT2D_rtlc5n1493_13_CYSELF,
      O => U_DCT2D_rtlc_389_add_65_ix65206z63358_O
    );
  U_DCT2D_rtlc5n1493_13_CYMUXF2_1256 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_13_CY0F,
      IB => U_DCT2D_rtlc5n1493_13_CY0F,
      SEL => U_DCT2D_rtlc5n1493_13_CYSELF,
      O => U_DCT2D_rtlc5n1493_13_CYMUXF2
    );
  U_DCT2D_rtlc5n1493_13_CYINIT_1257 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_389_add_65_ix65206z63362_O,
      O => U_DCT2D_rtlc5n1493_13_CYINIT
    );
  U_DCT2D_rtlc5n1493_13_CY0F_1258 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s(11),
      O => U_DCT2D_rtlc5n1493_13_CY0F
    );
  U_DCT2D_rtlc5n1493_13_CYSELF_1259 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z16,
      O => U_DCT2D_rtlc5n1493_13_CYSELF
    );
  U_DCT2D_rtlc5n1493_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_13_XORG,
      O => U_DCT2D_rtlc5n1493(14)
    );
  U_DCT2D_rtlc5n1493_13_XORG_1260 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_389_add_65_ix65206z63358_O,
      I1 => U_DCT2D_nx65206z13,
      O => U_DCT2D_rtlc5n1493_13_XORG
    );
  U_DCT2D_rtlc5n1493_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_13_CYMUXFAST,
      O => U_DCT2D_rtlc_389_add_65_ix65206z63355_O
    );
  U_DCT2D_rtlc5n1493_13_FASTCARRY_1261 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_389_add_65_ix65206z63362_O,
      O => U_DCT2D_rtlc5n1493_13_FASTCARRY
    );
  U_DCT2D_rtlc5n1493_13_CYAND_1262 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1493_13_CYSELG,
      I1 => U_DCT2D_rtlc5n1493_13_CYSELF,
      O => U_DCT2D_rtlc5n1493_13_CYAND
    );
  U_DCT2D_rtlc5n1493_13_CYMUXFAST_1263 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_13_CYMUXG2,
      IB => U_DCT2D_rtlc5n1493_13_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1493_13_CYAND,
      O => U_DCT2D_rtlc5n1493_13_CYMUXFAST
    );
  U_DCT2D_rtlc5n1493_13_CYMUXG2_1264 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_13_CY0G,
      IB => U_DCT2D_rtlc5n1493_13_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1493_13_CYSELG,
      O => U_DCT2D_rtlc5n1493_13_CYMUXG2
    );
  U_DCT2D_rtlc5n1493_13_CY0G_1265 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s(12),
      O => U_DCT2D_rtlc5n1493_13_CY0G
    );
  U_DCT2D_rtlc5n1493_13_CYSELG_1266 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z13,
      O => U_DCT2D_rtlc5n1493_13_CYSELG
    );
  U_DCT2D_rtlc5n1493_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_15_XORF,
      O => U_DCT2D_rtlc5n1493(15)
    );
  U_DCT2D_rtlc5n1493_15_XORF_1267 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1493_15_CYINIT,
      I1 => U_DCT2D_nx65206z10,
      O => U_DCT2D_rtlc5n1493_15_XORF
    );
  U_DCT2D_rtlc5n1493_15_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_15_CY0F,
      IB => U_DCT2D_rtlc5n1493_15_CYINIT,
      SEL => U_DCT2D_rtlc5n1493_15_CYSELF,
      O => U_DCT2D_rtlc_389_add_65_ix65206z63351_O
    );
  U_DCT2D_rtlc5n1493_15_CYMUXF2_1268 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_15_CY0F,
      IB => U_DCT2D_rtlc5n1493_15_CY0F,
      SEL => U_DCT2D_rtlc5n1493_15_CYSELF,
      O => U_DCT2D_rtlc5n1493_15_CYMUXF2
    );
  U_DCT2D_rtlc5n1493_15_CYINIT_1269 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_389_add_65_ix65206z63355_O,
      O => U_DCT2D_rtlc5n1493_15_CYINIT
    );
  U_DCT2D_rtlc5n1493_15_CY0F_1270 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s(13),
      O => U_DCT2D_rtlc5n1493_15_CY0F
    );
  U_DCT2D_rtlc5n1493_15_CYSELF_1271 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z10,
      O => U_DCT2D_rtlc5n1493_15_CYSELF
    );
  U_DCT2D_rtlc5n1493_15_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_15_XORG,
      O => U_DCT2D_rtlc5n1493(16)
    );
  U_DCT2D_rtlc5n1493_15_XORG_1272 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_389_add_65_ix65206z63351_O,
      I1 => U_DCT2D_nx65206z7,
      O => U_DCT2D_rtlc5n1493_15_XORG
    );
  U_DCT2D_rtlc5n1493_15_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_15_CYMUXFAST,
      O => U_DCT2D_rtlc_389_add_65_ix65206z63348_O
    );
  U_DCT2D_rtlc5n1493_15_FASTCARRY_1273 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_389_add_65_ix65206z63355_O,
      O => U_DCT2D_rtlc5n1493_15_FASTCARRY
    );
  U_DCT2D_rtlc5n1493_15_CYAND_1274 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1493_15_CYSELG,
      I1 => U_DCT2D_rtlc5n1493_15_CYSELF,
      O => U_DCT2D_rtlc5n1493_15_CYAND
    );
  U_DCT2D_rtlc5n1493_15_CYMUXFAST_1275 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_15_CYMUXG2,
      IB => U_DCT2D_rtlc5n1493_15_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1493_15_CYAND,
      O => U_DCT2D_rtlc5n1493_15_CYMUXFAST
    );
  U_DCT2D_rtlc5n1493_15_CYMUXG2_1276 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1493_15_CY0G,
      IB => U_DCT2D_rtlc5n1493_15_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1493_15_CYSELG,
      O => U_DCT2D_rtlc5n1493_15_CYMUXG2
    );
  U_DCT2D_rtlc5n1493_15_CY0G_1277 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s(13),
      O => U_DCT2D_rtlc5n1493_15_CY0G
    );
  U_DCT2D_rtlc5n1493_15_CYSELG_1278 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z7,
      O => U_DCT2D_rtlc5n1493_15_CYSELG
    );
  U_DCT2D_nx65206z5_rt_1279 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT2D_nx65206z5,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z5_rt
    );
  U_DCT2D_rtlc5n1493_17_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1493_17_XORF,
      O => U_DCT2D_rtlc5n1493(17)
    );
  U_DCT2D_rtlc5n1493_17_XORF_1280 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1493_17_CYINIT,
      I1 => U_DCT2D_nx65206z5_rt,
      O => U_DCT2D_rtlc5n1493_17_XORF
    );
  U_DCT2D_rtlc5n1493_17_CYINIT_1281 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_389_add_65_ix65206z63348_O,
      O => U_DCT2D_rtlc5n1493_17_CYINIT
    );
  U_DCT1D_rtlc5n1359_6_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_6_XORF,
      O => U_DCT1D_rtlc5n1359(6)
    );
  U_DCT1D_rtlc5n1359_6_XORF_1282 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1359_6_CYINIT,
      I1 => U_DCT1D_nx59700z431,
      O => U_DCT1D_rtlc5n1359_6_XORF
    );
  U_DCT1D_rtlc5n1359_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_6_CY0F,
      IB => U_DCT1D_rtlc5n1359_6_CYINIT,
      SEL => U_DCT1D_rtlc5n1359_6_CYSELF,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63921_O
    );
  U_DCT1D_rtlc5n1359_6_CYINIT_1283 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_6_BXINVNOT,
      O => U_DCT1D_rtlc5n1359_6_CYINIT
    );
  U_DCT1D_rtlc5n1359_6_CY0F_1284 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z432,
      O => U_DCT1D_rtlc5n1359_6_CY0F
    );
  U_DCT1D_rtlc5n1359_6_FAND : X_AND2
    port map (
      I0 => romodatao6_s(0),
      I1 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z432
    );
  U_DCT1D_rtlc5n1359_6_CYSELF_1285 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z431,
      O => U_DCT1D_rtlc5n1359_6_CYSELF
    );
  U_DCT1D_rtlc5n1359_6_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_9,
      O => U_DCT1D_rtlc5n1359_6_BXINVNOT
    );
  U_DCT1D_rtlc5n1359_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_6_XORG,
      O => U_DCT1D_rtlc5n1359(7)
    );
  U_DCT1D_rtlc5n1359_6_XORG_1286 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_522_add_32_ix59700z63921_O,
      I1 => U_DCT1D_nx59700z427,
      O => U_DCT1D_rtlc5n1359_6_XORG
    );
  U_DCT1D_rtlc5n1359_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_6_CYMUXG,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63916_O
    );
  U_DCT1D_rtlc5n1359_6_CYMUXG_1287 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_6_CY0G,
      IB => U_DCT1D_rtlc_522_add_32_ix59700z63921_O,
      SEL => U_DCT1D_rtlc5n1359_6_CYSELG,
      O => U_DCT1D_rtlc5n1359_6_CYMUXG
    );
  U_DCT1D_rtlc5n1359_6_CY0G_1288 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z428,
      O => U_DCT1D_rtlc5n1359_6_CY0G
    );
  U_DCT1D_rtlc5n1359_6_CYSELG_1289 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z427,
      O => U_DCT1D_rtlc5n1359_6_CYSELG
    );
  U_DCT1D_ix59700z1885 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z420,
      ADR1 => U_DCT1D_rtlc5n1347(9),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z419
    );
  U_DCT1D_rtlc5n1359_8_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_8_XORF,
      O => U_DCT1D_rtlc5n1359(8)
    );
  U_DCT1D_rtlc5n1359_8_XORF_1290 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1359_8_CYINIT,
      I1 => U_DCT1D_nx59700z423,
      O => U_DCT1D_rtlc5n1359_8_XORF
    );
  U_DCT1D_rtlc5n1359_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_8_CY0F,
      IB => U_DCT1D_rtlc5n1359_8_CYINIT,
      SEL => U_DCT1D_rtlc5n1359_8_CYSELF,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63910_O
    );
  U_DCT1D_rtlc5n1359_8_CYMUXF2_1291 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_8_CY0F,
      IB => U_DCT1D_rtlc5n1359_8_CY0F,
      SEL => U_DCT1D_rtlc5n1359_8_CYSELF,
      O => U_DCT1D_rtlc5n1359_8_CYMUXF2
    );
  U_DCT1D_rtlc5n1359_8_CYINIT_1292 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63916_O,
      O => U_DCT1D_rtlc5n1359_8_CYINIT
    );
  U_DCT1D_rtlc5n1359_8_CY0F_1293 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z424,
      O => U_DCT1D_rtlc5n1359_8_CY0F
    );
  U_DCT1D_rtlc5n1359_8_CYSELF_1294 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z423,
      O => U_DCT1D_rtlc5n1359_8_CYSELF
    );
  U_DCT1D_rtlc5n1359_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_8_XORG,
      O => U_DCT1D_rtlc5n1359(9)
    );
  U_DCT1D_rtlc5n1359_8_XORG_1295 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_522_add_32_ix59700z63910_O,
      I1 => U_DCT1D_nx59700z419,
      O => U_DCT1D_rtlc5n1359_8_XORG
    );
  U_DCT1D_rtlc5n1359_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_8_CYMUXFAST,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63904_O
    );
  U_DCT1D_rtlc5n1359_8_FASTCARRY_1296 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63916_O,
      O => U_DCT1D_rtlc5n1359_8_FASTCARRY
    );
  U_DCT1D_rtlc5n1359_8_CYAND_1297 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1359_8_CYSELG,
      I1 => U_DCT1D_rtlc5n1359_8_CYSELF,
      O => U_DCT1D_rtlc5n1359_8_CYAND
    );
  U_DCT1D_rtlc5n1359_8_CYMUXFAST_1298 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_8_CYMUXG2,
      IB => U_DCT1D_rtlc5n1359_8_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1359_8_CYAND,
      O => U_DCT1D_rtlc5n1359_8_CYMUXFAST
    );
  U_DCT1D_rtlc5n1359_8_CYMUXG2_1299 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_8_CY0G,
      IB => U_DCT1D_rtlc5n1359_8_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1359_8_CYSELG,
      O => U_DCT1D_rtlc5n1359_8_CYMUXG2
    );
  U_DCT1D_rtlc5n1359_8_CY0G_1300 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z420,
      O => U_DCT1D_rtlc5n1359_8_CY0G
    );
  U_DCT1D_rtlc5n1359_8_CYSELG_1301 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z419,
      O => U_DCT1D_rtlc5n1359_8_CYSELG
    );
  U_DCT1D_rtlc5n1359_10_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_10_XORF,
      O => U_DCT1D_rtlc5n1359(10)
    );
  U_DCT1D_rtlc5n1359_10_XORF_1302 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1359_10_CYINIT,
      I1 => U_DCT1D_nx59700z415,
      O => U_DCT1D_rtlc5n1359_10_XORF
    );
  U_DCT1D_rtlc5n1359_10_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_10_CY0F,
      IB => U_DCT1D_rtlc5n1359_10_CYINIT,
      SEL => U_DCT1D_rtlc5n1359_10_CYSELF,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63898_O
    );
  U_DCT1D_rtlc5n1359_10_CYMUXF2_1303 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_10_CY0F,
      IB => U_DCT1D_rtlc5n1359_10_CY0F,
      SEL => U_DCT1D_rtlc5n1359_10_CYSELF,
      O => U_DCT1D_rtlc5n1359_10_CYMUXF2
    );
  U_DCT1D_rtlc5n1359_10_CYINIT_1304 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63904_O,
      O => U_DCT1D_rtlc5n1359_10_CYINIT
    );
  U_DCT1D_rtlc5n1359_10_CY0F_1305 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z416,
      O => U_DCT1D_rtlc5n1359_10_CY0F
    );
  U_DCT1D_rtlc5n1359_10_CYSELF_1306 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z415,
      O => U_DCT1D_rtlc5n1359_10_CYSELF
    );
  U_DCT1D_rtlc5n1359_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_10_XORG,
      O => U_DCT1D_rtlc5n1359(11)
    );
  U_DCT1D_rtlc5n1359_10_XORG_1307 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_522_add_32_ix59700z63898_O,
      I1 => U_DCT1D_nx59700z411,
      O => U_DCT1D_rtlc5n1359_10_XORG
    );
  U_DCT1D_rtlc5n1359_10_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_10_CYMUXFAST,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63892_O
    );
  U_DCT1D_rtlc5n1359_10_FASTCARRY_1308 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63904_O,
      O => U_DCT1D_rtlc5n1359_10_FASTCARRY
    );
  U_DCT1D_rtlc5n1359_10_CYAND_1309 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1359_10_CYSELG,
      I1 => U_DCT1D_rtlc5n1359_10_CYSELF,
      O => U_DCT1D_rtlc5n1359_10_CYAND
    );
  U_DCT1D_rtlc5n1359_10_CYMUXFAST_1310 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_10_CYMUXG2,
      IB => U_DCT1D_rtlc5n1359_10_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1359_10_CYAND,
      O => U_DCT1D_rtlc5n1359_10_CYMUXFAST
    );
  U_DCT1D_rtlc5n1359_10_CYMUXG2_1311 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_10_CY0G,
      IB => U_DCT1D_rtlc5n1359_10_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1359_10_CYSELG,
      O => U_DCT1D_rtlc5n1359_10_CYMUXG2
    );
  U_DCT1D_rtlc5n1359_10_CY0G_1312 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z412,
      O => U_DCT1D_rtlc5n1359_10_CY0G
    );
  U_DCT1D_rtlc5n1359_10_CYSELG_1313 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z411,
      O => U_DCT1D_rtlc5n1359_10_CYSELG
    );
  U_DCT1D_rtlc5n1359_12_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_12_XORF,
      O => U_DCT1D_rtlc5n1359(12)
    );
  U_DCT1D_rtlc5n1359_12_XORF_1314 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1359_12_CYINIT,
      I1 => U_DCT1D_nx59700z407,
      O => U_DCT1D_rtlc5n1359_12_XORF
    );
  U_DCT1D_rtlc5n1359_12_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_12_CY0F,
      IB => U_DCT1D_rtlc5n1359_12_CYINIT,
      SEL => U_DCT1D_rtlc5n1359_12_CYSELF,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63886_O
    );
  U_DCT1D_rtlc5n1359_12_CYMUXF2_1315 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_12_CY0F,
      IB => U_DCT1D_rtlc5n1359_12_CY0F,
      SEL => U_DCT1D_rtlc5n1359_12_CYSELF,
      O => U_DCT1D_rtlc5n1359_12_CYMUXF2
    );
  U_DCT1D_rtlc5n1359_12_CYINIT_1316 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63892_O,
      O => U_DCT1D_rtlc5n1359_12_CYINIT
    );
  U_DCT1D_rtlc5n1359_12_CY0F_1317 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z408,
      O => U_DCT1D_rtlc5n1359_12_CY0F
    );
  U_DCT1D_rtlc5n1359_12_CYSELF_1318 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z407,
      O => U_DCT1D_rtlc5n1359_12_CYSELF
    );
  U_DCT1D_rtlc5n1359_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_12_XORG,
      O => U_DCT1D_rtlc5n1359(13)
    );
  U_DCT1D_rtlc5n1359_12_XORG_1319 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_522_add_32_ix59700z63886_O,
      I1 => U_DCT1D_nx59700z403,
      O => U_DCT1D_rtlc5n1359_12_XORG
    );
  U_DCT1D_rtlc5n1359_12_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_12_CYMUXFAST,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63880_O
    );
  U_DCT1D_rtlc5n1359_12_FASTCARRY_1320 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63892_O,
      O => U_DCT1D_rtlc5n1359_12_FASTCARRY
    );
  U_DCT1D_rtlc5n1359_12_CYAND_1321 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1359_12_CYSELG,
      I1 => U_DCT1D_rtlc5n1359_12_CYSELF,
      O => U_DCT1D_rtlc5n1359_12_CYAND
    );
  U_DCT1D_rtlc5n1359_12_CYMUXFAST_1322 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_12_CYMUXG2,
      IB => U_DCT1D_rtlc5n1359_12_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1359_12_CYAND,
      O => U_DCT1D_rtlc5n1359_12_CYMUXFAST
    );
  U_DCT1D_rtlc5n1359_12_CYMUXG2_1323 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_12_CY0G,
      IB => U_DCT1D_rtlc5n1359_12_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1359_12_CYSELG,
      O => U_DCT1D_rtlc5n1359_12_CYMUXG2
    );
  U_DCT1D_rtlc5n1359_12_CY0G_1324 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z404,
      O => U_DCT1D_rtlc5n1359_12_CY0G
    );
  U_DCT1D_rtlc5n1359_12_CYSELG_1325 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z403,
      O => U_DCT1D_rtlc5n1359_12_CYSELG
    );
  U_DCT1D_rtlc5n1359_14_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_14_XORF,
      O => U_DCT1D_rtlc5n1359(14)
    );
  U_DCT1D_rtlc5n1359_14_XORF_1326 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1359_14_CYINIT,
      I1 => U_DCT1D_nx59700z399,
      O => U_DCT1D_rtlc5n1359_14_XORF
    );
  U_DCT1D_rtlc5n1359_14_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_14_CY0F,
      IB => U_DCT1D_rtlc5n1359_14_CYINIT,
      SEL => U_DCT1D_rtlc5n1359_14_CYSELF,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63874_O
    );
  U_DCT1D_rtlc5n1359_14_CYMUXF2_1327 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_14_CY0F,
      IB => U_DCT1D_rtlc5n1359_14_CY0F,
      SEL => U_DCT1D_rtlc5n1359_14_CYSELF,
      O => U_DCT1D_rtlc5n1359_14_CYMUXF2
    );
  U_DCT1D_rtlc5n1359_14_CYINIT_1328 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63880_O,
      O => U_DCT1D_rtlc5n1359_14_CYINIT
    );
  U_DCT1D_rtlc5n1359_14_CY0F_1329 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z400,
      O => U_DCT1D_rtlc5n1359_14_CY0F
    );
  U_DCT1D_rtlc5n1359_14_CYSELF_1330 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z399,
      O => U_DCT1D_rtlc5n1359_14_CYSELF
    );
  U_DCT1D_rtlc5n1359_14_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_14_XORG,
      O => U_DCT1D_rtlc5n1359(15)
    );
  U_DCT1D_rtlc5n1359_14_XORG_1331 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_522_add_32_ix59700z63874_O,
      I1 => U_DCT1D_nx59700z395,
      O => U_DCT1D_rtlc5n1359_14_XORG
    );
  U_DCT1D_rtlc5n1359_14_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_14_CYMUXFAST,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63868_O
    );
  U_DCT1D_rtlc5n1359_14_FASTCARRY_1332 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63880_O,
      O => U_DCT1D_rtlc5n1359_14_FASTCARRY
    );
  U_DCT1D_rtlc5n1359_14_CYAND_1333 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1359_14_CYSELG,
      I1 => U_DCT1D_rtlc5n1359_14_CYSELF,
      O => U_DCT1D_rtlc5n1359_14_CYAND
    );
  U_DCT1D_rtlc5n1359_14_CYMUXFAST_1334 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_14_CYMUXG2,
      IB => U_DCT1D_rtlc5n1359_14_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1359_14_CYAND,
      O => U_DCT1D_rtlc5n1359_14_CYMUXFAST
    );
  U_DCT1D_rtlc5n1359_14_CYMUXG2_1335 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_14_CY0G,
      IB => U_DCT1D_rtlc5n1359_14_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1359_14_CYSELG,
      O => U_DCT1D_rtlc5n1359_14_CYMUXG2
    );
  U_DCT1D_rtlc5n1359_14_CY0G_1336 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z396,
      O => U_DCT1D_rtlc5n1359_14_CY0G
    );
  U_DCT1D_rtlc5n1359_14_CYSELG_1337 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z395,
      O => U_DCT1D_rtlc5n1359_14_CYSELG
    );
  U_DCT1D_rtlc5n1359_16_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_16_XORF,
      O => U_DCT1D_rtlc5n1359(16)
    );
  U_DCT1D_rtlc5n1359_16_XORF_1338 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1359_16_CYINIT,
      I1 => U_DCT1D_nx59700z391,
      O => U_DCT1D_rtlc5n1359_16_XORF
    );
  U_DCT1D_rtlc5n1359_16_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_16_CY0F,
      IB => U_DCT1D_rtlc5n1359_16_CYINIT,
      SEL => U_DCT1D_rtlc5n1359_16_CYSELF,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63862_O
    );
  U_DCT1D_rtlc5n1359_16_CYMUXF2_1339 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_16_CY0F,
      IB => U_DCT1D_rtlc5n1359_16_CY0F,
      SEL => U_DCT1D_rtlc5n1359_16_CYSELF,
      O => U_DCT1D_rtlc5n1359_16_CYMUXF2
    );
  U_DCT1D_rtlc5n1359_16_CYINIT_1340 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63868_O,
      O => U_DCT1D_rtlc5n1359_16_CYINIT
    );
  U_DCT1D_rtlc5n1359_16_CY0F_1341 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z392,
      O => U_DCT1D_rtlc5n1359_16_CY0F
    );
  U_DCT1D_rtlc5n1359_16_CYSELF_1342 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z391,
      O => U_DCT1D_rtlc5n1359_16_CYSELF
    );
  U_DCT1D_rtlc5n1359_16_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_16_XORG,
      O => U_DCT1D_rtlc5n1359(17)
    );
  U_DCT1D_rtlc5n1359_16_XORG_1343 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_522_add_32_ix59700z63862_O,
      I1 => U_DCT1D_nx59700z387,
      O => U_DCT1D_rtlc5n1359_16_XORG
    );
  U_DCT1D_rtlc5n1359_16_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_16_CYMUXFAST,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63856_O
    );
  U_DCT1D_rtlc5n1359_16_FASTCARRY_1344 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63868_O,
      O => U_DCT1D_rtlc5n1359_16_FASTCARRY
    );
  U_DCT1D_rtlc5n1359_16_CYAND_1345 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1359_16_CYSELG,
      I1 => U_DCT1D_rtlc5n1359_16_CYSELF,
      O => U_DCT1D_rtlc5n1359_16_CYAND
    );
  U_DCT1D_rtlc5n1359_16_CYMUXFAST_1346 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_16_CYMUXG2,
      IB => U_DCT1D_rtlc5n1359_16_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1359_16_CYAND,
      O => U_DCT1D_rtlc5n1359_16_CYMUXFAST
    );
  U_DCT1D_rtlc5n1359_16_CYMUXG2_1347 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_16_CY0G,
      IB => U_DCT1D_rtlc5n1359_16_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1359_16_CYSELG,
      O => U_DCT1D_rtlc5n1359_16_CYMUXG2
    );
  U_DCT1D_rtlc5n1359_16_CY0G_1348 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z388,
      O => U_DCT1D_rtlc5n1359_16_CY0G
    );
  U_DCT1D_rtlc5n1359_16_CYSELG_1349 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z387,
      O => U_DCT1D_rtlc5n1359_16_CYSELG
    );
  U_DCT1D_rtlc5n1359_18_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_18_XORF,
      O => U_DCT1D_rtlc5n1359(18)
    );
  U_DCT1D_rtlc5n1359_18_XORF_1350 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1359_18_CYINIT,
      I1 => U_DCT1D_nx59700z383,
      O => U_DCT1D_rtlc5n1359_18_XORF
    );
  U_DCT1D_rtlc5n1359_18_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_18_CY0F,
      IB => U_DCT1D_rtlc5n1359_18_CYINIT,
      SEL => U_DCT1D_rtlc5n1359_18_CYSELF,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63851_O
    );
  U_DCT1D_rtlc5n1359_18_CYMUXF2_1351 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_18_CY0F,
      IB => U_DCT1D_rtlc5n1359_18_CY0F,
      SEL => U_DCT1D_rtlc5n1359_18_CYSELF,
      O => U_DCT1D_rtlc5n1359_18_CYMUXF2
    );
  U_DCT1D_rtlc5n1359_18_CYINIT_1352 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63856_O,
      O => U_DCT1D_rtlc5n1359_18_CYINIT
    );
  U_DCT1D_rtlc5n1359_18_CY0F_1353 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z384,
      O => U_DCT1D_rtlc5n1359_18_CY0F
    );
  U_DCT1D_rtlc5n1359_18_CYSELF_1354 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z383,
      O => U_DCT1D_rtlc5n1359_18_CYSELF
    );
  U_DCT1D_rtlc5n1359_18_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_18_XORG,
      O => U_DCT1D_rtlc5n1359(19)
    );
  U_DCT1D_rtlc5n1359_18_XORG_1355 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_522_add_32_ix59700z63851_O,
      I1 => U_DCT1D_nx59700z380,
      O => U_DCT1D_rtlc5n1359_18_XORG
    );
  U_DCT1D_rtlc5n1359_18_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_18_CYMUXFAST,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63846_O
    );
  U_DCT1D_rtlc5n1359_18_FASTCARRY_1356 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63856_O,
      O => U_DCT1D_rtlc5n1359_18_FASTCARRY
    );
  U_DCT1D_rtlc5n1359_18_CYAND_1357 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1359_18_CYSELG,
      I1 => U_DCT1D_rtlc5n1359_18_CYSELF,
      O => U_DCT1D_rtlc5n1359_18_CYAND
    );
  U_DCT1D_rtlc5n1359_18_CYMUXFAST_1358 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_18_CYMUXG2,
      IB => U_DCT1D_rtlc5n1359_18_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1359_18_CYAND,
      O => U_DCT1D_rtlc5n1359_18_CYMUXFAST
    );
  U_DCT1D_rtlc5n1359_18_CYMUXG2_1359 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_18_CY0G,
      IB => U_DCT1D_rtlc5n1359_18_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1359_18_CYSELG,
      O => U_DCT1D_rtlc5n1359_18_CYMUXG2
    );
  U_DCT1D_rtlc5n1359_18_CY0G_1360 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z253,
      O => U_DCT1D_rtlc5n1359_18_CY0G
    );
  U_DCT1D_rtlc5n1359_18_CYSELG_1361 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z380,
      O => U_DCT1D_rtlc5n1359_18_CYSELG
    );
  U_DCT1D_ix59700z1675 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_rtlc5n1347(21),
      ADR2 => U_DCT1D_nx59700z253,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z252
    );
  U_DCT1D_rtlc5n1359_20_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_20_XORF,
      O => U_DCT1D_rtlc5n1359(20)
    );
  U_DCT1D_rtlc5n1359_20_XORF_1362 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1359_20_CYINIT,
      I1 => U_DCT1D_nx59700z377,
      O => U_DCT1D_rtlc5n1359_20_XORF
    );
  U_DCT1D_rtlc5n1359_20_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1359_20_CY0F,
      IB => U_DCT1D_rtlc5n1359_20_CYINIT,
      SEL => U_DCT1D_rtlc5n1359_20_CYSELF,
      O => U_DCT1D_rtlc_522_add_32_ix59700z63841_O
    );
  U_DCT1D_rtlc5n1359_20_CYINIT_1363 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_522_add_32_ix59700z63846_O,
      O => U_DCT1D_rtlc5n1359_20_CYINIT
    );
  U_DCT1D_rtlc5n1359_20_CY0F_1364 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z253,
      O => U_DCT1D_rtlc5n1359_20_CY0F
    );
  U_DCT1D_rtlc5n1359_20_CYSELF_1365 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z377,
      O => U_DCT1D_rtlc5n1359_20_CYSELF
    );
  U_DCT1D_rtlc5n1359_20_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1359_20_XORG,
      O => U_DCT1D_rtlc5n1359(21)
    );
  U_DCT1D_rtlc5n1359_20_XORG_1366 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_522_add_32_ix59700z63841_O,
      I1 => U_DCT1D_nx59700z252,
      O => U_DCT1D_rtlc5n1359_20_XORG
    );
  U_DCT1D_reg_databuf_reg_2_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_2_2_DXMUX,
      CE => U_DCT1D_databuf_reg_2_2_CEINV,
      CLK => U_DCT1D_databuf_reg_2_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_2_2_FFX_RST,
      O => U_DCT1D_databuf_reg_2_Q(2)
    );
  U_DCT1D_databuf_reg_2_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_2_2_FFX_RST
    );
  U_DCT2D_databuf_reg_6_0_DXMUX_1367 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_0_XORF,
      O => U_DCT2D_databuf_reg_6_0_DXMUX
    );
  U_DCT2D_databuf_reg_6_0_XORF_1368 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_0_CYINIT,
      I1 => U_DCT2D_nx39282z1,
      O => U_DCT2D_databuf_reg_6_0_XORF
    );
  U_DCT2D_databuf_reg_6_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_0_CY0F,
      IB => U_DCT2D_databuf_reg_6_0_CYINIT,
      SEL => U_DCT2D_databuf_reg_6_0_CYSELF,
      O => U_DCT2D_rtlc5_99_sub_43_ix40279z63342_O
    );
  U_DCT2D_databuf_reg_6_0_CYINIT_1369 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GLOBAL_LOGIC1_27,
      O => U_DCT2D_databuf_reg_6_0_CYINIT
    );
  U_DCT2D_databuf_reg_6_0_CY0F_1370 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_0_Q,
      O => U_DCT2D_databuf_reg_6_0_CY0F
    );
  U_DCT2D_databuf_reg_6_0_CYSELF_1371 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx39282z1,
      O => U_DCT2D_databuf_reg_6_0_CYSELF
    );
  U_DCT2D_databuf_reg_6_0_DYMUX_1372 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_0_XORG,
      O => U_DCT2D_databuf_reg_6_0_DYMUX
    );
  U_DCT2D_databuf_reg_6_0_XORG_1373 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_99_sub_43_ix40279z63342_O,
      I1 => U_DCT2D_nx40279z1,
      O => U_DCT2D_databuf_reg_6_0_XORG
    );
  U_DCT2D_databuf_reg_6_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_0_CYMUXG,
      O => U_DCT2D_rtlc5_99_sub_43_ix41276z63342_O
    );
  U_DCT2D_databuf_reg_6_0_CYMUXG_1374 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_0_CY0G,
      IB => U_DCT2D_rtlc5_99_sub_43_ix40279z63342_O,
      SEL => U_DCT2D_databuf_reg_6_0_CYSELG,
      O => U_DCT2D_databuf_reg_6_0_CYMUXG
    );
  U_DCT2D_databuf_reg_6_0_CY0G_1375 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_1_Q,
      O => U_DCT2D_databuf_reg_6_0_CY0G
    );
  U_DCT2D_databuf_reg_6_0_CYSELG_1376 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx40279z1,
      O => U_DCT2D_databuf_reg_6_0_CYSELG
    );
  U_DCT2D_databuf_reg_6_0_SRINV_1377 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_6_0_SRINV
    );
  U_DCT2D_databuf_reg_6_0_CLKINV_1378 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_6_0_CLKINV
    );
  U_DCT2D_databuf_reg_6_0_CEINV_1379 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_6_0_CEINV
    );
  U_DCT2D_databuf_reg_6_2_DXMUX_1380 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_2_XORF,
      O => U_DCT2D_databuf_reg_6_2_DXMUX
    );
  U_DCT2D_databuf_reg_6_2_XORF_1381 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_2_CYINIT,
      I1 => U_DCT2D_nx41276z1,
      O => U_DCT2D_databuf_reg_6_2_XORF
    );
  U_DCT2D_databuf_reg_6_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_2_CY0F,
      IB => U_DCT2D_databuf_reg_6_2_CYINIT,
      SEL => U_DCT2D_databuf_reg_6_2_CYSELF,
      O => U_DCT2D_rtlc5_99_sub_43_ix42273z63342_O
    );
  U_DCT2D_databuf_reg_6_2_CYMUXF2_1382 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_2_CY0F,
      IB => U_DCT2D_databuf_reg_6_2_CY0F,
      SEL => U_DCT2D_databuf_reg_6_2_CYSELF,
      O => U_DCT2D_databuf_reg_6_2_CYMUXF2
    );
  U_DCT2D_databuf_reg_6_2_CYINIT_1383 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_99_sub_43_ix41276z63342_O,
      O => U_DCT2D_databuf_reg_6_2_CYINIT
    );
  U_DCT2D_databuf_reg_6_2_CY0F_1384 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_2_Q,
      O => U_DCT2D_databuf_reg_6_2_CY0F
    );
  U_DCT2D_databuf_reg_6_2_CYSELF_1385 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx41276z1,
      O => U_DCT2D_databuf_reg_6_2_CYSELF
    );
  U_DCT2D_databuf_reg_6_2_DYMUX_1386 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_2_XORG,
      O => U_DCT2D_databuf_reg_6_2_DYMUX
    );
  U_DCT2D_databuf_reg_6_2_XORG_1387 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_99_sub_43_ix42273z63342_O,
      I1 => U_DCT2D_nx42273z1,
      O => U_DCT2D_databuf_reg_6_2_XORG
    );
  U_DCT2D_databuf_reg_6_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_2_CYMUXFAST,
      O => U_DCT2D_rtlc5_99_sub_43_ix43270z63342_O
    );
  U_DCT2D_databuf_reg_6_2_FASTCARRY_1388 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_99_sub_43_ix41276z63342_O,
      O => U_DCT2D_databuf_reg_6_2_FASTCARRY
    );
  U_DCT2D_databuf_reg_6_2_CYAND_1389 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_6_2_CYSELG,
      I1 => U_DCT2D_databuf_reg_6_2_CYSELF,
      O => U_DCT2D_databuf_reg_6_2_CYAND
    );
  U_DCT2D_databuf_reg_6_2_CYMUXFAST_1390 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_2_CYMUXG2,
      IB => U_DCT2D_databuf_reg_6_2_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_6_2_CYAND,
      O => U_DCT2D_databuf_reg_6_2_CYMUXFAST
    );
  U_DCT2D_databuf_reg_6_2_CYMUXG2_1391 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_2_CY0G,
      IB => U_DCT2D_databuf_reg_6_2_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_6_2_CYSELG,
      O => U_DCT2D_databuf_reg_6_2_CYMUXG2
    );
  U_DCT2D_databuf_reg_6_2_CY0G_1392 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_3_Q,
      O => U_DCT2D_databuf_reg_6_2_CY0G
    );
  U_DCT2D_databuf_reg_6_2_CYSELG_1393 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx42273z1,
      O => U_DCT2D_databuf_reg_6_2_CYSELG
    );
  U_DCT2D_databuf_reg_6_2_SRINV_1394 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_6_2_SRINV
    );
  U_DCT2D_databuf_reg_6_2_CLKINV_1395 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_6_2_CLKINV
    );
  U_DCT2D_databuf_reg_6_2_CEINV_1396 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_6_2_CEINV
    );
  U_DCT2D_databuf_reg_6_4_DXMUX_1397 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_4_XORF,
      O => U_DCT2D_databuf_reg_6_4_DXMUX
    );
  U_DCT2D_databuf_reg_6_4_XORF_1398 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_4_CYINIT,
      I1 => U_DCT2D_nx43270z1,
      O => U_DCT2D_databuf_reg_6_4_XORF
    );
  U_DCT2D_databuf_reg_6_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_4_CY0F,
      IB => U_DCT2D_databuf_reg_6_4_CYINIT,
      SEL => U_DCT2D_databuf_reg_6_4_CYSELF,
      O => U_DCT2D_rtlc5_99_sub_43_ix44267z63342_O
    );
  U_DCT2D_databuf_reg_6_4_CYMUXF2_1399 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_4_CY0F,
      IB => U_DCT2D_databuf_reg_6_4_CY0F,
      SEL => U_DCT2D_databuf_reg_6_4_CYSELF,
      O => U_DCT2D_databuf_reg_6_4_CYMUXF2
    );
  U_DCT2D_databuf_reg_6_4_CYINIT_1400 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_99_sub_43_ix43270z63342_O,
      O => U_DCT2D_databuf_reg_6_4_CYINIT
    );
  U_DCT2D_databuf_reg_6_4_CY0F_1401 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_4_Q,
      O => U_DCT2D_databuf_reg_6_4_CY0F
    );
  U_DCT2D_databuf_reg_6_4_CYSELF_1402 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx43270z1,
      O => U_DCT2D_databuf_reg_6_4_CYSELF
    );
  U_DCT2D_databuf_reg_6_4_DYMUX_1403 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_4_XORG,
      O => U_DCT2D_databuf_reg_6_4_DYMUX
    );
  U_DCT2D_databuf_reg_6_4_XORG_1404 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_99_sub_43_ix44267z63342_O,
      I1 => U_DCT2D_nx44267z1,
      O => U_DCT2D_databuf_reg_6_4_XORG
    );
  U_DCT2D_databuf_reg_6_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_4_CYMUXFAST,
      O => U_DCT2D_rtlc5_99_sub_43_ix45264z63342_O
    );
  U_DCT2D_databuf_reg_6_4_FASTCARRY_1405 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_99_sub_43_ix43270z63342_O,
      O => U_DCT2D_databuf_reg_6_4_FASTCARRY
    );
  U_DCT2D_databuf_reg_6_4_CYAND_1406 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_6_4_CYSELG,
      I1 => U_DCT2D_databuf_reg_6_4_CYSELF,
      O => U_DCT2D_databuf_reg_6_4_CYAND
    );
  U_DCT2D_databuf_reg_6_4_CYMUXFAST_1407 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_4_CYMUXG2,
      IB => U_DCT2D_databuf_reg_6_4_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_6_4_CYAND,
      O => U_DCT2D_databuf_reg_6_4_CYMUXFAST
    );
  U_DCT2D_databuf_reg_6_4_CYMUXG2_1408 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_4_CY0G,
      IB => U_DCT2D_databuf_reg_6_4_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_6_4_CYSELG,
      O => U_DCT2D_databuf_reg_6_4_CYMUXG2
    );
  U_DCT2D_databuf_reg_6_4_CY0G_1409 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_5_Q,
      O => U_DCT2D_databuf_reg_6_4_CY0G
    );
  U_DCT2D_databuf_reg_6_4_CYSELG_1410 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx44267z1,
      O => U_DCT2D_databuf_reg_6_4_CYSELG
    );
  U_DCT2D_databuf_reg_6_4_SRINV_1411 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_6_4_SRINV
    );
  U_DCT2D_databuf_reg_6_4_CLKINV_1412 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_6_4_CLKINV
    );
  U_DCT2D_databuf_reg_6_4_CEINV_1413 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_6_4_CEINV
    );
  U_DCT1D_ix64807z1321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_2_Q(5),
      ADR2 => U_DCT1D_latchbuf_reg_5_Q(5),
      ADR3 => VCC,
      O => U_DCT1D_nx64807z1
    );
  U_DCT2D_databuf_reg_6_6_DXMUX_1414 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_6_XORF,
      O => U_DCT2D_databuf_reg_6_6_DXMUX
    );
  U_DCT2D_databuf_reg_6_6_XORF_1415 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_6_CYINIT,
      I1 => U_DCT2D_nx45264z1,
      O => U_DCT2D_databuf_reg_6_6_XORF
    );
  U_DCT2D_databuf_reg_6_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_6_CY0F,
      IB => U_DCT2D_databuf_reg_6_6_CYINIT,
      SEL => U_DCT2D_databuf_reg_6_6_CYSELF,
      O => U_DCT2D_rtlc5_99_sub_43_ix46261z63342_O
    );
  U_DCT2D_databuf_reg_6_6_CYMUXF2_1416 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_6_CY0F,
      IB => U_DCT2D_databuf_reg_6_6_CY0F,
      SEL => U_DCT2D_databuf_reg_6_6_CYSELF,
      O => U_DCT2D_databuf_reg_6_6_CYMUXF2
    );
  U_DCT2D_databuf_reg_6_6_CYINIT_1417 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_99_sub_43_ix45264z63342_O,
      O => U_DCT2D_databuf_reg_6_6_CYINIT
    );
  U_DCT2D_databuf_reg_6_6_CY0F_1418 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_6_Q,
      O => U_DCT2D_databuf_reg_6_6_CY0F
    );
  U_DCT2D_databuf_reg_6_6_CYSELF_1419 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx45264z1,
      O => U_DCT2D_databuf_reg_6_6_CYSELF
    );
  U_DCT2D_databuf_reg_6_6_DYMUX_1420 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_6_XORG,
      O => U_DCT2D_databuf_reg_6_6_DYMUX
    );
  U_DCT2D_databuf_reg_6_6_XORG_1421 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_99_sub_43_ix46261z63342_O,
      I1 => U_DCT2D_nx46261z1,
      O => U_DCT2D_databuf_reg_6_6_XORG
    );
  U_DCT2D_databuf_reg_6_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_6_CYMUXFAST,
      O => U_DCT2D_rtlc5_99_sub_43_ix47258z63342_O
    );
  U_DCT2D_databuf_reg_6_6_FASTCARRY_1422 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_99_sub_43_ix45264z63342_O,
      O => U_DCT2D_databuf_reg_6_6_FASTCARRY
    );
  U_DCT2D_databuf_reg_6_6_CYAND_1423 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_6_6_CYSELG,
      I1 => U_DCT2D_databuf_reg_6_6_CYSELF,
      O => U_DCT2D_databuf_reg_6_6_CYAND
    );
  U_DCT2D_databuf_reg_6_6_CYMUXFAST_1424 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_6_CYMUXG2,
      IB => U_DCT2D_databuf_reg_6_6_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_6_6_CYAND,
      O => U_DCT2D_databuf_reg_6_6_CYMUXFAST
    );
  U_DCT2D_databuf_reg_6_6_CYMUXG2_1425 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_6_CY0G,
      IB => U_DCT2D_databuf_reg_6_6_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_6_6_CYSELG,
      O => U_DCT2D_databuf_reg_6_6_CYMUXG2
    );
  U_DCT2D_databuf_reg_6_6_CY0G_1426 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_7_Q,
      O => U_DCT2D_databuf_reg_6_6_CY0G
    );
  U_DCT2D_databuf_reg_6_6_CYSELG_1427 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx46261z1,
      O => U_DCT2D_databuf_reg_6_6_CYSELG
    );
  U_DCT2D_databuf_reg_6_6_SRINV_1428 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_6_6_SRINV
    );
  U_DCT2D_databuf_reg_6_6_CLKINV_1429 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_6_6_CLKINV
    );
  U_DCT2D_databuf_reg_6_6_CEINV_1430 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_6_6_CEINV
    );
  U_DCT2D_databuf_reg_6_8_DXMUX_1431 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_8_XORF,
      O => U_DCT2D_databuf_reg_6_8_DXMUX
    );
  U_DCT2D_databuf_reg_6_8_XORF_1432 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_8_CYINIT,
      I1 => U_DCT2D_nx47258z1,
      O => U_DCT2D_databuf_reg_6_8_XORF
    );
  U_DCT2D_databuf_reg_6_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_8_CY0F,
      IB => U_DCT2D_databuf_reg_6_8_CYINIT,
      SEL => U_DCT2D_databuf_reg_6_8_CYSELF,
      O => U_DCT2D_rtlc5_99_sub_43_ix48255z63342_O
    );
  U_DCT2D_databuf_reg_6_8_CYMUXF2_1433 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_8_CY0F,
      IB => U_DCT2D_databuf_reg_6_8_CY0F,
      SEL => U_DCT2D_databuf_reg_6_8_CYSELF,
      O => U_DCT2D_databuf_reg_6_8_CYMUXF2
    );
  U_DCT2D_databuf_reg_6_8_CYINIT_1434 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_99_sub_43_ix47258z63342_O,
      O => U_DCT2D_databuf_reg_6_8_CYINIT
    );
  U_DCT2D_databuf_reg_6_8_CY0F_1435 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_8_Q,
      O => U_DCT2D_databuf_reg_6_8_CY0F
    );
  U_DCT2D_databuf_reg_6_8_CYSELF_1436 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx47258z1,
      O => U_DCT2D_databuf_reg_6_8_CYSELF
    );
  U_DCT2D_databuf_reg_6_8_DYMUX_1437 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_8_XORG,
      O => U_DCT2D_databuf_reg_6_8_DYMUX
    );
  U_DCT2D_databuf_reg_6_8_XORG_1438 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_99_sub_43_ix48255z63342_O,
      I1 => U_DCT2D_nx48255z1,
      O => U_DCT2D_databuf_reg_6_8_XORG
    );
  U_DCT2D_databuf_reg_6_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_8_CYMUXFAST,
      O => U_DCT2D_rtlc5_99_sub_43_ix8385z63342_O
    );
  U_DCT2D_databuf_reg_6_8_FASTCARRY_1439 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_99_sub_43_ix47258z63342_O,
      O => U_DCT2D_databuf_reg_6_8_FASTCARRY
    );
  U_DCT2D_databuf_reg_6_8_CYAND_1440 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_6_8_CYSELG,
      I1 => U_DCT2D_databuf_reg_6_8_CYSELF,
      O => U_DCT2D_databuf_reg_6_8_CYAND
    );
  U_DCT2D_databuf_reg_6_8_CYMUXFAST_1441 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_8_CYMUXG2,
      IB => U_DCT2D_databuf_reg_6_8_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_6_8_CYAND,
      O => U_DCT2D_databuf_reg_6_8_CYMUXFAST
    );
  U_DCT2D_databuf_reg_6_8_CYMUXG2_1442 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_6_8_CY0G,
      IB => U_DCT2D_databuf_reg_6_8_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_6_8_CYSELG,
      O => U_DCT2D_databuf_reg_6_8_CYMUXG2
    );
  U_DCT2D_databuf_reg_6_8_CY0G_1443 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_10_Q,
      O => U_DCT2D_databuf_reg_6_8_CY0G
    );
  U_DCT2D_databuf_reg_6_8_CYSELG_1444 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx48255z1,
      O => U_DCT2D_databuf_reg_6_8_CYSELG
    );
  U_DCT2D_databuf_reg_6_8_SRINV_1445 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_6_8_SRINV
    );
  U_DCT2D_databuf_reg_6_8_CLKINV_1446 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_6_8_CLKINV
    );
  U_DCT2D_databuf_reg_6_8_CEINV_1447 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_6_8_CEINV
    );
  U_DCT2D_databuf_reg_6_10_DXMUX_1448 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_10_XORF,
      O => U_DCT2D_databuf_reg_6_10_DXMUX
    );
  U_DCT2D_databuf_reg_6_10_XORF_1449 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_10_CYINIT,
      I1 => U_DCT2D_nx8385z1_rt,
      O => U_DCT2D_databuf_reg_6_10_XORF
    );
  U_DCT2D_databuf_reg_6_10_CYINIT_1450 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_99_sub_43_ix8385z63342_O,
      O => U_DCT2D_databuf_reg_6_10_CYINIT
    );
  U_DCT2D_databuf_reg_6_10_CLKINV_1451 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_6_10_CLKINV
    );
  U_DCT2D_databuf_reg_6_10_CEINV_1452 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_6_10_CEINV
    );
  U_DCT1D_databuf_reg_0_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_0_0_FFX_RST
    );
  U_DCT1D_reg_databuf_reg_0_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_0_0_DXMUX,
      CE => U_DCT1D_databuf_reg_0_0_CEINV,
      CLK => U_DCT1D_databuf_reg_0_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_0_0_FFX_RST,
      O => U_DCT1D_databuf_reg_0_Q(0)
    );
  U_DCT1D_ix60980z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_0_Q(0),
      ADR1 => U_DCT1D_latchbuf_reg_7_Q(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx60980z1
    );
  U_DCT1D_databuf_reg_0_0_DXMUX_1453 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_0_XORF,
      O => U_DCT1D_databuf_reg_0_0_DXMUX
    );
  U_DCT1D_databuf_reg_0_0_XORF_1454 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_0_CYINIT,
      I1 => U_DCT1D_nx60980z1,
      O => U_DCT1D_databuf_reg_0_0_XORF
    );
  U_DCT1D_databuf_reg_0_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_0_CY0F,
      IB => U_DCT1D_databuf_reg_0_0_CYINIT,
      SEL => U_DCT1D_databuf_reg_0_0_CYSELF,
      O => U_DCT1D_rtlc5_1419_add_8_ix59983z63342_O
    );
  U_DCT1D_databuf_reg_0_0_CYINIT_1455 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_0_BXINVNOT,
      O => U_DCT1D_databuf_reg_0_0_CYINIT
    );
  U_DCT1D_databuf_reg_0_0_CY0F_1456 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(0),
      O => U_DCT1D_databuf_reg_0_0_CY0F
    );
  U_DCT1D_databuf_reg_0_0_CYSELF_1457 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx60980z1,
      O => U_DCT1D_databuf_reg_0_0_CYSELF
    );
  U_DCT1D_databuf_reg_0_0_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_5,
      O => U_DCT1D_databuf_reg_0_0_BXINVNOT
    );
  U_DCT1D_databuf_reg_0_0_DYMUX_1458 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_0_XORG,
      O => U_DCT1D_databuf_reg_0_0_DYMUX
    );
  U_DCT1D_databuf_reg_0_0_XORG_1459 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1419_add_8_ix59983z63342_O,
      I1 => U_DCT1D_nx59983z1,
      O => U_DCT1D_databuf_reg_0_0_XORG
    );
  U_DCT1D_databuf_reg_0_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_0_CYMUXG,
      O => U_DCT1D_rtlc5_1419_add_8_ix58986z63342_O
    );
  U_DCT1D_databuf_reg_0_0_CYMUXG_1460 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_0_CY0G,
      IB => U_DCT1D_rtlc5_1419_add_8_ix59983z63342_O,
      SEL => U_DCT1D_databuf_reg_0_0_CYSELG,
      O => U_DCT1D_databuf_reg_0_0_CYMUXG
    );
  U_DCT1D_databuf_reg_0_0_CY0G_1461 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(1),
      O => U_DCT1D_databuf_reg_0_0_CY0G
    );
  U_DCT1D_databuf_reg_0_0_CYSELG_1462 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59983z1,
      O => U_DCT1D_databuf_reg_0_0_CYSELG
    );
  U_DCT1D_databuf_reg_0_0_SRINV_1463 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_0_0_SRINV
    );
  U_DCT1D_databuf_reg_0_0_CLKINV_1464 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_0_0_CLKINV
    );
  U_DCT1D_databuf_reg_0_0_CEINV_1465 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_0_0_CEINV
    );
  U_DCT1D_ix58986z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_0_Q(2),
      ADR1 => U_DCT1D_latchbuf_reg_7_Q(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx58986z1
    );
  U_DCT1D_databuf_reg_0_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_0_2_FFY_RST
    );
  U_DCT1D_reg_databuf_reg_0_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_0_2_DYMUX,
      CE => U_DCT1D_databuf_reg_0_2_CEINV,
      CLK => U_DCT1D_databuf_reg_0_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_0_2_FFY_RST,
      O => U_DCT1D_databuf_reg_0_Q(3)
    );
  U_DCT1D_ix57989z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_7_Q(3),
      ADR1 => U_DCT1D_latchbuf_reg_0_Q(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx57989z1
    );
  U_DCT1D_databuf_reg_0_2_DXMUX_1466 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_2_XORF,
      O => U_DCT1D_databuf_reg_0_2_DXMUX
    );
  U_DCT1D_databuf_reg_0_2_XORF_1467 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_2_CYINIT,
      I1 => U_DCT1D_nx58986z1,
      O => U_DCT1D_databuf_reg_0_2_XORF
    );
  U_DCT1D_databuf_reg_0_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_2_CY0F,
      IB => U_DCT1D_databuf_reg_0_2_CYINIT,
      SEL => U_DCT1D_databuf_reg_0_2_CYSELF,
      O => U_DCT1D_rtlc5_1419_add_8_ix57989z63342_O
    );
  U_DCT1D_databuf_reg_0_2_CYMUXF2_1468 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_2_CY0F,
      IB => U_DCT1D_databuf_reg_0_2_CY0F,
      SEL => U_DCT1D_databuf_reg_0_2_CYSELF,
      O => U_DCT1D_databuf_reg_0_2_CYMUXF2
    );
  U_DCT1D_databuf_reg_0_2_CYINIT_1469 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1419_add_8_ix58986z63342_O,
      O => U_DCT1D_databuf_reg_0_2_CYINIT
    );
  U_DCT1D_databuf_reg_0_2_CY0F_1470 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(2),
      O => U_DCT1D_databuf_reg_0_2_CY0F
    );
  U_DCT1D_databuf_reg_0_2_CYSELF_1471 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx58986z1,
      O => U_DCT1D_databuf_reg_0_2_CYSELF
    );
  U_DCT1D_databuf_reg_0_2_DYMUX_1472 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_2_XORG,
      O => U_DCT1D_databuf_reg_0_2_DYMUX
    );
  U_DCT1D_databuf_reg_0_2_XORG_1473 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1419_add_8_ix57989z63342_O,
      I1 => U_DCT1D_nx57989z1,
      O => U_DCT1D_databuf_reg_0_2_XORG
    );
  U_DCT1D_databuf_reg_0_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_2_CYMUXFAST,
      O => U_DCT1D_rtlc5_1419_add_8_ix56992z63342_O
    );
  U_DCT1D_databuf_reg_0_2_FASTCARRY_1474 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1419_add_8_ix58986z63342_O,
      O => U_DCT1D_databuf_reg_0_2_FASTCARRY
    );
  U_DCT1D_databuf_reg_0_2_CYAND_1475 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_0_2_CYSELG,
      I1 => U_DCT1D_databuf_reg_0_2_CYSELF,
      O => U_DCT1D_databuf_reg_0_2_CYAND
    );
  U_DCT1D_databuf_reg_0_2_CYMUXFAST_1476 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_2_CYMUXG2,
      IB => U_DCT1D_databuf_reg_0_2_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_0_2_CYAND,
      O => U_DCT1D_databuf_reg_0_2_CYMUXFAST
    );
  U_DCT1D_databuf_reg_0_2_CYMUXG2_1477 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_2_CY0G,
      IB => U_DCT1D_databuf_reg_0_2_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_0_2_CYSELG,
      O => U_DCT1D_databuf_reg_0_2_CYMUXG2
    );
  U_DCT1D_databuf_reg_0_2_CY0G_1478 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(3),
      O => U_DCT1D_databuf_reg_0_2_CY0G
    );
  U_DCT1D_databuf_reg_0_2_CYSELG_1479 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx57989z1,
      O => U_DCT1D_databuf_reg_0_2_CYSELG
    );
  U_DCT1D_databuf_reg_0_2_SRINV_1480 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_0_2_SRINV
    );
  U_DCT1D_databuf_reg_0_2_CLKINV_1481 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_0_2_CLKINV
    );
  U_DCT1D_databuf_reg_0_2_CEINV_1482 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_0_2_CEINV
    );
  U_DCT1D_databuf_reg_0_4_DXMUX_1483 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_4_XORF,
      O => U_DCT1D_databuf_reg_0_4_DXMUX
    );
  U_DCT1D_databuf_reg_0_4_XORF_1484 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_4_CYINIT,
      I1 => U_DCT1D_nx56992z1,
      O => U_DCT1D_databuf_reg_0_4_XORF
    );
  U_DCT1D_databuf_reg_0_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_4_CY0F,
      IB => U_DCT1D_databuf_reg_0_4_CYINIT,
      SEL => U_DCT1D_databuf_reg_0_4_CYSELF,
      O => U_DCT1D_rtlc5_1419_add_8_ix55995z63342_O
    );
  U_DCT1D_databuf_reg_0_4_CYMUXF2_1485 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_4_CY0F,
      IB => U_DCT1D_databuf_reg_0_4_CY0F,
      SEL => U_DCT1D_databuf_reg_0_4_CYSELF,
      O => U_DCT1D_databuf_reg_0_4_CYMUXF2
    );
  U_DCT1D_databuf_reg_0_4_CYINIT_1486 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1419_add_8_ix56992z63342_O,
      O => U_DCT1D_databuf_reg_0_4_CYINIT
    );
  U_DCT1D_databuf_reg_0_4_CY0F_1487 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(4),
      O => U_DCT1D_databuf_reg_0_4_CY0F
    );
  U_DCT1D_databuf_reg_0_4_CYSELF_1488 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx56992z1,
      O => U_DCT1D_databuf_reg_0_4_CYSELF
    );
  U_DCT1D_databuf_reg_0_4_DYMUX_1489 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_4_XORG,
      O => U_DCT1D_databuf_reg_0_4_DYMUX
    );
  U_DCT1D_databuf_reg_0_4_XORG_1490 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1419_add_8_ix55995z63342_O,
      I1 => U_DCT1D_nx55995z1,
      O => U_DCT1D_databuf_reg_0_4_XORG
    );
  U_DCT1D_databuf_reg_0_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_4_CYMUXFAST,
      O => U_DCT1D_rtlc5_1419_add_8_ix54998z63342_O
    );
  U_DCT1D_databuf_reg_0_4_FASTCARRY_1491 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1419_add_8_ix56992z63342_O,
      O => U_DCT1D_databuf_reg_0_4_FASTCARRY
    );
  U_DCT1D_databuf_reg_0_4_CYAND_1492 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_0_4_CYSELG,
      I1 => U_DCT1D_databuf_reg_0_4_CYSELF,
      O => U_DCT1D_databuf_reg_0_4_CYAND
    );
  U_DCT1D_databuf_reg_0_4_CYMUXFAST_1493 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_4_CYMUXG2,
      IB => U_DCT1D_databuf_reg_0_4_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_0_4_CYAND,
      O => U_DCT1D_databuf_reg_0_4_CYMUXFAST
    );
  U_DCT1D_databuf_reg_0_4_CYMUXG2_1494 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_4_CY0G,
      IB => U_DCT1D_databuf_reg_0_4_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_0_4_CYSELG,
      O => U_DCT1D_databuf_reg_0_4_CYMUXG2
    );
  U_DCT1D_databuf_reg_0_4_CY0G_1495 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(5),
      O => U_DCT1D_databuf_reg_0_4_CY0G
    );
  U_DCT1D_databuf_reg_0_4_CYSELG_1496 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx55995z1,
      O => U_DCT1D_databuf_reg_0_4_CYSELG
    );
  U_DCT1D_databuf_reg_0_4_SRINV_1497 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_0_4_SRINV
    );
  U_DCT1D_databuf_reg_0_4_CLKINV_1498 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_0_4_CLKINV
    );
  U_DCT1D_databuf_reg_0_4_CEINV_1499 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_0_4_CEINV
    );
  U_DCT1D_databuf_reg_0_6_DXMUX_1500 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_6_XORF,
      O => U_DCT1D_databuf_reg_0_6_DXMUX
    );
  U_DCT1D_databuf_reg_0_6_XORF_1501 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_6_CYINIT,
      I1 => U_DCT1D_nx54998z1,
      O => U_DCT1D_databuf_reg_0_6_XORF
    );
  U_DCT1D_databuf_reg_0_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_6_CY0F,
      IB => U_DCT1D_databuf_reg_0_6_CYINIT,
      SEL => U_DCT1D_databuf_reg_0_6_CYSELF,
      O => U_DCT1D_rtlc5_1419_add_8_ix54001z63342_O
    );
  U_DCT1D_databuf_reg_0_6_CYMUXF2_1502 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_6_CY0F,
      IB => U_DCT1D_databuf_reg_0_6_CY0F,
      SEL => U_DCT1D_databuf_reg_0_6_CYSELF,
      O => U_DCT1D_databuf_reg_0_6_CYMUXF2
    );
  U_DCT1D_databuf_reg_0_6_CYINIT_1503 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1419_add_8_ix54998z63342_O,
      O => U_DCT1D_databuf_reg_0_6_CYINIT
    );
  U_DCT1D_databuf_reg_0_6_CY0F_1504 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(6),
      O => U_DCT1D_databuf_reg_0_6_CY0F
    );
  U_DCT1D_databuf_reg_0_6_CYSELF_1505 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx54998z1,
      O => U_DCT1D_databuf_reg_0_6_CYSELF
    );
  U_DCT1D_databuf_reg_0_6_DYMUX_1506 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_6_XORG,
      O => U_DCT1D_databuf_reg_0_6_DYMUX
    );
  U_DCT1D_databuf_reg_0_6_XORG_1507 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1419_add_8_ix54001z63342_O,
      I1 => U_DCT1D_nx54001z1,
      O => U_DCT1D_databuf_reg_0_6_XORG
    );
  U_DCT1D_databuf_reg_0_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_6_CYMUXFAST,
      O => U_DCT1D_rtlc5_1419_add_8_ix53004z63342_O
    );
  U_DCT1D_databuf_reg_0_6_FASTCARRY_1508 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1419_add_8_ix54998z63342_O,
      O => U_DCT1D_databuf_reg_0_6_FASTCARRY
    );
  U_DCT1D_databuf_reg_0_6_CYAND_1509 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_0_6_CYSELG,
      I1 => U_DCT1D_databuf_reg_0_6_CYSELF,
      O => U_DCT1D_databuf_reg_0_6_CYAND
    );
  U_DCT1D_databuf_reg_0_6_CYMUXFAST_1510 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_6_CYMUXG2,
      IB => U_DCT1D_databuf_reg_0_6_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_0_6_CYAND,
      O => U_DCT1D_databuf_reg_0_6_CYMUXFAST
    );
  U_DCT1D_databuf_reg_0_6_CYMUXG2_1511 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_0_6_CY0G,
      IB => U_DCT1D_databuf_reg_0_6_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_0_6_CYSELG,
      O => U_DCT1D_databuf_reg_0_6_CYMUXG2
    );
  U_DCT1D_databuf_reg_0_6_CY0G_1512 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_Q(7),
      O => U_DCT1D_databuf_reg_0_6_CY0G
    );
  U_DCT1D_databuf_reg_0_6_CYSELG_1513 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx54001z1,
      O => U_DCT1D_databuf_reg_0_6_CYSELG
    );
  U_DCT1D_databuf_reg_0_6_SRINV_1514 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_0_6_SRINV
    );
  U_DCT1D_databuf_reg_0_6_CLKINV_1515 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_0_6_CLKINV
    );
  U_DCT1D_databuf_reg_0_6_CEINV_1516 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_0_6_CEINV
    );
  U_DCT1D_databuf_reg_0_8_DXMUX_1517 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_8_XORF,
      O => U_DCT1D_databuf_reg_0_8_DXMUX
    );
  U_DCT1D_databuf_reg_0_8_XORF_1518 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_8_CYINIT,
      I1 => U_DCT1D_nx53004z1_rt,
      O => U_DCT1D_databuf_reg_0_8_XORF
    );
  U_DCT1D_databuf_reg_0_8_CYINIT_1519 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1419_add_8_ix53004z63342_O,
      O => U_DCT1D_databuf_reg_0_8_CYINIT
    );
  U_DCT1D_databuf_reg_0_8_CLKINV_1520 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_0_8_CLKINV
    );
  U_DCT1D_databuf_reg_0_8_CEINV_1521 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_0_8_CEINV
    );
  U_DCT1D_databuf_reg_5_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_5_0_FFX_RST
    );
  U_DCT1D_reg_databuf_reg_5_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_5_0_DXMUX,
      CE => U_DCT1D_databuf_reg_5_0_CEINV,
      CLK => U_DCT1D_databuf_reg_5_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_5_0_FFX_RST,
      O => U_DCT1D_databuf_reg_5_Q(0)
    );
  U_DCT1D_ix44417z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_6_Q(0),
      ADR1 => U_DCT1D_latchbuf_reg_1_Q(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx44417z1
    );
  U_DCT1D_databuf_reg_5_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_5_0_FFY_RST
    );
  U_DCT1D_reg_databuf_reg_5_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_5_0_DYMUX,
      CE => U_DCT1D_databuf_reg_5_0_CEINV,
      CLK => U_DCT1D_databuf_reg_5_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_5_0_FFY_RST,
      O => U_DCT1D_databuf_reg_5_Q(1)
    );
  U_DCT1D_databuf_reg_5_0_DXMUX_1522 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_0_XORF,
      O => U_DCT1D_databuf_reg_5_0_DXMUX
    );
  U_DCT1D_databuf_reg_5_0_XORF_1523 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_0_CYINIT,
      I1 => U_DCT1D_nx44417z1,
      O => U_DCT1D_databuf_reg_5_0_XORF
    );
  U_DCT1D_databuf_reg_5_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_0_CY0F,
      IB => U_DCT1D_databuf_reg_5_0_CYINIT,
      SEL => U_DCT1D_databuf_reg_5_0_CYSELF,
      O => U_DCT1D_rtlc5_84_sub_5_ix45414z63342_O
    );
  U_DCT1D_databuf_reg_5_0_CYINIT_1524 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GLOBAL_LOGIC1_8,
      O => U_DCT1D_databuf_reg_5_0_CYINIT
    );
  U_DCT1D_databuf_reg_5_0_CY0F_1525 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(0),
      O => U_DCT1D_databuf_reg_5_0_CY0F
    );
  U_DCT1D_databuf_reg_5_0_CYSELF_1526 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx44417z1,
      O => U_DCT1D_databuf_reg_5_0_CYSELF
    );
  U_DCT1D_databuf_reg_5_0_DYMUX_1527 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_0_XORG,
      O => U_DCT1D_databuf_reg_5_0_DYMUX
    );
  U_DCT1D_databuf_reg_5_0_XORG_1528 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_84_sub_5_ix45414z63342_O,
      I1 => U_DCT1D_nx45414z1,
      O => U_DCT1D_databuf_reg_5_0_XORG
    );
  U_DCT1D_databuf_reg_5_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_0_CYMUXG,
      O => U_DCT1D_rtlc5_84_sub_5_ix46411z63342_O
    );
  U_DCT1D_databuf_reg_5_0_CYMUXG_1529 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_0_CY0G,
      IB => U_DCT1D_rtlc5_84_sub_5_ix45414z63342_O,
      SEL => U_DCT1D_databuf_reg_5_0_CYSELG,
      O => U_DCT1D_databuf_reg_5_0_CYMUXG
    );
  U_DCT1D_databuf_reg_5_0_CY0G_1530 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(1),
      O => U_DCT1D_databuf_reg_5_0_CY0G
    );
  U_DCT1D_databuf_reg_5_0_CYSELG_1531 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx45414z1,
      O => U_DCT1D_databuf_reg_5_0_CYSELG
    );
  U_DCT1D_databuf_reg_5_0_SRINV_1532 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_5_0_SRINV
    );
  U_DCT1D_databuf_reg_5_0_CLKINV_1533 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_5_0_CLKINV
    );
  U_DCT1D_databuf_reg_5_0_CEINV_1534 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_5_0_CEINV
    );
  U_DCT1D_databuf_reg_5_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_5_2_FFY_RST
    );
  U_DCT1D_reg_databuf_reg_5_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_5_2_DYMUX,
      CE => U_DCT1D_databuf_reg_5_2_CEINV,
      CLK => U_DCT1D_databuf_reg_5_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_5_2_FFY_RST,
      O => U_DCT1D_databuf_reg_5_Q(3)
    );
  U_DCT1D_ix47408z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_1_Q(3),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_6_Q(3),
      ADR3 => VCC,
      O => U_DCT1D_nx47408z1
    );
  U_DCT1D_databuf_reg_5_2_DXMUX_1535 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_2_XORF,
      O => U_DCT1D_databuf_reg_5_2_DXMUX
    );
  U_DCT1D_databuf_reg_5_2_XORF_1536 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_2_CYINIT,
      I1 => U_DCT1D_nx46411z1,
      O => U_DCT1D_databuf_reg_5_2_XORF
    );
  U_DCT1D_databuf_reg_5_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_2_CY0F,
      IB => U_DCT1D_databuf_reg_5_2_CYINIT,
      SEL => U_DCT1D_databuf_reg_5_2_CYSELF,
      O => U_DCT1D_rtlc5_84_sub_5_ix47408z63342_O
    );
  U_DCT1D_databuf_reg_5_2_CYMUXF2_1537 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_2_CY0F,
      IB => U_DCT1D_databuf_reg_5_2_CY0F,
      SEL => U_DCT1D_databuf_reg_5_2_CYSELF,
      O => U_DCT1D_databuf_reg_5_2_CYMUXF2
    );
  U_DCT1D_databuf_reg_5_2_CYINIT_1538 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_84_sub_5_ix46411z63342_O,
      O => U_DCT1D_databuf_reg_5_2_CYINIT
    );
  U_DCT1D_databuf_reg_5_2_CY0F_1539 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(2),
      O => U_DCT1D_databuf_reg_5_2_CY0F
    );
  U_DCT1D_databuf_reg_5_2_CYSELF_1540 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx46411z1,
      O => U_DCT1D_databuf_reg_5_2_CYSELF
    );
  U_DCT1D_databuf_reg_5_2_DYMUX_1541 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_2_XORG,
      O => U_DCT1D_databuf_reg_5_2_DYMUX
    );
  U_DCT1D_databuf_reg_5_2_XORG_1542 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_84_sub_5_ix47408z63342_O,
      I1 => U_DCT1D_nx47408z1,
      O => U_DCT1D_databuf_reg_5_2_XORG
    );
  U_DCT1D_databuf_reg_5_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_2_CYMUXFAST,
      O => U_DCT1D_rtlc5_84_sub_5_ix48405z63342_O
    );
  U_DCT1D_databuf_reg_5_2_FASTCARRY_1543 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_84_sub_5_ix46411z63342_O,
      O => U_DCT1D_databuf_reg_5_2_FASTCARRY
    );
  U_DCT1D_databuf_reg_5_2_CYAND_1544 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_5_2_CYSELG,
      I1 => U_DCT1D_databuf_reg_5_2_CYSELF,
      O => U_DCT1D_databuf_reg_5_2_CYAND
    );
  U_DCT1D_databuf_reg_5_2_CYMUXFAST_1545 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_2_CYMUXG2,
      IB => U_DCT1D_databuf_reg_5_2_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_5_2_CYAND,
      O => U_DCT1D_databuf_reg_5_2_CYMUXFAST
    );
  U_DCT1D_databuf_reg_5_2_CYMUXG2_1546 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_2_CY0G,
      IB => U_DCT1D_databuf_reg_5_2_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_5_2_CYSELG,
      O => U_DCT1D_databuf_reg_5_2_CYMUXG2
    );
  U_DCT1D_databuf_reg_5_2_CY0G_1547 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(3),
      O => U_DCT1D_databuf_reg_5_2_CY0G
    );
  U_DCT1D_databuf_reg_5_2_CYSELG_1548 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx47408z1,
      O => U_DCT1D_databuf_reg_5_2_CYSELG
    );
  U_DCT1D_databuf_reg_5_2_SRINV_1549 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_5_2_SRINV
    );
  U_DCT1D_databuf_reg_5_2_CLKINV_1550 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_5_2_CLKINV
    );
  U_DCT1D_databuf_reg_5_2_CEINV_1551 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_5_2_CEINV
    );
  U_DCT1D_databuf_reg_5_4_DXMUX_1552 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_4_XORF,
      O => U_DCT1D_databuf_reg_5_4_DXMUX
    );
  U_DCT1D_databuf_reg_5_4_XORF_1553 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_4_CYINIT,
      I1 => U_DCT1D_nx48405z1,
      O => U_DCT1D_databuf_reg_5_4_XORF
    );
  U_DCT1D_databuf_reg_5_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_4_CY0F,
      IB => U_DCT1D_databuf_reg_5_4_CYINIT,
      SEL => U_DCT1D_databuf_reg_5_4_CYSELF,
      O => U_DCT1D_rtlc5_84_sub_5_ix49402z63342_O
    );
  U_DCT1D_databuf_reg_5_4_CYMUXF2_1554 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_4_CY0F,
      IB => U_DCT1D_databuf_reg_5_4_CY0F,
      SEL => U_DCT1D_databuf_reg_5_4_CYSELF,
      O => U_DCT1D_databuf_reg_5_4_CYMUXF2
    );
  U_DCT1D_databuf_reg_5_4_CYINIT_1555 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_84_sub_5_ix48405z63342_O,
      O => U_DCT1D_databuf_reg_5_4_CYINIT
    );
  U_DCT1D_databuf_reg_5_4_CY0F_1556 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(4),
      O => U_DCT1D_databuf_reg_5_4_CY0F
    );
  U_DCT1D_databuf_reg_5_4_CYSELF_1557 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx48405z1,
      O => U_DCT1D_databuf_reg_5_4_CYSELF
    );
  U_DCT1D_databuf_reg_5_4_DYMUX_1558 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_4_XORG,
      O => U_DCT1D_databuf_reg_5_4_DYMUX
    );
  U_DCT1D_databuf_reg_5_4_XORG_1559 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_84_sub_5_ix49402z63342_O,
      I1 => U_DCT1D_nx49402z1,
      O => U_DCT1D_databuf_reg_5_4_XORG
    );
  U_DCT1D_databuf_reg_5_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_4_CYMUXFAST,
      O => U_DCT1D_rtlc5_84_sub_5_ix50399z63342_O
    );
  U_DCT1D_databuf_reg_5_4_FASTCARRY_1560 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_84_sub_5_ix48405z63342_O,
      O => U_DCT1D_databuf_reg_5_4_FASTCARRY
    );
  U_DCT1D_databuf_reg_5_4_CYAND_1561 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_5_4_CYSELG,
      I1 => U_DCT1D_databuf_reg_5_4_CYSELF,
      O => U_DCT1D_databuf_reg_5_4_CYAND
    );
  U_DCT1D_databuf_reg_5_4_CYMUXFAST_1562 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_4_CYMUXG2,
      IB => U_DCT1D_databuf_reg_5_4_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_5_4_CYAND,
      O => U_DCT1D_databuf_reg_5_4_CYMUXFAST
    );
  U_DCT1D_databuf_reg_5_4_CYMUXG2_1563 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_4_CY0G,
      IB => U_DCT1D_databuf_reg_5_4_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_5_4_CYSELG,
      O => U_DCT1D_databuf_reg_5_4_CYMUXG2
    );
  U_DCT1D_databuf_reg_5_4_CY0G_1564 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(5),
      O => U_DCT1D_databuf_reg_5_4_CY0G
    );
  U_DCT1D_databuf_reg_5_4_CYSELG_1565 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx49402z1,
      O => U_DCT1D_databuf_reg_5_4_CYSELG
    );
  U_DCT1D_databuf_reg_5_4_SRINV_1566 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_5_4_SRINV
    );
  U_DCT1D_databuf_reg_5_4_CLKINV_1567 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_5_4_CLKINV
    );
  U_DCT1D_databuf_reg_5_4_CEINV_1568 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_5_4_CEINV
    );
  U_DCT1D_databuf_reg_5_6_DXMUX_1569 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_6_XORF,
      O => U_DCT1D_databuf_reg_5_6_DXMUX
    );
  U_DCT1D_databuf_reg_5_6_XORF_1570 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_6_CYINIT,
      I1 => U_DCT1D_nx50399z1,
      O => U_DCT1D_databuf_reg_5_6_XORF
    );
  U_DCT1D_databuf_reg_5_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_6_CY0F,
      IB => U_DCT1D_databuf_reg_5_6_CYINIT,
      SEL => U_DCT1D_databuf_reg_5_6_CYSELF,
      O => U_DCT1D_rtlc5_84_sub_5_ix51396z63342_O
    );
  U_DCT1D_databuf_reg_5_6_CYMUXF2_1571 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_6_CY0F,
      IB => U_DCT1D_databuf_reg_5_6_CY0F,
      SEL => U_DCT1D_databuf_reg_5_6_CYSELF,
      O => U_DCT1D_databuf_reg_5_6_CYMUXF2
    );
  U_DCT1D_databuf_reg_5_6_CYINIT_1572 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_84_sub_5_ix50399z63342_O,
      O => U_DCT1D_databuf_reg_5_6_CYINIT
    );
  U_DCT1D_databuf_reg_5_6_CY0F_1573 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(6),
      O => U_DCT1D_databuf_reg_5_6_CY0F
    );
  U_DCT1D_databuf_reg_5_6_CYSELF_1574 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx50399z1,
      O => U_DCT1D_databuf_reg_5_6_CYSELF
    );
  U_DCT1D_databuf_reg_5_6_DYMUX_1575 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_6_XORG,
      O => U_DCT1D_databuf_reg_5_6_DYMUX
    );
  U_DCT1D_databuf_reg_5_6_XORG_1576 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_84_sub_5_ix51396z63342_O,
      I1 => U_DCT1D_nx51396z1,
      O => U_DCT1D_databuf_reg_5_6_XORG
    );
  U_DCT1D_databuf_reg_5_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_6_CYMUXFAST,
      O => U_DCT1D_rtlc5_84_sub_5_ix52393z63342_O
    );
  U_DCT1D_databuf_reg_5_6_FASTCARRY_1577 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_84_sub_5_ix50399z63342_O,
      O => U_DCT1D_databuf_reg_5_6_FASTCARRY
    );
  U_DCT1D_databuf_reg_5_6_CYAND_1578 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_5_6_CYSELG,
      I1 => U_DCT1D_databuf_reg_5_6_CYSELF,
      O => U_DCT1D_databuf_reg_5_6_CYAND
    );
  U_DCT1D_databuf_reg_5_6_CYMUXFAST_1579 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_6_CYMUXG2,
      IB => U_DCT1D_databuf_reg_5_6_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_5_6_CYAND,
      O => U_DCT1D_databuf_reg_5_6_CYMUXFAST
    );
  U_DCT1D_databuf_reg_5_6_CYMUXG2_1580 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_5_6_CY0G,
      IB => U_DCT1D_databuf_reg_5_6_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_5_6_CYSELG,
      O => U_DCT1D_databuf_reg_5_6_CYMUXG2
    );
  U_DCT1D_databuf_reg_5_6_CY0G_1581 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(7),
      O => U_DCT1D_databuf_reg_5_6_CY0G
    );
  U_DCT1D_databuf_reg_5_6_CYSELG_1582 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx51396z1,
      O => U_DCT1D_databuf_reg_5_6_CYSELG
    );
  U_DCT1D_databuf_reg_5_6_SRINV_1583 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_5_6_SRINV
    );
  U_DCT1D_databuf_reg_5_6_CLKINV_1584 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_5_6_CLKINV
    );
  U_DCT1D_databuf_reg_5_6_CEINV_1585 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_5_6_CEINV
    );
  U_DCT1D_databuf_reg_5_8_DXMUX_1586 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_8_XORF,
      O => U_DCT1D_databuf_reg_5_8_DXMUX
    );
  U_DCT1D_databuf_reg_5_8_XORF_1587 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_8_CYINIT,
      I1 => U_DCT1D_nx52393z1_rt,
      O => U_DCT1D_databuf_reg_5_8_XORF
    );
  U_DCT1D_databuf_reg_5_8_CYINIT_1588 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_84_sub_5_ix52393z63342_O,
      O => U_DCT1D_databuf_reg_5_8_CYINIT
    );
  U_DCT1D_databuf_reg_5_8_CLKINV_1589 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_5_8_CLKINV
    );
  U_DCT1D_databuf_reg_5_8_CEINV_1590 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_5_8_CEINV
    );
  U_DCT2D_databuf_reg_5_0_DXMUX_1591 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_0_XORF,
      O => U_DCT2D_databuf_reg_5_0_DXMUX
    );
  U_DCT2D_databuf_reg_5_0_XORF_1592 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_0_CYINIT,
      I1 => U_DCT2D_nx44417z1,
      O => U_DCT2D_databuf_reg_5_0_XORF
    );
  U_DCT2D_databuf_reg_5_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_0_CY0F,
      IB => U_DCT2D_databuf_reg_5_0_CYINIT,
      SEL => U_DCT2D_databuf_reg_5_0_CYSELF,
      O => U_DCT2D_rtlc5_98_sub_42_ix45414z63342_O
    );
  U_DCT2D_databuf_reg_5_0_CYINIT_1593 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GLOBAL_LOGIC1_25,
      O => U_DCT2D_databuf_reg_5_0_CYINIT
    );
  U_DCT2D_databuf_reg_5_0_CY0F_1594 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_0_Q,
      O => U_DCT2D_databuf_reg_5_0_CY0F
    );
  U_DCT2D_databuf_reg_5_0_CYSELF_1595 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx44417z1,
      O => U_DCT2D_databuf_reg_5_0_CYSELF
    );
  U_DCT2D_databuf_reg_5_0_DYMUX_1596 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_0_XORG,
      O => U_DCT2D_databuf_reg_5_0_DYMUX
    );
  U_DCT2D_databuf_reg_5_0_XORG_1597 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_98_sub_42_ix45414z63342_O,
      I1 => U_DCT2D_nx45414z1,
      O => U_DCT2D_databuf_reg_5_0_XORG
    );
  U_DCT2D_databuf_reg_5_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_0_CYMUXG,
      O => U_DCT2D_rtlc5_98_sub_42_ix46411z63342_O
    );
  U_DCT2D_databuf_reg_5_0_CYMUXG_1598 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_0_CY0G,
      IB => U_DCT2D_rtlc5_98_sub_42_ix45414z63342_O,
      SEL => U_DCT2D_databuf_reg_5_0_CYSELG,
      O => U_DCT2D_databuf_reg_5_0_CYMUXG
    );
  U_DCT2D_databuf_reg_5_0_CY0G_1599 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_1_Q,
      O => U_DCT2D_databuf_reg_5_0_CY0G
    );
  U_DCT2D_databuf_reg_5_0_CYSELG_1600 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx45414z1,
      O => U_DCT2D_databuf_reg_5_0_CYSELG
    );
  U_DCT2D_databuf_reg_5_0_SRINV_1601 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_5_0_SRINV
    );
  U_DCT2D_databuf_reg_5_0_CLKINV_1602 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_5_0_CLKINV
    );
  U_DCT2D_databuf_reg_5_0_CEINV_1603 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_5_0_CEINV
    );
  U_DCT2D_databuf_reg_5_2_DXMUX_1604 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_2_XORF,
      O => U_DCT2D_databuf_reg_5_2_DXMUX
    );
  U_DCT2D_databuf_reg_5_2_XORF_1605 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_2_CYINIT,
      I1 => U_DCT2D_nx46411z1,
      O => U_DCT2D_databuf_reg_5_2_XORF
    );
  U_DCT2D_databuf_reg_5_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_2_CY0F,
      IB => U_DCT2D_databuf_reg_5_2_CYINIT,
      SEL => U_DCT2D_databuf_reg_5_2_CYSELF,
      O => U_DCT2D_rtlc5_98_sub_42_ix47408z63342_O
    );
  U_DCT2D_databuf_reg_5_2_CYMUXF2_1606 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_2_CY0F,
      IB => U_DCT2D_databuf_reg_5_2_CY0F,
      SEL => U_DCT2D_databuf_reg_5_2_CYSELF,
      O => U_DCT2D_databuf_reg_5_2_CYMUXF2
    );
  U_DCT2D_databuf_reg_5_2_CYINIT_1607 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_98_sub_42_ix46411z63342_O,
      O => U_DCT2D_databuf_reg_5_2_CYINIT
    );
  U_DCT2D_databuf_reg_5_2_CY0F_1608 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_2_Q,
      O => U_DCT2D_databuf_reg_5_2_CY0F
    );
  U_DCT2D_databuf_reg_5_2_CYSELF_1609 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx46411z1,
      O => U_DCT2D_databuf_reg_5_2_CYSELF
    );
  U_DCT2D_databuf_reg_5_2_DYMUX_1610 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_2_XORG,
      O => U_DCT2D_databuf_reg_5_2_DYMUX
    );
  U_DCT2D_databuf_reg_5_2_XORG_1611 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_98_sub_42_ix47408z63342_O,
      I1 => U_DCT2D_nx47408z1,
      O => U_DCT2D_databuf_reg_5_2_XORG
    );
  U_DCT2D_databuf_reg_5_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_2_CYMUXFAST,
      O => U_DCT2D_rtlc5_98_sub_42_ix48405z63342_O
    );
  U_DCT2D_databuf_reg_5_2_FASTCARRY_1612 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_98_sub_42_ix46411z63342_O,
      O => U_DCT2D_databuf_reg_5_2_FASTCARRY
    );
  U_DCT2D_databuf_reg_5_2_CYAND_1613 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_5_2_CYSELG,
      I1 => U_DCT2D_databuf_reg_5_2_CYSELF,
      O => U_DCT2D_databuf_reg_5_2_CYAND
    );
  U_DCT2D_databuf_reg_5_2_CYMUXFAST_1614 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_2_CYMUXG2,
      IB => U_DCT2D_databuf_reg_5_2_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_5_2_CYAND,
      O => U_DCT2D_databuf_reg_5_2_CYMUXFAST
    );
  U_DCT2D_databuf_reg_5_2_CYMUXG2_1615 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_2_CY0G,
      IB => U_DCT2D_databuf_reg_5_2_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_5_2_CYSELG,
      O => U_DCT2D_databuf_reg_5_2_CYMUXG2
    );
  U_DCT2D_databuf_reg_5_2_CY0G_1616 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_3_Q,
      O => U_DCT2D_databuf_reg_5_2_CY0G
    );
  U_DCT2D_databuf_reg_5_2_CYSELG_1617 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx47408z1,
      O => U_DCT2D_databuf_reg_5_2_CYSELG
    );
  U_DCT2D_databuf_reg_5_2_SRINV_1618 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_5_2_SRINV
    );
  U_DCT2D_databuf_reg_5_2_CLKINV_1619 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_5_2_CLKINV
    );
  U_DCT2D_databuf_reg_5_2_CEINV_1620 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_5_2_CEINV
    );
  U_DCT2D_databuf_reg_5_4_DXMUX_1621 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_4_XORF,
      O => U_DCT2D_databuf_reg_5_4_DXMUX
    );
  U_DCT2D_databuf_reg_5_4_XORF_1622 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_4_CYINIT,
      I1 => U_DCT2D_nx48405z1,
      O => U_DCT2D_databuf_reg_5_4_XORF
    );
  U_DCT2D_databuf_reg_5_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_4_CY0F,
      IB => U_DCT2D_databuf_reg_5_4_CYINIT,
      SEL => U_DCT2D_databuf_reg_5_4_CYSELF,
      O => U_DCT2D_rtlc5_98_sub_42_ix49402z63342_O
    );
  U_DCT2D_databuf_reg_5_4_CYMUXF2_1623 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_4_CY0F,
      IB => U_DCT2D_databuf_reg_5_4_CY0F,
      SEL => U_DCT2D_databuf_reg_5_4_CYSELF,
      O => U_DCT2D_databuf_reg_5_4_CYMUXF2
    );
  U_DCT2D_databuf_reg_5_4_CYINIT_1624 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_98_sub_42_ix48405z63342_O,
      O => U_DCT2D_databuf_reg_5_4_CYINIT
    );
  U_DCT2D_databuf_reg_5_4_CY0F_1625 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_4_Q,
      O => U_DCT2D_databuf_reg_5_4_CY0F
    );
  U_DCT2D_databuf_reg_5_4_CYSELF_1626 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx48405z1,
      O => U_DCT2D_databuf_reg_5_4_CYSELF
    );
  U_DCT2D_databuf_reg_5_4_DYMUX_1627 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_4_XORG,
      O => U_DCT2D_databuf_reg_5_4_DYMUX
    );
  U_DCT2D_databuf_reg_5_4_XORG_1628 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_98_sub_42_ix49402z63342_O,
      I1 => U_DCT2D_nx49402z1,
      O => U_DCT2D_databuf_reg_5_4_XORG
    );
  U_DCT2D_databuf_reg_5_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_4_CYMUXFAST,
      O => U_DCT2D_rtlc5_98_sub_42_ix50399z63342_O
    );
  U_DCT2D_databuf_reg_5_4_FASTCARRY_1629 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_98_sub_42_ix48405z63342_O,
      O => U_DCT2D_databuf_reg_5_4_FASTCARRY
    );
  U_DCT2D_databuf_reg_5_4_CYAND_1630 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_5_4_CYSELG,
      I1 => U_DCT2D_databuf_reg_5_4_CYSELF,
      O => U_DCT2D_databuf_reg_5_4_CYAND
    );
  U_DCT2D_databuf_reg_5_4_CYMUXFAST_1631 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_4_CYMUXG2,
      IB => U_DCT2D_databuf_reg_5_4_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_5_4_CYAND,
      O => U_DCT2D_databuf_reg_5_4_CYMUXFAST
    );
  U_DCT2D_databuf_reg_5_4_CYMUXG2_1632 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_4_CY0G,
      IB => U_DCT2D_databuf_reg_5_4_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_5_4_CYSELG,
      O => U_DCT2D_databuf_reg_5_4_CYMUXG2
    );
  U_DCT2D_databuf_reg_5_4_CY0G_1633 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_5_Q,
      O => U_DCT2D_databuf_reg_5_4_CY0G
    );
  U_DCT2D_databuf_reg_5_4_CYSELG_1634 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx49402z1,
      O => U_DCT2D_databuf_reg_5_4_CYSELG
    );
  U_DCT2D_databuf_reg_5_4_SRINV_1635 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_5_4_SRINV
    );
  U_DCT2D_databuf_reg_5_4_CLKINV_1636 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_5_4_CLKINV
    );
  U_DCT2D_databuf_reg_5_4_CEINV_1637 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_5_4_CEINV
    );
  U_DCT2D_databuf_reg_5_6_DXMUX_1638 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_6_XORF,
      O => U_DCT2D_databuf_reg_5_6_DXMUX
    );
  U_DCT2D_databuf_reg_5_6_XORF_1639 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_6_CYINIT,
      I1 => U_DCT2D_nx50399z1,
      O => U_DCT2D_databuf_reg_5_6_XORF
    );
  U_DCT2D_databuf_reg_5_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_6_CY0F,
      IB => U_DCT2D_databuf_reg_5_6_CYINIT,
      SEL => U_DCT2D_databuf_reg_5_6_CYSELF,
      O => U_DCT2D_rtlc5_98_sub_42_ix51396z63342_O
    );
  U_DCT2D_databuf_reg_5_6_CYMUXF2_1640 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_6_CY0F,
      IB => U_DCT2D_databuf_reg_5_6_CY0F,
      SEL => U_DCT2D_databuf_reg_5_6_CYSELF,
      O => U_DCT2D_databuf_reg_5_6_CYMUXF2
    );
  U_DCT2D_databuf_reg_5_6_CYINIT_1641 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_98_sub_42_ix50399z63342_O,
      O => U_DCT2D_databuf_reg_5_6_CYINIT
    );
  U_DCT2D_databuf_reg_5_6_CY0F_1642 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_6_Q,
      O => U_DCT2D_databuf_reg_5_6_CY0F
    );
  U_DCT2D_databuf_reg_5_6_CYSELF_1643 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx50399z1,
      O => U_DCT2D_databuf_reg_5_6_CYSELF
    );
  U_DCT2D_databuf_reg_5_6_DYMUX_1644 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_6_XORG,
      O => U_DCT2D_databuf_reg_5_6_DYMUX
    );
  U_DCT2D_databuf_reg_5_6_XORG_1645 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_98_sub_42_ix51396z63342_O,
      I1 => U_DCT2D_nx51396z1,
      O => U_DCT2D_databuf_reg_5_6_XORG
    );
  U_DCT2D_databuf_reg_5_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_6_CYMUXFAST,
      O => U_DCT2D_rtlc5_98_sub_42_ix52393z63342_O
    );
  U_DCT2D_databuf_reg_5_6_FASTCARRY_1646 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_98_sub_42_ix50399z63342_O,
      O => U_DCT2D_databuf_reg_5_6_FASTCARRY
    );
  U_DCT2D_databuf_reg_5_6_CYAND_1647 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_5_6_CYSELG,
      I1 => U_DCT2D_databuf_reg_5_6_CYSELF,
      O => U_DCT2D_databuf_reg_5_6_CYAND
    );
  U_DCT2D_databuf_reg_5_6_CYMUXFAST_1648 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_6_CYMUXG2,
      IB => U_DCT2D_databuf_reg_5_6_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_5_6_CYAND,
      O => U_DCT2D_databuf_reg_5_6_CYMUXFAST
    );
  U_DCT2D_databuf_reg_5_6_CYMUXG2_1649 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_6_CY0G,
      IB => U_DCT2D_databuf_reg_5_6_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_5_6_CYSELG,
      O => U_DCT2D_databuf_reg_5_6_CYMUXG2
    );
  U_DCT2D_databuf_reg_5_6_CY0G_1650 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_7_Q,
      O => U_DCT2D_databuf_reg_5_6_CY0G
    );
  U_DCT2D_databuf_reg_5_6_CYSELG_1651 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx51396z1,
      O => U_DCT2D_databuf_reg_5_6_CYSELG
    );
  U_DCT2D_databuf_reg_5_6_SRINV_1652 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_5_6_SRINV
    );
  U_DCT2D_databuf_reg_5_6_CLKINV_1653 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_5_6_CLKINV
    );
  U_DCT2D_databuf_reg_5_6_CEINV_1654 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_5_6_CEINV
    );
  U_DCT2D_databuf_reg_5_8_DXMUX_1655 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_8_XORF,
      O => U_DCT2D_databuf_reg_5_8_DXMUX
    );
  U_DCT2D_databuf_reg_5_8_XORF_1656 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_8_CYINIT,
      I1 => U_DCT2D_nx52393z1,
      O => U_DCT2D_databuf_reg_5_8_XORF
    );
  U_DCT2D_databuf_reg_5_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_8_CY0F,
      IB => U_DCT2D_databuf_reg_5_8_CYINIT,
      SEL => U_DCT2D_databuf_reg_5_8_CYSELF,
      O => U_DCT2D_rtlc5_98_sub_42_ix53390z63342_O
    );
  U_DCT2D_databuf_reg_5_8_CYMUXF2_1657 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_8_CY0F,
      IB => U_DCT2D_databuf_reg_5_8_CY0F,
      SEL => U_DCT2D_databuf_reg_5_8_CYSELF,
      O => U_DCT2D_databuf_reg_5_8_CYMUXF2
    );
  U_DCT2D_databuf_reg_5_8_CYINIT_1658 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_98_sub_42_ix52393z63342_O,
      O => U_DCT2D_databuf_reg_5_8_CYINIT
    );
  U_DCT2D_databuf_reg_5_8_CY0F_1659 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_8_Q,
      O => U_DCT2D_databuf_reg_5_8_CY0F
    );
  U_DCT2D_databuf_reg_5_8_CYSELF_1660 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx52393z1,
      O => U_DCT2D_databuf_reg_5_8_CYSELF
    );
  U_DCT2D_databuf_reg_5_8_DYMUX_1661 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_8_XORG,
      O => U_DCT2D_databuf_reg_5_8_DYMUX
    );
  U_DCT2D_databuf_reg_5_8_XORG_1662 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5_98_sub_42_ix53390z63342_O,
      I1 => U_DCT2D_nx53390z1,
      O => U_DCT2D_databuf_reg_5_8_XORG
    );
  U_DCT2D_databuf_reg_5_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_8_CYMUXFAST,
      O => U_DCT2D_rtlc5_98_sub_42_ix64938z63342_O
    );
  U_DCT2D_databuf_reg_5_8_FASTCARRY_1663 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_98_sub_42_ix52393z63342_O,
      O => U_DCT2D_databuf_reg_5_8_FASTCARRY
    );
  U_DCT2D_databuf_reg_5_8_CYAND_1664 : X_AND2
    port map (
      I0 => U_DCT2D_databuf_reg_5_8_CYSELG,
      I1 => U_DCT2D_databuf_reg_5_8_CYSELF,
      O => U_DCT2D_databuf_reg_5_8_CYAND
    );
  U_DCT2D_databuf_reg_5_8_CYMUXFAST_1665 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_8_CYMUXG2,
      IB => U_DCT2D_databuf_reg_5_8_FASTCARRY,
      SEL => U_DCT2D_databuf_reg_5_8_CYAND,
      O => U_DCT2D_databuf_reg_5_8_CYMUXFAST
    );
  U_DCT2D_databuf_reg_5_8_CYMUXG2_1666 : X_MUX2
    port map (
      IA => U_DCT2D_databuf_reg_5_8_CY0G,
      IB => U_DCT2D_databuf_reg_5_8_CYMUXF2,
      SEL => U_DCT2D_databuf_reg_5_8_CYSELG,
      O => U_DCT2D_databuf_reg_5_8_CYMUXG2
    );
  U_DCT2D_databuf_reg_5_8_CY0G_1667 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_10_Q,
      O => U_DCT2D_databuf_reg_5_8_CY0G
    );
  U_DCT2D_databuf_reg_5_8_CYSELG_1668 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx53390z1,
      O => U_DCT2D_databuf_reg_5_8_CYSELG
    );
  U_DCT2D_databuf_reg_5_8_SRINV_1669 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_5_8_SRINV
    );
  U_DCT2D_databuf_reg_5_8_CLKINV_1670 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_5_8_CLKINV
    );
  U_DCT2D_databuf_reg_5_8_CEINV_1671 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_5_8_CEINV
    );
  U_DCT2D_databuf_reg_5_10_DXMUX_1672 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_10_XORF,
      O => U_DCT2D_databuf_reg_5_10_DXMUX
    );
  U_DCT2D_databuf_reg_5_10_XORF_1673 : X_XOR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_10_CYINIT,
      I1 => U_DCT2D_nx64938z1_rt,
      O => U_DCT2D_databuf_reg_5_10_XORF
    );
  U_DCT2D_databuf_reg_5_10_CYINIT_1674 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_98_sub_42_ix64938z63342_O,
      O => U_DCT2D_databuf_reg_5_10_CYINIT
    );
  U_DCT2D_databuf_reg_5_10_CLKINV_1675 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_databuf_reg_5_10_CLKINV
    );
  U_DCT2D_databuf_reg_5_10_CEINV_1676 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702,
      O => U_DCT2D_databuf_reg_5_10_CEINV
    );
  U_DCT1D_databuf_reg_3_0_DXMUX_1677 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_0_XORF,
      O => U_DCT1D_databuf_reg_3_0_DXMUX
    );
  U_DCT1D_databuf_reg_3_0_XORF_1678 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_0_CYINIT,
      I1 => U_DCT1D_nx54687z1,
      O => U_DCT1D_databuf_reg_3_0_XORF
    );
  U_DCT1D_databuf_reg_3_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_0_CY0F,
      IB => U_DCT1D_databuf_reg_3_0_CYINIT,
      SEL => U_DCT1D_databuf_reg_3_0_CYSELF,
      O => U_DCT1D_rtlc5_1422_add_11_ix55684z63342_O
    );
  U_DCT1D_databuf_reg_3_0_CYINIT_1679 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_0_BXINVNOT,
      O => U_DCT1D_databuf_reg_3_0_CYINIT
    );
  U_DCT1D_databuf_reg_3_0_CY0F_1680 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(0),
      O => U_DCT1D_databuf_reg_3_0_CY0F
    );
  U_DCT1D_databuf_reg_3_0_CYSELF_1681 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx54687z1,
      O => U_DCT1D_databuf_reg_3_0_CYSELF
    );
  U_DCT1D_databuf_reg_3_0_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_11,
      O => U_DCT1D_databuf_reg_3_0_BXINVNOT
    );
  U_DCT1D_databuf_reg_3_0_DYMUX_1682 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_0_XORG,
      O => U_DCT1D_databuf_reg_3_0_DYMUX
    );
  U_DCT1D_databuf_reg_3_0_XORG_1683 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1422_add_11_ix55684z63342_O,
      I1 => U_DCT1D_nx55684z1,
      O => U_DCT1D_databuf_reg_3_0_XORG
    );
  U_DCT1D_databuf_reg_3_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_0_CYMUXG,
      O => U_DCT1D_rtlc5_1422_add_11_ix56681z63342_O
    );
  U_DCT1D_databuf_reg_3_0_CYMUXG_1684 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_0_CY0G,
      IB => U_DCT1D_rtlc5_1422_add_11_ix55684z63342_O,
      SEL => U_DCT1D_databuf_reg_3_0_CYSELG,
      O => U_DCT1D_databuf_reg_3_0_CYMUXG
    );
  U_DCT1D_databuf_reg_3_0_CY0G_1685 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(1),
      O => U_DCT1D_databuf_reg_3_0_CY0G
    );
  U_DCT1D_databuf_reg_3_0_CYSELG_1686 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx55684z1,
      O => U_DCT1D_databuf_reg_3_0_CYSELG
    );
  U_DCT1D_databuf_reg_3_0_SRINV_1687 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_3_0_SRINV
    );
  U_DCT1D_databuf_reg_3_0_CLKINV_1688 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_3_0_CLKINV
    );
  U_DCT1D_databuf_reg_3_0_CEINV_1689 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_3_0_CEINV
    );
  U_DCT1D_databuf_reg_3_2_DXMUX_1690 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_2_XORF,
      O => U_DCT1D_databuf_reg_3_2_DXMUX
    );
  U_DCT1D_databuf_reg_3_2_XORF_1691 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_2_CYINIT,
      I1 => U_DCT1D_nx56681z1,
      O => U_DCT1D_databuf_reg_3_2_XORF
    );
  U_DCT1D_databuf_reg_3_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_2_CY0F,
      IB => U_DCT1D_databuf_reg_3_2_CYINIT,
      SEL => U_DCT1D_databuf_reg_3_2_CYSELF,
      O => U_DCT1D_rtlc5_1422_add_11_ix57678z63342_O
    );
  U_DCT1D_databuf_reg_3_2_CYMUXF2_1692 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_2_CY0F,
      IB => U_DCT1D_databuf_reg_3_2_CY0F,
      SEL => U_DCT1D_databuf_reg_3_2_CYSELF,
      O => U_DCT1D_databuf_reg_3_2_CYMUXF2
    );
  U_DCT1D_databuf_reg_3_2_CYINIT_1693 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1422_add_11_ix56681z63342_O,
      O => U_DCT1D_databuf_reg_3_2_CYINIT
    );
  U_DCT1D_databuf_reg_3_2_CY0F_1694 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(2),
      O => U_DCT1D_databuf_reg_3_2_CY0F
    );
  U_DCT1D_databuf_reg_3_2_CYSELF_1695 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx56681z1,
      O => U_DCT1D_databuf_reg_3_2_CYSELF
    );
  U_DCT1D_databuf_reg_3_2_DYMUX_1696 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_2_XORG,
      O => U_DCT1D_databuf_reg_3_2_DYMUX
    );
  U_DCT1D_databuf_reg_3_2_XORG_1697 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1422_add_11_ix57678z63342_O,
      I1 => U_DCT1D_nx57678z1,
      O => U_DCT1D_databuf_reg_3_2_XORG
    );
  U_DCT1D_databuf_reg_3_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_2_CYMUXFAST,
      O => U_DCT1D_rtlc5_1422_add_11_ix58675z63342_O
    );
  U_DCT1D_databuf_reg_3_2_FASTCARRY_1698 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1422_add_11_ix56681z63342_O,
      O => U_DCT1D_databuf_reg_3_2_FASTCARRY
    );
  U_DCT1D_databuf_reg_3_2_CYAND_1699 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_3_2_CYSELG,
      I1 => U_DCT1D_databuf_reg_3_2_CYSELF,
      O => U_DCT1D_databuf_reg_3_2_CYAND
    );
  U_DCT1D_databuf_reg_3_2_CYMUXFAST_1700 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_2_CYMUXG2,
      IB => U_DCT1D_databuf_reg_3_2_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_3_2_CYAND,
      O => U_DCT1D_databuf_reg_3_2_CYMUXFAST
    );
  U_DCT1D_databuf_reg_3_2_CYMUXG2_1701 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_2_CY0G,
      IB => U_DCT1D_databuf_reg_3_2_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_3_2_CYSELG,
      O => U_DCT1D_databuf_reg_3_2_CYMUXG2
    );
  U_DCT1D_databuf_reg_3_2_CY0G_1702 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(3),
      O => U_DCT1D_databuf_reg_3_2_CY0G
    );
  U_DCT1D_databuf_reg_3_2_CYSELG_1703 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx57678z1,
      O => U_DCT1D_databuf_reg_3_2_CYSELG
    );
  U_DCT1D_databuf_reg_3_2_SRINV_1704 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_3_2_SRINV
    );
  U_DCT1D_databuf_reg_3_2_CLKINV_1705 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_3_2_CLKINV
    );
  U_DCT1D_databuf_reg_3_2_CEINV_1706 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_3_2_CEINV
    );
  U_DCT1D_databuf_reg_3_4_DXMUX_1707 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_4_XORF,
      O => U_DCT1D_databuf_reg_3_4_DXMUX
    );
  U_DCT1D_databuf_reg_3_4_XORF_1708 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_4_CYINIT,
      I1 => U_DCT1D_nx58675z1,
      O => U_DCT1D_databuf_reg_3_4_XORF
    );
  U_DCT1D_databuf_reg_3_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_4_CY0F,
      IB => U_DCT1D_databuf_reg_3_4_CYINIT,
      SEL => U_DCT1D_databuf_reg_3_4_CYSELF,
      O => U_DCT1D_rtlc5_1422_add_11_ix59672z63342_O
    );
  U_DCT1D_databuf_reg_3_4_CYMUXF2_1709 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_4_CY0F,
      IB => U_DCT1D_databuf_reg_3_4_CY0F,
      SEL => U_DCT1D_databuf_reg_3_4_CYSELF,
      O => U_DCT1D_databuf_reg_3_4_CYMUXF2
    );
  U_DCT1D_databuf_reg_3_4_CYINIT_1710 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1422_add_11_ix58675z63342_O,
      O => U_DCT1D_databuf_reg_3_4_CYINIT
    );
  U_DCT1D_databuf_reg_3_4_CY0F_1711 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(4),
      O => U_DCT1D_databuf_reg_3_4_CY0F
    );
  U_DCT1D_databuf_reg_3_4_CYSELF_1712 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx58675z1,
      O => U_DCT1D_databuf_reg_3_4_CYSELF
    );
  U_DCT1D_databuf_reg_3_4_DYMUX_1713 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_4_XORG,
      O => U_DCT1D_databuf_reg_3_4_DYMUX
    );
  U_DCT1D_databuf_reg_3_4_XORG_1714 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1422_add_11_ix59672z63342_O,
      I1 => U_DCT1D_nx59672z1,
      O => U_DCT1D_databuf_reg_3_4_XORG
    );
  U_DCT1D_databuf_reg_3_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_4_CYMUXFAST,
      O => U_DCT1D_rtlc5_1422_add_11_ix60669z63342_O
    );
  U_DCT1D_databuf_reg_3_4_FASTCARRY_1715 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1422_add_11_ix58675z63342_O,
      O => U_DCT1D_databuf_reg_3_4_FASTCARRY
    );
  U_DCT1D_databuf_reg_3_4_CYAND_1716 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_3_4_CYSELG,
      I1 => U_DCT1D_databuf_reg_3_4_CYSELF,
      O => U_DCT1D_databuf_reg_3_4_CYAND
    );
  U_DCT1D_databuf_reg_3_4_CYMUXFAST_1717 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_4_CYMUXG2,
      IB => U_DCT1D_databuf_reg_3_4_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_3_4_CYAND,
      O => U_DCT1D_databuf_reg_3_4_CYMUXFAST
    );
  U_DCT1D_databuf_reg_3_4_CYMUXG2_1718 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_4_CY0G,
      IB => U_DCT1D_databuf_reg_3_4_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_3_4_CYSELG,
      O => U_DCT1D_databuf_reg_3_4_CYMUXG2
    );
  U_DCT1D_databuf_reg_3_4_CY0G_1719 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(5),
      O => U_DCT1D_databuf_reg_3_4_CY0G
    );
  U_DCT1D_databuf_reg_3_4_CYSELG_1720 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59672z1,
      O => U_DCT1D_databuf_reg_3_4_CYSELG
    );
  U_DCT1D_databuf_reg_3_4_SRINV_1721 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_3_4_SRINV
    );
  U_DCT1D_databuf_reg_3_4_CLKINV_1722 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_3_4_CLKINV
    );
  U_DCT1D_databuf_reg_3_4_CEINV_1723 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_3_4_CEINV
    );
  U_DCT1D_databuf_reg_3_6_DXMUX_1724 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_6_XORF,
      O => U_DCT1D_databuf_reg_3_6_DXMUX
    );
  U_DCT1D_databuf_reg_3_6_XORF_1725 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_6_CYINIT,
      I1 => U_DCT1D_nx60669z1,
      O => U_DCT1D_databuf_reg_3_6_XORF
    );
  U_DCT1D_databuf_reg_3_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_6_CY0F,
      IB => U_DCT1D_databuf_reg_3_6_CYINIT,
      SEL => U_DCT1D_databuf_reg_3_6_CYSELF,
      O => U_DCT1D_rtlc5_1422_add_11_ix61666z63342_O
    );
  U_DCT1D_databuf_reg_3_6_CYMUXF2_1726 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_6_CY0F,
      IB => U_DCT1D_databuf_reg_3_6_CY0F,
      SEL => U_DCT1D_databuf_reg_3_6_CYSELF,
      O => U_DCT1D_databuf_reg_3_6_CYMUXF2
    );
  U_DCT1D_databuf_reg_3_6_CYINIT_1727 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1422_add_11_ix60669z63342_O,
      O => U_DCT1D_databuf_reg_3_6_CYINIT
    );
  U_DCT1D_databuf_reg_3_6_CY0F_1728 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(6),
      O => U_DCT1D_databuf_reg_3_6_CY0F
    );
  U_DCT1D_databuf_reg_3_6_CYSELF_1729 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx60669z1,
      O => U_DCT1D_databuf_reg_3_6_CYSELF
    );
  U_DCT1D_databuf_reg_3_6_DYMUX_1730 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_6_XORG,
      O => U_DCT1D_databuf_reg_3_6_DYMUX
    );
  U_DCT1D_databuf_reg_3_6_XORG_1731 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_1422_add_11_ix61666z63342_O,
      I1 => U_DCT1D_nx61666z1,
      O => U_DCT1D_databuf_reg_3_6_XORG
    );
  U_DCT1D_databuf_reg_3_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_6_CYMUXFAST,
      O => U_DCT1D_rtlc5_1422_add_11_ix62663z63342_O
    );
  U_DCT1D_databuf_reg_3_6_FASTCARRY_1732 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1422_add_11_ix60669z63342_O,
      O => U_DCT1D_databuf_reg_3_6_FASTCARRY
    );
  U_DCT1D_databuf_reg_3_6_CYAND_1733 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_3_6_CYSELG,
      I1 => U_DCT1D_databuf_reg_3_6_CYSELF,
      O => U_DCT1D_databuf_reg_3_6_CYAND
    );
  U_DCT1D_databuf_reg_3_6_CYMUXFAST_1734 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_6_CYMUXG2,
      IB => U_DCT1D_databuf_reg_3_6_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_3_6_CYAND,
      O => U_DCT1D_databuf_reg_3_6_CYMUXFAST
    );
  U_DCT1D_databuf_reg_3_6_CYMUXG2_1735 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_3_6_CY0G,
      IB => U_DCT1D_databuf_reg_3_6_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_3_6_CYSELG,
      O => U_DCT1D_databuf_reg_3_6_CYMUXG2
    );
  U_DCT1D_databuf_reg_3_6_CY0G_1736 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(7),
      O => U_DCT1D_databuf_reg_3_6_CY0G
    );
  U_DCT1D_databuf_reg_3_6_CYSELG_1737 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx61666z1,
      O => U_DCT1D_databuf_reg_3_6_CYSELG
    );
  U_DCT1D_databuf_reg_3_6_SRINV_1738 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_3_6_SRINV
    );
  U_DCT1D_databuf_reg_3_6_CLKINV_1739 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_3_6_CLKINV
    );
  U_DCT1D_databuf_reg_3_6_CEINV_1740 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_3_6_CEINV
    );
  U_DCT1D_databuf_reg_3_8_DXMUX_1741 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_8_XORF,
      O => U_DCT1D_databuf_reg_3_8_DXMUX
    );
  U_DCT1D_databuf_reg_3_8_XORF_1742 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_8_CYINIT,
      I1 => U_DCT1D_nx62663z1_rt,
      O => U_DCT1D_databuf_reg_3_8_XORF
    );
  U_DCT1D_databuf_reg_3_8_CYINIT_1743 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_1422_add_11_ix62663z63342_O,
      O => U_DCT1D_databuf_reg_3_8_CYINIT
    );
  U_DCT1D_databuf_reg_3_8_CLKINV_1744 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_3_8_CLKINV
    );
  U_DCT1D_databuf_reg_3_8_CEINV_1745 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_3_8_CEINV
    );
  U_DCT2D_rtlc5n1492_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_4_CY0F,
      IB => U_DCT2D_rtlc5n1492_4_CYINIT,
      SEL => U_DCT2D_rtlc5n1492_4_CYSELF,
      O => U_DCT2D_rtlc_387_add_64_ix65206z63433_O
    );
  U_DCT2D_rtlc5n1492_4_CYINIT_1746 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_4_BXINVNOT,
      O => U_DCT2D_rtlc5n1492_4_CYINIT
    );
  U_DCT2D_rtlc5n1492_4_CY0F_1747 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s(3),
      O => U_DCT2D_rtlc5n1492_4_CY0F
    );
  U_DCT2D_rtlc5n1492_4_CYSELF_1748 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z77,
      O => U_DCT2D_rtlc5n1492_4_CYSELF
    );
  U_DCT2D_rtlc5n1492_4_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_37,
      O => U_DCT2D_rtlc5n1492_4_BXINVNOT
    );
  U_DCT2D_rtlc5n1492_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_4_XORG,
      O => U_DCT2D_rtlc5n1492(4)
    );
  U_DCT2D_rtlc5n1492_4_XORG_1749 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_387_add_64_ix65206z63433_O,
      I1 => U_DCT2D_nx65206z74,
      O => U_DCT2D_rtlc5n1492_4_XORG
    );
  U_DCT2D_rtlc5n1492_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_4_CYMUXG,
      O => U_DCT2D_rtlc_387_add_64_ix65206z63429_O
    );
  U_DCT2D_rtlc5n1492_4_CYMUXG_1750 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_4_CY0G,
      IB => U_DCT2D_rtlc_387_add_64_ix65206z63433_O,
      SEL => U_DCT2D_rtlc5n1492_4_CYSELG,
      O => U_DCT2D_rtlc5n1492_4_CYMUXG
    );
  U_DCT2D_rtlc5n1492_4_CY0G_1751 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s(4),
      O => U_DCT2D_rtlc5n1492_4_CY0G
    );
  U_DCT2D_rtlc5n1492_4_CYSELG_1752 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z74,
      O => U_DCT2D_rtlc5n1492_4_CYSELG
    );
  U_DCT2D_rtlc5n1492_5_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_5_XORF,
      O => U_DCT2D_rtlc5n1492(5)
    );
  U_DCT2D_rtlc5n1492_5_XORF_1753 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1492_5_CYINIT,
      I1 => U_DCT2D_nx65206z71,
      O => U_DCT2D_rtlc5n1492_5_XORF
    );
  U_DCT2D_rtlc5n1492_5_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_5_CY0F,
      IB => U_DCT2D_rtlc5n1492_5_CYINIT,
      SEL => U_DCT2D_rtlc5n1492_5_CYSELF,
      O => U_DCT2D_rtlc_387_add_64_ix65206z63426_O
    );
  U_DCT2D_rtlc5n1492_5_CYMUXF2_1754 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_5_CY0F,
      IB => U_DCT2D_rtlc5n1492_5_CY0F,
      SEL => U_DCT2D_rtlc5n1492_5_CYSELF,
      O => U_DCT2D_rtlc5n1492_5_CYMUXF2
    );
  U_DCT2D_rtlc5n1492_5_CYINIT_1755 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_387_add_64_ix65206z63429_O,
      O => U_DCT2D_rtlc5n1492_5_CYINIT
    );
  U_DCT2D_rtlc5n1492_5_CY0F_1756 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s(5),
      O => U_DCT2D_rtlc5n1492_5_CY0F
    );
  U_DCT2D_rtlc5n1492_5_CYSELF_1757 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z71,
      O => U_DCT2D_rtlc5n1492_5_CYSELF
    );
  U_DCT2D_rtlc5n1492_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_5_XORG,
      O => U_DCT2D_rtlc5n1492(6)
    );
  U_DCT2D_rtlc5n1492_5_XORG_1758 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_387_add_64_ix65206z63426_O,
      I1 => U_DCT2D_nx65206z68,
      O => U_DCT2D_rtlc5n1492_5_XORG
    );
  U_DCT2D_rtlc5n1492_5_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_5_CYMUXFAST,
      O => U_DCT2D_rtlc_387_add_64_ix65206z63422_O
    );
  U_DCT2D_rtlc5n1492_5_FASTCARRY_1759 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_387_add_64_ix65206z63429_O,
      O => U_DCT2D_rtlc5n1492_5_FASTCARRY
    );
  U_DCT2D_rtlc5n1492_5_CYAND_1760 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1492_5_CYSELG,
      I1 => U_DCT2D_rtlc5n1492_5_CYSELF,
      O => U_DCT2D_rtlc5n1492_5_CYAND
    );
  U_DCT2D_rtlc5n1492_5_CYMUXFAST_1761 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_5_CYMUXG2,
      IB => U_DCT2D_rtlc5n1492_5_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1492_5_CYAND,
      O => U_DCT2D_rtlc5n1492_5_CYMUXFAST
    );
  U_DCT2D_rtlc5n1492_5_CYMUXG2_1762 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_5_CY0G,
      IB => U_DCT2D_rtlc5n1492_5_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1492_5_CYSELG,
      O => U_DCT2D_rtlc5n1492_5_CYMUXG2
    );
  U_DCT2D_rtlc5n1492_5_CY0G_1763 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s(6),
      O => U_DCT2D_rtlc5n1492_5_CY0G
    );
  U_DCT2D_rtlc5n1492_5_CYSELG_1764 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z68,
      O => U_DCT2D_rtlc5n1492_5_CYSELG
    );
  U_DCT2D_rtlc5n1492_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_7_XORF,
      O => U_DCT2D_rtlc5n1492(7)
    );
  U_DCT2D_rtlc5n1492_7_XORF_1765 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1492_7_CYINIT,
      I1 => U_DCT2D_nx65206z65,
      O => U_DCT2D_rtlc5n1492_7_XORF
    );
  U_DCT2D_rtlc5n1492_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_7_CY0F,
      IB => U_DCT2D_rtlc5n1492_7_CYINIT,
      SEL => U_DCT2D_rtlc5n1492_7_CYSELF,
      O => U_DCT2D_rtlc_387_add_64_ix65206z63419_O
    );
  U_DCT2D_rtlc5n1492_7_CYMUXF2_1766 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_7_CY0F,
      IB => U_DCT2D_rtlc5n1492_7_CY0F,
      SEL => U_DCT2D_rtlc5n1492_7_CYSELF,
      O => U_DCT2D_rtlc5n1492_7_CYMUXF2
    );
  U_DCT2D_rtlc5n1492_7_CYINIT_1767 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_387_add_64_ix65206z63422_O,
      O => U_DCT2D_rtlc5n1492_7_CYINIT
    );
  U_DCT2D_rtlc5n1492_7_CY0F_1768 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s(7),
      O => U_DCT2D_rtlc5n1492_7_CY0F
    );
  U_DCT2D_rtlc5n1492_7_CYSELF_1769 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z65,
      O => U_DCT2D_rtlc5n1492_7_CYSELF
    );
  U_DCT2D_rtlc5n1492_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_7_XORG,
      O => U_DCT2D_rtlc5n1492(8)
    );
  U_DCT2D_rtlc5n1492_7_XORG_1770 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_387_add_64_ix65206z63419_O,
      I1 => U_DCT2D_nx65206z62,
      O => U_DCT2D_rtlc5n1492_7_XORG
    );
  U_DCT2D_rtlc5n1492_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_7_CYMUXFAST,
      O => U_DCT2D_rtlc_387_add_64_ix65206z63415_O
    );
  U_DCT2D_rtlc5n1492_7_FASTCARRY_1771 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_387_add_64_ix65206z63422_O,
      O => U_DCT2D_rtlc5n1492_7_FASTCARRY
    );
  U_DCT2D_rtlc5n1492_7_CYAND_1772 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1492_7_CYSELG,
      I1 => U_DCT2D_rtlc5n1492_7_CYSELF,
      O => U_DCT2D_rtlc5n1492_7_CYAND
    );
  U_DCT2D_rtlc5n1492_7_CYMUXFAST_1773 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_7_CYMUXG2,
      IB => U_DCT2D_rtlc5n1492_7_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1492_7_CYAND,
      O => U_DCT2D_rtlc5n1492_7_CYMUXFAST
    );
  U_DCT2D_rtlc5n1492_7_CYMUXG2_1774 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_7_CY0G,
      IB => U_DCT2D_rtlc5n1492_7_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1492_7_CYSELG,
      O => U_DCT2D_rtlc5n1492_7_CYMUXG2
    );
  U_DCT2D_rtlc5n1492_7_CY0G_1775 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s(8),
      O => U_DCT2D_rtlc5n1492_7_CY0G
    );
  U_DCT2D_rtlc5n1492_7_CYSELG_1776 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z62,
      O => U_DCT2D_rtlc5n1492_7_CYSELG
    );
  U_DCT2D_rtlc5n1492_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_9_XORF,
      O => U_DCT2D_rtlc5n1492(9)
    );
  U_DCT2D_rtlc5n1492_9_XORF_1777 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1492_9_CYINIT,
      I1 => U_DCT2D_nx65206z59,
      O => U_DCT2D_rtlc5n1492_9_XORF
    );
  U_DCT2D_rtlc5n1492_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_9_CY0F,
      IB => U_DCT2D_rtlc5n1492_9_CYINIT,
      SEL => U_DCT2D_rtlc5n1492_9_CYSELF,
      O => U_DCT2D_rtlc_387_add_64_ix65206z63412_O
    );
  U_DCT2D_rtlc5n1492_9_CYMUXF2_1778 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_9_CY0F,
      IB => U_DCT2D_rtlc5n1492_9_CY0F,
      SEL => U_DCT2D_rtlc5n1492_9_CYSELF,
      O => U_DCT2D_rtlc5n1492_9_CYMUXF2
    );
  U_DCT2D_rtlc5n1492_9_CYINIT_1779 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_387_add_64_ix65206z63415_O,
      O => U_DCT2D_rtlc5n1492_9_CYINIT
    );
  U_DCT2D_rtlc5n1492_9_CY0F_1780 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s(9),
      O => U_DCT2D_rtlc5n1492_9_CY0F
    );
  U_DCT2D_rtlc5n1492_9_CYSELF_1781 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z59,
      O => U_DCT2D_rtlc5n1492_9_CYSELF
    );
  U_DCT2D_rtlc5n1492_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_9_XORG,
      O => U_DCT2D_rtlc5n1492(10)
    );
  U_DCT2D_rtlc5n1492_9_XORG_1782 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_387_add_64_ix65206z63412_O,
      I1 => U_DCT2D_nx65206z56,
      O => U_DCT2D_rtlc5n1492_9_XORG
    );
  U_DCT2D_rtlc5n1492_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_9_CYMUXFAST,
      O => U_DCT2D_rtlc_387_add_64_ix65206z63408_O
    );
  U_DCT2D_rtlc5n1492_9_FASTCARRY_1783 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_387_add_64_ix65206z63415_O,
      O => U_DCT2D_rtlc5n1492_9_FASTCARRY
    );
  U_DCT2D_rtlc5n1492_9_CYAND_1784 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1492_9_CYSELG,
      I1 => U_DCT2D_rtlc5n1492_9_CYSELF,
      O => U_DCT2D_rtlc5n1492_9_CYAND
    );
  U_DCT2D_rtlc5n1492_9_CYMUXFAST_1785 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_9_CYMUXG2,
      IB => U_DCT2D_rtlc5n1492_9_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1492_9_CYAND,
      O => U_DCT2D_rtlc5n1492_9_CYMUXFAST
    );
  U_DCT2D_rtlc5n1492_9_CYMUXG2_1786 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_9_CY0G,
      IB => U_DCT2D_rtlc5n1492_9_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1492_9_CYSELG,
      O => U_DCT2D_rtlc5n1492_9_CYMUXG2
    );
  U_DCT2D_rtlc5n1492_9_CY0G_1787 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s(10),
      O => U_DCT2D_rtlc5n1492_9_CY0G
    );
  U_DCT2D_rtlc5n1492_9_CYSELG_1788 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z56,
      O => U_DCT2D_rtlc5n1492_9_CYSELG
    );
  U_DCT2D_rtlc5n1492_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_11_XORF,
      O => U_DCT2D_rtlc5n1492(11)
    );
  U_DCT2D_rtlc5n1492_11_XORF_1789 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1492_11_CYINIT,
      I1 => U_DCT2D_nx65206z53,
      O => U_DCT2D_rtlc5n1492_11_XORF
    );
  U_DCT2D_rtlc5n1492_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_11_CY0F,
      IB => U_DCT2D_rtlc5n1492_11_CYINIT,
      SEL => U_DCT2D_rtlc5n1492_11_CYSELF,
      O => U_DCT2D_rtlc_387_add_64_ix65206z63405_O
    );
  U_DCT2D_rtlc5n1492_11_CYMUXF2_1790 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_11_CY0F,
      IB => U_DCT2D_rtlc5n1492_11_CY0F,
      SEL => U_DCT2D_rtlc5n1492_11_CYSELF,
      O => U_DCT2D_rtlc5n1492_11_CYMUXF2
    );
  U_DCT2D_rtlc5n1492_11_CYINIT_1791 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_387_add_64_ix65206z63408_O,
      O => U_DCT2D_rtlc5n1492_11_CYINIT
    );
  U_DCT2D_rtlc5n1492_11_CY0F_1792 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s(11),
      O => U_DCT2D_rtlc5n1492_11_CY0F
    );
  U_DCT2D_rtlc5n1492_11_CYSELF_1793 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z53,
      O => U_DCT2D_rtlc5n1492_11_CYSELF
    );
  U_DCT2D_rtlc5n1492_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_11_XORG,
      O => U_DCT2D_rtlc5n1492(12)
    );
  U_DCT2D_rtlc5n1492_11_XORG_1794 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_387_add_64_ix65206z63405_O,
      I1 => U_DCT2D_nx65206z50,
      O => U_DCT2D_rtlc5n1492_11_XORG
    );
  U_DCT2D_rtlc5n1492_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_11_CYMUXFAST,
      O => U_DCT2D_rtlc_387_add_64_ix65206z63401_O
    );
  U_DCT2D_rtlc5n1492_11_FASTCARRY_1795 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_387_add_64_ix65206z63408_O,
      O => U_DCT2D_rtlc5n1492_11_FASTCARRY
    );
  U_DCT2D_rtlc5n1492_11_CYAND_1796 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1492_11_CYSELG,
      I1 => U_DCT2D_rtlc5n1492_11_CYSELF,
      O => U_DCT2D_rtlc5n1492_11_CYAND
    );
  U_DCT2D_rtlc5n1492_11_CYMUXFAST_1797 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_11_CYMUXG2,
      IB => U_DCT2D_rtlc5n1492_11_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1492_11_CYAND,
      O => U_DCT2D_rtlc5n1492_11_CYMUXFAST
    );
  U_DCT2D_rtlc5n1492_11_CYMUXG2_1798 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_11_CY0G,
      IB => U_DCT2D_rtlc5n1492_11_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1492_11_CYSELG,
      O => U_DCT2D_rtlc5n1492_11_CYMUXG2
    );
  U_DCT2D_rtlc5n1492_11_CY0G_1799 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s(12),
      O => U_DCT2D_rtlc5n1492_11_CY0G
    );
  U_DCT2D_rtlc5n1492_11_CYSELG_1800 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z50,
      O => U_DCT2D_rtlc5n1492_11_CYSELG
    );
  U_DCT2D_rtlc5n1492_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_13_XORF,
      O => U_DCT2D_rtlc5n1492(13)
    );
  U_DCT2D_rtlc5n1492_13_XORF_1801 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1492_13_CYINIT,
      I1 => U_DCT2D_nx65206z47,
      O => U_DCT2D_rtlc5n1492_13_XORF
    );
  U_DCT2D_rtlc5n1492_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_13_CY0F,
      IB => U_DCT2D_rtlc5n1492_13_CYINIT,
      SEL => U_DCT2D_rtlc5n1492_13_CYSELF,
      O => U_DCT2D_rtlc_387_add_64_ix65206z63398_O
    );
  U_DCT2D_rtlc5n1492_13_CYMUXF2_1802 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_13_CY0F,
      IB => U_DCT2D_rtlc5n1492_13_CY0F,
      SEL => U_DCT2D_rtlc5n1492_13_CYSELF,
      O => U_DCT2D_rtlc5n1492_13_CYMUXF2
    );
  U_DCT2D_rtlc5n1492_13_CYINIT_1803 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_387_add_64_ix65206z63401_O,
      O => U_DCT2D_rtlc5n1492_13_CYINIT
    );
  U_DCT2D_rtlc5n1492_13_CY0F_1804 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s(13),
      O => U_DCT2D_rtlc5n1492_13_CY0F
    );
  U_DCT2D_rtlc5n1492_13_CYSELF_1805 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z47,
      O => U_DCT2D_rtlc5n1492_13_CYSELF
    );
  U_DCT2D_rtlc5n1492_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_13_XORG,
      O => U_DCT2D_rtlc5n1492(14)
    );
  U_DCT2D_rtlc5n1492_13_XORG_1806 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_387_add_64_ix65206z63398_O,
      I1 => U_DCT2D_nx65206z44,
      O => U_DCT2D_rtlc5n1492_13_XORG
    );
  U_DCT2D_rtlc5n1492_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_13_CYMUXFAST,
      O => U_DCT2D_rtlc_387_add_64_ix65206z63392_O
    );
  U_DCT2D_rtlc5n1492_13_FASTCARRY_1807 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_387_add_64_ix65206z63401_O,
      O => U_DCT2D_rtlc5n1492_13_FASTCARRY
    );
  U_DCT2D_rtlc5n1492_13_CYAND_1808 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1492_13_CYSELG,
      I1 => U_DCT2D_rtlc5n1492_13_CYSELF,
      O => U_DCT2D_rtlc5n1492_13_CYAND
    );
  U_DCT2D_rtlc5n1492_13_CYMUXFAST_1809 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_13_CYMUXG2,
      IB => U_DCT2D_rtlc5n1492_13_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1492_13_CYAND,
      O => U_DCT2D_rtlc5n1492_13_CYMUXFAST
    );
  U_DCT2D_rtlc5n1492_13_CYMUXG2_1810 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1492_13_CY0G,
      IB => U_DCT2D_rtlc5n1492_13_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1492_13_CYSELG,
      O => U_DCT2D_rtlc5n1492_13_CYMUXG2
    );
  U_DCT2D_rtlc5n1492_13_CY0G_1811 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s(13),
      O => U_DCT2D_rtlc5n1492_13_CY0G
    );
  U_DCT2D_rtlc5n1492_13_CYSELG_1812 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z44,
      O => U_DCT2D_rtlc5n1492_13_CYSELG
    );
  U_DCT2D_nx65206z42_rt_1813 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_nx65206z42,
      O => U_DCT2D_nx65206z42_rt
    );
  U_DCT2D_rtlc5n1492_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1492_15_XORF,
      O => U_DCT2D_rtlc5n1492(15)
    );
  U_DCT2D_rtlc5n1492_15_XORF_1814 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1492_15_CYINIT,
      I1 => U_DCT2D_nx65206z42_rt,
      O => U_DCT2D_rtlc5n1492_15_XORF
    );
  U_DCT2D_rtlc5n1492_15_CYINIT_1815 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_387_add_64_ix65206z63392_O,
      O => U_DCT2D_rtlc5n1492_15_CYINIT
    );
  U_DCT2D_rtlc5n1495_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_9_XORF,
      O => U_DCT2D_rtlc5n1495(9)
    );
  U_DCT2D_rtlc5n1495_9_XORF_1816 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1495_9_CYINIT,
      I1 => U_DCT2D_nx65206z369,
      O => U_DCT2D_rtlc5n1495_9_XORF
    );
  U_DCT2D_rtlc5n1495_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_9_CY0F,
      IB => U_DCT2D_rtlc5n1495_9_CYINIT,
      SEL => U_DCT2D_rtlc5n1495_9_CYSELF,
      O => U_DCT2D_rtlc_396_add_68_ix65206z63835_O
    );
  U_DCT2D_rtlc5n1495_9_CYINIT_1817 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_9_BXINVNOT,
      O => U_DCT2D_rtlc5n1495_9_CYINIT
    );
  U_DCT2D_rtlc5n1495_9_CY0F_1818 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s(3),
      O => U_DCT2D_rtlc5n1495_9_CY0F
    );
  U_DCT2D_rtlc5n1495_9_CYSELF_1819 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z369,
      O => U_DCT2D_rtlc5n1495_9_CYSELF
    );
  U_DCT2D_rtlc5n1495_9_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_4,
      O => U_DCT2D_rtlc5n1495_9_BXINVNOT
    );
  U_DCT2D_rtlc5n1495_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_9_XORG,
      O => U_DCT2D_rtlc5n1495(10)
    );
  U_DCT2D_rtlc5n1495_9_XORG_1820 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_396_add_68_ix65206z63835_O,
      I1 => U_DCT2D_nx65206z366,
      O => U_DCT2D_rtlc5n1495_9_XORG
    );
  U_DCT2D_rtlc5n1495_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_9_CYMUXG,
      O => U_DCT2D_rtlc_396_add_68_ix65206z63832_O
    );
  U_DCT2D_rtlc5n1495_9_CYMUXG_1821 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_9_CY0G,
      IB => U_DCT2D_rtlc_396_add_68_ix65206z63835_O,
      SEL => U_DCT2D_rtlc5n1495_9_CYSELG,
      O => U_DCT2D_rtlc5n1495_9_CYMUXG
    );
  U_DCT2D_rtlc5n1495_9_CY0G_1822 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s(4),
      O => U_DCT2D_rtlc5n1495_9_CY0G
    );
  U_DCT2D_rtlc5n1495_9_CYSELG_1823 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z366,
      O => U_DCT2D_rtlc5n1495_9_CYSELG
    );
  U_DCT2D_rtlc5n1495_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_11_XORF,
      O => U_DCT2D_rtlc5n1495(11)
    );
  U_DCT2D_rtlc5n1495_11_XORF_1824 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1495_11_CYINIT,
      I1 => U_DCT2D_nx65206z363,
      O => U_DCT2D_rtlc5n1495_11_XORF
    );
  U_DCT2D_rtlc5n1495_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_11_CY0F,
      IB => U_DCT2D_rtlc5n1495_11_CYINIT,
      SEL => U_DCT2D_rtlc5n1495_11_CYSELF,
      O => U_DCT2D_rtlc_396_add_68_ix65206z63828_O
    );
  U_DCT2D_rtlc5n1495_11_CYMUXF2_1825 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_11_CY0F,
      IB => U_DCT2D_rtlc5n1495_11_CY0F,
      SEL => U_DCT2D_rtlc5n1495_11_CYSELF,
      O => U_DCT2D_rtlc5n1495_11_CYMUXF2
    );
  U_DCT2D_rtlc5n1495_11_CYINIT_1826 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_396_add_68_ix65206z63832_O,
      O => U_DCT2D_rtlc5n1495_11_CYINIT
    );
  U_DCT2D_rtlc5n1495_11_CY0F_1827 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s(5),
      O => U_DCT2D_rtlc5n1495_11_CY0F
    );
  U_DCT2D_rtlc5n1495_11_CYSELF_1828 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z363,
      O => U_DCT2D_rtlc5n1495_11_CYSELF
    );
  U_DCT2D_rtlc5n1495_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_11_XORG,
      O => U_DCT2D_rtlc5n1495(12)
    );
  U_DCT2D_rtlc5n1495_11_XORG_1829 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_396_add_68_ix65206z63828_O,
      I1 => U_DCT2D_nx65206z360,
      O => U_DCT2D_rtlc5n1495_11_XORG
    );
  U_DCT2D_rtlc5n1495_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_11_CYMUXFAST,
      O => U_DCT2D_rtlc_396_add_68_ix65206z63825_O
    );
  U_DCT2D_rtlc5n1495_11_FASTCARRY_1830 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_396_add_68_ix65206z63832_O,
      O => U_DCT2D_rtlc5n1495_11_FASTCARRY
    );
  U_DCT2D_rtlc5n1495_11_CYAND_1831 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1495_11_CYSELG,
      I1 => U_DCT2D_rtlc5n1495_11_CYSELF,
      O => U_DCT2D_rtlc5n1495_11_CYAND
    );
  U_DCT2D_rtlc5n1495_11_CYMUXFAST_1832 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_11_CYMUXG2,
      IB => U_DCT2D_rtlc5n1495_11_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1495_11_CYAND,
      O => U_DCT2D_rtlc5n1495_11_CYMUXFAST
    );
  U_DCT2D_rtlc5n1495_11_CYMUXG2_1833 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_11_CY0G,
      IB => U_DCT2D_rtlc5n1495_11_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1495_11_CYSELG,
      O => U_DCT2D_rtlc5n1495_11_CYMUXG2
    );
  U_DCT2D_rtlc5n1495_11_CY0G_1834 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s(6),
      O => U_DCT2D_rtlc5n1495_11_CY0G
    );
  U_DCT2D_rtlc5n1495_11_CYSELG_1835 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z360,
      O => U_DCT2D_rtlc5n1495_11_CYSELG
    );
  U_DCT2D_rtlc5n1495_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_13_XORF,
      O => U_DCT2D_rtlc5n1495(13)
    );
  U_DCT2D_rtlc5n1495_13_XORF_1836 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1495_13_CYINIT,
      I1 => U_DCT2D_nx65206z357,
      O => U_DCT2D_rtlc5n1495_13_XORF
    );
  U_DCT2D_rtlc5n1495_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_13_CY0F,
      IB => U_DCT2D_rtlc5n1495_13_CYINIT,
      SEL => U_DCT2D_rtlc5n1495_13_CYSELF,
      O => U_DCT2D_rtlc_396_add_68_ix65206z63821_O
    );
  U_DCT2D_rtlc5n1495_13_CYMUXF2_1837 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_13_CY0F,
      IB => U_DCT2D_rtlc5n1495_13_CY0F,
      SEL => U_DCT2D_rtlc5n1495_13_CYSELF,
      O => U_DCT2D_rtlc5n1495_13_CYMUXF2
    );
  U_DCT2D_rtlc5n1495_13_CYINIT_1838 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_396_add_68_ix65206z63825_O,
      O => U_DCT2D_rtlc5n1495_13_CYINIT
    );
  U_DCT2D_rtlc5n1495_13_CY0F_1839 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s(7),
      O => U_DCT2D_rtlc5n1495_13_CY0F
    );
  U_DCT2D_rtlc5n1495_13_CYSELF_1840 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z357,
      O => U_DCT2D_rtlc5n1495_13_CYSELF
    );
  U_DCT2D_rtlc5n1495_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_13_XORG,
      O => U_DCT2D_rtlc5n1495(14)
    );
  U_DCT2D_rtlc5n1495_13_XORG_1841 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_396_add_68_ix65206z63821_O,
      I1 => U_DCT2D_nx65206z354,
      O => U_DCT2D_rtlc5n1495_13_XORG
    );
  U_DCT2D_rtlc5n1495_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_13_CYMUXFAST,
      O => U_DCT2D_rtlc_396_add_68_ix65206z63818_O
    );
  U_DCT2D_rtlc5n1495_13_FASTCARRY_1842 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_396_add_68_ix65206z63825_O,
      O => U_DCT2D_rtlc5n1495_13_FASTCARRY
    );
  U_DCT2D_rtlc5n1495_13_CYAND_1843 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1495_13_CYSELG,
      I1 => U_DCT2D_rtlc5n1495_13_CYSELF,
      O => U_DCT2D_rtlc5n1495_13_CYAND
    );
  U_DCT2D_rtlc5n1495_13_CYMUXFAST_1844 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_13_CYMUXG2,
      IB => U_DCT2D_rtlc5n1495_13_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1495_13_CYAND,
      O => U_DCT2D_rtlc5n1495_13_CYMUXFAST
    );
  U_DCT2D_rtlc5n1495_13_CYMUXG2_1845 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_13_CY0G,
      IB => U_DCT2D_rtlc5n1495_13_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1495_13_CYSELG,
      O => U_DCT2D_rtlc5n1495_13_CYMUXG2
    );
  U_DCT2D_rtlc5n1495_13_CY0G_1846 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s(8),
      O => U_DCT2D_rtlc5n1495_13_CY0G
    );
  U_DCT2D_rtlc5n1495_13_CYSELG_1847 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z354,
      O => U_DCT2D_rtlc5n1495_13_CYSELG
    );
  U_DCT2D_rtlc5n1495_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_15_XORF,
      O => U_DCT2D_rtlc5n1495(15)
    );
  U_DCT2D_rtlc5n1495_15_XORF_1848 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1495_15_CYINIT,
      I1 => U_DCT2D_nx65206z351,
      O => U_DCT2D_rtlc5n1495_15_XORF
    );
  U_DCT2D_rtlc5n1495_15_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_15_CY0F,
      IB => U_DCT2D_rtlc5n1495_15_CYINIT,
      SEL => U_DCT2D_rtlc5n1495_15_CYSELF,
      O => U_DCT2D_rtlc_396_add_68_ix65206z63814_O
    );
  U_DCT2D_rtlc5n1495_15_CYMUXF2_1849 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_15_CY0F,
      IB => U_DCT2D_rtlc5n1495_15_CY0F,
      SEL => U_DCT2D_rtlc5n1495_15_CYSELF,
      O => U_DCT2D_rtlc5n1495_15_CYMUXF2
    );
  U_DCT2D_rtlc5n1495_15_CYINIT_1850 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_396_add_68_ix65206z63818_O,
      O => U_DCT2D_rtlc5n1495_15_CYINIT
    );
  U_DCT2D_rtlc5n1495_15_CY0F_1851 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s(9),
      O => U_DCT2D_rtlc5n1495_15_CY0F
    );
  U_DCT2D_rtlc5n1495_15_CYSELF_1852 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z351,
      O => U_DCT2D_rtlc5n1495_15_CYSELF
    );
  U_DCT2D_rtlc5n1495_15_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_15_XORG,
      O => U_DCT2D_rtlc5n1495(16)
    );
  U_DCT2D_rtlc5n1495_15_XORG_1853 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_396_add_68_ix65206z63814_O,
      I1 => U_DCT2D_nx65206z348,
      O => U_DCT2D_rtlc5n1495_15_XORG
    );
  U_DCT2D_rtlc5n1495_15_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_15_CYMUXFAST,
      O => U_DCT2D_rtlc_396_add_68_ix65206z63811_O
    );
  U_DCT2D_rtlc5n1495_15_FASTCARRY_1854 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_396_add_68_ix65206z63818_O,
      O => U_DCT2D_rtlc5n1495_15_FASTCARRY
    );
  U_DCT2D_rtlc5n1495_15_CYAND_1855 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1495_15_CYSELG,
      I1 => U_DCT2D_rtlc5n1495_15_CYSELF,
      O => U_DCT2D_rtlc5n1495_15_CYAND
    );
  U_DCT2D_rtlc5n1495_15_CYMUXFAST_1856 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_15_CYMUXG2,
      IB => U_DCT2D_rtlc5n1495_15_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1495_15_CYAND,
      O => U_DCT2D_rtlc5n1495_15_CYMUXFAST
    );
  U_DCT2D_rtlc5n1495_15_CYMUXG2_1857 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_15_CY0G,
      IB => U_DCT2D_rtlc5n1495_15_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1495_15_CYSELG,
      O => U_DCT2D_rtlc5n1495_15_CYMUXG2
    );
  U_DCT2D_rtlc5n1495_15_CY0G_1858 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s(10),
      O => U_DCT2D_rtlc5n1495_15_CY0G
    );
  U_DCT2D_rtlc5n1495_15_CYSELG_1859 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z348,
      O => U_DCT2D_rtlc5n1495_15_CYSELG
    );
  U_DCT1D_reg_databuf_reg_2_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_2_4_DYMUX,
      CE => U_DCT1D_databuf_reg_2_4_CEINV,
      CLK => U_DCT1D_databuf_reg_2_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_2_4_FFY_RST,
      O => U_DCT1D_databuf_reg_2_Q(5)
    );
  U_DCT1D_databuf_reg_2_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_2_4_FFY_RST
    );
  U_DCT2D_rtlc5n1495_17_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_17_XORF,
      O => U_DCT2D_rtlc5n1495(17)
    );
  U_DCT2D_rtlc5n1495_17_XORF_1860 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1495_17_CYINIT,
      I1 => U_DCT2D_nx65206z345,
      O => U_DCT2D_rtlc5n1495_17_XORF
    );
  U_DCT2D_rtlc5n1495_17_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_17_CY0F,
      IB => U_DCT2D_rtlc5n1495_17_CYINIT,
      SEL => U_DCT2D_rtlc5n1495_17_CYSELF,
      O => U_DCT2D_rtlc_396_add_68_ix65206z63807_O
    );
  U_DCT2D_rtlc5n1495_17_CYMUXF2_1861 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_17_CY0F,
      IB => U_DCT2D_rtlc5n1495_17_CY0F,
      SEL => U_DCT2D_rtlc5n1495_17_CYSELF,
      O => U_DCT2D_rtlc5n1495_17_CYMUXF2
    );
  U_DCT2D_rtlc5n1495_17_CYINIT_1862 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_396_add_68_ix65206z63811_O,
      O => U_DCT2D_rtlc5n1495_17_CYINIT
    );
  U_DCT2D_rtlc5n1495_17_CY0F_1863 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s(11),
      O => U_DCT2D_rtlc5n1495_17_CY0F
    );
  U_DCT2D_rtlc5n1495_17_CYSELF_1864 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z345,
      O => U_DCT2D_rtlc5n1495_17_CYSELF
    );
  U_DCT2D_rtlc5n1495_17_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_17_XORG,
      O => U_DCT2D_rtlc5n1495(18)
    );
  U_DCT2D_rtlc5n1495_17_XORG_1865 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_396_add_68_ix65206z63807_O,
      I1 => U_DCT2D_nx65206z342,
      O => U_DCT2D_rtlc5n1495_17_XORG
    );
  U_DCT2D_rtlc5n1495_17_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_17_CYMUXFAST,
      O => U_DCT2D_rtlc_396_add_68_ix65206z63804_O
    );
  U_DCT2D_rtlc5n1495_17_FASTCARRY_1866 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_396_add_68_ix65206z63811_O,
      O => U_DCT2D_rtlc5n1495_17_FASTCARRY
    );
  U_DCT2D_rtlc5n1495_17_CYAND_1867 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1495_17_CYSELG,
      I1 => U_DCT2D_rtlc5n1495_17_CYSELF,
      O => U_DCT2D_rtlc5n1495_17_CYAND
    );
  U_DCT2D_rtlc5n1495_17_CYMUXFAST_1868 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_17_CYMUXG2,
      IB => U_DCT2D_rtlc5n1495_17_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1495_17_CYAND,
      O => U_DCT2D_rtlc5n1495_17_CYMUXFAST
    );
  U_DCT2D_rtlc5n1495_17_CYMUXG2_1869 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_17_CY0G,
      IB => U_DCT2D_rtlc5n1495_17_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1495_17_CYSELG,
      O => U_DCT2D_rtlc5n1495_17_CYMUXG2
    );
  U_DCT2D_rtlc5n1495_17_CY0G_1870 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s(12),
      O => U_DCT2D_rtlc5n1495_17_CY0G
    );
  U_DCT2D_rtlc5n1495_17_CYSELG_1871 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z342,
      O => U_DCT2D_rtlc5n1495_17_CYSELG
    );
  U_DCT2D_rtlc5n1495_19_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_19_XORF,
      O => U_DCT2D_rtlc5n1495(19)
    );
  U_DCT2D_rtlc5n1495_19_XORF_1872 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1495_19_CYINIT,
      I1 => U_DCT2D_nx65206z339,
      O => U_DCT2D_rtlc5n1495_19_XORF
    );
  U_DCT2D_rtlc5n1495_19_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_19_CY0F,
      IB => U_DCT2D_rtlc5n1495_19_CYINIT,
      SEL => U_DCT2D_rtlc5n1495_19_CYSELF,
      O => U_DCT2D_rtlc_396_add_68_ix65206z63800_O
    );
  U_DCT2D_rtlc5n1495_19_CYMUXF2_1873 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_19_CY0F,
      IB => U_DCT2D_rtlc5n1495_19_CY0F,
      SEL => U_DCT2D_rtlc5n1495_19_CYSELF,
      O => U_DCT2D_rtlc5n1495_19_CYMUXF2
    );
  U_DCT2D_rtlc5n1495_19_CYINIT_1874 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_396_add_68_ix65206z63804_O,
      O => U_DCT2D_rtlc5n1495_19_CYINIT
    );
  U_DCT2D_rtlc5n1495_19_CY0F_1875 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s(13),
      O => U_DCT2D_rtlc5n1495_19_CY0F
    );
  U_DCT2D_rtlc5n1495_19_CYSELF_1876 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z339,
      O => U_DCT2D_rtlc5n1495_19_CYSELF
    );
  U_DCT2D_rtlc5n1495_19_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_19_XORG,
      O => U_DCT2D_rtlc5n1495(20)
    );
  U_DCT2D_rtlc5n1495_19_XORG_1877 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_396_add_68_ix65206z63800_O,
      I1 => U_DCT2D_nx65206z336,
      O => U_DCT2D_rtlc5n1495_19_XORG
    );
  U_DCT2D_rtlc5n1495_19_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_19_CYMUXFAST,
      O => U_DCT2D_rtlc_396_add_68_ix65206z63797_O
    );
  U_DCT2D_rtlc5n1495_19_FASTCARRY_1878 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_396_add_68_ix65206z63804_O,
      O => U_DCT2D_rtlc5n1495_19_FASTCARRY
    );
  U_DCT2D_rtlc5n1495_19_CYAND_1879 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1495_19_CYSELG,
      I1 => U_DCT2D_rtlc5n1495_19_CYSELF,
      O => U_DCT2D_rtlc5n1495_19_CYAND
    );
  U_DCT2D_rtlc5n1495_19_CYMUXFAST_1880 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_19_CYMUXG2,
      IB => U_DCT2D_rtlc5n1495_19_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1495_19_CYAND,
      O => U_DCT2D_rtlc5n1495_19_CYMUXFAST
    );
  U_DCT2D_rtlc5n1495_19_CYMUXG2_1881 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1495_19_CY0G,
      IB => U_DCT2D_rtlc5n1495_19_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1495_19_CYSELG,
      O => U_DCT2D_rtlc5n1495_19_CYMUXG2
    );
  U_DCT2D_rtlc5n1495_19_CY0G_1882 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s(13),
      O => U_DCT2D_rtlc5n1495_19_CY0G
    );
  U_DCT2D_rtlc5n1495_19_CYSELG_1883 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z336,
      O => U_DCT2D_rtlc5n1495_19_CYSELG
    );
  U_DCT2D_nx65206z334_rt_1884 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT2D_nx65206z334,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z334_rt
    );
  U_DCT2D_rtlc5n1495_21_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1495_21_XORF,
      O => U_DCT2D_rtlc5n1495(21)
    );
  U_DCT2D_rtlc5n1495_21_XORF_1885 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1495_21_CYINIT,
      I1 => U_DCT2D_nx65206z334_rt,
      O => U_DCT2D_rtlc5n1495_21_XORF
    );
  U_DCT2D_rtlc5n1495_21_CYINIT_1886 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_396_add_68_ix65206z63797_O,
      O => U_DCT2D_rtlc5n1495_21_CYINIT
    );
  U_DCT1D_databuf_reg_6_0_DXMUX_1887 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_0_XORF,
      O => U_DCT1D_databuf_reg_6_0_DXMUX
    );
  U_DCT1D_databuf_reg_6_0_XORF_1888 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_0_CYINIT,
      I1 => U_DCT1D_nx39282z1,
      O => U_DCT1D_databuf_reg_6_0_XORF
    );
  U_DCT1D_databuf_reg_6_0_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_0_CY0F,
      IB => U_DCT1D_databuf_reg_6_0_CYINIT,
      SEL => U_DCT1D_databuf_reg_6_0_CYSELF,
      O => U_DCT1D_rtlc5_85_sub_6_ix40279z63342_O
    );
  U_DCT1D_databuf_reg_6_0_CYINIT_1889 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GLOBAL_LOGIC1_7,
      O => U_DCT1D_databuf_reg_6_0_CYINIT
    );
  U_DCT1D_databuf_reg_6_0_CY0F_1890 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(0),
      O => U_DCT1D_databuf_reg_6_0_CY0F
    );
  U_DCT1D_databuf_reg_6_0_CYSELF_1891 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx39282z1,
      O => U_DCT1D_databuf_reg_6_0_CYSELF
    );
  U_DCT1D_databuf_reg_6_0_DYMUX_1892 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_0_XORG,
      O => U_DCT1D_databuf_reg_6_0_DYMUX
    );
  U_DCT1D_databuf_reg_6_0_XORG_1893 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_85_sub_6_ix40279z63342_O,
      I1 => U_DCT1D_nx40279z1,
      O => U_DCT1D_databuf_reg_6_0_XORG
    );
  U_DCT1D_databuf_reg_6_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_0_CYMUXG,
      O => U_DCT1D_rtlc5_85_sub_6_ix41276z63342_O
    );
  U_DCT1D_databuf_reg_6_0_CYMUXG_1894 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_0_CY0G,
      IB => U_DCT1D_rtlc5_85_sub_6_ix40279z63342_O,
      SEL => U_DCT1D_databuf_reg_6_0_CYSELG,
      O => U_DCT1D_databuf_reg_6_0_CYMUXG
    );
  U_DCT1D_databuf_reg_6_0_CY0G_1895 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(1),
      O => U_DCT1D_databuf_reg_6_0_CY0G
    );
  U_DCT1D_databuf_reg_6_0_CYSELG_1896 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx40279z1,
      O => U_DCT1D_databuf_reg_6_0_CYSELG
    );
  U_DCT1D_databuf_reg_6_0_SRINV_1897 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_6_0_SRINV
    );
  U_DCT1D_databuf_reg_6_0_CLKINV_1898 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_6_0_CLKINV
    );
  U_DCT1D_databuf_reg_6_0_CEINV_1899 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_6_0_CEINV
    );
  U_DCT1D_databuf_reg_6_2_DXMUX_1900 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_2_XORF,
      O => U_DCT1D_databuf_reg_6_2_DXMUX
    );
  U_DCT1D_databuf_reg_6_2_XORF_1901 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_2_CYINIT,
      I1 => U_DCT1D_nx41276z1,
      O => U_DCT1D_databuf_reg_6_2_XORF
    );
  U_DCT1D_databuf_reg_6_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_2_CY0F,
      IB => U_DCT1D_databuf_reg_6_2_CYINIT,
      SEL => U_DCT1D_databuf_reg_6_2_CYSELF,
      O => U_DCT1D_rtlc5_85_sub_6_ix42273z63342_O
    );
  U_DCT1D_databuf_reg_6_2_CYMUXF2_1902 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_2_CY0F,
      IB => U_DCT1D_databuf_reg_6_2_CY0F,
      SEL => U_DCT1D_databuf_reg_6_2_CYSELF,
      O => U_DCT1D_databuf_reg_6_2_CYMUXF2
    );
  U_DCT1D_databuf_reg_6_2_CYINIT_1903 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_85_sub_6_ix41276z63342_O,
      O => U_DCT1D_databuf_reg_6_2_CYINIT
    );
  U_DCT1D_databuf_reg_6_2_CY0F_1904 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(2),
      O => U_DCT1D_databuf_reg_6_2_CY0F
    );
  U_DCT1D_databuf_reg_6_2_CYSELF_1905 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx41276z1,
      O => U_DCT1D_databuf_reg_6_2_CYSELF
    );
  U_DCT1D_databuf_reg_6_2_DYMUX_1906 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_2_XORG,
      O => U_DCT1D_databuf_reg_6_2_DYMUX
    );
  U_DCT1D_databuf_reg_6_2_XORG_1907 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_85_sub_6_ix42273z63342_O,
      I1 => U_DCT1D_nx42273z1,
      O => U_DCT1D_databuf_reg_6_2_XORG
    );
  U_DCT1D_databuf_reg_6_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_2_CYMUXFAST,
      O => U_DCT1D_rtlc5_85_sub_6_ix43270z63342_O
    );
  U_DCT1D_databuf_reg_6_2_FASTCARRY_1908 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_85_sub_6_ix41276z63342_O,
      O => U_DCT1D_databuf_reg_6_2_FASTCARRY
    );
  U_DCT1D_databuf_reg_6_2_CYAND_1909 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_6_2_CYSELG,
      I1 => U_DCT1D_databuf_reg_6_2_CYSELF,
      O => U_DCT1D_databuf_reg_6_2_CYAND
    );
  U_DCT1D_databuf_reg_6_2_CYMUXFAST_1910 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_2_CYMUXG2,
      IB => U_DCT1D_databuf_reg_6_2_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_6_2_CYAND,
      O => U_DCT1D_databuf_reg_6_2_CYMUXFAST
    );
  U_DCT1D_databuf_reg_6_2_CYMUXG2_1911 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_2_CY0G,
      IB => U_DCT1D_databuf_reg_6_2_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_6_2_CYSELG,
      O => U_DCT1D_databuf_reg_6_2_CYMUXG2
    );
  U_DCT1D_databuf_reg_6_2_CY0G_1912 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(3),
      O => U_DCT1D_databuf_reg_6_2_CY0G
    );
  U_DCT1D_databuf_reg_6_2_CYSELG_1913 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx42273z1,
      O => U_DCT1D_databuf_reg_6_2_CYSELG
    );
  U_DCT1D_databuf_reg_6_2_SRINV_1914 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_6_2_SRINV
    );
  U_DCT1D_databuf_reg_6_2_CLKINV_1915 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_6_2_CLKINV
    );
  U_DCT1D_databuf_reg_6_2_CEINV_1916 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_6_2_CEINV
    );
  U_DCT1D_databuf_reg_6_4_DXMUX_1917 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_4_XORF,
      O => U_DCT1D_databuf_reg_6_4_DXMUX
    );
  U_DCT1D_databuf_reg_6_4_XORF_1918 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_4_CYINIT,
      I1 => U_DCT1D_nx43270z1,
      O => U_DCT1D_databuf_reg_6_4_XORF
    );
  U_DCT1D_databuf_reg_6_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_4_CY0F,
      IB => U_DCT1D_databuf_reg_6_4_CYINIT,
      SEL => U_DCT1D_databuf_reg_6_4_CYSELF,
      O => U_DCT1D_rtlc5_85_sub_6_ix44267z63342_O
    );
  U_DCT1D_databuf_reg_6_4_CYMUXF2_1919 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_4_CY0F,
      IB => U_DCT1D_databuf_reg_6_4_CY0F,
      SEL => U_DCT1D_databuf_reg_6_4_CYSELF,
      O => U_DCT1D_databuf_reg_6_4_CYMUXF2
    );
  U_DCT1D_databuf_reg_6_4_CYINIT_1920 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_85_sub_6_ix43270z63342_O,
      O => U_DCT1D_databuf_reg_6_4_CYINIT
    );
  U_DCT1D_databuf_reg_6_4_CY0F_1921 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(4),
      O => U_DCT1D_databuf_reg_6_4_CY0F
    );
  U_DCT1D_databuf_reg_6_4_CYSELF_1922 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx43270z1,
      O => U_DCT1D_databuf_reg_6_4_CYSELF
    );
  U_DCT1D_databuf_reg_6_4_DYMUX_1923 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_4_XORG,
      O => U_DCT1D_databuf_reg_6_4_DYMUX
    );
  U_DCT1D_databuf_reg_6_4_XORG_1924 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_85_sub_6_ix44267z63342_O,
      I1 => U_DCT1D_nx44267z1,
      O => U_DCT1D_databuf_reg_6_4_XORG
    );
  U_DCT1D_databuf_reg_6_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_4_CYMUXFAST,
      O => U_DCT1D_rtlc5_85_sub_6_ix45264z63342_O
    );
  U_DCT1D_databuf_reg_6_4_FASTCARRY_1925 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_85_sub_6_ix43270z63342_O,
      O => U_DCT1D_databuf_reg_6_4_FASTCARRY
    );
  U_DCT1D_databuf_reg_6_4_CYAND_1926 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_6_4_CYSELG,
      I1 => U_DCT1D_databuf_reg_6_4_CYSELF,
      O => U_DCT1D_databuf_reg_6_4_CYAND
    );
  U_DCT1D_databuf_reg_6_4_CYMUXFAST_1927 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_4_CYMUXG2,
      IB => U_DCT1D_databuf_reg_6_4_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_6_4_CYAND,
      O => U_DCT1D_databuf_reg_6_4_CYMUXFAST
    );
  U_DCT1D_databuf_reg_6_4_CYMUXG2_1928 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_4_CY0G,
      IB => U_DCT1D_databuf_reg_6_4_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_6_4_CYSELG,
      O => U_DCT1D_databuf_reg_6_4_CYMUXG2
    );
  U_DCT1D_databuf_reg_6_4_CY0G_1929 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(5),
      O => U_DCT1D_databuf_reg_6_4_CY0G
    );
  U_DCT1D_databuf_reg_6_4_CYSELG_1930 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx44267z1,
      O => U_DCT1D_databuf_reg_6_4_CYSELG
    );
  U_DCT1D_databuf_reg_6_4_SRINV_1931 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_6_4_SRINV
    );
  U_DCT1D_databuf_reg_6_4_CLKINV_1932 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_6_4_CLKINV
    );
  U_DCT1D_databuf_reg_6_4_CEINV_1933 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_6_4_CEINV
    );
  U_DCT1D_databuf_reg_6_6_DXMUX_1934 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_6_XORF,
      O => U_DCT1D_databuf_reg_6_6_DXMUX
    );
  U_DCT1D_databuf_reg_6_6_XORF_1935 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_6_CYINIT,
      I1 => U_DCT1D_nx45264z1,
      O => U_DCT1D_databuf_reg_6_6_XORF
    );
  U_DCT1D_databuf_reg_6_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_6_CY0F,
      IB => U_DCT1D_databuf_reg_6_6_CYINIT,
      SEL => U_DCT1D_databuf_reg_6_6_CYSELF,
      O => U_DCT1D_rtlc5_85_sub_6_ix46261z63342_O
    );
  U_DCT1D_databuf_reg_6_6_CYMUXF2_1936 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_6_CY0F,
      IB => U_DCT1D_databuf_reg_6_6_CY0F,
      SEL => U_DCT1D_databuf_reg_6_6_CYSELF,
      O => U_DCT1D_databuf_reg_6_6_CYMUXF2
    );
  U_DCT1D_databuf_reg_6_6_CYINIT_1937 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_85_sub_6_ix45264z63342_O,
      O => U_DCT1D_databuf_reg_6_6_CYINIT
    );
  U_DCT1D_databuf_reg_6_6_CY0F_1938 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(6),
      O => U_DCT1D_databuf_reg_6_6_CY0F
    );
  U_DCT1D_databuf_reg_6_6_CYSELF_1939 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx45264z1,
      O => U_DCT1D_databuf_reg_6_6_CYSELF
    );
  U_DCT1D_databuf_reg_6_6_DYMUX_1940 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_6_XORG,
      O => U_DCT1D_databuf_reg_6_6_DYMUX
    );
  U_DCT1D_databuf_reg_6_6_XORG_1941 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5_85_sub_6_ix46261z63342_O,
      I1 => U_DCT1D_nx46261z1,
      O => U_DCT1D_databuf_reg_6_6_XORG
    );
  U_DCT1D_databuf_reg_6_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_6_CYMUXFAST,
      O => U_DCT1D_rtlc5_85_sub_6_ix47258z63342_O
    );
  U_DCT1D_databuf_reg_6_6_FASTCARRY_1942 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_85_sub_6_ix45264z63342_O,
      O => U_DCT1D_databuf_reg_6_6_FASTCARRY
    );
  U_DCT1D_databuf_reg_6_6_CYAND_1943 : X_AND2
    port map (
      I0 => U_DCT1D_databuf_reg_6_6_CYSELG,
      I1 => U_DCT1D_databuf_reg_6_6_CYSELF,
      O => U_DCT1D_databuf_reg_6_6_CYAND
    );
  U_DCT1D_databuf_reg_6_6_CYMUXFAST_1944 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_6_CYMUXG2,
      IB => U_DCT1D_databuf_reg_6_6_FASTCARRY,
      SEL => U_DCT1D_databuf_reg_6_6_CYAND,
      O => U_DCT1D_databuf_reg_6_6_CYMUXFAST
    );
  U_DCT1D_databuf_reg_6_6_CYMUXG2_1945 : X_MUX2
    port map (
      IA => U_DCT1D_databuf_reg_6_6_CY0G,
      IB => U_DCT1D_databuf_reg_6_6_CYMUXF2,
      SEL => U_DCT1D_databuf_reg_6_6_CYSELG,
      O => U_DCT1D_databuf_reg_6_6_CYMUXG2
    );
  U_DCT1D_databuf_reg_6_6_CY0G_1946 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(7),
      O => U_DCT1D_databuf_reg_6_6_CY0G
    );
  U_DCT1D_databuf_reg_6_6_CYSELG_1947 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx46261z1,
      O => U_DCT1D_databuf_reg_6_6_CYSELG
    );
  U_DCT1D_databuf_reg_6_6_SRINV_1948 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_6_6_SRINV
    );
  U_DCT1D_databuf_reg_6_6_CLKINV_1949 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_6_6_CLKINV
    );
  U_DCT1D_databuf_reg_6_6_CEINV_1950 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_6_6_CEINV
    );
  U_DCT1D_databuf_reg_6_8_DXMUX_1951 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_8_XORF,
      O => U_DCT1D_databuf_reg_6_8_DXMUX
    );
  U_DCT1D_databuf_reg_6_8_XORF_1952 : X_XOR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_8_CYINIT,
      I1 => U_DCT1D_nx47258z1_rt,
      O => U_DCT1D_databuf_reg_6_8_XORF
    );
  U_DCT1D_databuf_reg_6_8_CYINIT_1953 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_85_sub_6_ix47258z63342_O,
      O => U_DCT1D_databuf_reg_6_8_CYINIT
    );
  U_DCT1D_databuf_reg_6_8_CLKINV_1954 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_databuf_reg_6_8_CLKINV
    );
  U_DCT1D_databuf_reg_6_8_CEINV_1955 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558,
      O => U_DCT1D_databuf_reg_6_8_CEINV
    );
  U_DCT1D_rtlc5n1345_3_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_3_XORF,
      O => U_DCT1D_rtlc5n1345(3)
    );
  U_DCT1D_rtlc5n1345_3_XORF_1956 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1345_3_CYINIT,
      I1 => U_DCT1D_nx59700z162,
      O => U_DCT1D_rtlc5n1345_3_XORF
    );
  U_DCT1D_rtlc5n1345_3_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_3_CY0F,
      IB => U_DCT1D_rtlc5n1345_3_CYINIT,
      SEL => U_DCT1D_rtlc5n1345_3_CYSELF,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63535_O
    );
  U_DCT1D_rtlc5n1345_3_CYINIT_1957 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_3_BXINVNOT,
      O => U_DCT1D_rtlc5n1345_3_CYINIT
    );
  U_DCT1D_rtlc5n1345_3_CY0F_1958 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(1),
      O => U_DCT1D_rtlc5n1345_3_CY0F
    );
  U_DCT1D_rtlc5n1345_3_CYSELF_1959 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z162,
      O => U_DCT1D_rtlc5n1345_3_CYSELF
    );
  U_DCT1D_rtlc5n1345_3_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_1,
      O => U_DCT1D_rtlc5n1345_3_BXINVNOT
    );
  U_DCT1D_rtlc5n1345_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_3_XORG,
      O => U_DCT1D_rtlc5n1345(4)
    );
  U_DCT1D_rtlc5n1345_3_XORG_1960 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_493_add_21_ix59700z63535_O,
      I1 => U_DCT1D_nx59700z159,
      O => U_DCT1D_rtlc5n1345_3_XORG
    );
  U_DCT1D_rtlc5n1345_3_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_3_CYMUXG,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63531_O
    );
  U_DCT1D_rtlc5n1345_3_CYMUXG_1961 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_3_CY0G,
      IB => U_DCT1D_rtlc_493_add_21_ix59700z63535_O,
      SEL => U_DCT1D_rtlc5n1345_3_CYSELG,
      O => U_DCT1D_rtlc5n1345_3_CYMUXG
    );
  U_DCT1D_rtlc5n1345_3_CY0G_1962 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(2),
      O => U_DCT1D_rtlc5n1345_3_CY0G
    );
  U_DCT1D_rtlc5n1345_3_CYSELG_1963 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z159,
      O => U_DCT1D_rtlc5n1345_3_CYSELG
    );
  U_DCT1D_rtlc5n1345_5_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_5_XORF,
      O => U_DCT1D_rtlc5n1345(5)
    );
  U_DCT1D_rtlc5n1345_5_XORF_1964 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1345_5_CYINIT,
      I1 => U_DCT1D_nx59700z156,
      O => U_DCT1D_rtlc5n1345_5_XORF
    );
  U_DCT1D_rtlc5n1345_5_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_5_CY0F,
      IB => U_DCT1D_rtlc5n1345_5_CYINIT,
      SEL => U_DCT1D_rtlc5n1345_5_CYSELF,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63528_O
    );
  U_DCT1D_rtlc5n1345_5_CYMUXF2_1965 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_5_CY0F,
      IB => U_DCT1D_rtlc5n1345_5_CY0F,
      SEL => U_DCT1D_rtlc5n1345_5_CYSELF,
      O => U_DCT1D_rtlc5n1345_5_CYMUXF2
    );
  U_DCT1D_rtlc5n1345_5_CYINIT_1966 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63531_O,
      O => U_DCT1D_rtlc5n1345_5_CYINIT
    );
  U_DCT1D_rtlc5n1345_5_CY0F_1967 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(3),
      O => U_DCT1D_rtlc5n1345_5_CY0F
    );
  U_DCT1D_rtlc5n1345_5_CYSELF_1968 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z156,
      O => U_DCT1D_rtlc5n1345_5_CYSELF
    );
  U_DCT1D_rtlc5n1345_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_5_XORG,
      O => U_DCT1D_rtlc5n1345(6)
    );
  U_DCT1D_rtlc5n1345_5_XORG_1969 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_493_add_21_ix59700z63528_O,
      I1 => U_DCT1D_nx59700z153,
      O => U_DCT1D_rtlc5n1345_5_XORG
    );
  U_DCT1D_rtlc5n1345_5_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_5_CYMUXFAST,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63524_O
    );
  U_DCT1D_rtlc5n1345_5_FASTCARRY_1970 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63531_O,
      O => U_DCT1D_rtlc5n1345_5_FASTCARRY
    );
  U_DCT1D_rtlc5n1345_5_CYAND_1971 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1345_5_CYSELG,
      I1 => U_DCT1D_rtlc5n1345_5_CYSELF,
      O => U_DCT1D_rtlc5n1345_5_CYAND
    );
  U_DCT1D_rtlc5n1345_5_CYMUXFAST_1972 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_5_CYMUXG2,
      IB => U_DCT1D_rtlc5n1345_5_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1345_5_CYAND,
      O => U_DCT1D_rtlc5n1345_5_CYMUXFAST
    );
  U_DCT1D_rtlc5n1345_5_CYMUXG2_1973 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_5_CY0G,
      IB => U_DCT1D_rtlc5n1345_5_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1345_5_CYSELG,
      O => U_DCT1D_rtlc5n1345_5_CYMUXG2
    );
  U_DCT1D_rtlc5n1345_5_CY0G_1974 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(4),
      O => U_DCT1D_rtlc5n1345_5_CY0G
    );
  U_DCT1D_rtlc5n1345_5_CYSELG_1975 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z153,
      O => U_DCT1D_rtlc5n1345_5_CYSELG
    );
  U_DCT1D_ix63810z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_2_Q(4),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_5_Q(4),
      O => U_DCT1D_nx63810z1
    );
  U_DCT1D_rtlc5n1345_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_7_XORF,
      O => U_DCT1D_rtlc5n1345(7)
    );
  U_DCT1D_rtlc5n1345_7_XORF_1976 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1345_7_CYINIT,
      I1 => U_DCT1D_nx59700z150,
      O => U_DCT1D_rtlc5n1345_7_XORF
    );
  U_DCT1D_rtlc5n1345_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_7_CY0F,
      IB => U_DCT1D_rtlc5n1345_7_CYINIT,
      SEL => U_DCT1D_rtlc5n1345_7_CYSELF,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63521_O
    );
  U_DCT1D_rtlc5n1345_7_CYMUXF2_1977 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_7_CY0F,
      IB => U_DCT1D_rtlc5n1345_7_CY0F,
      SEL => U_DCT1D_rtlc5n1345_7_CYSELF,
      O => U_DCT1D_rtlc5n1345_7_CYMUXF2
    );
  U_DCT1D_rtlc5n1345_7_CYINIT_1978 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63524_O,
      O => U_DCT1D_rtlc5n1345_7_CYINIT
    );
  U_DCT1D_rtlc5n1345_7_CY0F_1979 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(5),
      O => U_DCT1D_rtlc5n1345_7_CY0F
    );
  U_DCT1D_rtlc5n1345_7_CYSELF_1980 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z150,
      O => U_DCT1D_rtlc5n1345_7_CYSELF
    );
  U_DCT1D_rtlc5n1345_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_7_XORG,
      O => U_DCT1D_rtlc5n1345(8)
    );
  U_DCT1D_rtlc5n1345_7_XORG_1981 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_493_add_21_ix59700z63521_O,
      I1 => U_DCT1D_nx59700z147,
      O => U_DCT1D_rtlc5n1345_7_XORG
    );
  U_DCT1D_rtlc5n1345_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_7_CYMUXFAST,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63517_O
    );
  U_DCT1D_rtlc5n1345_7_FASTCARRY_1982 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63524_O,
      O => U_DCT1D_rtlc5n1345_7_FASTCARRY
    );
  U_DCT1D_rtlc5n1345_7_CYAND_1983 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1345_7_CYSELG,
      I1 => U_DCT1D_rtlc5n1345_7_CYSELF,
      O => U_DCT1D_rtlc5n1345_7_CYAND
    );
  U_DCT1D_rtlc5n1345_7_CYMUXFAST_1984 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_7_CYMUXG2,
      IB => U_DCT1D_rtlc5n1345_7_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1345_7_CYAND,
      O => U_DCT1D_rtlc5n1345_7_CYMUXFAST
    );
  U_DCT1D_rtlc5n1345_7_CYMUXG2_1985 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_7_CY0G,
      IB => U_DCT1D_rtlc5n1345_7_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1345_7_CYSELG,
      O => U_DCT1D_rtlc5n1345_7_CYMUXG2
    );
  U_DCT1D_rtlc5n1345_7_CY0G_1986 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(6),
      O => U_DCT1D_rtlc5n1345_7_CY0G
    );
  U_DCT1D_rtlc5n1345_7_CYSELG_1987 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z147,
      O => U_DCT1D_rtlc5n1345_7_CYSELG
    );
  U_DCT1D_rtlc5n1345_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_9_XORF,
      O => U_DCT1D_rtlc5n1345(9)
    );
  U_DCT1D_rtlc5n1345_9_XORF_1988 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1345_9_CYINIT,
      I1 => U_DCT1D_nx59700z144,
      O => U_DCT1D_rtlc5n1345_9_XORF
    );
  U_DCT1D_rtlc5n1345_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_9_CY0F,
      IB => U_DCT1D_rtlc5n1345_9_CYINIT,
      SEL => U_DCT1D_rtlc5n1345_9_CYSELF,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63514_O
    );
  U_DCT1D_rtlc5n1345_9_CYMUXF2_1989 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_9_CY0F,
      IB => U_DCT1D_rtlc5n1345_9_CY0F,
      SEL => U_DCT1D_rtlc5n1345_9_CYSELF,
      O => U_DCT1D_rtlc5n1345_9_CYMUXF2
    );
  U_DCT1D_rtlc5n1345_9_CYINIT_1990 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63517_O,
      O => U_DCT1D_rtlc5n1345_9_CYINIT
    );
  U_DCT1D_rtlc5n1345_9_CY0F_1991 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(7),
      O => U_DCT1D_rtlc5n1345_9_CY0F
    );
  U_DCT1D_rtlc5n1345_9_CYSELF_1992 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z144,
      O => U_DCT1D_rtlc5n1345_9_CYSELF
    );
  U_DCT1D_rtlc5n1345_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_9_XORG,
      O => U_DCT1D_rtlc5n1345(10)
    );
  U_DCT1D_rtlc5n1345_9_XORG_1993 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_493_add_21_ix59700z63514_O,
      I1 => U_DCT1D_nx59700z141,
      O => U_DCT1D_rtlc5n1345_9_XORG
    );
  U_DCT1D_rtlc5n1345_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_9_CYMUXFAST,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63510_O
    );
  U_DCT1D_rtlc5n1345_9_FASTCARRY_1994 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63517_O,
      O => U_DCT1D_rtlc5n1345_9_FASTCARRY
    );
  U_DCT1D_rtlc5n1345_9_CYAND_1995 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1345_9_CYSELG,
      I1 => U_DCT1D_rtlc5n1345_9_CYSELF,
      O => U_DCT1D_rtlc5n1345_9_CYAND
    );
  U_DCT1D_rtlc5n1345_9_CYMUXFAST_1996 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_9_CYMUXG2,
      IB => U_DCT1D_rtlc5n1345_9_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1345_9_CYAND,
      O => U_DCT1D_rtlc5n1345_9_CYMUXFAST
    );
  U_DCT1D_rtlc5n1345_9_CYMUXG2_1997 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_9_CY0G,
      IB => U_DCT1D_rtlc5n1345_9_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1345_9_CYSELG,
      O => U_DCT1D_rtlc5n1345_9_CYMUXG2
    );
  U_DCT1D_rtlc5n1345_9_CY0G_1998 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(8),
      O => U_DCT1D_rtlc5n1345_9_CY0G
    );
  U_DCT1D_rtlc5n1345_9_CYSELG_1999 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z141,
      O => U_DCT1D_rtlc5n1345_9_CYSELG
    );
  U_DCT1D_rtlc5n1345_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_11_XORF,
      O => U_DCT1D_rtlc5n1345(11)
    );
  U_DCT1D_rtlc5n1345_11_XORF_2000 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1345_11_CYINIT,
      I1 => U_DCT1D_nx59700z138,
      O => U_DCT1D_rtlc5n1345_11_XORF
    );
  U_DCT1D_rtlc5n1345_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_11_CY0F,
      IB => U_DCT1D_rtlc5n1345_11_CYINIT,
      SEL => U_DCT1D_rtlc5n1345_11_CYSELF,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63506_O
    );
  U_DCT1D_rtlc5n1345_11_CYMUXF2_2001 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_11_CY0F,
      IB => U_DCT1D_rtlc5n1345_11_CY0F,
      SEL => U_DCT1D_rtlc5n1345_11_CYSELF,
      O => U_DCT1D_rtlc5n1345_11_CYMUXF2
    );
  U_DCT1D_rtlc5n1345_11_CYINIT_2002 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63510_O,
      O => U_DCT1D_rtlc5n1345_11_CYINIT
    );
  U_DCT1D_rtlc5n1345_11_CY0F_2003 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(9),
      O => U_DCT1D_rtlc5n1345_11_CY0F
    );
  U_DCT1D_rtlc5n1345_11_CYSELF_2004 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z138,
      O => U_DCT1D_rtlc5n1345_11_CYSELF
    );
  U_DCT1D_rtlc5n1345_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_11_XORG,
      O => U_DCT1D_rtlc5n1345(12)
    );
  U_DCT1D_rtlc5n1345_11_XORG_2005 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_493_add_21_ix59700z63506_O,
      I1 => U_DCT1D_nx59700z135,
      O => U_DCT1D_rtlc5n1345_11_XORG
    );
  U_DCT1D_rtlc5n1345_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_11_CYMUXFAST,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63503_O
    );
  U_DCT1D_rtlc5n1345_11_FASTCARRY_2006 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63510_O,
      O => U_DCT1D_rtlc5n1345_11_FASTCARRY
    );
  U_DCT1D_rtlc5n1345_11_CYAND_2007 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1345_11_CYSELG,
      I1 => U_DCT1D_rtlc5n1345_11_CYSELF,
      O => U_DCT1D_rtlc5n1345_11_CYAND
    );
  U_DCT1D_rtlc5n1345_11_CYMUXFAST_2008 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_11_CYMUXG2,
      IB => U_DCT1D_rtlc5n1345_11_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1345_11_CYAND,
      O => U_DCT1D_rtlc5n1345_11_CYMUXFAST
    );
  U_DCT1D_rtlc5n1345_11_CYMUXG2_2009 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_11_CY0G,
      IB => U_DCT1D_rtlc5n1345_11_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1345_11_CYSELG,
      O => U_DCT1D_rtlc5n1345_11_CYMUXG2
    );
  U_DCT1D_rtlc5n1345_11_CY0G_2010 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(10),
      O => U_DCT1D_rtlc5n1345_11_CY0G
    );
  U_DCT1D_rtlc5n1345_11_CYSELG_2011 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z135,
      O => U_DCT1D_rtlc5n1345_11_CYSELG
    );
  U_DCT1D_rtlc5n1345_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_13_XORF,
      O => U_DCT1D_rtlc5n1345(13)
    );
  U_DCT1D_rtlc5n1345_13_XORF_2012 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1345_13_CYINIT,
      I1 => U_DCT1D_nx59700z132,
      O => U_DCT1D_rtlc5n1345_13_XORF
    );
  U_DCT1D_rtlc5n1345_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_13_CY0F,
      IB => U_DCT1D_rtlc5n1345_13_CYINIT,
      SEL => U_DCT1D_rtlc5n1345_13_CYSELF,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63499_O
    );
  U_DCT1D_rtlc5n1345_13_CYMUXF2_2013 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_13_CY0F,
      IB => U_DCT1D_rtlc5n1345_13_CY0F,
      SEL => U_DCT1D_rtlc5n1345_13_CYSELF,
      O => U_DCT1D_rtlc5n1345_13_CYMUXF2
    );
  U_DCT1D_rtlc5n1345_13_CYINIT_2014 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63503_O,
      O => U_DCT1D_rtlc5n1345_13_CYINIT
    );
  U_DCT1D_rtlc5n1345_13_CY0F_2015 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(11),
      O => U_DCT1D_rtlc5n1345_13_CY0F
    );
  U_DCT1D_rtlc5n1345_13_CYSELF_2016 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z132,
      O => U_DCT1D_rtlc5n1345_13_CYSELF
    );
  U_DCT1D_rtlc5n1345_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_13_XORG,
      O => U_DCT1D_rtlc5n1345(14)
    );
  U_DCT1D_rtlc5n1345_13_XORG_2017 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_493_add_21_ix59700z63499_O,
      I1 => U_DCT1D_nx59700z129,
      O => U_DCT1D_rtlc5n1345_13_XORG
    );
  U_DCT1D_rtlc5n1345_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_13_CYMUXFAST,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63496_O
    );
  U_DCT1D_rtlc5n1345_13_FASTCARRY_2018 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63503_O,
      O => U_DCT1D_rtlc5n1345_13_FASTCARRY
    );
  U_DCT1D_rtlc5n1345_13_CYAND_2019 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1345_13_CYSELG,
      I1 => U_DCT1D_rtlc5n1345_13_CYSELF,
      O => U_DCT1D_rtlc5n1345_13_CYAND
    );
  U_DCT1D_rtlc5n1345_13_CYMUXFAST_2020 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_13_CYMUXG2,
      IB => U_DCT1D_rtlc5n1345_13_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1345_13_CYAND,
      O => U_DCT1D_rtlc5n1345_13_CYMUXFAST
    );
  U_DCT1D_rtlc5n1345_13_CYMUXG2_2021 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_13_CY0G,
      IB => U_DCT1D_rtlc5n1345_13_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1345_13_CYSELG,
      O => U_DCT1D_rtlc5n1345_13_CYMUXG2
    );
  U_DCT1D_rtlc5n1345_13_CY0G_2022 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(12),
      O => U_DCT1D_rtlc5n1345_13_CY0G
    );
  U_DCT1D_rtlc5n1345_13_CYSELG_2023 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z129,
      O => U_DCT1D_rtlc5n1345_13_CYSELG
    );
  U_DCT1D_rtlc5n1345_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_15_XORF,
      O => U_DCT1D_rtlc5n1345(15)
    );
  U_DCT1D_rtlc5n1345_15_XORF_2024 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1345_15_CYINIT,
      I1 => U_DCT1D_nx59700z126,
      O => U_DCT1D_rtlc5n1345_15_XORF
    );
  U_DCT1D_rtlc5n1345_15_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_15_CY0F,
      IB => U_DCT1D_rtlc5n1345_15_CYINIT,
      SEL => U_DCT1D_rtlc5n1345_15_CYSELF,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63492_O
    );
  U_DCT1D_rtlc5n1345_15_CYMUXF2_2025 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_15_CY0F,
      IB => U_DCT1D_rtlc5n1345_15_CY0F,
      SEL => U_DCT1D_rtlc5n1345_15_CYSELF,
      O => U_DCT1D_rtlc5n1345_15_CYMUXF2
    );
  U_DCT1D_rtlc5n1345_15_CYINIT_2026 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63496_O,
      O => U_DCT1D_rtlc5n1345_15_CYINIT
    );
  U_DCT1D_rtlc5n1345_15_CY0F_2027 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(13),
      O => U_DCT1D_rtlc5n1345_15_CY0F
    );
  U_DCT1D_rtlc5n1345_15_CYSELF_2028 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z126,
      O => U_DCT1D_rtlc5n1345_15_CYSELF
    );
  U_DCT1D_rtlc5n1345_15_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_15_XORG,
      O => U_DCT1D_rtlc5n1345(16)
    );
  U_DCT1D_rtlc5n1345_15_XORG_2029 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_493_add_21_ix59700z63492_O,
      I1 => U_DCT1D_nx59700z123,
      O => U_DCT1D_rtlc5n1345_15_XORG
    );
  U_DCT1D_rtlc5n1345_15_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_15_CYMUXFAST,
      O => U_DCT1D_rtlc_493_add_21_ix59700z63489_O
    );
  U_DCT1D_rtlc5n1345_15_FASTCARRY_2030 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63496_O,
      O => U_DCT1D_rtlc5n1345_15_FASTCARRY
    );
  U_DCT1D_rtlc5n1345_15_CYAND_2031 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1345_15_CYSELG,
      I1 => U_DCT1D_rtlc5n1345_15_CYSELF,
      O => U_DCT1D_rtlc5n1345_15_CYAND
    );
  U_DCT1D_rtlc5n1345_15_CYMUXFAST_2032 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_15_CYMUXG2,
      IB => U_DCT1D_rtlc5n1345_15_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1345_15_CYAND,
      O => U_DCT1D_rtlc5n1345_15_CYMUXFAST
    );
  U_DCT1D_rtlc5n1345_15_CYMUXG2_2033 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1345_15_CY0G,
      IB => U_DCT1D_rtlc5n1345_15_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1345_15_CYSELG,
      O => U_DCT1D_rtlc5n1345_15_CYMUXG2
    );
  U_DCT1D_rtlc5n1345_15_CY0G_2034 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s(13),
      O => U_DCT1D_rtlc5n1345_15_CY0G
    );
  U_DCT1D_rtlc5n1345_15_CYSELG_2035 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z123,
      O => U_DCT1D_rtlc5n1345_15_CYSELG
    );
  U_DCT1D_nx59700z121_rt_2036 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z121,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z121_rt
    );
  U_DCT1D_rtlc5n1345_17_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1345_17_XORF,
      O => U_DCT1D_rtlc5n1345(17)
    );
  U_DCT1D_rtlc5n1345_17_XORF_2037 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1345_17_CYINIT,
      I1 => U_DCT1D_nx59700z121_rt,
      O => U_DCT1D_rtlc5n1345_17_XORF
    );
  U_DCT1D_rtlc5n1345_17_CYINIT_2038 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_493_add_21_ix59700z63489_O,
      O => U_DCT1D_rtlc5n1345_17_CYINIT
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CY0F,
      IB => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYINIT,
      SEL => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYSELF,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64143_O
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYINIT_2039 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_BXINVNOT,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYINIT
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CY0F_2040 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z570,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CY0F
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYSELF_2041 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z569,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYSELF
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64139_O_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_35,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_BXINVNOT
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64139_O_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYMUXG,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64139_O
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYMUXG_2042 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CY0G,
      IB => U_DCT2D_rtlc_404_add_70_ix65206z64143_O,
      SEL => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYSELG,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYMUXG
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CY0G_2043 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z567,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CY0G
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYSELG_2044 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z566,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64139_O_CYSELG
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYMUXF2_2045 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CY0F,
      IB => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CY0F,
      SEL => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYSELF,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYMUXF2
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CY0F_2046 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z564,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CY0F
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYSELF_2047 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z563,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYSELF
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64131_O_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYMUXFAST,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64131_O
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64131_O_FASTCARRY_2048 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64139_O,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_FASTCARRY
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYAND_2049 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYSELG,
      I1 => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYSELF,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYAND
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYMUXFAST_2050 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYMUXG2,
      IB => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_FASTCARRY,
      SEL => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYAND,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYMUXFAST
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYMUXG2_2051 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CY0G,
      IB => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYMUXF2,
      SEL => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYSELG,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYMUXG2
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CY0G_2052 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z561,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CY0G
    );
  U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYSELG_2053 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z560,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64131_O_CYSELG
    );
  U_DCT2D_rtlc5n1499_8_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_8_XORF,
      O => U_DCT2D_rtlc5n1499(8)
    );
  U_DCT2D_rtlc5n1499_8_XORF_2054 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1499_8_CYINIT,
      I1 => U_DCT2D_nx65206z556,
      O => U_DCT2D_rtlc5n1499_8_XORF
    );
  U_DCT2D_rtlc5n1499_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_8_CY0F,
      IB => U_DCT2D_rtlc5n1499_8_CYINIT,
      SEL => U_DCT2D_rtlc5n1499_8_CYSELF,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64124_O
    );
  U_DCT2D_rtlc5n1499_8_CYMUXF2_2055 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_8_CY0F,
      IB => U_DCT2D_rtlc5n1499_8_CY0F,
      SEL => U_DCT2D_rtlc5n1499_8_CYSELF,
      O => U_DCT2D_rtlc5n1499_8_CYMUXF2
    );
  U_DCT2D_rtlc5n1499_8_CYINIT_2056 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64131_O,
      O => U_DCT2D_rtlc5n1499_8_CYINIT
    );
  U_DCT2D_rtlc5n1499_8_CY0F_2057 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z557,
      O => U_DCT2D_rtlc5n1499_8_CY0F
    );
  U_DCT2D_rtlc5n1499_8_CYSELF_2058 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z556,
      O => U_DCT2D_rtlc5n1499_8_CYSELF
    );
  U_DCT2D_rtlc5n1499_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_8_XORG,
      O => U_DCT2D_rtlc5n1499(9)
    );
  U_DCT2D_rtlc5n1499_8_XORG_2059 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_404_add_70_ix65206z64124_O,
      I1 => U_DCT2D_nx65206z552,
      O => U_DCT2D_rtlc5n1499_8_XORG
    );
  U_DCT2D_rtlc5n1499_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_8_CYMUXFAST,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64119_O
    );
  U_DCT2D_rtlc5n1499_8_FASTCARRY_2060 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64131_O,
      O => U_DCT2D_rtlc5n1499_8_FASTCARRY
    );
  U_DCT2D_rtlc5n1499_8_CYAND_2061 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1499_8_CYSELG,
      I1 => U_DCT2D_rtlc5n1499_8_CYSELF,
      O => U_DCT2D_rtlc5n1499_8_CYAND
    );
  U_DCT2D_rtlc5n1499_8_CYMUXFAST_2062 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_8_CYMUXG2,
      IB => U_DCT2D_rtlc5n1499_8_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1499_8_CYAND,
      O => U_DCT2D_rtlc5n1499_8_CYMUXFAST
    );
  U_DCT2D_rtlc5n1499_8_CYMUXG2_2063 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_8_CY0G,
      IB => U_DCT2D_rtlc5n1499_8_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1499_8_CYSELG,
      O => U_DCT2D_rtlc5n1499_8_CYMUXG2
    );
  U_DCT2D_rtlc5n1499_8_CY0G_2064 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z553,
      O => U_DCT2D_rtlc5n1499_8_CY0G
    );
  U_DCT2D_rtlc5n1499_8_CYSELG_2065 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z552,
      O => U_DCT2D_rtlc5n1499_8_CYSELG
    );
  U_DCT2D_rtlc5n1499_10_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_10_XORF,
      O => U_DCT2D_rtlc5n1499(10)
    );
  U_DCT2D_rtlc5n1499_10_XORF_2066 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1499_10_CYINIT,
      I1 => U_DCT2D_nx65206z548,
      O => U_DCT2D_rtlc5n1499_10_XORF
    );
  U_DCT2D_rtlc5n1499_10_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_10_CY0F,
      IB => U_DCT2D_rtlc5n1499_10_CYINIT,
      SEL => U_DCT2D_rtlc5n1499_10_CYSELF,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64113_O
    );
  U_DCT2D_rtlc5n1499_10_CYMUXF2_2067 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_10_CY0F,
      IB => U_DCT2D_rtlc5n1499_10_CY0F,
      SEL => U_DCT2D_rtlc5n1499_10_CYSELF,
      O => U_DCT2D_rtlc5n1499_10_CYMUXF2
    );
  U_DCT2D_rtlc5n1499_10_CYINIT_2068 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64119_O,
      O => U_DCT2D_rtlc5n1499_10_CYINIT
    );
  U_DCT2D_rtlc5n1499_10_CY0F_2069 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z549,
      O => U_DCT2D_rtlc5n1499_10_CY0F
    );
  U_DCT2D_rtlc5n1499_10_CYSELF_2070 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z548,
      O => U_DCT2D_rtlc5n1499_10_CYSELF
    );
  U_DCT2D_rtlc5n1499_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_10_XORG,
      O => U_DCT2D_rtlc5n1499(11)
    );
  U_DCT2D_rtlc5n1499_10_XORG_2071 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_404_add_70_ix65206z64113_O,
      I1 => U_DCT2D_nx65206z544,
      O => U_DCT2D_rtlc5n1499_10_XORG
    );
  U_DCT2D_rtlc5n1499_10_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_10_CYMUXFAST,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64108_O
    );
  U_DCT2D_rtlc5n1499_10_FASTCARRY_2072 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64119_O,
      O => U_DCT2D_rtlc5n1499_10_FASTCARRY
    );
  U_DCT2D_rtlc5n1499_10_CYAND_2073 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1499_10_CYSELG,
      I1 => U_DCT2D_rtlc5n1499_10_CYSELF,
      O => U_DCT2D_rtlc5n1499_10_CYAND
    );
  U_DCT2D_rtlc5n1499_10_CYMUXFAST_2074 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_10_CYMUXG2,
      IB => U_DCT2D_rtlc5n1499_10_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1499_10_CYAND,
      O => U_DCT2D_rtlc5n1499_10_CYMUXFAST
    );
  U_DCT2D_rtlc5n1499_10_CYMUXG2_2075 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_10_CY0G,
      IB => U_DCT2D_rtlc5n1499_10_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1499_10_CYSELG,
      O => U_DCT2D_rtlc5n1499_10_CYMUXG2
    );
  U_DCT2D_rtlc5n1499_10_CY0G_2076 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z545,
      O => U_DCT2D_rtlc5n1499_10_CY0G
    );
  U_DCT2D_rtlc5n1499_10_CYSELG_2077 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z544,
      O => U_DCT2D_rtlc5n1499_10_CYSELG
    );
  U_DCT2D_rtlc5n1499_12_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_12_XORF,
      O => U_DCT2D_rtlc5n1499(12)
    );
  U_DCT2D_rtlc5n1499_12_XORF_2078 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1499_12_CYINIT,
      I1 => U_DCT2D_nx65206z540,
      O => U_DCT2D_rtlc5n1499_12_XORF
    );
  U_DCT2D_rtlc5n1499_12_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_12_CY0F,
      IB => U_DCT2D_rtlc5n1499_12_CYINIT,
      SEL => U_DCT2D_rtlc5n1499_12_CYSELF,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64103_O
    );
  U_DCT2D_rtlc5n1499_12_CYMUXF2_2079 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_12_CY0F,
      IB => U_DCT2D_rtlc5n1499_12_CY0F,
      SEL => U_DCT2D_rtlc5n1499_12_CYSELF,
      O => U_DCT2D_rtlc5n1499_12_CYMUXF2
    );
  U_DCT2D_rtlc5n1499_12_CYINIT_2080 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64108_O,
      O => U_DCT2D_rtlc5n1499_12_CYINIT
    );
  U_DCT2D_rtlc5n1499_12_CY0F_2081 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z541,
      O => U_DCT2D_rtlc5n1499_12_CY0F
    );
  U_DCT2D_rtlc5n1499_12_CYSELF_2082 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z540,
      O => U_DCT2D_rtlc5n1499_12_CYSELF
    );
  U_DCT2D_rtlc5n1499_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_12_XORG,
      O => U_DCT2D_rtlc5n1499(13)
    );
  U_DCT2D_rtlc5n1499_12_XORG_2083 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_404_add_70_ix65206z64103_O,
      I1 => U_DCT2D_nx65206z536,
      O => U_DCT2D_rtlc5n1499_12_XORG
    );
  U_DCT2D_rtlc5n1499_12_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_12_CYMUXFAST,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64097_O
    );
  U_DCT2D_rtlc5n1499_12_FASTCARRY_2084 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64108_O,
      O => U_DCT2D_rtlc5n1499_12_FASTCARRY
    );
  U_DCT2D_rtlc5n1499_12_CYAND_2085 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1499_12_CYSELG,
      I1 => U_DCT2D_rtlc5n1499_12_CYSELF,
      O => U_DCT2D_rtlc5n1499_12_CYAND
    );
  U_DCT2D_rtlc5n1499_12_CYMUXFAST_2086 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_12_CYMUXG2,
      IB => U_DCT2D_rtlc5n1499_12_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1499_12_CYAND,
      O => U_DCT2D_rtlc5n1499_12_CYMUXFAST
    );
  U_DCT2D_rtlc5n1499_12_CYMUXG2_2087 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_12_CY0G,
      IB => U_DCT2D_rtlc5n1499_12_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1499_12_CYSELG,
      O => U_DCT2D_rtlc5n1499_12_CYMUXG2
    );
  U_DCT2D_rtlc5n1499_12_CY0G_2088 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z537,
      O => U_DCT2D_rtlc5n1499_12_CY0G
    );
  U_DCT2D_rtlc5n1499_12_CYSELG_2089 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z536,
      O => U_DCT2D_rtlc5n1499_12_CYSELG
    );
  U_DCT2D_rtlc5n1499_14_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_14_XORF,
      O => U_DCT2D_rtlc5n1499(14)
    );
  U_DCT2D_rtlc5n1499_14_XORF_2090 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1499_14_CYINIT,
      I1 => U_DCT2D_nx65206z532,
      O => U_DCT2D_rtlc5n1499_14_XORF
    );
  U_DCT2D_rtlc5n1499_14_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_14_CY0F,
      IB => U_DCT2D_rtlc5n1499_14_CYINIT,
      SEL => U_DCT2D_rtlc5n1499_14_CYSELF,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64092_O
    );
  U_DCT2D_rtlc5n1499_14_CYMUXF2_2091 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_14_CY0F,
      IB => U_DCT2D_rtlc5n1499_14_CY0F,
      SEL => U_DCT2D_rtlc5n1499_14_CYSELF,
      O => U_DCT2D_rtlc5n1499_14_CYMUXF2
    );
  U_DCT2D_rtlc5n1499_14_CYINIT_2092 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64097_O,
      O => U_DCT2D_rtlc5n1499_14_CYINIT
    );
  U_DCT2D_rtlc5n1499_14_CY0F_2093 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z533,
      O => U_DCT2D_rtlc5n1499_14_CY0F
    );
  U_DCT2D_rtlc5n1499_14_CYSELF_2094 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z532,
      O => U_DCT2D_rtlc5n1499_14_CYSELF
    );
  U_DCT2D_rtlc5n1499_14_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_14_XORG,
      O => U_DCT2D_rtlc5n1499(15)
    );
  U_DCT2D_rtlc5n1499_14_XORG_2095 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_404_add_70_ix65206z64092_O,
      I1 => U_DCT2D_nx65206z528,
      O => U_DCT2D_rtlc5n1499_14_XORG
    );
  U_DCT2D_rtlc5n1499_14_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_14_CYMUXFAST,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64087_O
    );
  U_DCT2D_rtlc5n1499_14_FASTCARRY_2096 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64097_O,
      O => U_DCT2D_rtlc5n1499_14_FASTCARRY
    );
  U_DCT2D_rtlc5n1499_14_CYAND_2097 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1499_14_CYSELG,
      I1 => U_DCT2D_rtlc5n1499_14_CYSELF,
      O => U_DCT2D_rtlc5n1499_14_CYAND
    );
  U_DCT2D_rtlc5n1499_14_CYMUXFAST_2098 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_14_CYMUXG2,
      IB => U_DCT2D_rtlc5n1499_14_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1499_14_CYAND,
      O => U_DCT2D_rtlc5n1499_14_CYMUXFAST
    );
  U_DCT2D_rtlc5n1499_14_CYMUXG2_2099 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_14_CY0G,
      IB => U_DCT2D_rtlc5n1499_14_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1499_14_CYSELG,
      O => U_DCT2D_rtlc5n1499_14_CYMUXG2
    );
  U_DCT2D_rtlc5n1499_14_CY0G_2100 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z529,
      O => U_DCT2D_rtlc5n1499_14_CY0G
    );
  U_DCT2D_rtlc5n1499_14_CYSELG_2101 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z528,
      O => U_DCT2D_rtlc5n1499_14_CYSELG
    );
  U_DCT2D_rtlc5n1499_16_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_16_XORF,
      O => U_DCT2D_rtlc5n1499(16)
    );
  U_DCT2D_rtlc5n1499_16_XORF_2102 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1499_16_CYINIT,
      I1 => U_DCT2D_nx65206z524,
      O => U_DCT2D_rtlc5n1499_16_XORF
    );
  U_DCT2D_rtlc5n1499_16_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_16_CY0F,
      IB => U_DCT2D_rtlc5n1499_16_CYINIT,
      SEL => U_DCT2D_rtlc5n1499_16_CYSELF,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64082_O
    );
  U_DCT2D_rtlc5n1499_16_CYMUXF2_2103 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_16_CY0F,
      IB => U_DCT2D_rtlc5n1499_16_CY0F,
      SEL => U_DCT2D_rtlc5n1499_16_CYSELF,
      O => U_DCT2D_rtlc5n1499_16_CYMUXF2
    );
  U_DCT2D_rtlc5n1499_16_CYINIT_2104 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64087_O,
      O => U_DCT2D_rtlc5n1499_16_CYINIT
    );
  U_DCT2D_rtlc5n1499_16_CY0F_2105 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z525,
      O => U_DCT2D_rtlc5n1499_16_CY0F
    );
  U_DCT2D_rtlc5n1499_16_CYSELF_2106 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z524,
      O => U_DCT2D_rtlc5n1499_16_CYSELF
    );
  U_DCT2D_rtlc5n1499_16_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_16_XORG,
      O => U_DCT2D_rtlc5n1499(17)
    );
  U_DCT2D_rtlc5n1499_16_XORG_2107 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_404_add_70_ix65206z64082_O,
      I1 => U_DCT2D_nx65206z520,
      O => U_DCT2D_rtlc5n1499_16_XORG
    );
  U_DCT2D_rtlc5n1499_16_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_16_CYMUXFAST,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64077_O
    );
  U_DCT2D_rtlc5n1499_16_FASTCARRY_2108 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64087_O,
      O => U_DCT2D_rtlc5n1499_16_FASTCARRY
    );
  U_DCT2D_rtlc5n1499_16_CYAND_2109 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1499_16_CYSELG,
      I1 => U_DCT2D_rtlc5n1499_16_CYSELF,
      O => U_DCT2D_rtlc5n1499_16_CYAND
    );
  U_DCT2D_rtlc5n1499_16_CYMUXFAST_2110 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_16_CYMUXG2,
      IB => U_DCT2D_rtlc5n1499_16_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1499_16_CYAND,
      O => U_DCT2D_rtlc5n1499_16_CYMUXFAST
    );
  U_DCT2D_rtlc5n1499_16_CYMUXG2_2111 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_16_CY0G,
      IB => U_DCT2D_rtlc5n1499_16_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1499_16_CYSELG,
      O => U_DCT2D_rtlc5n1499_16_CYMUXG2
    );
  U_DCT2D_rtlc5n1499_16_CY0G_2112 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z521,
      O => U_DCT2D_rtlc5n1499_16_CY0G
    );
  U_DCT2D_rtlc5n1499_16_CYSELG_2113 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z520,
      O => U_DCT2D_rtlc5n1499_16_CYSELG
    );
  U_DCT2D_rtlc5n1499_18_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_18_XORF,
      O => U_DCT2D_rtlc5n1499(18)
    );
  U_DCT2D_rtlc5n1499_18_XORF_2114 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1499_18_CYINIT,
      I1 => U_DCT2D_nx65206z517,
      O => U_DCT2D_rtlc5n1499_18_XORF
    );
  U_DCT2D_rtlc5n1499_18_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_18_CY0F,
      IB => U_DCT2D_rtlc5n1499_18_CYINIT,
      SEL => U_DCT2D_rtlc5n1499_18_CYSELF,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64073_O
    );
  U_DCT2D_rtlc5n1499_18_CYMUXF2_2115 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_18_CY0F,
      IB => U_DCT2D_rtlc5n1499_18_CY0F,
      SEL => U_DCT2D_rtlc5n1499_18_CYSELF,
      O => U_DCT2D_rtlc5n1499_18_CYMUXF2
    );
  U_DCT2D_rtlc5n1499_18_CYINIT_2116 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64077_O,
      O => U_DCT2D_rtlc5n1499_18_CYINIT
    );
  U_DCT2D_rtlc5n1499_18_CY0F_2117 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z3,
      O => U_DCT2D_rtlc5n1499_18_CY0F
    );
  U_DCT2D_rtlc5n1499_18_CYSELF_2118 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z517,
      O => U_DCT2D_rtlc5n1499_18_CYSELF
    );
  U_DCT2D_rtlc5n1499_18_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_18_XORG,
      O => U_DCT2D_rtlc5n1499(19)
    );
  U_DCT2D_rtlc5n1499_18_XORG_2119 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_404_add_70_ix65206z64073_O,
      I1 => U_DCT2D_nx65206z514,
      O => U_DCT2D_rtlc5n1499_18_XORG
    );
  U_DCT2D_rtlc5n1499_18_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_18_CYMUXFAST,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64069_O
    );
  U_DCT2D_rtlc5n1499_18_FASTCARRY_2120 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64077_O,
      O => U_DCT2D_rtlc5n1499_18_FASTCARRY
    );
  U_DCT2D_rtlc5n1499_18_CYAND_2121 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1499_18_CYSELG,
      I1 => U_DCT2D_rtlc5n1499_18_CYSELF,
      O => U_DCT2D_rtlc5n1499_18_CYAND
    );
  U_DCT2D_rtlc5n1499_18_CYMUXFAST_2122 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_18_CYMUXG2,
      IB => U_DCT2D_rtlc5n1499_18_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1499_18_CYAND,
      O => U_DCT2D_rtlc5n1499_18_CYMUXFAST
    );
  U_DCT2D_rtlc5n1499_18_CYMUXG2_2123 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_18_CY0G,
      IB => U_DCT2D_rtlc5n1499_18_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1499_18_CYSELG,
      O => U_DCT2D_rtlc5n1499_18_CYMUXG2
    );
  U_DCT2D_rtlc5n1499_18_CY0G_2124 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z3,
      O => U_DCT2D_rtlc5n1499_18_CY0G
    );
  U_DCT2D_rtlc5n1499_18_CYSELG_2125 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z514,
      O => U_DCT2D_rtlc5n1499_18_CYSELG
    );
  U_DCT2D_rtlc5n1499_20_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_20_XORF,
      O => U_DCT2D_rtlc5n1499(20)
    );
  U_DCT2D_rtlc5n1499_20_XORF_2126 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1499_20_CYINIT,
      I1 => U_DCT2D_nx65206z511,
      O => U_DCT2D_rtlc5n1499_20_XORF
    );
  U_DCT2D_rtlc5n1499_20_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_20_CY0F,
      IB => U_DCT2D_rtlc5n1499_20_CYINIT,
      SEL => U_DCT2D_rtlc5n1499_20_CYSELF,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64065_O
    );
  U_DCT2D_rtlc5n1499_20_CYMUXF2_2127 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_20_CY0F,
      IB => U_DCT2D_rtlc5n1499_20_CY0F,
      SEL => U_DCT2D_rtlc5n1499_20_CYSELF,
      O => U_DCT2D_rtlc5n1499_20_CYMUXF2
    );
  U_DCT2D_rtlc5n1499_20_CYINIT_2128 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64069_O,
      O => U_DCT2D_rtlc5n1499_20_CYINIT
    );
  U_DCT2D_rtlc5n1499_20_CY0F_2129 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z3,
      O => U_DCT2D_rtlc5n1499_20_CY0F
    );
  U_DCT2D_rtlc5n1499_20_CYSELF_2130 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z511,
      O => U_DCT2D_rtlc5n1499_20_CYSELF
    );
  U_DCT2D_rtlc5n1499_20_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_20_XORG,
      O => U_DCT2D_rtlc5n1499(21)
    );
  U_DCT2D_rtlc5n1499_20_XORG_2131 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_404_add_70_ix65206z64065_O,
      I1 => U_DCT2D_nx65206z508,
      O => U_DCT2D_rtlc5n1499_20_XORG
    );
  U_DCT2D_rtlc5n1499_20_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_20_CYMUXFAST,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64060_O
    );
  U_DCT2D_rtlc5n1499_20_FASTCARRY_2132 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64069_O,
      O => U_DCT2D_rtlc5n1499_20_FASTCARRY
    );
  U_DCT2D_rtlc5n1499_20_CYAND_2133 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1499_20_CYSELG,
      I1 => U_DCT2D_rtlc5n1499_20_CYSELF,
      O => U_DCT2D_rtlc5n1499_20_CYAND
    );
  U_DCT2D_rtlc5n1499_20_CYMUXFAST_2134 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_20_CYMUXG2,
      IB => U_DCT2D_rtlc5n1499_20_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1499_20_CYAND,
      O => U_DCT2D_rtlc5n1499_20_CYMUXFAST
    );
  U_DCT2D_rtlc5n1499_20_CYMUXG2_2135 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_20_CY0G,
      IB => U_DCT2D_rtlc5n1499_20_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1499_20_CYSELG,
      O => U_DCT2D_rtlc5n1499_20_CYMUXG2
    );
  U_DCT2D_rtlc5n1499_20_CY0G_2136 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z3,
      O => U_DCT2D_rtlc5n1499_20_CY0G
    );
  U_DCT2D_rtlc5n1499_20_CYSELG_2137 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z508,
      O => U_DCT2D_rtlc5n1499_20_CYSELG
    );
  U_DCT2D_ix65206z1323 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_nx115_bus(18),
      ADR2 => U_DCT2D_nx65206z3,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z2
    );
  U_DCT2D_rtlc5n1499_22_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_22_XORF,
      O => U_DCT2D_rtlc5n1499(22)
    );
  U_DCT2D_rtlc5n1499_22_XORF_2138 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1499_22_CYINIT,
      I1 => U_DCT2D_nx65206z505,
      O => U_DCT2D_rtlc5n1499_22_XORF
    );
  U_DCT2D_rtlc5n1499_22_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1499_22_CY0F,
      IB => U_DCT2D_rtlc5n1499_22_CYINIT,
      SEL => U_DCT2D_rtlc5n1499_22_CYSELF,
      O => U_DCT2D_rtlc_404_add_70_ix65206z64056_O
    );
  U_DCT2D_rtlc5n1499_22_CYINIT_2139 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_404_add_70_ix65206z64060_O,
      O => U_DCT2D_rtlc5n1499_22_CYINIT
    );
  U_DCT2D_rtlc5n1499_22_CY0F_2140 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z3,
      O => U_DCT2D_rtlc5n1499_22_CY0F
    );
  U_DCT2D_rtlc5n1499_22_CYSELF_2141 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z505,
      O => U_DCT2D_rtlc5n1499_22_CYSELF
    );
  U_DCT2D_rtlc5n1499_22_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499_22_XORG,
      O => U_DCT2D_rtlc5n1499(23)
    );
  U_DCT2D_rtlc5n1499_22_XORG_2142 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_404_add_70_ix65206z64056_O,
      I1 => U_DCT2D_nx65206z2,
      O => U_DCT2D_rtlc5n1499_22_XORG
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CY0F,
      IB => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYINIT,
      SEL => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYSELF,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64314_O
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYINIT_2143 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_BXINVNOT,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYINIT
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CY0F_2144 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(8),
      O => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CY0F
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYSELF_2145 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z693,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYSELF
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64310_O_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_38,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_BXINVNOT
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64310_O_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYMUXG,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64310_O
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYMUXG_2146 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CY0G,
      IB => U_DCT2D_rtlc_385_add_63_ix65206z64314_O,
      SEL => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYSELG,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYMUXG
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CY0G_2147 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(9),
      O => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CY0G
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYSELG_2148 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z691,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64310_O_CYSELG
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYMUXF2_2149 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CY0F,
      IB => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CY0F,
      SEL => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYSELF,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYMUXF2
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CY0F_2150 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(10),
      O => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CY0F
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYSELF_2151 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z689,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYSELF
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64302_O_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYMUXFAST,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64302_O
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64302_O_FASTCARRY_2152 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64310_O,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_FASTCARRY
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYAND_2153 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYSELG,
      I1 => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYSELF,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYAND
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYMUXFAST_2154 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYMUXG2,
      IB => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_FASTCARRY,
      SEL => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYAND,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYMUXFAST
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYMUXG2_2155 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CY0G,
      IB => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYMUXF2,
      SEL => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYSELG,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYMUXG2
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CY0G_2156 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(11),
      O => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CY0G
    );
  U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYSELG_2157 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z687,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64302_O_CYSELG
    );
  U_DCT2D_rtlc5n1491_12_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_12_XORF,
      O => U_DCT2D_rtlc5n1491(12)
    );
  U_DCT2D_rtlc5n1491_12_XORF_2158 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1491_12_CYINIT,
      I1 => U_DCT2D_nx65206z684,
      O => U_DCT2D_rtlc5n1491_12_XORF
    );
  U_DCT2D_rtlc5n1491_12_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_12_CY0F,
      IB => U_DCT2D_rtlc5n1491_12_CYINIT,
      SEL => U_DCT2D_rtlc5n1491_12_CYSELF,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64297_O
    );
  U_DCT2D_rtlc5n1491_12_CYMUXF2_2159 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_12_CY0F,
      IB => U_DCT2D_rtlc5n1491_12_CY0F,
      SEL => U_DCT2D_rtlc5n1491_12_CYSELF,
      O => U_DCT2D_rtlc5n1491_12_CYMUXF2
    );
  U_DCT2D_rtlc5n1491_12_CYINIT_2160 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64302_O,
      O => U_DCT2D_rtlc5n1491_12_CYINIT
    );
  U_DCT2D_rtlc5n1491_12_CY0F_2161 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(12),
      O => U_DCT2D_rtlc5n1491_12_CY0F
    );
  U_DCT2D_rtlc5n1491_12_CYSELF_2162 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z684,
      O => U_DCT2D_rtlc5n1491_12_CYSELF
    );
  U_DCT2D_rtlc5n1491_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_12_XORG,
      O => U_DCT2D_rtlc5n1491(13)
    );
  U_DCT2D_rtlc5n1491_12_XORG_2163 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_385_add_63_ix65206z64297_O,
      I1 => U_DCT2D_nx65206z681,
      O => U_DCT2D_rtlc5n1491_12_XORG
    );
  U_DCT2D_rtlc5n1491_12_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_12_CYMUXFAST,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64290_O
    );
  U_DCT2D_rtlc5n1491_12_FASTCARRY_2164 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64302_O,
      O => U_DCT2D_rtlc5n1491_12_FASTCARRY
    );
  U_DCT2D_rtlc5n1491_12_CYAND_2165 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1491_12_CYSELG,
      I1 => U_DCT2D_rtlc5n1491_12_CYSELF,
      O => U_DCT2D_rtlc5n1491_12_CYAND
    );
  U_DCT2D_rtlc5n1491_12_CYMUXFAST_2166 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_12_CYMUXG2,
      IB => U_DCT2D_rtlc5n1491_12_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1491_12_CYAND,
      O => U_DCT2D_rtlc5n1491_12_CYMUXFAST
    );
  U_DCT2D_rtlc5n1491_12_CYMUXG2_2167 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_12_CY0G,
      IB => U_DCT2D_rtlc5n1491_12_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1491_12_CYSELG,
      O => U_DCT2D_rtlc5n1491_12_CYMUXG2
    );
  U_DCT2D_rtlc5n1491_12_CY0G_2168 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(13),
      O => U_DCT2D_rtlc5n1491_12_CY0G
    );
  U_DCT2D_rtlc5n1491_12_CYSELG_2169 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z681,
      O => U_DCT2D_rtlc5n1491_12_CYSELG
    );
  U_DCT2D_rtlc5n1491_14_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_14_XORF,
      O => U_DCT2D_rtlc5n1491(14)
    );
  U_DCT2D_rtlc5n1491_14_XORF_2170 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1491_14_CYINIT,
      I1 => U_DCT2D_nx65206z678,
      O => U_DCT2D_rtlc5n1491_14_XORF
    );
  U_DCT2D_rtlc5n1491_14_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_14_CY0F,
      IB => U_DCT2D_rtlc5n1491_14_CYINIT,
      SEL => U_DCT2D_rtlc5n1491_14_CYSELF,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64285_O
    );
  U_DCT2D_rtlc5n1491_14_CYMUXF2_2171 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_14_CY0F,
      IB => U_DCT2D_rtlc5n1491_14_CY0F,
      SEL => U_DCT2D_rtlc5n1491_14_CYSELF,
      O => U_DCT2D_rtlc5n1491_14_CYMUXF2
    );
  U_DCT2D_rtlc5n1491_14_CYINIT_2172 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64290_O,
      O => U_DCT2D_rtlc5n1491_14_CYINIT
    );
  U_DCT2D_rtlc5n1491_14_CY0F_2173 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(14),
      O => U_DCT2D_rtlc5n1491_14_CY0F
    );
  U_DCT2D_rtlc5n1491_14_CYSELF_2174 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z678,
      O => U_DCT2D_rtlc5n1491_14_CYSELF
    );
  U_DCT2D_rtlc5n1491_14_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_14_XORG,
      O => U_DCT2D_rtlc5n1491(15)
    );
  U_DCT2D_rtlc5n1491_14_XORG_2175 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_385_add_63_ix65206z64285_O,
      I1 => U_DCT2D_nx65206z675,
      O => U_DCT2D_rtlc5n1491_14_XORG
    );
  U_DCT2D_rtlc5n1491_14_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_14_CYMUXFAST,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64280_O
    );
  U_DCT2D_rtlc5n1491_14_FASTCARRY_2176 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64290_O,
      O => U_DCT2D_rtlc5n1491_14_FASTCARRY
    );
  U_DCT2D_rtlc5n1491_14_CYAND_2177 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1491_14_CYSELG,
      I1 => U_DCT2D_rtlc5n1491_14_CYSELF,
      O => U_DCT2D_rtlc5n1491_14_CYAND
    );
  U_DCT2D_rtlc5n1491_14_CYMUXFAST_2178 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_14_CYMUXG2,
      IB => U_DCT2D_rtlc5n1491_14_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1491_14_CYAND,
      O => U_DCT2D_rtlc5n1491_14_CYMUXFAST
    );
  U_DCT2D_rtlc5n1491_14_CYMUXG2_2179 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_14_CY0G,
      IB => U_DCT2D_rtlc5n1491_14_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1491_14_CYSELG,
      O => U_DCT2D_rtlc5n1491_14_CYMUXG2
    );
  U_DCT2D_rtlc5n1491_14_CY0G_2180 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(15),
      O => U_DCT2D_rtlc5n1491_14_CY0G
    );
  U_DCT2D_rtlc5n1491_14_CYSELG_2181 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z675,
      O => U_DCT2D_rtlc5n1491_14_CYSELG
    );
  U_DCT1D_reg_databuf_reg_2_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_2_4_DXMUX,
      CE => U_DCT1D_databuf_reg_2_4_CEINV,
      CLK => U_DCT1D_databuf_reg_2_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_2_4_FFX_RST,
      O => U_DCT1D_databuf_reg_2_Q(4)
    );
  U_DCT1D_databuf_reg_2_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_2_4_FFX_RST
    );
  U_DCT2D_rtlc5n1491_16_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_16_XORF,
      O => U_DCT2D_rtlc5n1491(16)
    );
  U_DCT2D_rtlc5n1491_16_XORF_2182 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1491_16_CYINIT,
      I1 => U_DCT2D_nx65206z672,
      O => U_DCT2D_rtlc5n1491_16_XORF
    );
  U_DCT2D_rtlc5n1491_16_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_16_CY0F,
      IB => U_DCT2D_rtlc5n1491_16_CYINIT,
      SEL => U_DCT2D_rtlc5n1491_16_CYSELF,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64275_O
    );
  U_DCT2D_rtlc5n1491_16_CYMUXF2_2183 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_16_CY0F,
      IB => U_DCT2D_rtlc5n1491_16_CY0F,
      SEL => U_DCT2D_rtlc5n1491_16_CYSELF,
      O => U_DCT2D_rtlc5n1491_16_CYMUXF2
    );
  U_DCT2D_rtlc5n1491_16_CYINIT_2184 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64280_O,
      O => U_DCT2D_rtlc5n1491_16_CYINIT
    );
  U_DCT2D_rtlc5n1491_16_CY0F_2185 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(16),
      O => U_DCT2D_rtlc5n1491_16_CY0F
    );
  U_DCT2D_rtlc5n1491_16_CYSELF_2186 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z672,
      O => U_DCT2D_rtlc5n1491_16_CYSELF
    );
  U_DCT2D_rtlc5n1491_16_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_16_XORG,
      O => U_DCT2D_rtlc5n1491(17)
    );
  U_DCT2D_rtlc5n1491_16_XORG_2187 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_385_add_63_ix65206z64275_O,
      I1 => U_DCT2D_nx65206z669,
      O => U_DCT2D_rtlc5n1491_16_XORG
    );
  U_DCT2D_rtlc5n1491_16_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_16_CYMUXFAST,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64270_O
    );
  U_DCT2D_rtlc5n1491_16_FASTCARRY_2188 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64280_O,
      O => U_DCT2D_rtlc5n1491_16_FASTCARRY
    );
  U_DCT2D_rtlc5n1491_16_CYAND_2189 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1491_16_CYSELG,
      I1 => U_DCT2D_rtlc5n1491_16_CYSELF,
      O => U_DCT2D_rtlc5n1491_16_CYAND
    );
  U_DCT2D_rtlc5n1491_16_CYMUXFAST_2190 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_16_CYMUXG2,
      IB => U_DCT2D_rtlc5n1491_16_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1491_16_CYAND,
      O => U_DCT2D_rtlc5n1491_16_CYMUXFAST
    );
  U_DCT2D_rtlc5n1491_16_CYMUXG2_2191 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_16_CY0G,
      IB => U_DCT2D_rtlc5n1491_16_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1491_16_CYSELG,
      O => U_DCT2D_rtlc5n1491_16_CYMUXG2
    );
  U_DCT2D_rtlc5n1491_16_CY0G_2192 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(17),
      O => U_DCT2D_rtlc5n1491_16_CY0G
    );
  U_DCT2D_rtlc5n1491_16_CYSELG_2193 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z669,
      O => U_DCT2D_rtlc5n1491_16_CYSELG
    );
  U_DCT2D_rtlc5n1491_18_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_18_XORF,
      O => U_DCT2D_rtlc5n1491(18)
    );
  U_DCT2D_rtlc5n1491_18_XORF_2194 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1491_18_CYINIT,
      I1 => U_DCT2D_nx65206z666,
      O => U_DCT2D_rtlc5n1491_18_XORF
    );
  U_DCT2D_rtlc5n1491_18_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_18_CY0F,
      IB => U_DCT2D_rtlc5n1491_18_CYINIT,
      SEL => U_DCT2D_rtlc5n1491_18_CYSELF,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64265_O
    );
  U_DCT2D_rtlc5n1491_18_CYMUXF2_2195 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_18_CY0F,
      IB => U_DCT2D_rtlc5n1491_18_CY0F,
      SEL => U_DCT2D_rtlc5n1491_18_CYSELF,
      O => U_DCT2D_rtlc5n1491_18_CYMUXF2
    );
  U_DCT2D_rtlc5n1491_18_CYINIT_2196 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64270_O,
      O => U_DCT2D_rtlc5n1491_18_CYINIT
    );
  U_DCT2D_rtlc5n1491_18_CY0F_2197 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(18),
      O => U_DCT2D_rtlc5n1491_18_CY0F
    );
  U_DCT2D_rtlc5n1491_18_CYSELF_2198 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z666,
      O => U_DCT2D_rtlc5n1491_18_CYSELF
    );
  U_DCT2D_rtlc5n1491_18_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_18_XORG,
      O => U_DCT2D_rtlc5n1491(19)
    );
  U_DCT2D_rtlc5n1491_18_XORG_2199 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_385_add_63_ix65206z64265_O,
      I1 => U_DCT2D_nx65206z663,
      O => U_DCT2D_rtlc5n1491_18_XORG
    );
  U_DCT2D_rtlc5n1491_18_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_18_CYMUXFAST,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64260_O
    );
  U_DCT2D_rtlc5n1491_18_FASTCARRY_2200 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64270_O,
      O => U_DCT2D_rtlc5n1491_18_FASTCARRY
    );
  U_DCT2D_rtlc5n1491_18_CYAND_2201 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1491_18_CYSELG,
      I1 => U_DCT2D_rtlc5n1491_18_CYSELF,
      O => U_DCT2D_rtlc5n1491_18_CYAND
    );
  U_DCT2D_rtlc5n1491_18_CYMUXFAST_2202 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_18_CYMUXG2,
      IB => U_DCT2D_rtlc5n1491_18_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1491_18_CYAND,
      O => U_DCT2D_rtlc5n1491_18_CYMUXFAST
    );
  U_DCT2D_rtlc5n1491_18_CYMUXG2_2203 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_18_CY0G,
      IB => U_DCT2D_rtlc5n1491_18_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1491_18_CYSELG,
      O => U_DCT2D_rtlc5n1491_18_CYMUXG2
    );
  U_DCT2D_rtlc5n1491_18_CY0G_2204 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(19),
      O => U_DCT2D_rtlc5n1491_18_CY0G
    );
  U_DCT2D_rtlc5n1491_18_CYSELG_2205 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z663,
      O => U_DCT2D_rtlc5n1491_18_CYSELG
    );
  U_DCT2D_rtlc5n1491_20_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_20_XORF,
      O => U_DCT2D_rtlc5n1491(20)
    );
  U_DCT2D_rtlc5n1491_20_XORF_2206 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1491_20_CYINIT,
      I1 => U_DCT2D_nx65206z660,
      O => U_DCT2D_rtlc5n1491_20_XORF
    );
  U_DCT2D_rtlc5n1491_20_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_20_CY0F,
      IB => U_DCT2D_rtlc5n1491_20_CYINIT,
      SEL => U_DCT2D_rtlc5n1491_20_CYSELF,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64253_O
    );
  U_DCT2D_rtlc5n1491_20_CYMUXF2_2207 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_20_CY0F,
      IB => U_DCT2D_rtlc5n1491_20_CY0F,
      SEL => U_DCT2D_rtlc5n1491_20_CYSELF,
      O => U_DCT2D_rtlc5n1491_20_CYMUXF2
    );
  U_DCT2D_rtlc5n1491_20_CYINIT_2208 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64260_O,
      O => U_DCT2D_rtlc5n1491_20_CYINIT
    );
  U_DCT2D_rtlc5n1491_20_CY0F_2209 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(20),
      O => U_DCT2D_rtlc5n1491_20_CY0F
    );
  U_DCT2D_rtlc5n1491_20_CYSELF_2210 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z660,
      O => U_DCT2D_rtlc5n1491_20_CYSELF
    );
  U_DCT2D_rtlc5n1491_20_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_20_XORG,
      O => U_DCT2D_rtlc5n1491(21)
    );
  U_DCT2D_rtlc5n1491_20_XORG_2211 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_385_add_63_ix65206z64253_O,
      I1 => U_DCT2D_nx65206z657,
      O => U_DCT2D_rtlc5n1491_20_XORG
    );
  U_DCT2D_rtlc5n1491_20_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_20_CYMUXFAST,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64248_O
    );
  U_DCT2D_rtlc5n1491_20_FASTCARRY_2212 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64260_O,
      O => U_DCT2D_rtlc5n1491_20_FASTCARRY
    );
  U_DCT2D_rtlc5n1491_20_CYAND_2213 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1491_20_CYSELG,
      I1 => U_DCT2D_rtlc5n1491_20_CYSELF,
      O => U_DCT2D_rtlc5n1491_20_CYAND
    );
  U_DCT2D_rtlc5n1491_20_CYMUXFAST_2214 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_20_CYMUXG2,
      IB => U_DCT2D_rtlc5n1491_20_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1491_20_CYAND,
      O => U_DCT2D_rtlc5n1491_20_CYMUXFAST
    );
  U_DCT2D_rtlc5n1491_20_CYMUXG2_2215 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_20_CY0G,
      IB => U_DCT2D_rtlc5n1491_20_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1491_20_CYSELG,
      O => U_DCT2D_rtlc5n1491_20_CYMUXG2
    );
  U_DCT2D_rtlc5n1491_20_CY0G_2216 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(21),
      O => U_DCT2D_rtlc5n1491_20_CY0G
    );
  U_DCT2D_rtlc5n1491_20_CYSELG_2217 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z657,
      O => U_DCT2D_rtlc5n1491_20_CYSELG
    );
  U_DCT2D_rtlc5n1491_22_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_22_XORF,
      O => U_DCT2D_rtlc5n1491(22)
    );
  U_DCT2D_rtlc5n1491_22_XORF_2218 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1491_22_CYINIT,
      I1 => U_DCT2D_nx65206z654,
      O => U_DCT2D_rtlc5n1491_22_XORF
    );
  U_DCT2D_rtlc5n1491_22_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1491_22_CY0F,
      IB => U_DCT2D_rtlc5n1491_22_CYINIT,
      SEL => U_DCT2D_rtlc5n1491_22_CYSELF,
      O => U_DCT2D_rtlc_385_add_63_ix65206z64243_O
    );
  U_DCT2D_rtlc5n1491_22_CYINIT_2219 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_385_add_63_ix65206z64248_O,
      O => U_DCT2D_rtlc5n1491_22_CYINIT
    );
  U_DCT2D_rtlc5n1491_22_CY0F_2220 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1499(22),
      O => U_DCT2D_rtlc5n1491_22_CY0F
    );
  U_DCT2D_rtlc5n1491_22_CYSELF_2221 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z654,
      O => U_DCT2D_rtlc5n1491_22_CYSELF
    );
  U_DCT2D_rtlc5n1491_22_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491_22_XORG,
      O => U_DCT2D_rtlc5n1491(23)
    );
  U_DCT2D_rtlc5n1491_22_XORG_2222 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_385_add_63_ix65206z64243_O,
      I1 => U_DCT2D_nx65206z1_rt,
      O => U_DCT2D_rtlc5n1491_22_XORG
    );
  U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CY0F,
      IB => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYINIT,
      SEL => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYSELF,
      O => U_DCT1D_rtlc_508_add_26_ix59700z64004_O
    );
  U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYINIT_2223 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_BXINVNOT,
      O => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYINIT
    );
  U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CY0F_2224 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z493,
      O => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CY0F
    );
  U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYSELF_2225 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z492,
      O => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYSELF
    );
  U_DCT1D_rtlc_508_add_26_ix59700z64000_O_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_15,
      O => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_BXINVNOT
    );
  U_DCT1D_rtlc_508_add_26_ix59700z64000_O_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYMUXG,
      O => U_DCT1D_rtlc_508_add_26_ix59700z64000_O
    );
  U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYMUXG_2226 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CY0G,
      IB => U_DCT1D_rtlc_508_add_26_ix59700z64004_O,
      SEL => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYSELG,
      O => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYMUXG
    );
  U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CY0G_2227 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z490,
      O => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CY0G
    );
  U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYSELG_2228 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z489,
      O => U_DCT1D_rtlc_508_add_26_ix59700z64000_O_CYSELG
    );
  U_DCT1D_ix59700z1973 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1359(7),
      ADR1 => U_DCT1D_nx59700z484,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z483
    );
  U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYMUXF2_2229 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CY0F,
      IB => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CY0F,
      SEL => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYSELF,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYMUXF2
    );
  U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CY0F_2230 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z487,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CY0F
    );
  U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYSELF_2231 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z486,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYSELF
    );
  U_DCT1D_rtlc_508_add_26_ix59700z63992_O_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYMUXFAST,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63992_O
    );
  U_DCT1D_rtlc_508_add_26_ix59700z63992_O_FASTCARRY_2232 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z64000_O,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_FASTCARRY
    );
  U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYAND_2233 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYSELG,
      I1 => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYSELF,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYAND
    );
  U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYMUXFAST_2234 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYMUXG2,
      IB => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_FASTCARRY,
      SEL => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYAND,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYMUXFAST
    );
  U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYMUXG2_2235 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CY0G,
      IB => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYMUXF2,
      SEL => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYSELG,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYMUXG2
    );
  U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CY0G_2236 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z484,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CY0G
    );
  U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYSELG_2237 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z483,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63992_O_CYSELG
    );
  U_DCT1D_rtlc5n1350_8_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_8_XORF,
      O => U_DCT1D_rtlc5n1350(8)
    );
  U_DCT1D_rtlc5n1350_8_XORF_2238 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1350_8_CYINIT,
      I1 => U_DCT1D_nx59700z479,
      O => U_DCT1D_rtlc5n1350_8_XORF
    );
  U_DCT1D_rtlc5n1350_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_8_CY0F,
      IB => U_DCT1D_rtlc5n1350_8_CYINIT,
      SEL => U_DCT1D_rtlc5n1350_8_CYSELF,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63985_O
    );
  U_DCT1D_rtlc5n1350_8_CYMUXF2_2239 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_8_CY0F,
      IB => U_DCT1D_rtlc5n1350_8_CY0F,
      SEL => U_DCT1D_rtlc5n1350_8_CYSELF,
      O => U_DCT1D_rtlc5n1350_8_CYMUXF2
    );
  U_DCT1D_rtlc5n1350_8_CYINIT_2240 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63992_O,
      O => U_DCT1D_rtlc5n1350_8_CYINIT
    );
  U_DCT1D_rtlc5n1350_8_CY0F_2241 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z480,
      O => U_DCT1D_rtlc5n1350_8_CY0F
    );
  U_DCT1D_rtlc5n1350_8_CYSELF_2242 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z479,
      O => U_DCT1D_rtlc5n1350_8_CYSELF
    );
  U_DCT1D_rtlc5n1350_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_8_XORG,
      O => U_DCT1D_rtlc5n1350(9)
    );
  U_DCT1D_rtlc5n1350_8_XORG_2243 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_508_add_26_ix59700z63985_O,
      I1 => U_DCT1D_nx59700z475,
      O => U_DCT1D_rtlc5n1350_8_XORG
    );
  U_DCT1D_rtlc5n1350_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_8_CYMUXFAST,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63980_O
    );
  U_DCT1D_rtlc5n1350_8_FASTCARRY_2244 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63992_O,
      O => U_DCT1D_rtlc5n1350_8_FASTCARRY
    );
  U_DCT1D_rtlc5n1350_8_CYAND_2245 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1350_8_CYSELG,
      I1 => U_DCT1D_rtlc5n1350_8_CYSELF,
      O => U_DCT1D_rtlc5n1350_8_CYAND
    );
  U_DCT1D_rtlc5n1350_8_CYMUXFAST_2246 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_8_CYMUXG2,
      IB => U_DCT1D_rtlc5n1350_8_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1350_8_CYAND,
      O => U_DCT1D_rtlc5n1350_8_CYMUXFAST
    );
  U_DCT1D_rtlc5n1350_8_CYMUXG2_2247 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_8_CY0G,
      IB => U_DCT1D_rtlc5n1350_8_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1350_8_CYSELG,
      O => U_DCT1D_rtlc5n1350_8_CYMUXG2
    );
  U_DCT1D_rtlc5n1350_8_CY0G_2248 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z476,
      O => U_DCT1D_rtlc5n1350_8_CY0G
    );
  U_DCT1D_rtlc5n1350_8_CYSELG_2249 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z475,
      O => U_DCT1D_rtlc5n1350_8_CYSELG
    );
  U_DCT1D_rtlc5n1350_10_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_10_XORF,
      O => U_DCT1D_rtlc5n1350(10)
    );
  U_DCT1D_rtlc5n1350_10_XORF_2250 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1350_10_CYINIT,
      I1 => U_DCT1D_nx59700z471,
      O => U_DCT1D_rtlc5n1350_10_XORF
    );
  U_DCT1D_rtlc5n1350_10_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_10_CY0F,
      IB => U_DCT1D_rtlc5n1350_10_CYINIT,
      SEL => U_DCT1D_rtlc5n1350_10_CYSELF,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63973_O
    );
  U_DCT1D_rtlc5n1350_10_CYMUXF2_2251 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_10_CY0F,
      IB => U_DCT1D_rtlc5n1350_10_CY0F,
      SEL => U_DCT1D_rtlc5n1350_10_CYSELF,
      O => U_DCT1D_rtlc5n1350_10_CYMUXF2
    );
  U_DCT1D_rtlc5n1350_10_CYINIT_2252 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63980_O,
      O => U_DCT1D_rtlc5n1350_10_CYINIT
    );
  U_DCT1D_rtlc5n1350_10_CY0F_2253 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z472,
      O => U_DCT1D_rtlc5n1350_10_CY0F
    );
  U_DCT1D_rtlc5n1350_10_CYSELF_2254 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z471,
      O => U_DCT1D_rtlc5n1350_10_CYSELF
    );
  U_DCT1D_rtlc5n1350_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_10_XORG,
      O => U_DCT1D_rtlc5n1350(11)
    );
  U_DCT1D_rtlc5n1350_10_XORG_2255 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_508_add_26_ix59700z63973_O,
      I1 => U_DCT1D_nx59700z467,
      O => U_DCT1D_rtlc5n1350_10_XORG
    );
  U_DCT1D_rtlc5n1350_10_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_10_CYMUXFAST,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63968_O
    );
  U_DCT1D_rtlc5n1350_10_FASTCARRY_2256 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63980_O,
      O => U_DCT1D_rtlc5n1350_10_FASTCARRY
    );
  U_DCT1D_rtlc5n1350_10_CYAND_2257 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1350_10_CYSELG,
      I1 => U_DCT1D_rtlc5n1350_10_CYSELF,
      O => U_DCT1D_rtlc5n1350_10_CYAND
    );
  U_DCT1D_rtlc5n1350_10_CYMUXFAST_2258 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_10_CYMUXG2,
      IB => U_DCT1D_rtlc5n1350_10_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1350_10_CYAND,
      O => U_DCT1D_rtlc5n1350_10_CYMUXFAST
    );
  U_DCT1D_rtlc5n1350_10_CYMUXG2_2259 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_10_CY0G,
      IB => U_DCT1D_rtlc5n1350_10_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1350_10_CYSELG,
      O => U_DCT1D_rtlc5n1350_10_CYMUXG2
    );
  U_DCT1D_rtlc5n1350_10_CY0G_2260 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z468,
      O => U_DCT1D_rtlc5n1350_10_CY0G
    );
  U_DCT1D_rtlc5n1350_10_CYSELG_2261 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z467,
      O => U_DCT1D_rtlc5n1350_10_CYSELG
    );
  U_DCT1D_rtlc5n1350_12_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_12_XORF,
      O => U_DCT1D_rtlc5n1350(12)
    );
  U_DCT1D_rtlc5n1350_12_XORF_2262 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1350_12_CYINIT,
      I1 => U_DCT1D_nx59700z463,
      O => U_DCT1D_rtlc5n1350_12_XORF
    );
  U_DCT1D_rtlc5n1350_12_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_12_CY0F,
      IB => U_DCT1D_rtlc5n1350_12_CYINIT,
      SEL => U_DCT1D_rtlc5n1350_12_CYSELF,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63962_O
    );
  U_DCT1D_rtlc5n1350_12_CYMUXF2_2263 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_12_CY0F,
      IB => U_DCT1D_rtlc5n1350_12_CY0F,
      SEL => U_DCT1D_rtlc5n1350_12_CYSELF,
      O => U_DCT1D_rtlc5n1350_12_CYMUXF2
    );
  U_DCT1D_rtlc5n1350_12_CYINIT_2264 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63968_O,
      O => U_DCT1D_rtlc5n1350_12_CYINIT
    );
  U_DCT1D_rtlc5n1350_12_CY0F_2265 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z464,
      O => U_DCT1D_rtlc5n1350_12_CY0F
    );
  U_DCT1D_rtlc5n1350_12_CYSELF_2266 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z463,
      O => U_DCT1D_rtlc5n1350_12_CYSELF
    );
  U_DCT1D_rtlc5n1350_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_12_XORG,
      O => U_DCT1D_rtlc5n1350(13)
    );
  U_DCT1D_rtlc5n1350_12_XORG_2267 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_508_add_26_ix59700z63962_O,
      I1 => U_DCT1D_nx59700z459,
      O => U_DCT1D_rtlc5n1350_12_XORG
    );
  U_DCT1D_rtlc5n1350_12_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_12_CYMUXFAST,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63957_O
    );
  U_DCT1D_rtlc5n1350_12_FASTCARRY_2268 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63968_O,
      O => U_DCT1D_rtlc5n1350_12_FASTCARRY
    );
  U_DCT1D_rtlc5n1350_12_CYAND_2269 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1350_12_CYSELG,
      I1 => U_DCT1D_rtlc5n1350_12_CYSELF,
      O => U_DCT1D_rtlc5n1350_12_CYAND
    );
  U_DCT1D_rtlc5n1350_12_CYMUXFAST_2270 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_12_CYMUXG2,
      IB => U_DCT1D_rtlc5n1350_12_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1350_12_CYAND,
      O => U_DCT1D_rtlc5n1350_12_CYMUXFAST
    );
  U_DCT1D_rtlc5n1350_12_CYMUXG2_2271 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_12_CY0G,
      IB => U_DCT1D_rtlc5n1350_12_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1350_12_CYSELG,
      O => U_DCT1D_rtlc5n1350_12_CYMUXG2
    );
  U_DCT1D_rtlc5n1350_12_CY0G_2272 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z460,
      O => U_DCT1D_rtlc5n1350_12_CY0G
    );
  U_DCT1D_rtlc5n1350_12_CYSELG_2273 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z459,
      O => U_DCT1D_rtlc5n1350_12_CYSELG
    );
  U_DCT1D_rtlc5n1350_14_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_14_XORF,
      O => U_DCT1D_rtlc5n1350(14)
    );
  U_DCT1D_rtlc5n1350_14_XORF_2274 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1350_14_CYINIT,
      I1 => U_DCT1D_nx59700z455,
      O => U_DCT1D_rtlc5n1350_14_XORF
    );
  U_DCT1D_rtlc5n1350_14_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_14_CY0F,
      IB => U_DCT1D_rtlc5n1350_14_CYINIT,
      SEL => U_DCT1D_rtlc5n1350_14_CYSELF,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63952_O
    );
  U_DCT1D_rtlc5n1350_14_CYMUXF2_2275 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_14_CY0F,
      IB => U_DCT1D_rtlc5n1350_14_CY0F,
      SEL => U_DCT1D_rtlc5n1350_14_CYSELF,
      O => U_DCT1D_rtlc5n1350_14_CYMUXF2
    );
  U_DCT1D_rtlc5n1350_14_CYINIT_2276 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63957_O,
      O => U_DCT1D_rtlc5n1350_14_CYINIT
    );
  U_DCT1D_rtlc5n1350_14_CY0F_2277 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z456,
      O => U_DCT1D_rtlc5n1350_14_CY0F
    );
  U_DCT1D_rtlc5n1350_14_CYSELF_2278 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z455,
      O => U_DCT1D_rtlc5n1350_14_CYSELF
    );
  U_DCT1D_rtlc5n1350_14_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_14_XORG,
      O => U_DCT1D_rtlc5n1350(15)
    );
  U_DCT1D_rtlc5n1350_14_XORG_2279 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_508_add_26_ix59700z63952_O,
      I1 => U_DCT1D_nx59700z451,
      O => U_DCT1D_rtlc5n1350_14_XORG
    );
  U_DCT1D_rtlc5n1350_14_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_14_CYMUXFAST,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63947_O
    );
  U_DCT1D_rtlc5n1350_14_FASTCARRY_2280 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63957_O,
      O => U_DCT1D_rtlc5n1350_14_FASTCARRY
    );
  U_DCT1D_rtlc5n1350_14_CYAND_2281 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1350_14_CYSELG,
      I1 => U_DCT1D_rtlc5n1350_14_CYSELF,
      O => U_DCT1D_rtlc5n1350_14_CYAND
    );
  U_DCT1D_rtlc5n1350_14_CYMUXFAST_2282 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_14_CYMUXG2,
      IB => U_DCT1D_rtlc5n1350_14_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1350_14_CYAND,
      O => U_DCT1D_rtlc5n1350_14_CYMUXFAST
    );
  U_DCT1D_rtlc5n1350_14_CYMUXG2_2283 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_14_CY0G,
      IB => U_DCT1D_rtlc5n1350_14_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1350_14_CYSELG,
      O => U_DCT1D_rtlc5n1350_14_CYMUXG2
    );
  U_DCT1D_rtlc5n1350_14_CY0G_2284 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z452,
      O => U_DCT1D_rtlc5n1350_14_CY0G
    );
  U_DCT1D_rtlc5n1350_14_CYSELG_2285 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z451,
      O => U_DCT1D_rtlc5n1350_14_CYSELG
    );
  U_DCT1D_rtlc5n1350_16_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_16_XORF,
      O => U_DCT1D_rtlc5n1350(16)
    );
  U_DCT1D_rtlc5n1350_16_XORF_2286 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1350_16_CYINIT,
      I1 => U_DCT1D_nx59700z447,
      O => U_DCT1D_rtlc5n1350_16_XORF
    );
  U_DCT1D_rtlc5n1350_16_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_16_CY0F,
      IB => U_DCT1D_rtlc5n1350_16_CYINIT,
      SEL => U_DCT1D_rtlc5n1350_16_CYSELF,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63942_O
    );
  U_DCT1D_rtlc5n1350_16_CYMUXF2_2287 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_16_CY0F,
      IB => U_DCT1D_rtlc5n1350_16_CY0F,
      SEL => U_DCT1D_rtlc5n1350_16_CYSELF,
      O => U_DCT1D_rtlc5n1350_16_CYMUXF2
    );
  U_DCT1D_rtlc5n1350_16_CYINIT_2288 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63947_O,
      O => U_DCT1D_rtlc5n1350_16_CYINIT
    );
  U_DCT1D_rtlc5n1350_16_CY0F_2289 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z448,
      O => U_DCT1D_rtlc5n1350_16_CY0F
    );
  U_DCT1D_rtlc5n1350_16_CYSELF_2290 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z447,
      O => U_DCT1D_rtlc5n1350_16_CYSELF
    );
  U_DCT1D_rtlc5n1350_16_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_16_XORG,
      O => U_DCT1D_rtlc5n1350(17)
    );
  U_DCT1D_rtlc5n1350_16_XORG_2291 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_508_add_26_ix59700z63942_O,
      I1 => U_DCT1D_nx59700z443,
      O => U_DCT1D_rtlc5n1350_16_XORG
    );
  U_DCT1D_rtlc5n1350_16_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_16_CYMUXFAST,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63937_O
    );
  U_DCT1D_rtlc5n1350_16_FASTCARRY_2292 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63947_O,
      O => U_DCT1D_rtlc5n1350_16_FASTCARRY
    );
  U_DCT1D_rtlc5n1350_16_CYAND_2293 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1350_16_CYSELG,
      I1 => U_DCT1D_rtlc5n1350_16_CYSELF,
      O => U_DCT1D_rtlc5n1350_16_CYAND
    );
  U_DCT1D_rtlc5n1350_16_CYMUXFAST_2294 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_16_CYMUXG2,
      IB => U_DCT1D_rtlc5n1350_16_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1350_16_CYAND,
      O => U_DCT1D_rtlc5n1350_16_CYMUXFAST
    );
  U_DCT1D_rtlc5n1350_16_CYMUXG2_2295 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_16_CY0G,
      IB => U_DCT1D_rtlc5n1350_16_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1350_16_CYSELG,
      O => U_DCT1D_rtlc5n1350_16_CYMUXG2
    );
  U_DCT1D_rtlc5n1350_16_CY0G_2296 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z444,
      O => U_DCT1D_rtlc5n1350_16_CY0G
    );
  U_DCT1D_rtlc5n1350_16_CYSELG_2297 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z443,
      O => U_DCT1D_rtlc5n1350_16_CYSELG
    );
  U_DCT1D_rtlc5n1350_18_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_18_XORF,
      O => U_DCT1D_rtlc5n1350(18)
    );
  U_DCT1D_rtlc5n1350_18_XORF_2298 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1350_18_CYINIT,
      I1 => U_DCT1D_nx59700z440,
      O => U_DCT1D_rtlc5n1350_18_XORF
    );
  U_DCT1D_rtlc5n1350_18_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_18_CY0F,
      IB => U_DCT1D_rtlc5n1350_18_CYINIT,
      SEL => U_DCT1D_rtlc5n1350_18_CYSELF,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63933_O
    );
  U_DCT1D_rtlc5n1350_18_CYMUXF2_2299 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_18_CY0F,
      IB => U_DCT1D_rtlc5n1350_18_CY0F,
      SEL => U_DCT1D_rtlc5n1350_18_CYSELF,
      O => U_DCT1D_rtlc5n1350_18_CYMUXF2
    );
  U_DCT1D_rtlc5n1350_18_CYINIT_2300 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63937_O,
      O => U_DCT1D_rtlc5n1350_18_CYINIT
    );
  U_DCT1D_rtlc5n1350_18_CY0F_2301 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z3,
      O => U_DCT1D_rtlc5n1350_18_CY0F
    );
  U_DCT1D_rtlc5n1350_18_CYSELF_2302 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z440,
      O => U_DCT1D_rtlc5n1350_18_CYSELF
    );
  U_DCT1D_rtlc5n1350_18_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_18_XORG,
      O => U_DCT1D_rtlc5n1350(19)
    );
  U_DCT1D_rtlc5n1350_18_XORG_2303 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_508_add_26_ix59700z63933_O,
      I1 => U_DCT1D_nx59700z437,
      O => U_DCT1D_rtlc5n1350_18_XORG
    );
  U_DCT1D_rtlc5n1350_18_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_18_CYMUXFAST,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63929_O
    );
  U_DCT1D_rtlc5n1350_18_FASTCARRY_2304 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63937_O,
      O => U_DCT1D_rtlc5n1350_18_FASTCARRY
    );
  U_DCT1D_rtlc5n1350_18_CYAND_2305 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1350_18_CYSELG,
      I1 => U_DCT1D_rtlc5n1350_18_CYSELF,
      O => U_DCT1D_rtlc5n1350_18_CYAND
    );
  U_DCT1D_rtlc5n1350_18_CYMUXFAST_2306 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_18_CYMUXG2,
      IB => U_DCT1D_rtlc5n1350_18_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1350_18_CYAND,
      O => U_DCT1D_rtlc5n1350_18_CYMUXFAST
    );
  U_DCT1D_rtlc5n1350_18_CYMUXG2_2307 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_18_CY0G,
      IB => U_DCT1D_rtlc5n1350_18_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1350_18_CYSELG,
      O => U_DCT1D_rtlc5n1350_18_CYMUXG2
    );
  U_DCT1D_rtlc5n1350_18_CY0G_2308 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z3,
      O => U_DCT1D_rtlc5n1350_18_CY0G
    );
  U_DCT1D_rtlc5n1350_18_CYSELG_2309 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z437,
      O => U_DCT1D_rtlc5n1350_18_CYSELG
    );
  U_DCT1D_ix1265z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_2_Q(7),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_5_Q(7),
      O => U_DCT1D_nx1265z1
    );
  U_DCT1D_rtlc5n1350_20_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_20_XORF,
      O => U_DCT1D_rtlc5n1350(20)
    );
  U_DCT1D_rtlc5n1350_20_XORF_2310 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1350_20_CYINIT,
      I1 => U_DCT1D_nx59700z434,
      O => U_DCT1D_rtlc5n1350_20_XORF
    );
  U_DCT1D_rtlc5n1350_20_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1350_20_CY0F,
      IB => U_DCT1D_rtlc5n1350_20_CYINIT,
      SEL => U_DCT1D_rtlc5n1350_20_CYSELF,
      O => U_DCT1D_rtlc_508_add_26_ix59700z63925_O
    );
  U_DCT1D_rtlc5n1350_20_CYINIT_2311 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_508_add_26_ix59700z63929_O,
      O => U_DCT1D_rtlc5n1350_20_CYINIT
    );
  U_DCT1D_rtlc5n1350_20_CY0F_2312 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z3,
      O => U_DCT1D_rtlc5n1350_20_CY0F
    );
  U_DCT1D_rtlc5n1350_20_CYSELF_2313 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z434,
      O => U_DCT1D_rtlc5n1350_20_CYSELF
    );
  U_DCT1D_rtlc5n1350_20_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350_20_XORG,
      O => U_DCT1D_rtlc5n1350(21)
    );
  U_DCT1D_rtlc5n1350_20_XORG_2314 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_508_add_26_ix59700z63925_O,
      I1 => U_DCT1D_nx59700z2,
      O => U_DCT1D_rtlc5n1350_20_XORG
    );
  U_DCT1D_rtlc5n1355_5_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_5_XORF,
      O => U_DCT1D_rtlc5n1355(5)
    );
  U_DCT1D_rtlc5n1355_5_XORF_2315 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1355_5_CYINIT,
      I1 => U_DCT1D_nx59700z40,
      O => U_DCT1D_rtlc5n1355_5_XORF
    );
  U_DCT1D_rtlc5n1355_5_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_5_CY0F,
      IB => U_DCT1D_rtlc5n1355_5_CYINIT,
      SEL => U_DCT1D_rtlc5n1355_5_CYSELF,
      O => U_DCT1D_rtlc_512_add_28_ix59700z63386_O
    );
  U_DCT1D_rtlc5n1355_5_CYINIT_2316 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_5_BXINVNOT,
      O => U_DCT1D_rtlc5n1355_5_CYINIT
    );
  U_DCT1D_rtlc5n1355_5_CY0F_2317 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s(3),
      O => U_DCT1D_rtlc5n1355_5_CY0F
    );
  U_DCT1D_rtlc5n1355_5_CYSELF_2318 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z40,
      O => U_DCT1D_rtlc5n1355_5_CYSELF
    );
  U_DCT1D_rtlc5n1355_5_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_14,
      O => U_DCT1D_rtlc5n1355_5_BXINVNOT
    );
  U_DCT1D_rtlc5n1355_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_5_XORG,
      O => U_DCT1D_rtlc5n1355(6)
    );
  U_DCT1D_rtlc5n1355_5_XORG_2319 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_512_add_28_ix59700z63386_O,
      I1 => U_DCT1D_nx59700z37,
      O => U_DCT1D_rtlc5n1355_5_XORG
    );
  U_DCT1D_rtlc5n1355_5_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_5_CYMUXG,
      O => U_DCT1D_rtlc_512_add_28_ix59700z63383_O
    );
  U_DCT1D_rtlc5n1355_5_CYMUXG_2320 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_5_CY0G,
      IB => U_DCT1D_rtlc_512_add_28_ix59700z63386_O,
      SEL => U_DCT1D_rtlc5n1355_5_CYSELG,
      O => U_DCT1D_rtlc5n1355_5_CYMUXG
    );
  U_DCT1D_rtlc5n1355_5_CY0G_2321 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s(4),
      O => U_DCT1D_rtlc5n1355_5_CY0G
    );
  U_DCT1D_rtlc5n1355_5_CYSELG_2322 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z37,
      O => U_DCT1D_rtlc5n1355_5_CYSELG
    );
  U_DCT1D_rtlc5n1355_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_7_XORF,
      O => U_DCT1D_rtlc5n1355(7)
    );
  U_DCT1D_rtlc5n1355_7_XORF_2323 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1355_7_CYINIT,
      I1 => U_DCT1D_nx59700z34,
      O => U_DCT1D_rtlc5n1355_7_XORF
    );
  U_DCT1D_rtlc5n1355_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_7_CY0F,
      IB => U_DCT1D_rtlc5n1355_7_CYINIT,
      SEL => U_DCT1D_rtlc5n1355_7_CYSELF,
      O => U_DCT1D_rtlc_512_add_28_ix59700z63379_O
    );
  U_DCT1D_rtlc5n1355_7_CYMUXF2_2324 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_7_CY0F,
      IB => U_DCT1D_rtlc5n1355_7_CY0F,
      SEL => U_DCT1D_rtlc5n1355_7_CYSELF,
      O => U_DCT1D_rtlc5n1355_7_CYMUXF2
    );
  U_DCT1D_rtlc5n1355_7_CYINIT_2325 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_512_add_28_ix59700z63383_O,
      O => U_DCT1D_rtlc5n1355_7_CYINIT
    );
  U_DCT1D_rtlc5n1355_7_CY0F_2326 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s(5),
      O => U_DCT1D_rtlc5n1355_7_CY0F
    );
  U_DCT1D_rtlc5n1355_7_CYSELF_2327 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z34,
      O => U_DCT1D_rtlc5n1355_7_CYSELF
    );
  U_DCT1D_rtlc5n1355_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_7_XORG,
      O => U_DCT1D_rtlc5n1355(8)
    );
  U_DCT1D_rtlc5n1355_7_XORG_2328 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_512_add_28_ix59700z63379_O,
      I1 => U_DCT1D_nx59700z31,
      O => U_DCT1D_rtlc5n1355_7_XORG
    );
  U_DCT1D_rtlc5n1355_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_7_CYMUXFAST,
      O => U_DCT1D_rtlc_512_add_28_ix59700z63376_O
    );
  U_DCT1D_rtlc5n1355_7_FASTCARRY_2329 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_512_add_28_ix59700z63383_O,
      O => U_DCT1D_rtlc5n1355_7_FASTCARRY
    );
  U_DCT1D_rtlc5n1355_7_CYAND_2330 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1355_7_CYSELG,
      I1 => U_DCT1D_rtlc5n1355_7_CYSELF,
      O => U_DCT1D_rtlc5n1355_7_CYAND
    );
  U_DCT1D_rtlc5n1355_7_CYMUXFAST_2331 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_7_CYMUXG2,
      IB => U_DCT1D_rtlc5n1355_7_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1355_7_CYAND,
      O => U_DCT1D_rtlc5n1355_7_CYMUXFAST
    );
  U_DCT1D_rtlc5n1355_7_CYMUXG2_2332 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_7_CY0G,
      IB => U_DCT1D_rtlc5n1355_7_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1355_7_CYSELG,
      O => U_DCT1D_rtlc5n1355_7_CYMUXG2
    );
  U_DCT1D_rtlc5n1355_7_CY0G_2333 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s(6),
      O => U_DCT1D_rtlc5n1355_7_CY0G
    );
  U_DCT1D_rtlc5n1355_7_CYSELG_2334 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z31,
      O => U_DCT1D_rtlc5n1355_7_CYSELG
    );
  U_DCT1D_rtlc5n1355_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_9_XORF,
      O => U_DCT1D_rtlc5n1355(9)
    );
  U_DCT1D_rtlc5n1355_9_XORF_2335 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1355_9_CYINIT,
      I1 => U_DCT1D_nx59700z28,
      O => U_DCT1D_rtlc5n1355_9_XORF
    );
  U_DCT1D_rtlc5n1355_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_9_CY0F,
      IB => U_DCT1D_rtlc5n1355_9_CYINIT,
      SEL => U_DCT1D_rtlc5n1355_9_CYSELF,
      O => U_DCT1D_rtlc_512_add_28_ix59700z63372_O
    );
  U_DCT1D_rtlc5n1355_9_CYMUXF2_2336 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_9_CY0F,
      IB => U_DCT1D_rtlc5n1355_9_CY0F,
      SEL => U_DCT1D_rtlc5n1355_9_CYSELF,
      O => U_DCT1D_rtlc5n1355_9_CYMUXF2
    );
  U_DCT1D_rtlc5n1355_9_CYINIT_2337 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_512_add_28_ix59700z63376_O,
      O => U_DCT1D_rtlc5n1355_9_CYINIT
    );
  U_DCT1D_rtlc5n1355_9_CY0F_2338 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s(7),
      O => U_DCT1D_rtlc5n1355_9_CY0F
    );
  U_DCT1D_rtlc5n1355_9_CYSELF_2339 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z28,
      O => U_DCT1D_rtlc5n1355_9_CYSELF
    );
  U_DCT1D_rtlc5n1355_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_9_XORG,
      O => U_DCT1D_rtlc5n1355(10)
    );
  U_DCT1D_rtlc5n1355_9_XORG_2340 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_512_add_28_ix59700z63372_O,
      I1 => U_DCT1D_nx59700z25,
      O => U_DCT1D_rtlc5n1355_9_XORG
    );
  U_DCT1D_rtlc5n1355_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_9_CYMUXFAST,
      O => U_DCT1D_rtlc_512_add_28_ix59700z63369_O
    );
  U_DCT1D_rtlc5n1355_9_FASTCARRY_2341 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_512_add_28_ix59700z63376_O,
      O => U_DCT1D_rtlc5n1355_9_FASTCARRY
    );
  U_DCT1D_rtlc5n1355_9_CYAND_2342 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1355_9_CYSELG,
      I1 => U_DCT1D_rtlc5n1355_9_CYSELF,
      O => U_DCT1D_rtlc5n1355_9_CYAND
    );
  U_DCT1D_rtlc5n1355_9_CYMUXFAST_2343 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_9_CYMUXG2,
      IB => U_DCT1D_rtlc5n1355_9_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1355_9_CYAND,
      O => U_DCT1D_rtlc5n1355_9_CYMUXFAST
    );
  U_DCT1D_rtlc5n1355_9_CYMUXG2_2344 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_9_CY0G,
      IB => U_DCT1D_rtlc5n1355_9_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1355_9_CYSELG,
      O => U_DCT1D_rtlc5n1355_9_CYMUXG2
    );
  U_DCT1D_rtlc5n1355_9_CY0G_2345 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s(8),
      O => U_DCT1D_rtlc5n1355_9_CY0G
    );
  U_DCT1D_rtlc5n1355_9_CYSELG_2346 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z25,
      O => U_DCT1D_rtlc5n1355_9_CYSELG
    );
  U_DCT1D_rtlc5n1355_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_11_XORF,
      O => U_DCT1D_rtlc5n1355(11)
    );
  U_DCT1D_rtlc5n1355_11_XORF_2347 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1355_11_CYINIT,
      I1 => U_DCT1D_nx59700z22,
      O => U_DCT1D_rtlc5n1355_11_XORF
    );
  U_DCT1D_rtlc5n1355_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_11_CY0F,
      IB => U_DCT1D_rtlc5n1355_11_CYINIT,
      SEL => U_DCT1D_rtlc5n1355_11_CYSELF,
      O => U_DCT1D_rtlc_512_add_28_ix59700z63365_O
    );
  U_DCT1D_rtlc5n1355_11_CYMUXF2_2348 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_11_CY0F,
      IB => U_DCT1D_rtlc5n1355_11_CY0F,
      SEL => U_DCT1D_rtlc5n1355_11_CYSELF,
      O => U_DCT1D_rtlc5n1355_11_CYMUXF2
    );
  U_DCT1D_rtlc5n1355_11_CYINIT_2349 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_512_add_28_ix59700z63369_O,
      O => U_DCT1D_rtlc5n1355_11_CYINIT
    );
  U_DCT1D_rtlc5n1355_11_CY0F_2350 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s(9),
      O => U_DCT1D_rtlc5n1355_11_CY0F
    );
  U_DCT1D_rtlc5n1355_11_CYSELF_2351 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z22,
      O => U_DCT1D_rtlc5n1355_11_CYSELF
    );
  U_DCT1D_rtlc5n1355_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_11_XORG,
      O => U_DCT1D_rtlc5n1355(12)
    );
  U_DCT1D_rtlc5n1355_11_XORG_2352 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_512_add_28_ix59700z63365_O,
      I1 => U_DCT1D_nx59700z19,
      O => U_DCT1D_rtlc5n1355_11_XORG
    );
  U_DCT1D_rtlc5n1355_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_11_CYMUXFAST,
      O => U_DCT1D_rtlc_512_add_28_ix59700z63362_O
    );
  U_DCT1D_rtlc5n1355_11_FASTCARRY_2353 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_512_add_28_ix59700z63369_O,
      O => U_DCT1D_rtlc5n1355_11_FASTCARRY
    );
  U_DCT1D_rtlc5n1355_11_CYAND_2354 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1355_11_CYSELG,
      I1 => U_DCT1D_rtlc5n1355_11_CYSELF,
      O => U_DCT1D_rtlc5n1355_11_CYAND
    );
  U_DCT1D_rtlc5n1355_11_CYMUXFAST_2355 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_11_CYMUXG2,
      IB => U_DCT1D_rtlc5n1355_11_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1355_11_CYAND,
      O => U_DCT1D_rtlc5n1355_11_CYMUXFAST
    );
  U_DCT1D_rtlc5n1355_11_CYMUXG2_2356 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_11_CY0G,
      IB => U_DCT1D_rtlc5n1355_11_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1355_11_CYSELG,
      O => U_DCT1D_rtlc5n1355_11_CYMUXG2
    );
  U_DCT1D_rtlc5n1355_11_CY0G_2357 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s(10),
      O => U_DCT1D_rtlc5n1355_11_CY0G
    );
  U_DCT1D_rtlc5n1355_11_CYSELG_2358 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z19,
      O => U_DCT1D_rtlc5n1355_11_CYSELG
    );
  U_DCT1D_rtlc5n1355_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_13_XORF,
      O => U_DCT1D_rtlc5n1355(13)
    );
  U_DCT1D_rtlc5n1355_13_XORF_2359 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1355_13_CYINIT,
      I1 => U_DCT1D_nx59700z16,
      O => U_DCT1D_rtlc5n1355_13_XORF
    );
  U_DCT1D_rtlc5n1355_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_13_CY0F,
      IB => U_DCT1D_rtlc5n1355_13_CYINIT,
      SEL => U_DCT1D_rtlc5n1355_13_CYSELF,
      O => U_DCT1D_rtlc_512_add_28_ix59700z63358_O
    );
  U_DCT1D_rtlc5n1355_13_CYMUXF2_2360 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_13_CY0F,
      IB => U_DCT1D_rtlc5n1355_13_CY0F,
      SEL => U_DCT1D_rtlc5n1355_13_CYSELF,
      O => U_DCT1D_rtlc5n1355_13_CYMUXF2
    );
  U_DCT1D_rtlc5n1355_13_CYINIT_2361 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_512_add_28_ix59700z63362_O,
      O => U_DCT1D_rtlc5n1355_13_CYINIT
    );
  U_DCT1D_rtlc5n1355_13_CY0F_2362 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s(11),
      O => U_DCT1D_rtlc5n1355_13_CY0F
    );
  U_DCT1D_rtlc5n1355_13_CYSELF_2363 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z16,
      O => U_DCT1D_rtlc5n1355_13_CYSELF
    );
  U_DCT1D_rtlc5n1355_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_13_XORG,
      O => U_DCT1D_rtlc5n1355(14)
    );
  U_DCT1D_rtlc5n1355_13_XORG_2364 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_512_add_28_ix59700z63358_O,
      I1 => U_DCT1D_nx59700z13,
      O => U_DCT1D_rtlc5n1355_13_XORG
    );
  U_DCT1D_rtlc5n1355_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_13_CYMUXFAST,
      O => U_DCT1D_rtlc_512_add_28_ix59700z63355_O
    );
  U_DCT1D_rtlc5n1355_13_FASTCARRY_2365 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_512_add_28_ix59700z63362_O,
      O => U_DCT1D_rtlc5n1355_13_FASTCARRY
    );
  U_DCT1D_rtlc5n1355_13_CYAND_2366 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1355_13_CYSELG,
      I1 => U_DCT1D_rtlc5n1355_13_CYSELF,
      O => U_DCT1D_rtlc5n1355_13_CYAND
    );
  U_DCT1D_rtlc5n1355_13_CYMUXFAST_2367 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_13_CYMUXG2,
      IB => U_DCT1D_rtlc5n1355_13_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1355_13_CYAND,
      O => U_DCT1D_rtlc5n1355_13_CYMUXFAST
    );
  U_DCT1D_rtlc5n1355_13_CYMUXG2_2368 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_13_CY0G,
      IB => U_DCT1D_rtlc5n1355_13_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1355_13_CYSELG,
      O => U_DCT1D_rtlc5n1355_13_CYMUXG2
    );
  U_DCT1D_rtlc5n1355_13_CY0G_2369 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s(12),
      O => U_DCT1D_rtlc5n1355_13_CY0G
    );
  U_DCT1D_rtlc5n1355_13_CYSELG_2370 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z13,
      O => U_DCT1D_rtlc5n1355_13_CYSELG
    );
  U_DCT1D_rtlc5n1355_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_15_XORF,
      O => U_DCT1D_rtlc5n1355(15)
    );
  U_DCT1D_rtlc5n1355_15_XORF_2371 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1355_15_CYINIT,
      I1 => U_DCT1D_nx59700z10,
      O => U_DCT1D_rtlc5n1355_15_XORF
    );
  U_DCT1D_rtlc5n1355_15_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_15_CY0F,
      IB => U_DCT1D_rtlc5n1355_15_CYINIT,
      SEL => U_DCT1D_rtlc5n1355_15_CYSELF,
      O => U_DCT1D_rtlc_512_add_28_ix59700z63351_O
    );
  U_DCT1D_rtlc5n1355_15_CYMUXF2_2372 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_15_CY0F,
      IB => U_DCT1D_rtlc5n1355_15_CY0F,
      SEL => U_DCT1D_rtlc5n1355_15_CYSELF,
      O => U_DCT1D_rtlc5n1355_15_CYMUXF2
    );
  U_DCT1D_rtlc5n1355_15_CYINIT_2373 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_512_add_28_ix59700z63355_O,
      O => U_DCT1D_rtlc5n1355_15_CYINIT
    );
  U_DCT1D_rtlc5n1355_15_CY0F_2374 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s(13),
      O => U_DCT1D_rtlc5n1355_15_CY0F
    );
  U_DCT1D_rtlc5n1355_15_CYSELF_2375 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z10,
      O => U_DCT1D_rtlc5n1355_15_CYSELF
    );
  U_DCT1D_rtlc5n1355_15_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_15_XORG,
      O => U_DCT1D_rtlc5n1355(16)
    );
  U_DCT1D_rtlc5n1355_15_XORG_2376 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_512_add_28_ix59700z63351_O,
      I1 => U_DCT1D_nx59700z7,
      O => U_DCT1D_rtlc5n1355_15_XORG
    );
  U_DCT1D_rtlc5n1355_15_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_15_CYMUXFAST,
      O => U_DCT1D_rtlc_512_add_28_ix59700z63348_O
    );
  U_DCT1D_rtlc5n1355_15_FASTCARRY_2377 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_512_add_28_ix59700z63355_O,
      O => U_DCT1D_rtlc5n1355_15_FASTCARRY
    );
  U_DCT1D_rtlc5n1355_15_CYAND_2378 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1355_15_CYSELG,
      I1 => U_DCT1D_rtlc5n1355_15_CYSELF,
      O => U_DCT1D_rtlc5n1355_15_CYAND
    );
  U_DCT1D_rtlc5n1355_15_CYMUXFAST_2379 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_15_CYMUXG2,
      IB => U_DCT1D_rtlc5n1355_15_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1355_15_CYAND,
      O => U_DCT1D_rtlc5n1355_15_CYMUXFAST
    );
  U_DCT1D_rtlc5n1355_15_CYMUXG2_2380 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1355_15_CY0G,
      IB => U_DCT1D_rtlc5n1355_15_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1355_15_CYSELG,
      O => U_DCT1D_rtlc5n1355_15_CYMUXG2
    );
  U_DCT1D_rtlc5n1355_15_CY0G_2381 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s(13),
      O => U_DCT1D_rtlc5n1355_15_CY0G
    );
  U_DCT1D_rtlc5n1355_15_CYSELG_2382 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z7,
      O => U_DCT1D_rtlc5n1355_15_CYSELG
    );
  U_DCT1D_nx59700z5_rt_2383 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z5,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z5_rt
    );
  U_DCT1D_rtlc5n1355_17_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1355_17_XORF,
      O => U_DCT1D_rtlc5n1355(17)
    );
  U_DCT1D_rtlc5n1355_17_XORF_2384 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1355_17_CYINIT,
      I1 => U_DCT1D_nx59700z5_rt,
      O => U_DCT1D_rtlc5n1355_17_XORF
    );
  U_DCT1D_rtlc5n1355_17_CYINIT_2385 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_512_add_28_ix59700z63348_O,
      O => U_DCT1D_rtlc5n1355_17_CYINIT
    );
  U_DCT2D_nx115_bus_2_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_2_XORF,
      O => U_DCT2D_nx115_bus(2)
    );
  U_DCT2D_nx115_bus_2_XORF_2386 : X_XOR2
    port map (
      I0 => U_DCT2D_nx115_bus_2_CYINIT,
      I1 => U_DCT2D_nx65206z502,
      O => U_DCT2D_nx115_bus_2_XORF
    );
  U_DCT2D_nx115_bus_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_2_CY0F,
      IB => U_DCT2D_nx115_bus_2_CYINIT,
      SEL => U_DCT2D_nx115_bus_2_CYSELF,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z64052_O
    );
  U_DCT2D_nx115_bus_2_CYINIT_2387 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_2_BXINVNOT,
      O => U_DCT2D_nx115_bus_2_CYINIT
    );
  U_DCT2D_nx115_bus_2_CY0F_2388 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z503,
      O => U_DCT2D_nx115_bus_2_CY0F
    );
  U_DCT2D_nx115_bus_2_FAND : X_AND2
    port map (
      I0 => romo2datao6_s(0),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z503
    );
  U_DCT2D_nx115_bus_2_CYSELF_2389 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z502,
      O => U_DCT2D_nx115_bus_2_CYSELF
    );
  U_DCT2D_nx115_bus_2_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_18,
      O => U_DCT2D_nx115_bus_2_BXINVNOT
    );
  U_DCT2D_nx115_bus_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_2_XORG,
      O => U_DCT2D_nx115_bus(3)
    );
  U_DCT2D_nx115_bus_2_XORG_2390 : X_XOR2
    port map (
      I0 => U_DCT2D_ix946_modgen_add_293_ix65206z64052_O,
      I1 => U_DCT2D_nx65206z499,
      O => U_DCT2D_nx115_bus_2_XORG
    );
  U_DCT2D_nx115_bus_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_2_CYMUXG,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z64046_O
    );
  U_DCT2D_nx115_bus_2_CYMUXG_2391 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_2_CY0G,
      IB => U_DCT2D_ix946_modgen_add_293_ix65206z64052_O,
      SEL => U_DCT2D_nx115_bus_2_CYSELG,
      O => U_DCT2D_nx115_bus_2_CYMUXG
    );
  U_DCT2D_nx115_bus_2_CY0G_2392 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z500,
      O => U_DCT2D_nx115_bus_2_CY0G
    );
  U_DCT2D_nx115_bus_2_GAND : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483(7),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z500
    );
  U_DCT2D_nx115_bus_2_CYSELG_2393 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z499,
      O => U_DCT2D_nx115_bus_2_CYSELG
    );
  U_DCT2D_ix65206z31409 : X_LUT4
    generic map(
      INIT => X"74B8"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1483(9),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1498(9),
      ADR3 => U_DCT2D_rtlc5n1482(9),
      O => U_DCT2D_nx65206z493
    );
  U_DCT2D_nx115_bus_4_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_4_XORF,
      O => U_DCT2D_nx115_bus(4)
    );
  U_DCT2D_nx115_bus_4_XORF_2394 : X_XOR2
    port map (
      I0 => U_DCT2D_nx115_bus_4_CYINIT,
      I1 => U_DCT2D_nx65206z496,
      O => U_DCT2D_nx115_bus_4_XORF
    );
  U_DCT2D_nx115_bus_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_4_CY0F,
      IB => U_DCT2D_nx115_bus_4_CYINIT,
      SEL => U_DCT2D_nx115_bus_4_CYSELF,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z64040_O
    );
  U_DCT2D_nx115_bus_4_CYMUXF2_2395 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_4_CY0F,
      IB => U_DCT2D_nx115_bus_4_CY0F,
      SEL => U_DCT2D_nx115_bus_4_CYSELF,
      O => U_DCT2D_nx115_bus_4_CYMUXF2
    );
  U_DCT2D_nx115_bus_4_CYINIT_2396 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z64046_O,
      O => U_DCT2D_nx115_bus_4_CYINIT
    );
  U_DCT2D_nx115_bus_4_CY0F_2397 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z497,
      O => U_DCT2D_nx115_bus_4_CY0F
    );
  U_DCT2D_nx115_bus_4_FAND : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483(8),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z497
    );
  U_DCT2D_nx115_bus_4_CYSELF_2398 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z496,
      O => U_DCT2D_nx115_bus_4_CYSELF
    );
  U_DCT2D_nx115_bus_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_4_XORG,
      O => U_DCT2D_nx115_bus(5)
    );
  U_DCT2D_nx115_bus_4_XORG_2399 : X_XOR2
    port map (
      I0 => U_DCT2D_ix946_modgen_add_293_ix65206z64040_O,
      I1 => U_DCT2D_nx65206z493,
      O => U_DCT2D_nx115_bus_4_XORG
    );
  U_DCT2D_nx115_bus_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_4_CYMUXFAST,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z64034_O
    );
  U_DCT2D_nx115_bus_4_FASTCARRY_2400 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z64046_O,
      O => U_DCT2D_nx115_bus_4_FASTCARRY
    );
  U_DCT2D_nx115_bus_4_CYAND_2401 : X_AND2
    port map (
      I0 => U_DCT2D_nx115_bus_4_CYSELG,
      I1 => U_DCT2D_nx115_bus_4_CYSELF,
      O => U_DCT2D_nx115_bus_4_CYAND
    );
  U_DCT2D_nx115_bus_4_CYMUXFAST_2402 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_4_CYMUXG2,
      IB => U_DCT2D_nx115_bus_4_FASTCARRY,
      SEL => U_DCT2D_nx115_bus_4_CYAND,
      O => U_DCT2D_nx115_bus_4_CYMUXFAST
    );
  U_DCT2D_nx115_bus_4_CYMUXG2_2403 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_4_CY0G,
      IB => U_DCT2D_nx115_bus_4_CYMUXF2,
      SEL => U_DCT2D_nx115_bus_4_CYSELG,
      O => U_DCT2D_nx115_bus_4_CYMUXG2
    );
  U_DCT2D_nx115_bus_4_CY0G_2404 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z494,
      O => U_DCT2D_nx115_bus_4_CY0G
    );
  U_DCT2D_nx115_bus_4_GAND : X_AND2
    port map (
      I0 => U_DCT2D_state_reg(0),
      I1 => U_DCT2D_rtlc5n1483(9),
      O => U_DCT2D_nx65206z494
    );
  U_DCT2D_nx115_bus_4_CYSELG_2405 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z493,
      O => U_DCT2D_nx115_bus_4_CYSELG
    );
  U_DCT2D_nx115_bus_6_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_6_XORF,
      O => U_DCT2D_nx115_bus(6)
    );
  U_DCT2D_nx115_bus_6_XORF_2406 : X_XOR2
    port map (
      I0 => U_DCT2D_nx115_bus_6_CYINIT,
      I1 => U_DCT2D_nx65206z490,
      O => U_DCT2D_nx115_bus_6_XORF
    );
  U_DCT2D_nx115_bus_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_6_CY0F,
      IB => U_DCT2D_nx115_bus_6_CYINIT,
      SEL => U_DCT2D_nx115_bus_6_CYSELF,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z64028_O
    );
  U_DCT2D_nx115_bus_6_CYMUXF2_2407 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_6_CY0F,
      IB => U_DCT2D_nx115_bus_6_CY0F,
      SEL => U_DCT2D_nx115_bus_6_CYSELF,
      O => U_DCT2D_nx115_bus_6_CYMUXF2
    );
  U_DCT2D_nx115_bus_6_CYINIT_2408 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z64034_O,
      O => U_DCT2D_nx115_bus_6_CYINIT
    );
  U_DCT2D_nx115_bus_6_CY0F_2409 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z491,
      O => U_DCT2D_nx115_bus_6_CY0F
    );
  U_DCT2D_nx115_bus_6_FAND : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483(10),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z491
    );
  U_DCT2D_nx115_bus_6_CYSELF_2410 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z490,
      O => U_DCT2D_nx115_bus_6_CYSELF
    );
  U_DCT2D_nx115_bus_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_6_XORG,
      O => U_DCT2D_nx115_bus(7)
    );
  U_DCT2D_nx115_bus_6_XORG_2411 : X_XOR2
    port map (
      I0 => U_DCT2D_ix946_modgen_add_293_ix65206z64028_O,
      I1 => U_DCT2D_nx65206z487,
      O => U_DCT2D_nx115_bus_6_XORG
    );
  U_DCT2D_nx115_bus_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_6_CYMUXFAST,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z64022_O
    );
  U_DCT2D_nx115_bus_6_FASTCARRY_2412 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z64034_O,
      O => U_DCT2D_nx115_bus_6_FASTCARRY
    );
  U_DCT2D_nx115_bus_6_CYAND_2413 : X_AND2
    port map (
      I0 => U_DCT2D_nx115_bus_6_CYSELG,
      I1 => U_DCT2D_nx115_bus_6_CYSELF,
      O => U_DCT2D_nx115_bus_6_CYAND
    );
  U_DCT2D_nx115_bus_6_CYMUXFAST_2414 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_6_CYMUXG2,
      IB => U_DCT2D_nx115_bus_6_FASTCARRY,
      SEL => U_DCT2D_nx115_bus_6_CYAND,
      O => U_DCT2D_nx115_bus_6_CYMUXFAST
    );
  U_DCT2D_nx115_bus_6_CYMUXG2_2415 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_6_CY0G,
      IB => U_DCT2D_nx115_bus_6_CYMUXF2,
      SEL => U_DCT2D_nx115_bus_6_CYSELG,
      O => U_DCT2D_nx115_bus_6_CYMUXG2
    );
  U_DCT2D_nx115_bus_6_CY0G_2416 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z488,
      O => U_DCT2D_nx115_bus_6_CY0G
    );
  U_DCT2D_nx115_bus_6_GAND : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483(11),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z488
    );
  U_DCT2D_nx115_bus_6_CYSELG_2417 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z487,
      O => U_DCT2D_nx115_bus_6_CYSELG
    );
  U_DCT2D_ix65206z31385 : X_LUT4
    generic map(
      INIT => X"74B8"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1483(13),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1498(13),
      ADR3 => U_DCT2D_rtlc5n1482(13),
      O => U_DCT2D_nx65206z481
    );
  U_DCT2D_nx115_bus_8_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_8_XORF,
      O => U_DCT2D_nx115_bus(8)
    );
  U_DCT2D_nx115_bus_8_XORF_2418 : X_XOR2
    port map (
      I0 => U_DCT2D_nx115_bus_8_CYINIT,
      I1 => U_DCT2D_nx65206z484,
      O => U_DCT2D_nx115_bus_8_XORF
    );
  U_DCT2D_nx115_bus_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_8_CY0F,
      IB => U_DCT2D_nx115_bus_8_CYINIT,
      SEL => U_DCT2D_nx115_bus_8_CYSELF,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z64016_O
    );
  U_DCT2D_nx115_bus_8_CYMUXF2_2419 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_8_CY0F,
      IB => U_DCT2D_nx115_bus_8_CY0F,
      SEL => U_DCT2D_nx115_bus_8_CYSELF,
      O => U_DCT2D_nx115_bus_8_CYMUXF2
    );
  U_DCT2D_nx115_bus_8_CYINIT_2420 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z64022_O,
      O => U_DCT2D_nx115_bus_8_CYINIT
    );
  U_DCT2D_nx115_bus_8_CY0F_2421 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z485,
      O => U_DCT2D_nx115_bus_8_CY0F
    );
  U_DCT2D_nx115_bus_8_FAND : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483(12),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z485
    );
  U_DCT2D_nx115_bus_8_CYSELF_2422 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z484,
      O => U_DCT2D_nx115_bus_8_CYSELF
    );
  U_DCT2D_nx115_bus_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_8_XORG,
      O => U_DCT2D_nx115_bus(9)
    );
  U_DCT2D_nx115_bus_8_XORG_2423 : X_XOR2
    port map (
      I0 => U_DCT2D_ix946_modgen_add_293_ix65206z64016_O,
      I1 => U_DCT2D_nx65206z481,
      O => U_DCT2D_nx115_bus_8_XORG
    );
  U_DCT2D_nx115_bus_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_8_CYMUXFAST,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z64010_O
    );
  U_DCT2D_nx115_bus_8_FASTCARRY_2424 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z64022_O,
      O => U_DCT2D_nx115_bus_8_FASTCARRY
    );
  U_DCT2D_nx115_bus_8_CYAND_2425 : X_AND2
    port map (
      I0 => U_DCT2D_nx115_bus_8_CYSELG,
      I1 => U_DCT2D_nx115_bus_8_CYSELF,
      O => U_DCT2D_nx115_bus_8_CYAND
    );
  U_DCT2D_nx115_bus_8_CYMUXFAST_2426 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_8_CYMUXG2,
      IB => U_DCT2D_nx115_bus_8_FASTCARRY,
      SEL => U_DCT2D_nx115_bus_8_CYAND,
      O => U_DCT2D_nx115_bus_8_CYMUXFAST
    );
  U_DCT2D_nx115_bus_8_CYMUXG2_2427 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_8_CY0G,
      IB => U_DCT2D_nx115_bus_8_CYMUXF2,
      SEL => U_DCT2D_nx115_bus_8_CYSELG,
      O => U_DCT2D_nx115_bus_8_CYMUXG2
    );
  U_DCT2D_nx115_bus_8_CY0G_2428 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z482,
      O => U_DCT2D_nx115_bus_8_CY0G
    );
  U_DCT2D_nx115_bus_8_GAND : X_AND2
    port map (
      I0 => U_DCT2D_state_reg(0),
      I1 => U_DCT2D_rtlc5n1483(13),
      O => U_DCT2D_nx65206z482
    );
  U_DCT2D_nx115_bus_8_CYSELG_2429 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z481,
      O => U_DCT2D_nx115_bus_8_CYSELG
    );
  U_DCT2D_nx115_bus_10_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_10_XORF,
      O => U_DCT2D_nx115_bus(10)
    );
  U_DCT2D_nx115_bus_10_XORF_2430 : X_XOR2
    port map (
      I0 => U_DCT2D_nx115_bus_10_CYINIT,
      I1 => U_DCT2D_nx65206z478,
      O => U_DCT2D_nx115_bus_10_XORF
    );
  U_DCT2D_nx115_bus_10_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_10_CY0F,
      IB => U_DCT2D_nx115_bus_10_CYINIT,
      SEL => U_DCT2D_nx115_bus_10_CYSELF,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z64004_O
    );
  U_DCT2D_nx115_bus_10_CYMUXF2_2431 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_10_CY0F,
      IB => U_DCT2D_nx115_bus_10_CY0F,
      SEL => U_DCT2D_nx115_bus_10_CYSELF,
      O => U_DCT2D_nx115_bus_10_CYMUXF2
    );
  U_DCT2D_nx115_bus_10_CYINIT_2432 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z64010_O,
      O => U_DCT2D_nx115_bus_10_CYINIT
    );
  U_DCT2D_nx115_bus_10_CY0F_2433 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z479,
      O => U_DCT2D_nx115_bus_10_CY0F
    );
  U_DCT2D_nx115_bus_10_FAND : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483(14),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z479
    );
  U_DCT2D_nx115_bus_10_CYSELF_2434 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z478,
      O => U_DCT2D_nx115_bus_10_CYSELF
    );
  U_DCT2D_nx115_bus_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_10_XORG,
      O => U_DCT2D_nx115_bus(11)
    );
  U_DCT2D_nx115_bus_10_XORG_2435 : X_XOR2
    port map (
      I0 => U_DCT2D_ix946_modgen_add_293_ix65206z64004_O,
      I1 => U_DCT2D_nx65206z475,
      O => U_DCT2D_nx115_bus_10_XORG
    );
  U_DCT2D_nx115_bus_10_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_10_CYMUXFAST,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z63998_O
    );
  U_DCT2D_nx115_bus_10_FASTCARRY_2436 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z64010_O,
      O => U_DCT2D_nx115_bus_10_FASTCARRY
    );
  U_DCT2D_nx115_bus_10_CYAND_2437 : X_AND2
    port map (
      I0 => U_DCT2D_nx115_bus_10_CYSELG,
      I1 => U_DCT2D_nx115_bus_10_CYSELF,
      O => U_DCT2D_nx115_bus_10_CYAND
    );
  U_DCT2D_nx115_bus_10_CYMUXFAST_2438 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_10_CYMUXG2,
      IB => U_DCT2D_nx115_bus_10_FASTCARRY,
      SEL => U_DCT2D_nx115_bus_10_CYAND,
      O => U_DCT2D_nx115_bus_10_CYMUXFAST
    );
  U_DCT2D_nx115_bus_10_CYMUXG2_2439 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_10_CY0G,
      IB => U_DCT2D_nx115_bus_10_CYMUXF2,
      SEL => U_DCT2D_nx115_bus_10_CYSELG,
      O => U_DCT2D_nx115_bus_10_CYMUXG2
    );
  U_DCT2D_nx115_bus_10_CY0G_2440 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z476,
      O => U_DCT2D_nx115_bus_10_CY0G
    );
  U_DCT2D_nx115_bus_10_GAND : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483(15),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z476
    );
  U_DCT2D_nx115_bus_10_CYSELG_2441 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z475,
      O => U_DCT2D_nx115_bus_10_CYSELG
    );
  U_DCT2D_ix65206z31361 : X_LUT4
    generic map(
      INIT => X"74B8"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1483(17),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1498(17),
      ADR3 => U_DCT2D_rtlc5n1482(17),
      O => U_DCT2D_nx65206z469
    );
  U_DCT2D_nx115_bus_12_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_12_XORF,
      O => U_DCT2D_nx115_bus(12)
    );
  U_DCT2D_nx115_bus_12_XORF_2442 : X_XOR2
    port map (
      I0 => U_DCT2D_nx115_bus_12_CYINIT,
      I1 => U_DCT2D_nx65206z472,
      O => U_DCT2D_nx115_bus_12_XORF
    );
  U_DCT2D_nx115_bus_12_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_12_CY0F,
      IB => U_DCT2D_nx115_bus_12_CYINIT,
      SEL => U_DCT2D_nx115_bus_12_CYSELF,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z63992_O
    );
  U_DCT2D_nx115_bus_12_CYMUXF2_2443 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_12_CY0F,
      IB => U_DCT2D_nx115_bus_12_CY0F,
      SEL => U_DCT2D_nx115_bus_12_CYSELF,
      O => U_DCT2D_nx115_bus_12_CYMUXF2
    );
  U_DCT2D_nx115_bus_12_CYINIT_2444 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z63998_O,
      O => U_DCT2D_nx115_bus_12_CYINIT
    );
  U_DCT2D_nx115_bus_12_CY0F_2445 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z473,
      O => U_DCT2D_nx115_bus_12_CY0F
    );
  U_DCT2D_nx115_bus_12_FAND : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483(16),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z473
    );
  U_DCT2D_nx115_bus_12_CYSELF_2446 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z472,
      O => U_DCT2D_nx115_bus_12_CYSELF
    );
  U_DCT2D_nx115_bus_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_12_XORG,
      O => U_DCT2D_nx115_bus(13)
    );
  U_DCT2D_nx115_bus_12_XORG_2447 : X_XOR2
    port map (
      I0 => U_DCT2D_ix946_modgen_add_293_ix65206z63992_O,
      I1 => U_DCT2D_nx65206z469,
      O => U_DCT2D_nx115_bus_12_XORG
    );
  U_DCT2D_nx115_bus_12_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_12_CYMUXFAST,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z63986_O
    );
  U_DCT2D_nx115_bus_12_FASTCARRY_2448 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z63998_O,
      O => U_DCT2D_nx115_bus_12_FASTCARRY
    );
  U_DCT2D_nx115_bus_12_CYAND_2449 : X_AND2
    port map (
      I0 => U_DCT2D_nx115_bus_12_CYSELG,
      I1 => U_DCT2D_nx115_bus_12_CYSELF,
      O => U_DCT2D_nx115_bus_12_CYAND
    );
  U_DCT2D_nx115_bus_12_CYMUXFAST_2450 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_12_CYMUXG2,
      IB => U_DCT2D_nx115_bus_12_FASTCARRY,
      SEL => U_DCT2D_nx115_bus_12_CYAND,
      O => U_DCT2D_nx115_bus_12_CYMUXFAST
    );
  U_DCT2D_nx115_bus_12_CYMUXG2_2451 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_12_CY0G,
      IB => U_DCT2D_nx115_bus_12_CYMUXF2,
      SEL => U_DCT2D_nx115_bus_12_CYSELG,
      O => U_DCT2D_nx115_bus_12_CYMUXG2
    );
  U_DCT2D_nx115_bus_12_CY0G_2452 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z470,
      O => U_DCT2D_nx115_bus_12_CY0G
    );
  U_DCT2D_nx115_bus_12_GAND : X_AND2
    port map (
      I0 => U_DCT2D_state_reg(0),
      I1 => U_DCT2D_rtlc5n1483(17),
      O => U_DCT2D_nx65206z470
    );
  U_DCT2D_nx115_bus_12_CYSELG_2453 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z469,
      O => U_DCT2D_nx115_bus_12_CYSELG
    );
  U_DCT2D_nx115_bus_14_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_14_XORF,
      O => U_DCT2D_nx115_bus(14)
    );
  U_DCT2D_nx115_bus_14_XORF_2454 : X_XOR2
    port map (
      I0 => U_DCT2D_nx115_bus_14_CYINIT,
      I1 => U_DCT2D_nx65206z466,
      O => U_DCT2D_nx115_bus_14_XORF
    );
  U_DCT2D_nx115_bus_14_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_14_CY0F,
      IB => U_DCT2D_nx115_bus_14_CYINIT,
      SEL => U_DCT2D_nx115_bus_14_CYSELF,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z63980_O
    );
  U_DCT2D_nx115_bus_14_CYMUXF2_2455 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_14_CY0F,
      IB => U_DCT2D_nx115_bus_14_CY0F,
      SEL => U_DCT2D_nx115_bus_14_CYSELF,
      O => U_DCT2D_nx115_bus_14_CYMUXF2
    );
  U_DCT2D_nx115_bus_14_CYINIT_2456 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z63986_O,
      O => U_DCT2D_nx115_bus_14_CYINIT
    );
  U_DCT2D_nx115_bus_14_CY0F_2457 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z467,
      O => U_DCT2D_nx115_bus_14_CY0F
    );
  U_DCT2D_nx115_bus_14_FAND : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483(18),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z467
    );
  U_DCT2D_nx115_bus_14_CYSELF_2458 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z466,
      O => U_DCT2D_nx115_bus_14_CYSELF
    );
  U_DCT2D_nx115_bus_14_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_14_XORG,
      O => U_DCT2D_nx115_bus(15)
    );
  U_DCT2D_nx115_bus_14_XORG_2459 : X_XOR2
    port map (
      I0 => U_DCT2D_ix946_modgen_add_293_ix65206z63980_O,
      I1 => U_DCT2D_nx65206z463,
      O => U_DCT2D_nx115_bus_14_XORG
    );
  U_DCT2D_nx115_bus_14_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_14_CYMUXFAST,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z63975_O
    );
  U_DCT2D_nx115_bus_14_FASTCARRY_2460 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z63986_O,
      O => U_DCT2D_nx115_bus_14_FASTCARRY
    );
  U_DCT2D_nx115_bus_14_CYAND_2461 : X_AND2
    port map (
      I0 => U_DCT2D_nx115_bus_14_CYSELG,
      I1 => U_DCT2D_nx115_bus_14_CYSELF,
      O => U_DCT2D_nx115_bus_14_CYAND
    );
  U_DCT2D_nx115_bus_14_CYMUXFAST_2462 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_14_CYMUXG2,
      IB => U_DCT2D_nx115_bus_14_FASTCARRY,
      SEL => U_DCT2D_nx115_bus_14_CYAND,
      O => U_DCT2D_nx115_bus_14_CYMUXFAST
    );
  U_DCT2D_nx115_bus_14_CYMUXG2_2463 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_14_CY0G,
      IB => U_DCT2D_nx115_bus_14_CYMUXF2,
      SEL => U_DCT2D_nx115_bus_14_CYSELG,
      O => U_DCT2D_nx115_bus_14_CYMUXG2
    );
  U_DCT2D_nx115_bus_14_CY0G_2464 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z464,
      O => U_DCT2D_nx115_bus_14_CY0G
    );
  U_DCT2D_nx115_bus_14_GAND : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483(19),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z464
    );
  U_DCT2D_nx115_bus_14_CYSELG_2465 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z463,
      O => U_DCT2D_nx115_bus_14_CYSELG
    );
  U_DCT2D_ix65206z31341 : X_LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1483(21),
      ADR2 => U_DCT2D_rtlc5n1482(19),
      ADR3 => U_DCT2D_rtlc5n1498(21),
      O => U_DCT2D_nx65206z457
    );
  U_DCT2D_nx115_bus_16_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_16_XORF,
      O => U_DCT2D_nx115_bus(16)
    );
  U_DCT2D_nx115_bus_16_XORF_2466 : X_XOR2
    port map (
      I0 => U_DCT2D_nx115_bus_16_CYINIT,
      I1 => U_DCT2D_nx65206z460,
      O => U_DCT2D_nx115_bus_16_XORF
    );
  U_DCT2D_nx115_bus_16_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_16_CY0F,
      IB => U_DCT2D_nx115_bus_16_CYINIT,
      SEL => U_DCT2D_nx115_bus_16_CYSELF,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z63970_O
    );
  U_DCT2D_nx115_bus_16_CYMUXF2_2467 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_16_CY0F,
      IB => U_DCT2D_nx115_bus_16_CY0F,
      SEL => U_DCT2D_nx115_bus_16_CYSELF,
      O => U_DCT2D_nx115_bus_16_CYMUXF2
    );
  U_DCT2D_nx115_bus_16_CYINIT_2468 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z63975_O,
      O => U_DCT2D_nx115_bus_16_CYINIT
    );
  U_DCT2D_nx115_bus_16_CY0F_2469 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z461,
      O => U_DCT2D_nx115_bus_16_CY0F
    );
  U_DCT2D_nx115_bus_16_FAND : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483(20),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z461
    );
  U_DCT2D_nx115_bus_16_CYSELF_2470 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z460,
      O => U_DCT2D_nx115_bus_16_CYSELF
    );
  U_DCT2D_nx115_bus_16_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_16_XORG,
      O => U_DCT2D_nx115_bus(17)
    );
  U_DCT2D_nx115_bus_16_XORG_2471 : X_XOR2
    port map (
      I0 => U_DCT2D_ix946_modgen_add_293_ix65206z63970_O,
      I1 => U_DCT2D_nx65206z457,
      O => U_DCT2D_nx115_bus_16_XORG
    );
  U_DCT2D_nx115_bus_16_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_16_CYMUXFAST,
      O => U_DCT2D_ix946_modgen_add_293_ix65206z63966_O
    );
  U_DCT2D_nx115_bus_16_FASTCARRY_2472 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z63975_O,
      O => U_DCT2D_nx115_bus_16_FASTCARRY
    );
  U_DCT2D_nx115_bus_16_CYAND_2473 : X_AND2
    port map (
      I0 => U_DCT2D_nx115_bus_16_CYSELG,
      I1 => U_DCT2D_nx115_bus_16_CYSELF,
      O => U_DCT2D_nx115_bus_16_CYAND
    );
  U_DCT2D_nx115_bus_16_CYMUXFAST_2474 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_16_CYMUXG2,
      IB => U_DCT2D_nx115_bus_16_FASTCARRY,
      SEL => U_DCT2D_nx115_bus_16_CYAND,
      O => U_DCT2D_nx115_bus_16_CYMUXFAST
    );
  U_DCT2D_nx115_bus_16_CYMUXG2_2475 : X_MUX2
    port map (
      IA => U_DCT2D_nx115_bus_16_CY0G,
      IB => U_DCT2D_nx115_bus_16_CYMUXF2,
      SEL => U_DCT2D_nx115_bus_16_CYSELG,
      O => U_DCT2D_nx115_bus_16_CYMUXG2
    );
  U_DCT2D_nx115_bus_16_CY0G_2476 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z458,
      O => U_DCT2D_nx115_bus_16_CY0G
    );
  U_DCT2D_nx115_bus_16_GAND : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1483(21),
      I1 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z458
    );
  U_DCT2D_nx115_bus_16_CYSELG_2477 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z457,
      O => U_DCT2D_nx115_bus_16_CYSELG
    );
  U_DCT1D_nx2262z1_rt_2478 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => U_DCT1D_nx2262z1,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx2262z1_rt
    );
  U_DCT2D_nx65206z252_rt_2479 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z252,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z252_rt
    );
  U_DCT2D_nx115_bus_18_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx115_bus_18_XORF,
      O => U_DCT2D_nx115_bus(18)
    );
  U_DCT2D_nx115_bus_18_XORF_2480 : X_XOR2
    port map (
      I0 => U_DCT2D_nx115_bus_18_CYINIT,
      I1 => U_DCT2D_nx65206z252_rt,
      O => U_DCT2D_nx115_bus_18_XORF
    );
  U_DCT2D_nx115_bus_18_CYINIT_2481 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix946_modgen_add_293_ix65206z63966_O,
      O => U_DCT2D_nx115_bus_18_CYINIT
    );
  U_DCT1D_rtlc5n1346_5_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_5_XORF,
      O => U_DCT1D_rtlc5n1346(5)
    );
  U_DCT1D_rtlc5n1346_5_XORF_2482 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1346_5_CYINIT,
      I1 => U_DCT1D_nx59700z296,
      O => U_DCT1D_rtlc5n1346_5_XORF
    );
  U_DCT1D_rtlc5n1346_5_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_5_CY0F,
      IB => U_DCT1D_rtlc5n1346_5_CYINIT,
      SEL => U_DCT1D_rtlc5n1346_5_CYSELF,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63745_O
    );
  U_DCT1D_rtlc5n1346_5_CYINIT_2483 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_5_BXINVNOT,
      O => U_DCT1D_rtlc5n1346_5_CYINIT
    );
  U_DCT1D_rtlc5n1346_5_CY0F_2484 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(1),
      O => U_DCT1D_rtlc5n1346_5_CY0F
    );
  U_DCT1D_rtlc5n1346_5_CYSELF_2485 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z296,
      O => U_DCT1D_rtlc5n1346_5_CYSELF
    );
  U_DCT1D_rtlc5n1346_5_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1,
      O => U_DCT1D_rtlc5n1346_5_BXINVNOT
    );
  U_DCT1D_rtlc5n1346_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_5_XORG,
      O => U_DCT1D_rtlc5n1346(6)
    );
  U_DCT1D_rtlc5n1346_5_XORG_2486 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_498_add_23_ix59700z63745_O,
      I1 => U_DCT1D_nx59700z293,
      O => U_DCT1D_rtlc5n1346_5_XORG
    );
  U_DCT1D_rtlc5n1346_5_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_5_CYMUXG,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63742_O
    );
  U_DCT1D_rtlc5n1346_5_CYMUXG_2487 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_5_CY0G,
      IB => U_DCT1D_rtlc_498_add_23_ix59700z63745_O,
      SEL => U_DCT1D_rtlc5n1346_5_CYSELG,
      O => U_DCT1D_rtlc5n1346_5_CYMUXG
    );
  U_DCT1D_rtlc5n1346_5_CY0G_2488 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(2),
      O => U_DCT1D_rtlc5n1346_5_CY0G
    );
  U_DCT1D_rtlc5n1346_5_CYSELG_2489 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z293,
      O => U_DCT1D_rtlc5n1346_5_CYSELG
    );
  U_DCT1D_rtlc5n1346_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_7_XORF,
      O => U_DCT1D_rtlc5n1346(7)
    );
  U_DCT1D_rtlc5n1346_7_XORF_2490 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1346_7_CYINIT,
      I1 => U_DCT1D_nx59700z290,
      O => U_DCT1D_rtlc5n1346_7_XORF
    );
  U_DCT1D_rtlc5n1346_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_7_CY0F,
      IB => U_DCT1D_rtlc5n1346_7_CYINIT,
      SEL => U_DCT1D_rtlc5n1346_7_CYSELF,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63738_O
    );
  U_DCT1D_rtlc5n1346_7_CYMUXF2_2491 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_7_CY0F,
      IB => U_DCT1D_rtlc5n1346_7_CY0F,
      SEL => U_DCT1D_rtlc5n1346_7_CYSELF,
      O => U_DCT1D_rtlc5n1346_7_CYMUXF2
    );
  U_DCT1D_rtlc5n1346_7_CYINIT_2492 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63742_O,
      O => U_DCT1D_rtlc5n1346_7_CYINIT
    );
  U_DCT1D_rtlc5n1346_7_CY0F_2493 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(3),
      O => U_DCT1D_rtlc5n1346_7_CY0F
    );
  U_DCT1D_rtlc5n1346_7_CYSELF_2494 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z290,
      O => U_DCT1D_rtlc5n1346_7_CYSELF
    );
  U_DCT1D_rtlc5n1346_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_7_XORG,
      O => U_DCT1D_rtlc5n1346(8)
    );
  U_DCT1D_rtlc5n1346_7_XORG_2495 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_498_add_23_ix59700z63738_O,
      I1 => U_DCT1D_nx59700z287,
      O => U_DCT1D_rtlc5n1346_7_XORG
    );
  U_DCT1D_rtlc5n1346_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_7_CYMUXFAST,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63735_O
    );
  U_DCT1D_rtlc5n1346_7_FASTCARRY_2496 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63742_O,
      O => U_DCT1D_rtlc5n1346_7_FASTCARRY
    );
  U_DCT1D_rtlc5n1346_7_CYAND_2497 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1346_7_CYSELG,
      I1 => U_DCT1D_rtlc5n1346_7_CYSELF,
      O => U_DCT1D_rtlc5n1346_7_CYAND
    );
  U_DCT1D_rtlc5n1346_7_CYMUXFAST_2498 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_7_CYMUXG2,
      IB => U_DCT1D_rtlc5n1346_7_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1346_7_CYAND,
      O => U_DCT1D_rtlc5n1346_7_CYMUXFAST
    );
  U_DCT1D_rtlc5n1346_7_CYMUXG2_2499 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_7_CY0G,
      IB => U_DCT1D_rtlc5n1346_7_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1346_7_CYSELG,
      O => U_DCT1D_rtlc5n1346_7_CYMUXG2
    );
  U_DCT1D_rtlc5n1346_7_CY0G_2500 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(4),
      O => U_DCT1D_rtlc5n1346_7_CY0G
    );
  U_DCT1D_rtlc5n1346_7_CYSELG_2501 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z287,
      O => U_DCT1D_rtlc5n1346_7_CYSELG
    );
  U_DCT1D_rtlc5n1346_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_9_XORF,
      O => U_DCT1D_rtlc5n1346(9)
    );
  U_DCT1D_rtlc5n1346_9_XORF_2502 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1346_9_CYINIT,
      I1 => U_DCT1D_nx59700z284,
      O => U_DCT1D_rtlc5n1346_9_XORF
    );
  U_DCT1D_rtlc5n1346_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_9_CY0F,
      IB => U_DCT1D_rtlc5n1346_9_CYINIT,
      SEL => U_DCT1D_rtlc5n1346_9_CYSELF,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63731_O
    );
  U_DCT1D_rtlc5n1346_9_CYMUXF2_2503 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_9_CY0F,
      IB => U_DCT1D_rtlc5n1346_9_CY0F,
      SEL => U_DCT1D_rtlc5n1346_9_CYSELF,
      O => U_DCT1D_rtlc5n1346_9_CYMUXF2
    );
  U_DCT1D_rtlc5n1346_9_CYINIT_2504 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63735_O,
      O => U_DCT1D_rtlc5n1346_9_CYINIT
    );
  U_DCT1D_rtlc5n1346_9_CY0F_2505 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(5),
      O => U_DCT1D_rtlc5n1346_9_CY0F
    );
  U_DCT1D_rtlc5n1346_9_CYSELF_2506 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z284,
      O => U_DCT1D_rtlc5n1346_9_CYSELF
    );
  U_DCT1D_rtlc5n1346_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_9_XORG,
      O => U_DCT1D_rtlc5n1346(10)
    );
  U_DCT1D_rtlc5n1346_9_XORG_2507 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_498_add_23_ix59700z63731_O,
      I1 => U_DCT1D_nx59700z281,
      O => U_DCT1D_rtlc5n1346_9_XORG
    );
  U_DCT1D_rtlc5n1346_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_9_CYMUXFAST,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63728_O
    );
  U_DCT1D_rtlc5n1346_9_FASTCARRY_2508 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63735_O,
      O => U_DCT1D_rtlc5n1346_9_FASTCARRY
    );
  U_DCT1D_rtlc5n1346_9_CYAND_2509 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1346_9_CYSELG,
      I1 => U_DCT1D_rtlc5n1346_9_CYSELF,
      O => U_DCT1D_rtlc5n1346_9_CYAND
    );
  U_DCT1D_rtlc5n1346_9_CYMUXFAST_2510 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_9_CYMUXG2,
      IB => U_DCT1D_rtlc5n1346_9_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1346_9_CYAND,
      O => U_DCT1D_rtlc5n1346_9_CYMUXFAST
    );
  U_DCT1D_rtlc5n1346_9_CYMUXG2_2511 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_9_CY0G,
      IB => U_DCT1D_rtlc5n1346_9_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1346_9_CYSELG,
      O => U_DCT1D_rtlc5n1346_9_CYMUXG2
    );
  U_DCT1D_rtlc5n1346_9_CY0G_2512 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(6),
      O => U_DCT1D_rtlc5n1346_9_CY0G
    );
  U_DCT1D_rtlc5n1346_9_CYSELG_2513 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z281,
      O => U_DCT1D_rtlc5n1346_9_CYSELG
    );
  U_DCT1D_rtlc5n1346_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_11_XORF,
      O => U_DCT1D_rtlc5n1346(11)
    );
  U_DCT1D_rtlc5n1346_11_XORF_2514 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1346_11_CYINIT,
      I1 => U_DCT1D_nx59700z278,
      O => U_DCT1D_rtlc5n1346_11_XORF
    );
  U_DCT1D_rtlc5n1346_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_11_CY0F,
      IB => U_DCT1D_rtlc5n1346_11_CYINIT,
      SEL => U_DCT1D_rtlc5n1346_11_CYSELF,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63724_O
    );
  U_DCT1D_rtlc5n1346_11_CYMUXF2_2515 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_11_CY0F,
      IB => U_DCT1D_rtlc5n1346_11_CY0F,
      SEL => U_DCT1D_rtlc5n1346_11_CYSELF,
      O => U_DCT1D_rtlc5n1346_11_CYMUXF2
    );
  U_DCT1D_rtlc5n1346_11_CYINIT_2516 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63728_O,
      O => U_DCT1D_rtlc5n1346_11_CYINIT
    );
  U_DCT1D_rtlc5n1346_11_CY0F_2517 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(7),
      O => U_DCT1D_rtlc5n1346_11_CY0F
    );
  U_DCT1D_rtlc5n1346_11_CYSELF_2518 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z278,
      O => U_DCT1D_rtlc5n1346_11_CYSELF
    );
  U_DCT1D_rtlc5n1346_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_11_XORG,
      O => U_DCT1D_rtlc5n1346(12)
    );
  U_DCT1D_rtlc5n1346_11_XORG_2519 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_498_add_23_ix59700z63724_O,
      I1 => U_DCT1D_nx59700z275,
      O => U_DCT1D_rtlc5n1346_11_XORG
    );
  U_DCT1D_rtlc5n1346_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_11_CYMUXFAST,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63721_O
    );
  U_DCT1D_rtlc5n1346_11_FASTCARRY_2520 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63728_O,
      O => U_DCT1D_rtlc5n1346_11_FASTCARRY
    );
  U_DCT1D_rtlc5n1346_11_CYAND_2521 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1346_11_CYSELG,
      I1 => U_DCT1D_rtlc5n1346_11_CYSELF,
      O => U_DCT1D_rtlc5n1346_11_CYAND
    );
  U_DCT1D_rtlc5n1346_11_CYMUXFAST_2522 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_11_CYMUXG2,
      IB => U_DCT1D_rtlc5n1346_11_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1346_11_CYAND,
      O => U_DCT1D_rtlc5n1346_11_CYMUXFAST
    );
  U_DCT1D_rtlc5n1346_11_CYMUXG2_2523 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_11_CY0G,
      IB => U_DCT1D_rtlc5n1346_11_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1346_11_CYSELG,
      O => U_DCT1D_rtlc5n1346_11_CYMUXG2
    );
  U_DCT1D_rtlc5n1346_11_CY0G_2524 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(8),
      O => U_DCT1D_rtlc5n1346_11_CY0G
    );
  U_DCT1D_rtlc5n1346_11_CYSELG_2525 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z275,
      O => U_DCT1D_rtlc5n1346_11_CYSELG
    );
  U_DCT1D_rtlc5n1346_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_13_XORF,
      O => U_DCT1D_rtlc5n1346(13)
    );
  U_DCT1D_rtlc5n1346_13_XORF_2526 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1346_13_CYINIT,
      I1 => U_DCT1D_nx59700z272,
      O => U_DCT1D_rtlc5n1346_13_XORF
    );
  U_DCT1D_rtlc5n1346_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_13_CY0F,
      IB => U_DCT1D_rtlc5n1346_13_CYINIT,
      SEL => U_DCT1D_rtlc5n1346_13_CYSELF,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63717_O
    );
  U_DCT1D_rtlc5n1346_13_CYMUXF2_2527 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_13_CY0F,
      IB => U_DCT1D_rtlc5n1346_13_CY0F,
      SEL => U_DCT1D_rtlc5n1346_13_CYSELF,
      O => U_DCT1D_rtlc5n1346_13_CYMUXF2
    );
  U_DCT1D_rtlc5n1346_13_CYINIT_2528 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63721_O,
      O => U_DCT1D_rtlc5n1346_13_CYINIT
    );
  U_DCT1D_rtlc5n1346_13_CY0F_2529 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(9),
      O => U_DCT1D_rtlc5n1346_13_CY0F
    );
  U_DCT1D_rtlc5n1346_13_CYSELF_2530 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z272,
      O => U_DCT1D_rtlc5n1346_13_CYSELF
    );
  U_DCT1D_rtlc5n1346_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_13_XORG,
      O => U_DCT1D_rtlc5n1346(14)
    );
  U_DCT1D_rtlc5n1346_13_XORG_2531 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_498_add_23_ix59700z63717_O,
      I1 => U_DCT1D_nx59700z269,
      O => U_DCT1D_rtlc5n1346_13_XORG
    );
  U_DCT1D_rtlc5n1346_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_13_CYMUXFAST,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63714_O
    );
  U_DCT1D_rtlc5n1346_13_FASTCARRY_2532 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63721_O,
      O => U_DCT1D_rtlc5n1346_13_FASTCARRY
    );
  U_DCT1D_rtlc5n1346_13_CYAND_2533 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1346_13_CYSELG,
      I1 => U_DCT1D_rtlc5n1346_13_CYSELF,
      O => U_DCT1D_rtlc5n1346_13_CYAND
    );
  U_DCT1D_rtlc5n1346_13_CYMUXFAST_2534 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_13_CYMUXG2,
      IB => U_DCT1D_rtlc5n1346_13_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1346_13_CYAND,
      O => U_DCT1D_rtlc5n1346_13_CYMUXFAST
    );
  U_DCT1D_rtlc5n1346_13_CYMUXG2_2535 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_13_CY0G,
      IB => U_DCT1D_rtlc5n1346_13_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1346_13_CYSELG,
      O => U_DCT1D_rtlc5n1346_13_CYMUXG2
    );
  U_DCT1D_rtlc5n1346_13_CY0G_2536 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(10),
      O => U_DCT1D_rtlc5n1346_13_CY0G
    );
  U_DCT1D_rtlc5n1346_13_CYSELG_2537 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z269,
      O => U_DCT1D_rtlc5n1346_13_CYSELG
    );
  U_DCT1D_rtlc5n1346_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_15_XORF,
      O => U_DCT1D_rtlc5n1346(15)
    );
  U_DCT1D_rtlc5n1346_15_XORF_2538 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1346_15_CYINIT,
      I1 => U_DCT1D_nx59700z266,
      O => U_DCT1D_rtlc5n1346_15_XORF
    );
  U_DCT1D_rtlc5n1346_15_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_15_CY0F,
      IB => U_DCT1D_rtlc5n1346_15_CYINIT,
      SEL => U_DCT1D_rtlc5n1346_15_CYSELF,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63710_O
    );
  U_DCT1D_rtlc5n1346_15_CYMUXF2_2539 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_15_CY0F,
      IB => U_DCT1D_rtlc5n1346_15_CY0F,
      SEL => U_DCT1D_rtlc5n1346_15_CYSELF,
      O => U_DCT1D_rtlc5n1346_15_CYMUXF2
    );
  U_DCT1D_rtlc5n1346_15_CYINIT_2540 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63714_O,
      O => U_DCT1D_rtlc5n1346_15_CYINIT
    );
  U_DCT1D_rtlc5n1346_15_CY0F_2541 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(11),
      O => U_DCT1D_rtlc5n1346_15_CY0F
    );
  U_DCT1D_rtlc5n1346_15_CYSELF_2542 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z266,
      O => U_DCT1D_rtlc5n1346_15_CYSELF
    );
  U_DCT1D_rtlc5n1346_15_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_15_XORG,
      O => U_DCT1D_rtlc5n1346(16)
    );
  U_DCT1D_rtlc5n1346_15_XORG_2543 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_498_add_23_ix59700z63710_O,
      I1 => U_DCT1D_nx59700z263,
      O => U_DCT1D_rtlc5n1346_15_XORG
    );
  U_DCT1D_rtlc5n1346_15_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_15_CYMUXFAST,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63707_O
    );
  U_DCT1D_rtlc5n1346_15_FASTCARRY_2544 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63714_O,
      O => U_DCT1D_rtlc5n1346_15_FASTCARRY
    );
  U_DCT1D_rtlc5n1346_15_CYAND_2545 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1346_15_CYSELG,
      I1 => U_DCT1D_rtlc5n1346_15_CYSELF,
      O => U_DCT1D_rtlc5n1346_15_CYAND
    );
  U_DCT1D_rtlc5n1346_15_CYMUXFAST_2546 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_15_CYMUXG2,
      IB => U_DCT1D_rtlc5n1346_15_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1346_15_CYAND,
      O => U_DCT1D_rtlc5n1346_15_CYMUXFAST
    );
  U_DCT1D_rtlc5n1346_15_CYMUXG2_2547 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_15_CY0G,
      IB => U_DCT1D_rtlc5n1346_15_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1346_15_CYSELG,
      O => U_DCT1D_rtlc5n1346_15_CYMUXG2
    );
  U_DCT1D_rtlc5n1346_15_CY0G_2548 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(12),
      O => U_DCT1D_rtlc5n1346_15_CY0G
    );
  U_DCT1D_rtlc5n1346_15_CYSELG_2549 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z263,
      O => U_DCT1D_rtlc5n1346_15_CYSELG
    );
  U_DCT1D_rtlc5n1346_17_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_17_XORF,
      O => U_DCT1D_rtlc5n1346(17)
    );
  U_DCT1D_rtlc5n1346_17_XORF_2550 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1346_17_CYINIT,
      I1 => U_DCT1D_nx59700z260,
      O => U_DCT1D_rtlc5n1346_17_XORF
    );
  U_DCT1D_rtlc5n1346_17_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_17_CY0F,
      IB => U_DCT1D_rtlc5n1346_17_CYINIT,
      SEL => U_DCT1D_rtlc5n1346_17_CYSELF,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63703_O
    );
  U_DCT1D_rtlc5n1346_17_CYMUXF2_2551 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_17_CY0F,
      IB => U_DCT1D_rtlc5n1346_17_CY0F,
      SEL => U_DCT1D_rtlc5n1346_17_CYSELF,
      O => U_DCT1D_rtlc5n1346_17_CYMUXF2
    );
  U_DCT1D_rtlc5n1346_17_CYINIT_2552 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63707_O,
      O => U_DCT1D_rtlc5n1346_17_CYINIT
    );
  U_DCT1D_rtlc5n1346_17_CY0F_2553 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(13),
      O => U_DCT1D_rtlc5n1346_17_CY0F
    );
  U_DCT1D_rtlc5n1346_17_CYSELF_2554 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z260,
      O => U_DCT1D_rtlc5n1346_17_CYSELF
    );
  U_DCT1D_rtlc5n1346_17_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_17_XORG,
      O => U_DCT1D_rtlc5n1346(18)
    );
  U_DCT1D_rtlc5n1346_17_XORG_2555 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_498_add_23_ix59700z63703_O,
      I1 => U_DCT1D_nx59700z257,
      O => U_DCT1D_rtlc5n1346_17_XORG
    );
  U_DCT1D_rtlc5n1346_17_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_17_CYMUXFAST,
      O => U_DCT1D_rtlc_498_add_23_ix59700z63700_O
    );
  U_DCT1D_rtlc5n1346_17_FASTCARRY_2556 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63707_O,
      O => U_DCT1D_rtlc5n1346_17_FASTCARRY
    );
  U_DCT1D_rtlc5n1346_17_CYAND_2557 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1346_17_CYSELG,
      I1 => U_DCT1D_rtlc5n1346_17_CYSELF,
      O => U_DCT1D_rtlc5n1346_17_CYAND
    );
  U_DCT1D_rtlc5n1346_17_CYMUXFAST_2558 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_17_CYMUXG2,
      IB => U_DCT1D_rtlc5n1346_17_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1346_17_CYAND,
      O => U_DCT1D_rtlc5n1346_17_CYMUXFAST
    );
  U_DCT1D_rtlc5n1346_17_CYMUXG2_2559 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1346_17_CY0G,
      IB => U_DCT1D_rtlc5n1346_17_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1346_17_CYSELG,
      O => U_DCT1D_rtlc5n1346_17_CYMUXG2
    );
  U_DCT1D_rtlc5n1346_17_CY0G_2560 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s(13),
      O => U_DCT1D_rtlc5n1346_17_CY0G
    );
  U_DCT1D_rtlc5n1346_17_CYSELG_2561 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z257,
      O => U_DCT1D_rtlc5n1346_17_CYSELG
    );
  U_DCT1D_nx59700z255_rt_2562 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z255,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z255_rt
    );
  U_DCT1D_rtlc5n1346_19_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1346_19_XORF,
      O => U_DCT1D_rtlc5n1346(19)
    );
  U_DCT1D_rtlc5n1346_19_XORF_2563 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1346_19_CYINIT,
      I1 => U_DCT1D_nx59700z255_rt,
      O => U_DCT1D_rtlc5n1346_19_XORF
    );
  U_DCT1D_rtlc5n1346_19_CYINIT_2564 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_498_add_23_ix59700z63700_O,
      O => U_DCT1D_rtlc5n1346_19_CYINIT
    );
  romodatao4_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_6_F5MUX,
      O => nx54672z943
    );
  romodatao4_s_6_F5MUX_2565 : X_MUX2
    port map (
      IA => nx54672z944,
      IB => nx54672z945,
      SEL => romodatao4_s_6_BXINV,
      O => romodatao4_s_6_F5MUX
    );
  romodatao4_s_6_BXINV_2566 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_6_BXINV
    );
  romodatao4_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_6_F6MUX,
      O => romodatao4_s(6)
    );
  romodatao4_s_6_F6MUX_2567 : X_MUX2
    port map (
      IA => nx54672z940,
      IB => nx54672z943,
      SEL => romodatao4_s_6_BYINV,
      O => romodatao4_s_6_F6MUX
    );
  romodatao4_s_6_BYINV_2568 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_6_BYINV
    );
  ix54672z22871 : X_LUT4
    generic map(
      INIT => X"08CE"
    )
    port map (
      ADR0 => romoaddro4_s(1),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(0),
      ADR3 => romoaddro4_s(2),
      O => nx54672z941
    );
  nx54672z940_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z940_F5MUX,
      O => nx54672z940
    );
  nx54672z940_F5MUX_2569 : X_MUX2
    port map (
      IA => nx54672z941,
      IB => nx54672z942,
      SEL => nx54672z940_BXINV,
      O => nx54672z940_F5MUX
    );
  nx54672z940_BXINV_2570 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z940_BXINV
    );
  U_DCT2D_reg_databuf_reg_7_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_7_0_DYMUX,
      CE => U_DCT2D_databuf_reg_7_0_CEINV,
      CLK => U_DCT2D_databuf_reg_7_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_7_0_FFY_RST,
      O => U_DCT2D_databuf_reg_7_Q(1)
    );
  U_DCT2D_databuf_reg_7_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_7_0_FFY_RST
    );
  romodatao4_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_5_F5MUX,
      O => nx54672z949
    );
  romodatao4_s_5_F5MUX_2571 : X_MUX2
    port map (
      IA => nx54672z950,
      IB => nx54672z951,
      SEL => romodatao4_s_5_BXINV,
      O => romodatao4_s_5_F5MUX
    );
  romodatao4_s_5_BXINV_2572 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_5_BXINV
    );
  romodatao4_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_5_F6MUX,
      O => romodatao4_s(5)
    );
  romodatao4_s_5_F6MUX_2573 : X_MUX2
    port map (
      IA => nx54672z946,
      IB => nx54672z949,
      SEL => romodatao4_s_5_BYINV,
      O => romodatao4_s_5_F6MUX
    );
  romodatao4_s_5_BYINV_2574 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_5_BYINV
    );
  nx54672z946_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z946_F5MUX,
      O => nx54672z946
    );
  nx54672z946_F5MUX_2575 : X_MUX2
    port map (
      IA => nx54672z947,
      IB => nx54672z948,
      SEL => nx54672z946_BXINV,
      O => nx54672z946_F5MUX
    );
  nx54672z946_BXINV_2576 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z946_BXINV
    );
  romodatao4_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_4_F5MUX,
      O => nx54672z955
    );
  romodatao4_s_4_F5MUX_2577 : X_MUX2
    port map (
      IA => nx54672z956,
      IB => nx54672z957,
      SEL => romodatao4_s_4_BXINV,
      O => romodatao4_s_4_F5MUX
    );
  romodatao4_s_4_BXINV_2578 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_4_BXINV
    );
  romodatao4_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_4_F6MUX,
      O => romodatao4_s(4)
    );
  romodatao4_s_4_F6MUX_2579 : X_MUX2
    port map (
      IA => nx54672z952,
      IB => nx54672z955,
      SEL => romodatao4_s_4_BYINV,
      O => romodatao4_s_4_F6MUX
    );
  romodatao4_s_4_BYINV_2580 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_4_BYINV
    );
  nx54672z952_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z952_F5MUX,
      O => nx54672z952
    );
  nx54672z952_F5MUX_2581 : X_MUX2
    port map (
      IA => nx54672z953,
      IB => nx54672z954,
      SEL => nx54672z952_BXINV,
      O => nx54672z952_F5MUX
    );
  nx54672z952_BXINV_2582 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z952_BXINV
    );
  romodatao3_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_12_F5MUX,
      O => nx54672z828
    );
  romodatao3_s_12_F5MUX_2583 : X_MUX2
    port map (
      IA => nx54672z829,
      IB => nx54672z830,
      SEL => romodatao3_s_12_BXINV,
      O => romodatao3_s_12_F5MUX
    );
  romodatao3_s_12_BXINV_2584 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_12_BXINV
    );
  romodatao3_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_12_F6MUX,
      O => romodatao3_s(12)
    );
  romodatao3_s_12_F6MUX_2585 : X_MUX2
    port map (
      IA => nx54672z825,
      IB => nx54672z828,
      SEL => romodatao3_s_12_BYINV,
      O => romodatao3_s_12_F6MUX
    );
  romodatao3_s_12_BYINV_2586 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_12_BYINV
    );
  ix54672z59827 : X_LUT4
    generic map(
      INIT => X"8880"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(1),
      ADR3 => romoaddro3_s(0),
      O => nx54672z826
    );
  nx54672z825_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z825_F5MUX,
      O => nx54672z825
    );
  nx54672z825_F5MUX_2587 : X_MUX2
    port map (
      IA => nx54672z826,
      IB => nx54672z827,
      SEL => nx54672z825_BXINV,
      O => nx54672z825_F5MUX
    );
  nx54672z825_BXINV_2588 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z825_BXINV
    );
  romodatao3_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_10_F5MUX,
      O => nx54672z840
    );
  romodatao3_s_10_F5MUX_2589 : X_MUX2
    port map (
      IA => nx54672z841,
      IB => nx54672z842,
      SEL => romodatao3_s_10_BXINV,
      O => romodatao3_s_10_F5MUX
    );
  romodatao3_s_10_BXINV_2590 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_10_BXINV
    );
  romodatao3_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_10_F6MUX,
      O => romodatao3_s(10)
    );
  romodatao3_s_10_F6MUX_2591 : X_MUX2
    port map (
      IA => nx54672z837,
      IB => nx54672z840,
      SEL => romodatao3_s_10_BYINV,
      O => romodatao3_s_10_F6MUX
    );
  romodatao3_s_10_BYINV_2592 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_10_BYINV
    );
  nx54672z837_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z837_F5MUX,
      O => nx54672z837
    );
  nx54672z837_F5MUX_2593 : X_MUX2
    port map (
      IA => nx54672z838,
      IB => nx54672z839,
      SEL => nx54672z837_BXINV,
      O => nx54672z837_F5MUX
    );
  nx54672z837_BXINV_2594 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z837_BXINV
    );
  romodatao3_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_4_F5MUX,
      O => nx54672z876
    );
  romodatao3_s_4_F5MUX_2595 : X_MUX2
    port map (
      IA => nx54672z877,
      IB => nx54672z878,
      SEL => romodatao3_s_4_BXINV,
      O => romodatao3_s_4_F5MUX
    );
  romodatao3_s_4_BXINV_2596 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_4_BXINV
    );
  romodatao3_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_4_F6MUX,
      O => romodatao3_s(4)
    );
  romodatao3_s_4_F6MUX_2597 : X_MUX2
    port map (
      IA => nx54672z873,
      IB => nx54672z876,
      SEL => romodatao3_s_4_BYINV,
      O => romodatao3_s_4_F6MUX
    );
  romodatao3_s_4_BYINV_2598 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_4_BYINV
    );
  nx54672z873_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z873_F5MUX,
      O => nx54672z873
    );
  nx54672z873_F5MUX_2599 : X_MUX2
    port map (
      IA => nx54672z874,
      IB => nx54672z875,
      SEL => nx54672z873_BXINV,
      O => nx54672z873_F5MUX
    );
  nx54672z873_BXINV_2600 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z873_BXINV
    );
  romodatao3_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_2_F5MUX,
      O => nx54672z888
    );
  romodatao3_s_2_F5MUX_2601 : X_MUX2
    port map (
      IA => nx54672z889,
      IB => nx54672z890,
      SEL => romodatao3_s_2_BXINV,
      O => romodatao3_s_2_F5MUX
    );
  romodatao3_s_2_BXINV_2602 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_2_BXINV
    );
  romodatao3_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_2_F6MUX,
      O => romodatao3_s(2)
    );
  romodatao3_s_2_F6MUX_2603 : X_MUX2
    port map (
      IA => nx54672z885,
      IB => nx54672z888,
      SEL => romodatao3_s_2_BYINV,
      O => romodatao3_s_2_F6MUX
    );
  romodatao3_s_2_BYINV_2604 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_2_BYINV
    );
  nx54672z885_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z885_F5MUX,
      O => nx54672z885
    );
  nx54672z885_F5MUX_2605 : X_MUX2
    port map (
      IA => nx54672z886,
      IB => nx54672z887,
      SEL => nx54672z885_BXINV,
      O => nx54672z885_F5MUX
    );
  nx54672z885_BXINV_2606 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z885_BXINV
    );
  romodatao3_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_0_F5MUX,
      O => U1_ROMO3_modgen_rom_ix0_nx_ro64_32_l
    );
  romodatao3_s_0_F5MUX_2607 : X_MUX2
    port map (
      IA => nx54672z897,
      IB => nx54672z898,
      SEL => romodatao3_s_0_BXINV,
      O => romodatao3_s_0_F5MUX
    );
  romodatao3_s_0_BXINV_2608 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_0_BXINV
    );
  romodatao3_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_0_F6MUX,
      O => romodatao3_s(0)
    );
  romodatao3_s_0_F6MUX_2609 : X_MUX2
    port map (
      IA => U1_ROMO3_modgen_rom_ix0_nx_ro64_32_u,
      IB => U1_ROMO3_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romodatao3_s_0_BYINV,
      O => romodatao3_s_0_F6MUX
    );
  romodatao3_s_0_BYINV_2610 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_0_BYINV
    );
  U1_ROMO3_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROMO3_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U1_ROMO3_modgen_rom_ix0_nx_ro64_32_u
    );
  U1_ROMO3_modgen_rom_ix0_nx_ro64_32_u_F5MUX_2611 : X_MUX2
    port map (
      IA => U1_ROMO3_modgen_rom_ix0_nx_rm64_16_u,
      IB => U1_ROMO3_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U1_ROMO3_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U1_ROMO3_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U1_ROMO3_modgen_rom_ix0_nx_ro64_32_u_BXINV_2612 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => U1_ROMO3_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romodatao2_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_10_F5MUX,
      O => nx54672z761
    );
  romodatao2_s_10_F5MUX_2613 : X_MUX2
    port map (
      IA => nx54672z762,
      IB => nx54672z763,
      SEL => romodatao2_s_10_BXINV,
      O => romodatao2_s_10_F5MUX
    );
  romodatao2_s_10_BXINV_2614 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_10_BXINV
    );
  romodatao2_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_10_F6MUX,
      O => romodatao2_s(10)
    );
  romodatao2_s_10_F6MUX_2615 : X_MUX2
    port map (
      IA => nx54672z758,
      IB => nx54672z761,
      SEL => romodatao2_s_10_BYINV,
      O => romodatao2_s_10_F6MUX
    );
  romodatao2_s_10_BYINV_2616 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_10_BYINV
    );
  U_DCT2D_ix34147z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_3_0_Q,
      ADR1 => U_DCT2D_latchbuf_reg_4_0_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx34147z1
    );
  nx54672z758_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z758_F5MUX,
      O => nx54672z758
    );
  nx54672z758_F5MUX_2617 : X_MUX2
    port map (
      IA => nx54672z759,
      IB => nx54672z760,
      SEL => nx54672z758_BXINV,
      O => nx54672z758_F5MUX
    );
  nx54672z758_BXINV_2618 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z758_BXINV
    );
  romodatao2_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_9_F5MUX,
      O => nx54672z767
    );
  romodatao2_s_9_F5MUX_2619 : X_MUX2
    port map (
      IA => nx54672z768,
      IB => nx54672z769,
      SEL => romodatao2_s_9_BXINV,
      O => romodatao2_s_9_F5MUX
    );
  romodatao2_s_9_BXINV_2620 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_9_BXINV
    );
  romodatao2_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_9_F6MUX,
      O => romodatao2_s(9)
    );
  romodatao2_s_9_F6MUX_2621 : X_MUX2
    port map (
      IA => nx54672z764,
      IB => nx54672z767,
      SEL => romodatao2_s_9_BYINV,
      O => romodatao2_s_9_F6MUX
    );
  romodatao2_s_9_BYINV_2622 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_9_BYINV
    );
  nx54672z764_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z764_F5MUX,
      O => nx54672z764
    );
  nx54672z764_F5MUX_2623 : X_MUX2
    port map (
      IA => nx54672z765,
      IB => nx54672z766,
      SEL => nx54672z764_BXINV,
      O => nx54672z764_F5MUX
    );
  nx54672z764_BXINV_2624 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z764_BXINV
    );
  romodatao2_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_8_F5MUX,
      O => nx54672z773
    );
  romodatao2_s_8_F5MUX_2625 : X_MUX2
    port map (
      IA => nx54672z774,
      IB => nx54672z775,
      SEL => romodatao2_s_8_BXINV,
      O => romodatao2_s_8_F5MUX
    );
  romodatao2_s_8_BXINV_2626 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_8_BXINV
    );
  romodatao2_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_8_F6MUX,
      O => romodatao2_s(8)
    );
  romodatao2_s_8_F6MUX_2627 : X_MUX2
    port map (
      IA => nx54672z770,
      IB => nx54672z773,
      SEL => romodatao2_s_8_BYINV,
      O => romodatao2_s_8_F6MUX
    );
  romodatao2_s_8_BYINV_2628 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_8_BYINV
    );
  nx54672z770_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z770_F5MUX,
      O => nx54672z770
    );
  nx54672z770_F5MUX_2629 : X_MUX2
    port map (
      IA => nx54672z771,
      IB => nx54672z772,
      SEL => nx54672z770_BXINV,
      O => nx54672z770_F5MUX
    );
  nx54672z770_BXINV_2630 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z770_BXINV
    );
  romodatao2_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_7_F5MUX,
      O => nx54672z779
    );
  romodatao2_s_7_F5MUX_2631 : X_MUX2
    port map (
      IA => nx54672z780,
      IB => nx54672z781,
      SEL => romodatao2_s_7_BXINV,
      O => romodatao2_s_7_F5MUX
    );
  romodatao2_s_7_BXINV_2632 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_7_BXINV
    );
  romodatao2_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_7_F6MUX,
      O => romodatao2_s(7)
    );
  romodatao2_s_7_F6MUX_2633 : X_MUX2
    port map (
      IA => nx54672z776,
      IB => nx54672z779,
      SEL => romodatao2_s_7_BYINV,
      O => romodatao2_s_7_F6MUX
    );
  romodatao2_s_7_BYINV_2634 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_7_BYINV
    );
  nx54672z776_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z776_F5MUX,
      O => nx54672z776
    );
  nx54672z776_F5MUX_2635 : X_MUX2
    port map (
      IA => nx54672z777,
      IB => nx54672z778,
      SEL => nx54672z776_BXINV,
      O => nx54672z776_F5MUX
    );
  nx54672z776_BXINV_2636 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z776_BXINV
    );
  romodatao2_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_6_F5MUX,
      O => nx54672z785
    );
  romodatao2_s_6_F5MUX_2637 : X_MUX2
    port map (
      IA => nx54672z786,
      IB => nx54672z787,
      SEL => romodatao2_s_6_BXINV,
      O => romodatao2_s_6_F5MUX
    );
  romodatao2_s_6_BXINV_2638 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_6_BXINV
    );
  romodatao2_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_6_F6MUX,
      O => romodatao2_s(6)
    );
  romodatao2_s_6_F6MUX_2639 : X_MUX2
    port map (
      IA => nx54672z782,
      IB => nx54672z785,
      SEL => romodatao2_s_6_BYINV,
      O => romodatao2_s_6_F6MUX
    );
  romodatao2_s_6_BYINV_2640 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_6_BYINV
    );
  nx54672z782_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z782_F5MUX,
      O => nx54672z782
    );
  nx54672z782_F5MUX_2641 : X_MUX2
    port map (
      IA => nx54672z783,
      IB => nx54672z784,
      SEL => nx54672z782_BXINV,
      O => nx54672z782_F5MUX
    );
  nx54672z782_BXINV_2642 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z782_BXINV
    );
  romodatao4_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_13_F5MUX,
      O => nx54672z901
    );
  romodatao4_s_13_F5MUX_2643 : X_MUX2
    port map (
      IA => nx54672z902,
      IB => nx54672z903,
      SEL => romodatao4_s_13_BXINV,
      O => romodatao4_s_13_F5MUX
    );
  romodatao4_s_13_BXINV_2644 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_13_BXINV
    );
  romodatao4_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_13_F6MUX,
      O => romodatao4_s(13)
    );
  romodatao4_s_13_F6MUX_2645 : X_MUX2
    port map (
      IA => nx54672z899,
      IB => nx54672z901,
      SEL => romodatao4_s_13_BYINV,
      O => romodatao4_s_13_F6MUX
    );
  romodatao4_s_13_BYINV_2646 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_13_BYINV
    );
  nx54672z899_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z899_F5MUX,
      O => nx54672z899
    );
  nx54672z899_F5MUX_2647 : X_MUX2
    port map (
      IA => nx54672z899_G,
      IB => nx54672z900,
      SEL => nx54672z899_BXINV,
      O => nx54672z899_F5MUX
    );
  nx54672z899_BXINV_2648 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z899_BXINV
    );
  romodatao3_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_13_F5MUX,
      O => nx54672z822
    );
  romodatao3_s_13_F5MUX_2649 : X_MUX2
    port map (
      IA => nx54672z823,
      IB => nx54672z824,
      SEL => romodatao3_s_13_BXINV,
      O => romodatao3_s_13_F5MUX
    );
  romodatao3_s_13_BXINV_2650 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_13_BXINV
    );
  romodatao3_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_13_F6MUX,
      O => romodatao3_s(13)
    );
  romodatao3_s_13_F6MUX_2651 : X_MUX2
    port map (
      IA => nx54672z820,
      IB => nx54672z822,
      SEL => romodatao3_s_13_BYINV,
      O => romodatao3_s_13_F6MUX
    );
  romodatao3_s_13_BYINV_2652 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_13_BYINV
    );
  nx54672z820_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z820_F5MUX,
      O => nx54672z820
    );
  nx54672z820_F5MUX_2653 : X_MUX2
    port map (
      IA => nx54672z820_G,
      IB => nx54672z821,
      SEL => nx54672z820_BXINV,
      O => nx54672z820_F5MUX
    );
  nx54672z820_BXINV_2654 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z820_BXINV
    );
  romodatao1_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_5_F5MUX,
      O => nx54672z712
    );
  romodatao1_s_5_F5MUX_2655 : X_MUX2
    port map (
      IA => nx54672z713,
      IB => nx54672z714,
      SEL => romodatao1_s_5_BXINV,
      O => romodatao1_s_5_F5MUX
    );
  romodatao1_s_5_BXINV_2656 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_5_BXINV
    );
  romodatao1_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_5_F6MUX,
      O => romodatao1_s(5)
    );
  romodatao1_s_5_F6MUX_2657 : X_MUX2
    port map (
      IA => nx54672z709,
      IB => nx54672z712,
      SEL => romodatao1_s_5_BYINV,
      O => romodatao1_s_5_F6MUX
    );
  romodatao1_s_5_BYINV_2658 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_5_BYINV
    );
  nx54672z709_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z709_F5MUX,
      O => nx54672z709
    );
  nx54672z709_F5MUX_2659 : X_MUX2
    port map (
      IA => nx54672z710,
      IB => nx54672z711,
      SEL => nx54672z709_BXINV,
      O => nx54672z709_F5MUX
    );
  nx54672z709_BXINV_2660 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z709_BXINV
    );
  romodatao1_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_4_F5MUX,
      O => nx54672z718
    );
  romodatao1_s_4_F5MUX_2661 : X_MUX2
    port map (
      IA => nx54672z719,
      IB => nx54672z720,
      SEL => romodatao1_s_4_BXINV,
      O => romodatao1_s_4_F5MUX
    );
  romodatao1_s_4_BXINV_2662 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_4_BXINV
    );
  romodatao1_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_4_F6MUX,
      O => romodatao1_s(4)
    );
  romodatao1_s_4_F6MUX_2663 : X_MUX2
    port map (
      IA => nx54672z715,
      IB => nx54672z718,
      SEL => romodatao1_s_4_BYINV,
      O => romodatao1_s_4_F6MUX
    );
  romodatao1_s_4_BYINV_2664 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_4_BYINV
    );
  nx54672z715_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z715_F5MUX,
      O => nx54672z715
    );
  nx54672z715_F5MUX_2665 : X_MUX2
    port map (
      IA => nx54672z716,
      IB => nx54672z717,
      SEL => nx54672z715_BXINV,
      O => nx54672z715_F5MUX
    );
  nx54672z715_BXINV_2666 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z715_BXINV
    );
  romodatao1_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_3_F5MUX,
      O => nx54672z724
    );
  romodatao1_s_3_F5MUX_2667 : X_MUX2
    port map (
      IA => nx54672z725,
      IB => nx54672z726,
      SEL => romodatao1_s_3_BXINV,
      O => romodatao1_s_3_F5MUX
    );
  romodatao1_s_3_BXINV_2668 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_3_BXINV
    );
  romodatao1_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_3_F6MUX,
      O => romodatao1_s(3)
    );
  romodatao1_s_3_F6MUX_2669 : X_MUX2
    port map (
      IA => nx54672z721,
      IB => nx54672z724,
      SEL => romodatao1_s_3_BYINV,
      O => romodatao1_s_3_F6MUX
    );
  romodatao1_s_3_BYINV_2670 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_3_BYINV
    );
  U_DCT2D_reg_databuf_reg_7_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_7_0_DXMUX,
      CE => U_DCT2D_databuf_reg_7_0_CEINV,
      CLK => U_DCT2D_databuf_reg_7_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_7_0_FFX_RST,
      O => U_DCT2D_databuf_reg_7_Q(0)
    );
  U_DCT2D_databuf_reg_7_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_7_0_FFX_RST
    );
  nx54672z721_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z721_F5MUX,
      O => nx54672z721
    );
  nx54672z721_F5MUX_2671 : X_MUX2
    port map (
      IA => nx54672z722,
      IB => nx54672z723,
      SEL => nx54672z721_BXINV,
      O => nx54672z721_F5MUX
    );
  nx54672z721_BXINV_2672 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z721_BXINV
    );
  romedatao6_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_13_F5MUX,
      O => nx54672z392
    );
  romedatao6_s_13_F5MUX_2673 : X_MUX2
    port map (
      IA => nx54672z393,
      IB => nx54672z394,
      SEL => romedatao6_s_13_BXINV,
      O => romedatao6_s_13_F5MUX
    );
  romedatao6_s_13_BXINV_2674 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao6_s_13_BXINV
    );
  romedatao6_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_13_F6MUX,
      O => romedatao6_s(13)
    );
  romedatao6_s_13_F6MUX_2675 : X_MUX2
    port map (
      IA => nx54672z390,
      IB => nx54672z392,
      SEL => romedatao6_s_13_BYINV,
      O => romedatao6_s_13_F6MUX
    );
  romedatao6_s_13_BYINV_2676 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao6_s_13_BYINV
    );
  nx54672z390_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z390_F5MUX,
      O => nx54672z390
    );
  nx54672z390_F5MUX_2677 : X_MUX2
    port map (
      IA => nx54672z390_G,
      IB => nx54672z391,
      SEL => nx54672z390_BXINV,
      O => nx54672z390_F5MUX
    );
  nx54672z390_BXINV_2678 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z390_BXINV
    );
  romedatao4_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_12_F5MUX,
      O => nx54672z268
    );
  romedatao4_s_12_F5MUX_2679 : X_MUX2
    port map (
      IA => nx54672z269,
      IB => nx54672z270,
      SEL => romedatao4_s_12_BXINV,
      O => romedatao4_s_12_F5MUX
    );
  romedatao4_s_12_BXINV_2680 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao4_s_12_BXINV
    );
  romedatao4_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_12_F6MUX,
      O => romedatao4_s(12)
    );
  romedatao4_s_12_F6MUX_2681 : X_MUX2
    port map (
      IA => nx54672z265,
      IB => nx54672z268,
      SEL => romedatao4_s_12_BYINV,
      O => romedatao4_s_12_F6MUX
    );
  romedatao4_s_12_BYINV_2682 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao4_s_12_BYINV
    );
  nx54672z265_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z265_F5MUX,
      O => nx54672z265
    );
  nx54672z265_F5MUX_2683 : X_MUX2
    port map (
      IA => nx54672z266,
      IB => nx54672z267,
      SEL => nx54672z265_BXINV,
      O => nx54672z265_F5MUX
    );
  nx54672z265_BXINV_2684 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z265_BXINV
    );
  romedatao4_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_11_F5MUX,
      O => nx54672z274
    );
  romedatao4_s_11_F5MUX_2685 : X_MUX2
    port map (
      IA => nx54672z275,
      IB => nx54672z276,
      SEL => romedatao4_s_11_BXINV,
      O => romedatao4_s_11_F5MUX
    );
  romedatao4_s_11_BXINV_2686 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao4_s_11_BXINV
    );
  romedatao4_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_11_F6MUX,
      O => romedatao4_s(11)
    );
  romedatao4_s_11_F6MUX_2687 : X_MUX2
    port map (
      IA => nx54672z271,
      IB => nx54672z274,
      SEL => romedatao4_s_11_BYINV,
      O => romedatao4_s_11_F6MUX
    );
  romedatao4_s_11_BYINV_2688 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao4_s_11_BYINV
    );
  nx54672z271_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z271_F5MUX,
      O => nx54672z271
    );
  nx54672z271_F5MUX_2689 : X_MUX2
    port map (
      IA => nx54672z272,
      IB => nx54672z273,
      SEL => nx54672z271_BXINV,
      O => nx54672z271_F5MUX
    );
  nx54672z271_BXINV_2690 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z271_BXINV
    );
  romedatao4_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_10_F5MUX,
      O => nx54672z280
    );
  romedatao4_s_10_F5MUX_2691 : X_MUX2
    port map (
      IA => nx54672z281,
      IB => nx54672z282,
      SEL => romedatao4_s_10_BXINV,
      O => romedatao4_s_10_F5MUX
    );
  romedatao4_s_10_BXINV_2692 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao4_s_10_BXINV
    );
  romedatao4_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_10_F6MUX,
      O => romedatao4_s(10)
    );
  romedatao4_s_10_F6MUX_2693 : X_MUX2
    port map (
      IA => nx54672z277,
      IB => nx54672z280,
      SEL => romedatao4_s_10_BYINV,
      O => romedatao4_s_10_F6MUX
    );
  romedatao4_s_10_BYINV_2694 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao4_s_10_BYINV
    );
  nx54672z277_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z277_F5MUX,
      O => nx54672z277
    );
  nx54672z277_F5MUX_2695 : X_MUX2
    port map (
      IA => nx54672z278,
      IB => nx54672z279,
      SEL => nx54672z277_BXINV,
      O => nx54672z277_F5MUX
    );
  nx54672z277_BXINV_2696 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z277_BXINV
    );
  romedatao4_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_4_F5MUX,
      O => nx54672z316
    );
  romedatao4_s_4_F5MUX_2697 : X_MUX2
    port map (
      IA => nx54672z317,
      IB => nx54672z318,
      SEL => romedatao4_s_4_BXINV,
      O => romedatao4_s_4_F5MUX
    );
  romedatao4_s_4_BXINV_2698 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao4_s_4_BXINV
    );
  romedatao4_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_4_F6MUX,
      O => romedatao4_s(4)
    );
  romedatao4_s_4_F6MUX_2699 : X_MUX2
    port map (
      IA => nx54672z313,
      IB => nx54672z316,
      SEL => romedatao4_s_4_BYINV,
      O => romedatao4_s_4_F6MUX
    );
  romedatao4_s_4_BYINV_2700 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao4_s_4_BYINV
    );
  U_DCT2D_ix37138z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_3_3_Q,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_4_3_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx37138z1
    );
  U_DCT1D_nx59700z428_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z428_XORF,
      O => U_DCT1D_nx59700z428
    );
  U_DCT1D_nx59700z428_XORF_2701 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z428_CYINIT,
      I1 => U_DCT1D_nx59700z428_F,
      O => U_DCT1D_nx59700z428_XORF
    );
  U_DCT1D_nx59700z428_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z428_CY0F,
      IB => U_DCT1D_nx59700z428_CYINIT,
      SEL => U_DCT1D_nx59700z428_CYSELF,
      O => U_DCT1D_ix740_modgen_add_290_ix59700z63793_O
    );
  U_DCT1D_nx59700z428_CYINIT_2702 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z428_BXINVNOT,
      O => U_DCT1D_nx59700z428_CYINIT
    );
  U_DCT1D_nx59700z428_CY0F_2703 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z333,
      O => U_DCT1D_nx59700z428_CY0F
    );
  U_DCT1D_nx59700z428_CYSELF_2704 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z428_F,
      O => U_DCT1D_nx59700z428_CYSELF
    );
  U_DCT1D_nx59700z428_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_2,
      O => U_DCT1D_nx59700z428_BXINVNOT
    );
  U_DCT1D_nx59700z428_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z428_XORG,
      O => U_DCT1D_nx59700z424
    );
  U_DCT1D_nx59700z428_XORG_2705 : X_XOR2
    port map (
      I0 => U_DCT1D_ix740_modgen_add_290_ix59700z63793_O,
      I1 => U_DCT1D_nx59700z329,
      O => U_DCT1D_nx59700z428_XORG
    );
  U_DCT1D_nx59700z428_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z428_CYMUXG,
      O => U_DCT1D_ix740_modgen_add_290_ix59700z63789_O
    );
  U_DCT1D_nx59700z428_CYMUXG_2706 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z428_CY0G,
      IB => U_DCT1D_ix740_modgen_add_290_ix59700z63793_O,
      SEL => U_DCT1D_nx59700z428_CYSELG,
      O => U_DCT1D_nx59700z428_CYMUXG
    );
  U_DCT1D_nx59700z428_CY0G_2707 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z330,
      O => U_DCT1D_nx59700z428_CY0G
    );
  U_DCT1D_nx59700z428_CYSELG_2708 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z329,
      O => U_DCT1D_nx59700z428_CYSELG
    );
  U_DCT1D_reg_databuf_reg_2_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_2_6_DYMUX,
      CE => U_DCT1D_databuf_reg_2_6_CEINV,
      CLK => U_DCT1D_databuf_reg_2_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_2_6_FFY_RST,
      O => U_DCT1D_databuf_reg_2_Q(7)
    );
  U_DCT1D_databuf_reg_2_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_2_6_FFY_RST
    );
  U_DCT1D_nx59700z420_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z420_XORF,
      O => U_DCT1D_nx59700z420
    );
  U_DCT1D_nx59700z420_XORF_2709 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z420_CYINIT,
      I1 => U_DCT1D_nx59700z326,
      O => U_DCT1D_nx59700z420_XORF
    );
  U_DCT1D_nx59700z420_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z420_CY0F,
      IB => U_DCT1D_nx59700z420_CYINIT,
      SEL => U_DCT1D_nx59700z420_CYSELF,
      O => U_DCT1D_ix740_modgen_add_290_ix59700z63785_O
    );
  U_DCT1D_nx59700z420_CYMUXF2_2710 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z420_CY0F,
      IB => U_DCT1D_nx59700z420_CY0F,
      SEL => U_DCT1D_nx59700z420_CYSELF,
      O => U_DCT1D_nx59700z420_CYMUXF2
    );
  U_DCT1D_nx59700z420_CYINIT_2711 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix740_modgen_add_290_ix59700z63789_O,
      O => U_DCT1D_nx59700z420_CYINIT
    );
  U_DCT1D_nx59700z420_CY0F_2712 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z327,
      O => U_DCT1D_nx59700z420_CY0F
    );
  U_DCT1D_nx59700z420_CYSELF_2713 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z326,
      O => U_DCT1D_nx59700z420_CYSELF
    );
  U_DCT1D_nx59700z420_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z420_XORG,
      O => U_DCT1D_nx59700z416
    );
  U_DCT1D_nx59700z420_XORG_2714 : X_XOR2
    port map (
      I0 => U_DCT1D_ix740_modgen_add_290_ix59700z63785_O,
      I1 => U_DCT1D_nx59700z323,
      O => U_DCT1D_nx59700z420_XORG
    );
  U_DCT1D_nx59700z420_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z420_CYMUXFAST,
      O => U_DCT1D_ix740_modgen_add_290_ix59700z63781_O
    );
  U_DCT1D_nx59700z420_FASTCARRY_2715 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix740_modgen_add_290_ix59700z63789_O,
      O => U_DCT1D_nx59700z420_FASTCARRY
    );
  U_DCT1D_nx59700z420_CYAND_2716 : X_AND2
    port map (
      I0 => U_DCT1D_nx59700z420_CYSELG,
      I1 => U_DCT1D_nx59700z420_CYSELF,
      O => U_DCT1D_nx59700z420_CYAND
    );
  U_DCT1D_nx59700z420_CYMUXFAST_2717 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z420_CYMUXG2,
      IB => U_DCT1D_nx59700z420_FASTCARRY,
      SEL => U_DCT1D_nx59700z420_CYAND,
      O => U_DCT1D_nx59700z420_CYMUXFAST
    );
  U_DCT1D_nx59700z420_CYMUXG2_2718 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z420_CY0G,
      IB => U_DCT1D_nx59700z420_CYMUXF2,
      SEL => U_DCT1D_nx59700z420_CYSELG,
      O => U_DCT1D_nx59700z420_CYMUXG2
    );
  U_DCT1D_nx59700z420_CY0G_2719 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z324,
      O => U_DCT1D_nx59700z420_CY0G
    );
  U_DCT1D_nx59700z420_CYSELG_2720 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z323,
      O => U_DCT1D_nx59700z420_CYSELG
    );
  U_DCT1D_nx59700z412_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z412_XORF,
      O => U_DCT1D_nx59700z412
    );
  U_DCT1D_nx59700z412_XORF_2721 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z412_CYINIT,
      I1 => U_DCT1D_nx59700z320,
      O => U_DCT1D_nx59700z412_XORF
    );
  U_DCT1D_nx59700z412_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z412_CY0F,
      IB => U_DCT1D_nx59700z412_CYINIT,
      SEL => U_DCT1D_nx59700z412_CYSELF,
      O => U_DCT1D_ix740_modgen_add_290_ix59700z63777_O
    );
  U_DCT1D_nx59700z412_CYMUXF2_2722 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z412_CY0F,
      IB => U_DCT1D_nx59700z412_CY0F,
      SEL => U_DCT1D_nx59700z412_CYSELF,
      O => U_DCT1D_nx59700z412_CYMUXF2
    );
  U_DCT1D_nx59700z412_CYINIT_2723 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix740_modgen_add_290_ix59700z63781_O,
      O => U_DCT1D_nx59700z412_CYINIT
    );
  U_DCT1D_nx59700z412_CY0F_2724 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z321,
      O => U_DCT1D_nx59700z412_CY0F
    );
  U_DCT1D_nx59700z412_CYSELF_2725 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z320,
      O => U_DCT1D_nx59700z412_CYSELF
    );
  U_DCT1D_nx59700z412_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z412_XORG,
      O => U_DCT1D_nx59700z408
    );
  U_DCT1D_nx59700z412_XORG_2726 : X_XOR2
    port map (
      I0 => U_DCT1D_ix740_modgen_add_290_ix59700z63777_O,
      I1 => U_DCT1D_nx59700z317,
      O => U_DCT1D_nx59700z412_XORG
    );
  U_DCT1D_nx59700z412_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z412_CYMUXFAST,
      O => U_DCT1D_ix740_modgen_add_290_ix59700z63773_O
    );
  U_DCT1D_nx59700z412_FASTCARRY_2727 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix740_modgen_add_290_ix59700z63781_O,
      O => U_DCT1D_nx59700z412_FASTCARRY
    );
  U_DCT1D_nx59700z412_CYAND_2728 : X_AND2
    port map (
      I0 => U_DCT1D_nx59700z412_CYSELG,
      I1 => U_DCT1D_nx59700z412_CYSELF,
      O => U_DCT1D_nx59700z412_CYAND
    );
  U_DCT1D_nx59700z412_CYMUXFAST_2729 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z412_CYMUXG2,
      IB => U_DCT1D_nx59700z412_FASTCARRY,
      SEL => U_DCT1D_nx59700z412_CYAND,
      O => U_DCT1D_nx59700z412_CYMUXFAST
    );
  U_DCT1D_nx59700z412_CYMUXG2_2730 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z412_CY0G,
      IB => U_DCT1D_nx59700z412_CYMUXF2,
      SEL => U_DCT1D_nx59700z412_CYSELG,
      O => U_DCT1D_nx59700z412_CYMUXG2
    );
  U_DCT1D_nx59700z412_CY0G_2731 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z318,
      O => U_DCT1D_nx59700z412_CY0G
    );
  U_DCT1D_nx59700z412_CYSELG_2732 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z317,
      O => U_DCT1D_nx59700z412_CYSELG
    );
  U_DCT1D_nx59700z404_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z404_XORF,
      O => U_DCT1D_nx59700z404
    );
  U_DCT1D_nx59700z404_XORF_2733 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z404_CYINIT,
      I1 => U_DCT1D_nx59700z314,
      O => U_DCT1D_nx59700z404_XORF
    );
  U_DCT1D_nx59700z404_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z404_CY0F,
      IB => U_DCT1D_nx59700z404_CYINIT,
      SEL => U_DCT1D_nx59700z404_CYSELF,
      O => U_DCT1D_ix740_modgen_add_290_ix59700z63769_O
    );
  U_DCT1D_nx59700z404_CYMUXF2_2734 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z404_CY0F,
      IB => U_DCT1D_nx59700z404_CY0F,
      SEL => U_DCT1D_nx59700z404_CYSELF,
      O => U_DCT1D_nx59700z404_CYMUXF2
    );
  U_DCT1D_nx59700z404_CYINIT_2735 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix740_modgen_add_290_ix59700z63773_O,
      O => U_DCT1D_nx59700z404_CYINIT
    );
  U_DCT1D_nx59700z404_CY0F_2736 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z315,
      O => U_DCT1D_nx59700z404_CY0F
    );
  U_DCT1D_nx59700z404_CYSELF_2737 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z314,
      O => U_DCT1D_nx59700z404_CYSELF
    );
  U_DCT1D_nx59700z404_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z404_XORG,
      O => U_DCT1D_nx59700z400
    );
  U_DCT1D_nx59700z404_XORG_2738 : X_XOR2
    port map (
      I0 => U_DCT1D_ix740_modgen_add_290_ix59700z63769_O,
      I1 => U_DCT1D_nx59700z311,
      O => U_DCT1D_nx59700z404_XORG
    );
  U_DCT1D_nx59700z404_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z404_CYMUXFAST,
      O => U_DCT1D_ix740_modgen_add_290_ix59700z63765_O
    );
  U_DCT1D_nx59700z404_FASTCARRY_2739 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix740_modgen_add_290_ix59700z63773_O,
      O => U_DCT1D_nx59700z404_FASTCARRY
    );
  U_DCT1D_nx59700z404_CYAND_2740 : X_AND2
    port map (
      I0 => U_DCT1D_nx59700z404_CYSELG,
      I1 => U_DCT1D_nx59700z404_CYSELF,
      O => U_DCT1D_nx59700z404_CYAND
    );
  U_DCT1D_nx59700z404_CYMUXFAST_2741 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z404_CYMUXG2,
      IB => U_DCT1D_nx59700z404_FASTCARRY,
      SEL => U_DCT1D_nx59700z404_CYAND,
      O => U_DCT1D_nx59700z404_CYMUXFAST
    );
  U_DCT1D_nx59700z404_CYMUXG2_2742 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z404_CY0G,
      IB => U_DCT1D_nx59700z404_CYMUXF2,
      SEL => U_DCT1D_nx59700z404_CYSELG,
      O => U_DCT1D_nx59700z404_CYMUXG2
    );
  U_DCT1D_nx59700z404_CY0G_2743 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z312,
      O => U_DCT1D_nx59700z404_CY0G
    );
  U_DCT1D_nx59700z404_CYSELG_2744 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z311,
      O => U_DCT1D_nx59700z404_CYSELG
    );
  U_DCT1D_nx59700z396_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z396_XORF,
      O => U_DCT1D_nx59700z396
    );
  U_DCT1D_nx59700z396_XORF_2745 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z396_CYINIT,
      I1 => U_DCT1D_nx59700z308,
      O => U_DCT1D_nx59700z396_XORF
    );
  U_DCT1D_nx59700z396_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z396_CY0F,
      IB => U_DCT1D_nx59700z396_CYINIT,
      SEL => U_DCT1D_nx59700z396_CYSELF,
      O => U_DCT1D_ix740_modgen_add_290_ix59700z63761_O
    );
  U_DCT1D_nx59700z396_CYMUXF2_2746 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z396_CY0F,
      IB => U_DCT1D_nx59700z396_CY0F,
      SEL => U_DCT1D_nx59700z396_CYSELF,
      O => U_DCT1D_nx59700z396_CYMUXF2
    );
  U_DCT1D_nx59700z396_CYINIT_2747 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix740_modgen_add_290_ix59700z63765_O,
      O => U_DCT1D_nx59700z396_CYINIT
    );
  U_DCT1D_nx59700z396_CY0F_2748 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z309,
      O => U_DCT1D_nx59700z396_CY0F
    );
  U_DCT1D_nx59700z396_CYSELF_2749 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z308,
      O => U_DCT1D_nx59700z396_CYSELF
    );
  U_DCT1D_nx59700z396_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z396_XORG,
      O => U_DCT1D_nx59700z392
    );
  U_DCT1D_nx59700z396_XORG_2750 : X_XOR2
    port map (
      I0 => U_DCT1D_ix740_modgen_add_290_ix59700z63761_O,
      I1 => U_DCT1D_nx59700z305,
      O => U_DCT1D_nx59700z396_XORG
    );
  U_DCT1D_nx59700z396_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z396_CYMUXFAST,
      O => U_DCT1D_ix740_modgen_add_290_ix59700z63757_O
    );
  U_DCT1D_nx59700z396_FASTCARRY_2751 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix740_modgen_add_290_ix59700z63765_O,
      O => U_DCT1D_nx59700z396_FASTCARRY
    );
  U_DCT1D_nx59700z396_CYAND_2752 : X_AND2
    port map (
      I0 => U_DCT1D_nx59700z396_CYSELG,
      I1 => U_DCT1D_nx59700z396_CYSELF,
      O => U_DCT1D_nx59700z396_CYAND
    );
  U_DCT1D_nx59700z396_CYMUXFAST_2753 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z396_CYMUXG2,
      IB => U_DCT1D_nx59700z396_FASTCARRY,
      SEL => U_DCT1D_nx59700z396_CYAND,
      O => U_DCT1D_nx59700z396_CYMUXFAST
    );
  U_DCT1D_nx59700z396_CYMUXG2_2754 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z396_CY0G,
      IB => U_DCT1D_nx59700z396_CYMUXF2,
      SEL => U_DCT1D_nx59700z396_CYSELG,
      O => U_DCT1D_nx59700z396_CYMUXG2
    );
  U_DCT1D_nx59700z396_CY0G_2755 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z306,
      O => U_DCT1D_nx59700z396_CY0G
    );
  U_DCT1D_nx59700z396_CYSELG_2756 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z305,
      O => U_DCT1D_nx59700z396_CYSELG
    );
  U_DCT1D_nx59700z388_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z388_XORF,
      O => U_DCT1D_nx59700z388
    );
  U_DCT1D_nx59700z388_XORF_2757 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z388_CYINIT,
      I1 => U_DCT1D_nx59700z302,
      O => U_DCT1D_nx59700z388_XORF
    );
  U_DCT1D_nx59700z388_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z388_CY0F,
      IB => U_DCT1D_nx59700z388_CYINIT,
      SEL => U_DCT1D_nx59700z388_CYSELF,
      O => U_DCT1D_ix740_modgen_add_290_ix59700z63753_O
    );
  U_DCT1D_nx59700z388_CYMUXF2_2758 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z388_CY0F,
      IB => U_DCT1D_nx59700z388_CY0F,
      SEL => U_DCT1D_nx59700z388_CYSELF,
      O => U_DCT1D_nx59700z388_CYMUXF2
    );
  U_DCT1D_nx59700z388_CYINIT_2759 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix740_modgen_add_290_ix59700z63757_O,
      O => U_DCT1D_nx59700z388_CYINIT
    );
  U_DCT1D_nx59700z388_CY0F_2760 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z303,
      O => U_DCT1D_nx59700z388_CY0F
    );
  U_DCT1D_nx59700z388_CYSELF_2761 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z302,
      O => U_DCT1D_nx59700z388_CYSELF
    );
  U_DCT1D_nx59700z388_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z388_XORG,
      O => U_DCT1D_nx59700z384
    );
  U_DCT1D_nx59700z388_XORG_2762 : X_XOR2
    port map (
      I0 => U_DCT1D_ix740_modgen_add_290_ix59700z63753_O,
      I1 => U_DCT1D_nx59700z299,
      O => U_DCT1D_nx59700z388_XORG
    );
  U_DCT1D_nx59700z388_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z388_CYMUXFAST,
      O => U_DCT1D_ix740_modgen_add_290_ix59700z63749_O
    );
  U_DCT1D_nx59700z388_FASTCARRY_2763 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix740_modgen_add_290_ix59700z63757_O,
      O => U_DCT1D_nx59700z388_FASTCARRY
    );
  U_DCT1D_nx59700z388_CYAND_2764 : X_AND2
    port map (
      I0 => U_DCT1D_nx59700z388_CYSELG,
      I1 => U_DCT1D_nx59700z388_CYSELF,
      O => U_DCT1D_nx59700z388_CYAND
    );
  U_DCT1D_nx59700z388_CYMUXFAST_2765 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z388_CYMUXG2,
      IB => U_DCT1D_nx59700z388_FASTCARRY,
      SEL => U_DCT1D_nx59700z388_CYAND,
      O => U_DCT1D_nx59700z388_CYMUXFAST
    );
  U_DCT1D_nx59700z388_CYMUXG2_2766 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z388_CY0G,
      IB => U_DCT1D_nx59700z388_CYMUXF2,
      SEL => U_DCT1D_nx59700z388_CYSELG,
      O => U_DCT1D_nx59700z388_CYMUXG2
    );
  U_DCT1D_nx59700z388_CY0G_2767 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z300,
      O => U_DCT1D_nx59700z388_CY0G
    );
  U_DCT1D_nx59700z388_CYSELG_2768 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z299,
      O => U_DCT1D_nx59700z388_CYSELG
    );
  U_DCT1D_nx59700z254_rt_2769 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z254,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z254_rt
    );
  U_DCT1D_nx59700z253_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z253_XORF,
      O => U_DCT1D_nx59700z253
    );
  U_DCT1D_nx59700z253_XORF_2770 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z253_CYINIT,
      I1 => U_DCT1D_nx59700z254_rt,
      O => U_DCT1D_nx59700z253_XORF
    );
  U_DCT1D_nx59700z253_CYINIT_2771 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix740_modgen_add_290_ix59700z63749_O,
      O => U_DCT1D_nx59700z253_CYINIT
    );
  U_DCT2D_rtlc5n1494_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_7_XORF,
      O => U_DCT2D_rtlc5n1494(7)
    );
  U_DCT2D_rtlc5n1494_7_XORF_2772 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1494_7_CYINIT,
      I1 => U_DCT2D_nx65206z332,
      O => U_DCT2D_rtlc5n1494_7_XORF
    );
  U_DCT2D_rtlc5n1494_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_7_CY0F,
      IB => U_DCT2D_rtlc5n1494_7_CYINIT,
      SEL => U_DCT2D_rtlc5n1494_7_CYSELF,
      O => U_DCT2D_rtlc_394_add_67_ix65206z63792_O
    );
  U_DCT2D_rtlc5n1494_7_CYINIT_2773 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_7_BXINVNOT,
      O => U_DCT2D_rtlc5n1494_7_CYINIT
    );
  U_DCT2D_rtlc5n1494_7_CY0F_2774 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s(3),
      O => U_DCT2D_rtlc5n1494_7_CY0F
    );
  U_DCT2D_rtlc5n1494_7_CYSELF_2775 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z332,
      O => U_DCT2D_rtlc5n1494_7_CYSELF
    );
  U_DCT2D_rtlc5n1494_7_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_3,
      O => U_DCT2D_rtlc5n1494_7_BXINVNOT
    );
  U_DCT2D_rtlc5n1494_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_7_XORG,
      O => U_DCT2D_rtlc5n1494(8)
    );
  U_DCT2D_rtlc5n1494_7_XORG_2776 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_394_add_67_ix65206z63792_O,
      I1 => U_DCT2D_nx65206z329,
      O => U_DCT2D_rtlc5n1494_7_XORG
    );
  U_DCT2D_rtlc5n1494_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_7_CYMUXG,
      O => U_DCT2D_rtlc_394_add_67_ix65206z63788_O
    );
  U_DCT2D_rtlc5n1494_7_CYMUXG_2777 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_7_CY0G,
      IB => U_DCT2D_rtlc_394_add_67_ix65206z63792_O,
      SEL => U_DCT2D_rtlc5n1494_7_CYSELG,
      O => U_DCT2D_rtlc5n1494_7_CYMUXG
    );
  U_DCT2D_rtlc5n1494_7_CY0G_2778 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s(4),
      O => U_DCT2D_rtlc5n1494_7_CY0G
    );
  U_DCT2D_rtlc5n1494_7_CYSELG_2779 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z329,
      O => U_DCT2D_rtlc5n1494_7_CYSELG
    );
  U_DCT2D_rtlc5n1494_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_9_XORF,
      O => U_DCT2D_rtlc5n1494(9)
    );
  U_DCT2D_rtlc5n1494_9_XORF_2780 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1494_9_CYINIT,
      I1 => U_DCT2D_nx65206z326,
      O => U_DCT2D_rtlc5n1494_9_XORF
    );
  U_DCT2D_rtlc5n1494_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_9_CY0F,
      IB => U_DCT2D_rtlc5n1494_9_CYINIT,
      SEL => U_DCT2D_rtlc5n1494_9_CYSELF,
      O => U_DCT2D_rtlc_394_add_67_ix65206z63784_O
    );
  U_DCT2D_rtlc5n1494_9_CYMUXF2_2781 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_9_CY0F,
      IB => U_DCT2D_rtlc5n1494_9_CY0F,
      SEL => U_DCT2D_rtlc5n1494_9_CYSELF,
      O => U_DCT2D_rtlc5n1494_9_CYMUXF2
    );
  U_DCT2D_rtlc5n1494_9_CYINIT_2782 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_394_add_67_ix65206z63788_O,
      O => U_DCT2D_rtlc5n1494_9_CYINIT
    );
  U_DCT2D_rtlc5n1494_9_CY0F_2783 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s(5),
      O => U_DCT2D_rtlc5n1494_9_CY0F
    );
  U_DCT2D_rtlc5n1494_9_CYSELF_2784 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z326,
      O => U_DCT2D_rtlc5n1494_9_CYSELF
    );
  U_DCT2D_rtlc5n1494_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_9_XORG,
      O => U_DCT2D_rtlc5n1494(10)
    );
  U_DCT2D_rtlc5n1494_9_XORG_2785 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_394_add_67_ix65206z63784_O,
      I1 => U_DCT2D_nx65206z323,
      O => U_DCT2D_rtlc5n1494_9_XORG
    );
  U_DCT2D_rtlc5n1494_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_9_CYMUXFAST,
      O => U_DCT2D_rtlc_394_add_67_ix65206z63781_O
    );
  U_DCT2D_rtlc5n1494_9_FASTCARRY_2786 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_394_add_67_ix65206z63788_O,
      O => U_DCT2D_rtlc5n1494_9_FASTCARRY
    );
  U_DCT2D_rtlc5n1494_9_CYAND_2787 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1494_9_CYSELG,
      I1 => U_DCT2D_rtlc5n1494_9_CYSELF,
      O => U_DCT2D_rtlc5n1494_9_CYAND
    );
  U_DCT2D_rtlc5n1494_9_CYMUXFAST_2788 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_9_CYMUXG2,
      IB => U_DCT2D_rtlc5n1494_9_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1494_9_CYAND,
      O => U_DCT2D_rtlc5n1494_9_CYMUXFAST
    );
  U_DCT2D_rtlc5n1494_9_CYMUXG2_2789 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_9_CY0G,
      IB => U_DCT2D_rtlc5n1494_9_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1494_9_CYSELG,
      O => U_DCT2D_rtlc5n1494_9_CYMUXG2
    );
  U_DCT2D_rtlc5n1494_9_CY0G_2790 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s(6),
      O => U_DCT2D_rtlc5n1494_9_CY0G
    );
  U_DCT2D_rtlc5n1494_9_CYSELG_2791 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z323,
      O => U_DCT2D_rtlc5n1494_9_CYSELG
    );
  U_DCT2D_rtlc5n1494_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_11_XORF,
      O => U_DCT2D_rtlc5n1494(11)
    );
  U_DCT2D_rtlc5n1494_11_XORF_2792 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1494_11_CYINIT,
      I1 => U_DCT2D_nx65206z320,
      O => U_DCT2D_rtlc5n1494_11_XORF
    );
  U_DCT2D_rtlc5n1494_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_11_CY0F,
      IB => U_DCT2D_rtlc5n1494_11_CYINIT,
      SEL => U_DCT2D_rtlc5n1494_11_CYSELF,
      O => U_DCT2D_rtlc_394_add_67_ix65206z63777_O
    );
  U_DCT2D_rtlc5n1494_11_CYMUXF2_2793 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_11_CY0F,
      IB => U_DCT2D_rtlc5n1494_11_CY0F,
      SEL => U_DCT2D_rtlc5n1494_11_CYSELF,
      O => U_DCT2D_rtlc5n1494_11_CYMUXF2
    );
  U_DCT2D_rtlc5n1494_11_CYINIT_2794 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_394_add_67_ix65206z63781_O,
      O => U_DCT2D_rtlc5n1494_11_CYINIT
    );
  U_DCT2D_rtlc5n1494_11_CY0F_2795 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s(7),
      O => U_DCT2D_rtlc5n1494_11_CY0F
    );
  U_DCT2D_rtlc5n1494_11_CYSELF_2796 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z320,
      O => U_DCT2D_rtlc5n1494_11_CYSELF
    );
  U_DCT2D_rtlc5n1494_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_11_XORG,
      O => U_DCT2D_rtlc5n1494(12)
    );
  U_DCT2D_rtlc5n1494_11_XORG_2797 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_394_add_67_ix65206z63777_O,
      I1 => U_DCT2D_nx65206z317,
      O => U_DCT2D_rtlc5n1494_11_XORG
    );
  U_DCT2D_rtlc5n1494_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_11_CYMUXFAST,
      O => U_DCT2D_rtlc_394_add_67_ix65206z63774_O
    );
  U_DCT2D_rtlc5n1494_11_FASTCARRY_2798 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_394_add_67_ix65206z63781_O,
      O => U_DCT2D_rtlc5n1494_11_FASTCARRY
    );
  U_DCT2D_rtlc5n1494_11_CYAND_2799 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1494_11_CYSELG,
      I1 => U_DCT2D_rtlc5n1494_11_CYSELF,
      O => U_DCT2D_rtlc5n1494_11_CYAND
    );
  U_DCT2D_rtlc5n1494_11_CYMUXFAST_2800 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_11_CYMUXG2,
      IB => U_DCT2D_rtlc5n1494_11_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1494_11_CYAND,
      O => U_DCT2D_rtlc5n1494_11_CYMUXFAST
    );
  U_DCT2D_rtlc5n1494_11_CYMUXG2_2801 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_11_CY0G,
      IB => U_DCT2D_rtlc5n1494_11_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1494_11_CYSELG,
      O => U_DCT2D_rtlc5n1494_11_CYMUXG2
    );
  U_DCT2D_rtlc5n1494_11_CY0G_2802 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s(8),
      O => U_DCT2D_rtlc5n1494_11_CY0G
    );
  U_DCT2D_rtlc5n1494_11_CYSELG_2803 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z317,
      O => U_DCT2D_rtlc5n1494_11_CYSELG
    );
  U_DCT2D_rtlc5n1494_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_13_XORF,
      O => U_DCT2D_rtlc5n1494(13)
    );
  U_DCT2D_rtlc5n1494_13_XORF_2804 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1494_13_CYINIT,
      I1 => U_DCT2D_nx65206z314,
      O => U_DCT2D_rtlc5n1494_13_XORF
    );
  U_DCT2D_rtlc5n1494_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_13_CY0F,
      IB => U_DCT2D_rtlc5n1494_13_CYINIT,
      SEL => U_DCT2D_rtlc5n1494_13_CYSELF,
      O => U_DCT2D_rtlc_394_add_67_ix65206z63770_O
    );
  U_DCT2D_rtlc5n1494_13_CYMUXF2_2805 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_13_CY0F,
      IB => U_DCT2D_rtlc5n1494_13_CY0F,
      SEL => U_DCT2D_rtlc5n1494_13_CYSELF,
      O => U_DCT2D_rtlc5n1494_13_CYMUXF2
    );
  U_DCT2D_rtlc5n1494_13_CYINIT_2806 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_394_add_67_ix65206z63774_O,
      O => U_DCT2D_rtlc5n1494_13_CYINIT
    );
  U_DCT2D_rtlc5n1494_13_CY0F_2807 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s(9),
      O => U_DCT2D_rtlc5n1494_13_CY0F
    );
  U_DCT2D_rtlc5n1494_13_CYSELF_2808 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z314,
      O => U_DCT2D_rtlc5n1494_13_CYSELF
    );
  U_DCT2D_rtlc5n1494_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_13_XORG,
      O => U_DCT2D_rtlc5n1494(14)
    );
  U_DCT2D_rtlc5n1494_13_XORG_2809 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_394_add_67_ix65206z63770_O,
      I1 => U_DCT2D_nx65206z311,
      O => U_DCT2D_rtlc5n1494_13_XORG
    );
  U_DCT2D_rtlc5n1494_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_13_CYMUXFAST,
      O => U_DCT2D_rtlc_394_add_67_ix65206z63767_O
    );
  U_DCT2D_rtlc5n1494_13_FASTCARRY_2810 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_394_add_67_ix65206z63774_O,
      O => U_DCT2D_rtlc5n1494_13_FASTCARRY
    );
  U_DCT2D_rtlc5n1494_13_CYAND_2811 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1494_13_CYSELG,
      I1 => U_DCT2D_rtlc5n1494_13_CYSELF,
      O => U_DCT2D_rtlc5n1494_13_CYAND
    );
  U_DCT2D_rtlc5n1494_13_CYMUXFAST_2812 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_13_CYMUXG2,
      IB => U_DCT2D_rtlc5n1494_13_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1494_13_CYAND,
      O => U_DCT2D_rtlc5n1494_13_CYMUXFAST
    );
  U_DCT2D_rtlc5n1494_13_CYMUXG2_2813 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_13_CY0G,
      IB => U_DCT2D_rtlc5n1494_13_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1494_13_CYSELG,
      O => U_DCT2D_rtlc5n1494_13_CYMUXG2
    );
  U_DCT2D_rtlc5n1494_13_CY0G_2814 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s(10),
      O => U_DCT2D_rtlc5n1494_13_CY0G
    );
  U_DCT2D_rtlc5n1494_13_CYSELG_2815 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z311,
      O => U_DCT2D_rtlc5n1494_13_CYSELG
    );
  U_DCT1D_ix268z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_2_Q(6),
      ADR1 => U_DCT1D_latchbuf_reg_5_Q(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx268z1
    );
  U_DCT2D_rtlc5n1494_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_15_XORF,
      O => U_DCT2D_rtlc5n1494(15)
    );
  U_DCT2D_rtlc5n1494_15_XORF_2816 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1494_15_CYINIT,
      I1 => U_DCT2D_nx65206z308,
      O => U_DCT2D_rtlc5n1494_15_XORF
    );
  U_DCT2D_rtlc5n1494_15_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_15_CY0F,
      IB => U_DCT2D_rtlc5n1494_15_CYINIT,
      SEL => U_DCT2D_rtlc5n1494_15_CYSELF,
      O => U_DCT2D_rtlc_394_add_67_ix65206z63763_O
    );
  U_DCT2D_rtlc5n1494_15_CYMUXF2_2817 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_15_CY0F,
      IB => U_DCT2D_rtlc5n1494_15_CY0F,
      SEL => U_DCT2D_rtlc5n1494_15_CYSELF,
      O => U_DCT2D_rtlc5n1494_15_CYMUXF2
    );
  U_DCT2D_rtlc5n1494_15_CYINIT_2818 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_394_add_67_ix65206z63767_O,
      O => U_DCT2D_rtlc5n1494_15_CYINIT
    );
  U_DCT2D_rtlc5n1494_15_CY0F_2819 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s(11),
      O => U_DCT2D_rtlc5n1494_15_CY0F
    );
  U_DCT2D_rtlc5n1494_15_CYSELF_2820 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z308,
      O => U_DCT2D_rtlc5n1494_15_CYSELF
    );
  U_DCT2D_rtlc5n1494_15_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_15_XORG,
      O => U_DCT2D_rtlc5n1494(16)
    );
  U_DCT2D_rtlc5n1494_15_XORG_2821 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_394_add_67_ix65206z63763_O,
      I1 => U_DCT2D_nx65206z305,
      O => U_DCT2D_rtlc5n1494_15_XORG
    );
  U_DCT2D_rtlc5n1494_15_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_15_CYMUXFAST,
      O => U_DCT2D_rtlc_394_add_67_ix65206z63760_O
    );
  U_DCT2D_rtlc5n1494_15_FASTCARRY_2822 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_394_add_67_ix65206z63767_O,
      O => U_DCT2D_rtlc5n1494_15_FASTCARRY
    );
  U_DCT2D_rtlc5n1494_15_CYAND_2823 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1494_15_CYSELG,
      I1 => U_DCT2D_rtlc5n1494_15_CYSELF,
      O => U_DCT2D_rtlc5n1494_15_CYAND
    );
  U_DCT2D_rtlc5n1494_15_CYMUXFAST_2824 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_15_CYMUXG2,
      IB => U_DCT2D_rtlc5n1494_15_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1494_15_CYAND,
      O => U_DCT2D_rtlc5n1494_15_CYMUXFAST
    );
  U_DCT2D_rtlc5n1494_15_CYMUXG2_2825 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_15_CY0G,
      IB => U_DCT2D_rtlc5n1494_15_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1494_15_CYSELG,
      O => U_DCT2D_rtlc5n1494_15_CYMUXG2
    );
  U_DCT2D_rtlc5n1494_15_CY0G_2826 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s(12),
      O => U_DCT2D_rtlc5n1494_15_CY0G
    );
  U_DCT2D_rtlc5n1494_15_CYSELG_2827 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z305,
      O => U_DCT2D_rtlc5n1494_15_CYSELG
    );
  U_DCT2D_rtlc5n1494_17_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_17_XORF,
      O => U_DCT2D_rtlc5n1494(17)
    );
  U_DCT2D_rtlc5n1494_17_XORF_2828 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1494_17_CYINIT,
      I1 => U_DCT2D_nx65206z302,
      O => U_DCT2D_rtlc5n1494_17_XORF
    );
  U_DCT2D_rtlc5n1494_17_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_17_CY0F,
      IB => U_DCT2D_rtlc5n1494_17_CYINIT,
      SEL => U_DCT2D_rtlc5n1494_17_CYSELF,
      O => U_DCT2D_rtlc_394_add_67_ix65206z63756_O
    );
  U_DCT2D_rtlc5n1494_17_CYMUXF2_2829 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_17_CY0F,
      IB => U_DCT2D_rtlc5n1494_17_CY0F,
      SEL => U_DCT2D_rtlc5n1494_17_CYSELF,
      O => U_DCT2D_rtlc5n1494_17_CYMUXF2
    );
  U_DCT2D_rtlc5n1494_17_CYINIT_2830 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_394_add_67_ix65206z63760_O,
      O => U_DCT2D_rtlc5n1494_17_CYINIT
    );
  U_DCT2D_rtlc5n1494_17_CY0F_2831 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s(13),
      O => U_DCT2D_rtlc5n1494_17_CY0F
    );
  U_DCT2D_rtlc5n1494_17_CYSELF_2832 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z302,
      O => U_DCT2D_rtlc5n1494_17_CYSELF
    );
  U_DCT2D_rtlc5n1494_17_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_17_XORG,
      O => U_DCT2D_rtlc5n1494(18)
    );
  U_DCT2D_rtlc5n1494_17_XORG_2833 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_394_add_67_ix65206z63756_O,
      I1 => U_DCT2D_nx65206z299,
      O => U_DCT2D_rtlc5n1494_17_XORG
    );
  U_DCT2D_rtlc5n1494_17_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_17_CYMUXFAST,
      O => U_DCT2D_rtlc_394_add_67_ix65206z63753_O
    );
  U_DCT2D_rtlc5n1494_17_FASTCARRY_2834 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_394_add_67_ix65206z63760_O,
      O => U_DCT2D_rtlc5n1494_17_FASTCARRY
    );
  U_DCT2D_rtlc5n1494_17_CYAND_2835 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1494_17_CYSELG,
      I1 => U_DCT2D_rtlc5n1494_17_CYSELF,
      O => U_DCT2D_rtlc5n1494_17_CYAND
    );
  U_DCT2D_rtlc5n1494_17_CYMUXFAST_2836 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_17_CYMUXG2,
      IB => U_DCT2D_rtlc5n1494_17_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1494_17_CYAND,
      O => U_DCT2D_rtlc5n1494_17_CYMUXFAST
    );
  U_DCT2D_rtlc5n1494_17_CYMUXG2_2837 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1494_17_CY0G,
      IB => U_DCT2D_rtlc5n1494_17_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1494_17_CYSELG,
      O => U_DCT2D_rtlc5n1494_17_CYMUXG2
    );
  U_DCT2D_rtlc5n1494_17_CY0G_2838 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s(13),
      O => U_DCT2D_rtlc5n1494_17_CY0G
    );
  U_DCT2D_rtlc5n1494_17_CYSELG_2839 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z299,
      O => U_DCT2D_rtlc5n1494_17_CYSELG
    );
  U_DCT2D_nx65206z297_rt_2840 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT2D_nx65206z297,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z297_rt
    );
  U_DCT2D_rtlc5n1494_19_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494_19_XORF,
      O => U_DCT2D_rtlc5n1494(19)
    );
  U_DCT2D_rtlc5n1494_19_XORF_2841 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1494_19_CYINIT,
      I1 => U_DCT2D_nx65206z297_rt,
      O => U_DCT2D_rtlc5n1494_19_XORF
    );
  U_DCT2D_rtlc5n1494_19_CYINIT_2842 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_394_add_67_ix65206z63753_O,
      O => U_DCT2D_rtlc5n1494_19_CYINIT
    );
  U_DCT2D_nx65206z570_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z570_XORF,
      O => U_DCT2D_nx65206z570
    );
  U_DCT2D_nx65206z570_XORF_2843 : X_XOR2
    port map (
      I0 => U_DCT2D_nx65206z570_CYINIT,
      I1 => U_DCT2D_nx65206z570_F,
      O => U_DCT2D_nx65206z570_XORF
    );
  U_DCT2D_nx65206z570_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z570_CY0F,
      IB => U_DCT2D_nx65206z570_CYINIT,
      SEL => U_DCT2D_nx65206z570_CYSELF,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63689_O
    );
  U_DCT2D_nx65206z570_CYINIT_2844 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z570_BXINVNOT,
      O => U_DCT2D_nx65206z570_CYINIT
    );
  U_DCT2D_nx65206z570_CY0F_2845 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z251,
      O => U_DCT2D_nx65206z570_CY0F
    );
  U_DCT2D_nx65206z570_CYSELF_2846 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z570_F,
      O => U_DCT2D_nx65206z570_CYSELF
    );
  U_DCT2D_nx65206z570_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_34,
      O => U_DCT2D_nx65206z570_BXINVNOT
    );
  U_DCT2D_nx65206z570_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z570_XORG,
      O => U_DCT2D_nx65206z567
    );
  U_DCT2D_nx65206z570_XORG_2847 : X_XOR2
    port map (
      I0 => U_DCT2D_ix959_modgen_add_291_ix65206z63689_O,
      I1 => U_DCT2D_nx65206z247,
      O => U_DCT2D_nx65206z570_XORG
    );
  U_DCT2D_nx65206z570_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z570_CYMUXG,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63683_O
    );
  U_DCT2D_nx65206z570_CYMUXG_2848 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z570_CY0G,
      IB => U_DCT2D_ix959_modgen_add_291_ix65206z63689_O,
      SEL => U_DCT2D_nx65206z570_CYSELG,
      O => U_DCT2D_nx65206z570_CYMUXG
    );
  U_DCT2D_nx65206z570_CY0G_2849 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z248,
      O => U_DCT2D_nx65206z570_CY0G
    );
  U_DCT2D_nx65206z570_CYSELG_2850 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z247,
      O => U_DCT2D_nx65206z570_CYSELG
    );
  U_DCT2D_nx65206z564_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z564_XORF,
      O => U_DCT2D_nx65206z564
    );
  U_DCT2D_nx65206z564_XORF_2851 : X_XOR2
    port map (
      I0 => U_DCT2D_nx65206z564_CYINIT,
      I1 => U_DCT2D_nx65206z244,
      O => U_DCT2D_nx65206z564_XORF
    );
  U_DCT2D_nx65206z564_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z564_CY0F,
      IB => U_DCT2D_nx65206z564_CYINIT,
      SEL => U_DCT2D_nx65206z564_CYSELF,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63677_O
    );
  U_DCT2D_nx65206z564_CYMUXF2_2852 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z564_CY0F,
      IB => U_DCT2D_nx65206z564_CY0F,
      SEL => U_DCT2D_nx65206z564_CYSELF,
      O => U_DCT2D_nx65206z564_CYMUXF2
    );
  U_DCT2D_nx65206z564_CYINIT_2853 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63683_O,
      O => U_DCT2D_nx65206z564_CYINIT
    );
  U_DCT2D_nx65206z564_CY0F_2854 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z245,
      O => U_DCT2D_nx65206z564_CY0F
    );
  U_DCT2D_nx65206z564_CYSELF_2855 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z244,
      O => U_DCT2D_nx65206z564_CYSELF
    );
  U_DCT2D_nx65206z564_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z564_XORG,
      O => U_DCT2D_nx65206z561
    );
  U_DCT2D_nx65206z564_XORG_2856 : X_XOR2
    port map (
      I0 => U_DCT2D_ix959_modgen_add_291_ix65206z63677_O,
      I1 => U_DCT2D_nx65206z241,
      O => U_DCT2D_nx65206z564_XORG
    );
  U_DCT2D_nx65206z564_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z564_CYMUXFAST,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63671_O
    );
  U_DCT2D_nx65206z564_FASTCARRY_2857 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63683_O,
      O => U_DCT2D_nx65206z564_FASTCARRY
    );
  U_DCT2D_nx65206z564_CYAND_2858 : X_AND2
    port map (
      I0 => U_DCT2D_nx65206z564_CYSELG,
      I1 => U_DCT2D_nx65206z564_CYSELF,
      O => U_DCT2D_nx65206z564_CYAND
    );
  U_DCT2D_nx65206z564_CYMUXFAST_2859 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z564_CYMUXG2,
      IB => U_DCT2D_nx65206z564_FASTCARRY,
      SEL => U_DCT2D_nx65206z564_CYAND,
      O => U_DCT2D_nx65206z564_CYMUXFAST
    );
  U_DCT2D_nx65206z564_CYMUXG2_2860 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z564_CY0G,
      IB => U_DCT2D_nx65206z564_CYMUXF2,
      SEL => U_DCT2D_nx65206z564_CYSELG,
      O => U_DCT2D_nx65206z564_CYMUXG2
    );
  U_DCT2D_nx65206z564_CY0G_2861 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z242,
      O => U_DCT2D_nx65206z564_CY0G
    );
  U_DCT2D_nx65206z564_CYSELG_2862 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z241,
      O => U_DCT2D_nx65206z564_CYSELG
    );
  U_DCT2D_nx65206z557_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z557_XORF,
      O => U_DCT2D_nx65206z557
    );
  U_DCT2D_nx65206z557_XORF_2863 : X_XOR2
    port map (
      I0 => U_DCT2D_nx65206z557_CYINIT,
      I1 => U_DCT2D_nx65206z238,
      O => U_DCT2D_nx65206z557_XORF
    );
  U_DCT2D_nx65206z557_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z557_CY0F,
      IB => U_DCT2D_nx65206z557_CYINIT,
      SEL => U_DCT2D_nx65206z557_CYSELF,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63665_O
    );
  U_DCT2D_nx65206z557_CYMUXF2_2864 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z557_CY0F,
      IB => U_DCT2D_nx65206z557_CY0F,
      SEL => U_DCT2D_nx65206z557_CYSELF,
      O => U_DCT2D_nx65206z557_CYMUXF2
    );
  U_DCT2D_nx65206z557_CYINIT_2865 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63671_O,
      O => U_DCT2D_nx65206z557_CYINIT
    );
  U_DCT2D_nx65206z557_CY0F_2866 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z239,
      O => U_DCT2D_nx65206z557_CY0F
    );
  U_DCT2D_nx65206z557_CYSELF_2867 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z238,
      O => U_DCT2D_nx65206z557_CYSELF
    );
  U_DCT2D_nx65206z557_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z557_XORG,
      O => U_DCT2D_nx65206z553
    );
  U_DCT2D_nx65206z557_XORG_2868 : X_XOR2
    port map (
      I0 => U_DCT2D_ix959_modgen_add_291_ix65206z63665_O,
      I1 => U_DCT2D_nx65206z235,
      O => U_DCT2D_nx65206z557_XORG
    );
  U_DCT2D_nx65206z557_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z557_CYMUXFAST,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63659_O
    );
  U_DCT2D_nx65206z557_FASTCARRY_2869 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63671_O,
      O => U_DCT2D_nx65206z557_FASTCARRY
    );
  U_DCT2D_nx65206z557_CYAND_2870 : X_AND2
    port map (
      I0 => U_DCT2D_nx65206z557_CYSELG,
      I1 => U_DCT2D_nx65206z557_CYSELF,
      O => U_DCT2D_nx65206z557_CYAND
    );
  U_DCT2D_nx65206z557_CYMUXFAST_2871 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z557_CYMUXG2,
      IB => U_DCT2D_nx65206z557_FASTCARRY,
      SEL => U_DCT2D_nx65206z557_CYAND,
      O => U_DCT2D_nx65206z557_CYMUXFAST
    );
  U_DCT2D_nx65206z557_CYMUXG2_2872 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z557_CY0G,
      IB => U_DCT2D_nx65206z557_CYMUXF2,
      SEL => U_DCT2D_nx65206z557_CYSELG,
      O => U_DCT2D_nx65206z557_CYMUXG2
    );
  U_DCT2D_nx65206z557_CY0G_2873 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z236,
      O => U_DCT2D_nx65206z557_CY0G
    );
  U_DCT2D_nx65206z557_CYSELG_2874 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z235,
      O => U_DCT2D_nx65206z557_CYSELG
    );
  U_DCT2D_nx65206z549_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z549_XORF,
      O => U_DCT2D_nx65206z549
    );
  U_DCT2D_nx65206z549_XORF_2875 : X_XOR2
    port map (
      I0 => U_DCT2D_nx65206z549_CYINIT,
      I1 => U_DCT2D_nx65206z232,
      O => U_DCT2D_nx65206z549_XORF
    );
  U_DCT2D_nx65206z549_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z549_CY0F,
      IB => U_DCT2D_nx65206z549_CYINIT,
      SEL => U_DCT2D_nx65206z549_CYSELF,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63653_O
    );
  U_DCT2D_nx65206z549_CYMUXF2_2876 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z549_CY0F,
      IB => U_DCT2D_nx65206z549_CY0F,
      SEL => U_DCT2D_nx65206z549_CYSELF,
      O => U_DCT2D_nx65206z549_CYMUXF2
    );
  U_DCT2D_nx65206z549_CYINIT_2877 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63659_O,
      O => U_DCT2D_nx65206z549_CYINIT
    );
  U_DCT2D_nx65206z549_CY0F_2878 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z233,
      O => U_DCT2D_nx65206z549_CY0F
    );
  U_DCT2D_nx65206z549_CYSELF_2879 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z232,
      O => U_DCT2D_nx65206z549_CYSELF
    );
  U_DCT2D_nx65206z549_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z549_XORG,
      O => U_DCT2D_nx65206z545
    );
  U_DCT2D_nx65206z549_XORG_2880 : X_XOR2
    port map (
      I0 => U_DCT2D_ix959_modgen_add_291_ix65206z63653_O,
      I1 => U_DCT2D_nx65206z229,
      O => U_DCT2D_nx65206z549_XORG
    );
  U_DCT2D_nx65206z549_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z549_CYMUXFAST,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63647_O
    );
  U_DCT2D_nx65206z549_FASTCARRY_2881 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63659_O,
      O => U_DCT2D_nx65206z549_FASTCARRY
    );
  U_DCT2D_nx65206z549_CYAND_2882 : X_AND2
    port map (
      I0 => U_DCT2D_nx65206z549_CYSELG,
      I1 => U_DCT2D_nx65206z549_CYSELF,
      O => U_DCT2D_nx65206z549_CYAND
    );
  U_DCT2D_nx65206z549_CYMUXFAST_2883 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z549_CYMUXG2,
      IB => U_DCT2D_nx65206z549_FASTCARRY,
      SEL => U_DCT2D_nx65206z549_CYAND,
      O => U_DCT2D_nx65206z549_CYMUXFAST
    );
  U_DCT2D_nx65206z549_CYMUXG2_2884 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z549_CY0G,
      IB => U_DCT2D_nx65206z549_CYMUXF2,
      SEL => U_DCT2D_nx65206z549_CYSELG,
      O => U_DCT2D_nx65206z549_CYMUXG2
    );
  U_DCT2D_nx65206z549_CY0G_2885 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z230,
      O => U_DCT2D_nx65206z549_CY0G
    );
  U_DCT2D_nx65206z549_CYSELG_2886 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z229,
      O => U_DCT2D_nx65206z549_CYSELG
    );
  U_DCT2D_nx65206z541_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z541_XORF,
      O => U_DCT2D_nx65206z541
    );
  U_DCT2D_nx65206z541_XORF_2887 : X_XOR2
    port map (
      I0 => U_DCT2D_nx65206z541_CYINIT,
      I1 => U_DCT2D_nx65206z226,
      O => U_DCT2D_nx65206z541_XORF
    );
  U_DCT2D_nx65206z541_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z541_CY0F,
      IB => U_DCT2D_nx65206z541_CYINIT,
      SEL => U_DCT2D_nx65206z541_CYSELF,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63641_O
    );
  U_DCT2D_nx65206z541_CYMUXF2_2888 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z541_CY0F,
      IB => U_DCT2D_nx65206z541_CY0F,
      SEL => U_DCT2D_nx65206z541_CYSELF,
      O => U_DCT2D_nx65206z541_CYMUXF2
    );
  U_DCT2D_nx65206z541_CYINIT_2889 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63647_O,
      O => U_DCT2D_nx65206z541_CYINIT
    );
  U_DCT2D_nx65206z541_CY0F_2890 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z227,
      O => U_DCT2D_nx65206z541_CY0F
    );
  U_DCT2D_nx65206z541_CYSELF_2891 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z226,
      O => U_DCT2D_nx65206z541_CYSELF
    );
  U_DCT2D_nx65206z541_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z541_XORG,
      O => U_DCT2D_nx65206z537
    );
  U_DCT2D_nx65206z541_XORG_2892 : X_XOR2
    port map (
      I0 => U_DCT2D_ix959_modgen_add_291_ix65206z63641_O,
      I1 => U_DCT2D_nx65206z223,
      O => U_DCT2D_nx65206z541_XORG
    );
  U_DCT2D_nx65206z541_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z541_CYMUXFAST,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63635_O
    );
  U_DCT2D_nx65206z541_FASTCARRY_2893 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63647_O,
      O => U_DCT2D_nx65206z541_FASTCARRY
    );
  U_DCT2D_nx65206z541_CYAND_2894 : X_AND2
    port map (
      I0 => U_DCT2D_nx65206z541_CYSELG,
      I1 => U_DCT2D_nx65206z541_CYSELF,
      O => U_DCT2D_nx65206z541_CYAND
    );
  U_DCT2D_nx65206z541_CYMUXFAST_2895 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z541_CYMUXG2,
      IB => U_DCT2D_nx65206z541_FASTCARRY,
      SEL => U_DCT2D_nx65206z541_CYAND,
      O => U_DCT2D_nx65206z541_CYMUXFAST
    );
  U_DCT2D_nx65206z541_CYMUXG2_2896 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z541_CY0G,
      IB => U_DCT2D_nx65206z541_CYMUXF2,
      SEL => U_DCT2D_nx65206z541_CYSELG,
      O => U_DCT2D_nx65206z541_CYMUXG2
    );
  U_DCT2D_nx65206z541_CY0G_2897 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z224,
      O => U_DCT2D_nx65206z541_CY0G
    );
  U_DCT2D_nx65206z541_CYSELG_2898 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z223,
      O => U_DCT2D_nx65206z541_CYSELG
    );
  U_DCT2D_nx65206z533_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z533_XORF,
      O => U_DCT2D_nx65206z533
    );
  U_DCT2D_nx65206z533_XORF_2899 : X_XOR2
    port map (
      I0 => U_DCT2D_nx65206z533_CYINIT,
      I1 => U_DCT2D_nx65206z220,
      O => U_DCT2D_nx65206z533_XORF
    );
  U_DCT2D_nx65206z533_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z533_CY0F,
      IB => U_DCT2D_nx65206z533_CYINIT,
      SEL => U_DCT2D_nx65206z533_CYSELF,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63629_O
    );
  U_DCT2D_nx65206z533_CYMUXF2_2900 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z533_CY0F,
      IB => U_DCT2D_nx65206z533_CY0F,
      SEL => U_DCT2D_nx65206z533_CYSELF,
      O => U_DCT2D_nx65206z533_CYMUXF2
    );
  U_DCT2D_nx65206z533_CYINIT_2901 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63635_O,
      O => U_DCT2D_nx65206z533_CYINIT
    );
  U_DCT2D_nx65206z533_CY0F_2902 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z221,
      O => U_DCT2D_nx65206z533_CY0F
    );
  U_DCT2D_nx65206z533_CYSELF_2903 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z220,
      O => U_DCT2D_nx65206z533_CYSELF
    );
  U_DCT2D_nx65206z533_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z533_XORG,
      O => U_DCT2D_nx65206z529
    );
  U_DCT2D_nx65206z533_XORG_2904 : X_XOR2
    port map (
      I0 => U_DCT2D_ix959_modgen_add_291_ix65206z63629_O,
      I1 => U_DCT2D_nx65206z217,
      O => U_DCT2D_nx65206z533_XORG
    );
  U_DCT2D_nx65206z533_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z533_CYMUXFAST,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63624_O
    );
  U_DCT2D_nx65206z533_FASTCARRY_2905 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63635_O,
      O => U_DCT2D_nx65206z533_FASTCARRY
    );
  U_DCT2D_nx65206z533_CYAND_2906 : X_AND2
    port map (
      I0 => U_DCT2D_nx65206z533_CYSELG,
      I1 => U_DCT2D_nx65206z533_CYSELF,
      O => U_DCT2D_nx65206z533_CYAND
    );
  U_DCT2D_nx65206z533_CYMUXFAST_2907 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z533_CYMUXG2,
      IB => U_DCT2D_nx65206z533_FASTCARRY,
      SEL => U_DCT2D_nx65206z533_CYAND,
      O => U_DCT2D_nx65206z533_CYMUXFAST
    );
  U_DCT2D_nx65206z533_CYMUXG2_2908 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z533_CY0G,
      IB => U_DCT2D_nx65206z533_CYMUXF2,
      SEL => U_DCT2D_nx65206z533_CYSELG,
      O => U_DCT2D_nx65206z533_CYMUXG2
    );
  U_DCT2D_nx65206z533_CY0G_2909 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z218,
      O => U_DCT2D_nx65206z533_CY0G
    );
  U_DCT2D_nx65206z533_CYSELG_2910 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z217,
      O => U_DCT2D_nx65206z533_CYSELG
    );
  U_DCT2D_nx65206z525_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z525_XORF,
      O => U_DCT2D_nx65206z525
    );
  U_DCT2D_nx65206z525_XORF_2911 : X_XOR2
    port map (
      I0 => U_DCT2D_nx65206z525_CYINIT,
      I1 => U_DCT2D_nx65206z214,
      O => U_DCT2D_nx65206z525_XORF
    );
  U_DCT2D_nx65206z525_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z525_CY0F,
      IB => U_DCT2D_nx65206z525_CYINIT,
      SEL => U_DCT2D_nx65206z525_CYSELF,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63619_O
    );
  U_DCT2D_nx65206z525_CYMUXF2_2912 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z525_CY0F,
      IB => U_DCT2D_nx65206z525_CY0F,
      SEL => U_DCT2D_nx65206z525_CYSELF,
      O => U_DCT2D_nx65206z525_CYMUXF2
    );
  U_DCT2D_nx65206z525_CYINIT_2913 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63624_O,
      O => U_DCT2D_nx65206z525_CYINIT
    );
  U_DCT2D_nx65206z525_CY0F_2914 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z215,
      O => U_DCT2D_nx65206z525_CY0F
    );
  U_DCT2D_nx65206z525_CYSELF_2915 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z214,
      O => U_DCT2D_nx65206z525_CYSELF
    );
  U_DCT2D_nx65206z525_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z525_XORG,
      O => U_DCT2D_nx65206z521
    );
  U_DCT2D_nx65206z525_XORG_2916 : X_XOR2
    port map (
      I0 => U_DCT2D_ix959_modgen_add_291_ix65206z63619_O,
      I1 => U_DCT2D_nx65206z211,
      O => U_DCT2D_nx65206z525_XORG
    );
  U_DCT2D_nx65206z525_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z525_CYMUXFAST,
      O => U_DCT2D_ix959_modgen_add_291_ix65206z63615_O
    );
  U_DCT2D_nx65206z525_FASTCARRY_2917 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63624_O,
      O => U_DCT2D_nx65206z525_FASTCARRY
    );
  U_DCT2D_nx65206z525_CYAND_2918 : X_AND2
    port map (
      I0 => U_DCT2D_nx65206z525_CYSELG,
      I1 => U_DCT2D_nx65206z525_CYSELF,
      O => U_DCT2D_nx65206z525_CYAND
    );
  U_DCT2D_nx65206z525_CYMUXFAST_2919 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z525_CYMUXG2,
      IB => U_DCT2D_nx65206z525_FASTCARRY,
      SEL => U_DCT2D_nx65206z525_CYAND,
      O => U_DCT2D_nx65206z525_CYMUXFAST
    );
  U_DCT2D_nx65206z525_CYMUXG2_2920 : X_MUX2
    port map (
      IA => U_DCT2D_nx65206z525_CY0G,
      IB => U_DCT2D_nx65206z525_CYMUXF2,
      SEL => U_DCT2D_nx65206z525_CYSELG,
      O => U_DCT2D_nx65206z525_CYMUXG2
    );
  U_DCT2D_nx65206z525_CY0G_2921 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z212,
      O => U_DCT2D_nx65206z525_CY0G
    );
  U_DCT2D_nx65206z525_CYSELG_2922 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z211,
      O => U_DCT2D_nx65206z525_CYSELG
    );
  U_DCT2D_nx65206z3_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z3_XORF,
      O => U_DCT2D_nx65206z3
    );
  U_DCT2D_nx65206z3_XORF_2923 : X_XOR2
    port map (
      I0 => U_DCT2D_nx65206z3_CYINIT,
      I1 => U_DCT2D_nx65206z4_rt,
      O => U_DCT2D_nx65206z3_XORF
    );
  U_DCT2D_nx65206z3_CYINIT_2924 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_ix959_modgen_add_291_ix65206z63615_O,
      O => U_DCT2D_nx65206z3_CYINIT
    );
  U_DCT1D_rtlc5n1344_2_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_2_CY0F,
      IB => U_DCT1D_rtlc5n1344_2_CYINIT,
      SEL => U_DCT1D_rtlc5n1344_2_CYSELF,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63485_O
    );
  U_DCT1D_rtlc5n1344_2_CYINIT_2925 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_2_BXINVNOT,
      O => U_DCT1D_rtlc5n1344_2_CYINIT
    );
  U_DCT1D_rtlc5n1344_2_CY0F_2926 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(1),
      O => U_DCT1D_rtlc5n1344_2_CY0F
    );
  U_DCT1D_rtlc5n1344_2_CYSELF_2927 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z120,
      O => U_DCT1D_rtlc5n1344_2_CYSELF
    );
  U_DCT1D_rtlc5n1344_2_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_0,
      O => U_DCT1D_rtlc5n1344_2_BXINVNOT
    );
  U_DCT1D_rtlc5n1344_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_2_XORG,
      O => U_DCT1D_rtlc5n1344(2)
    );
  U_DCT1D_rtlc5n1344_2_XORG_2928 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_491_add_20_ix59700z63485_O,
      I1 => U_DCT1D_nx59700z117,
      O => U_DCT1D_rtlc5n1344_2_XORG
    );
  U_DCT1D_rtlc5n1344_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_2_CYMUXG,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63482_O
    );
  U_DCT1D_rtlc5n1344_2_CYMUXG_2929 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_2_CY0G,
      IB => U_DCT1D_rtlc_491_add_20_ix59700z63485_O,
      SEL => U_DCT1D_rtlc5n1344_2_CYSELG,
      O => U_DCT1D_rtlc5n1344_2_CYMUXG
    );
  U_DCT1D_rtlc5n1344_2_CY0G_2930 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(2),
      O => U_DCT1D_rtlc5n1344_2_CY0G
    );
  U_DCT1D_rtlc5n1344_2_CYSELG_2931 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z117,
      O => U_DCT1D_rtlc5n1344_2_CYSELG
    );
  U_DCT1D_rtlc5n1344_3_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_3_XORF,
      O => U_DCT1D_rtlc5n1344(3)
    );
  U_DCT1D_rtlc5n1344_3_XORF_2932 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1344_3_CYINIT,
      I1 => U_DCT1D_nx59700z114,
      O => U_DCT1D_rtlc5n1344_3_XORF
    );
  U_DCT1D_rtlc5n1344_3_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_3_CY0F,
      IB => U_DCT1D_rtlc5n1344_3_CYINIT,
      SEL => U_DCT1D_rtlc5n1344_3_CYSELF,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63478_O
    );
  U_DCT1D_rtlc5n1344_3_CYMUXF2_2933 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_3_CY0F,
      IB => U_DCT1D_rtlc5n1344_3_CY0F,
      SEL => U_DCT1D_rtlc5n1344_3_CYSELF,
      O => U_DCT1D_rtlc5n1344_3_CYMUXF2
    );
  U_DCT1D_rtlc5n1344_3_CYINIT_2934 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63482_O,
      O => U_DCT1D_rtlc5n1344_3_CYINIT
    );
  U_DCT1D_rtlc5n1344_3_CY0F_2935 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(3),
      O => U_DCT1D_rtlc5n1344_3_CY0F
    );
  U_DCT1D_rtlc5n1344_3_CYSELF_2936 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z114,
      O => U_DCT1D_rtlc5n1344_3_CYSELF
    );
  U_DCT1D_rtlc5n1344_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_3_XORG,
      O => U_DCT1D_rtlc5n1344(4)
    );
  U_DCT1D_rtlc5n1344_3_XORG_2937 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_491_add_20_ix59700z63478_O,
      I1 => U_DCT1D_nx59700z111,
      O => U_DCT1D_rtlc5n1344_3_XORG
    );
  U_DCT1D_rtlc5n1344_3_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_3_CYMUXFAST,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63474_O
    );
  U_DCT1D_rtlc5n1344_3_FASTCARRY_2938 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63482_O,
      O => U_DCT1D_rtlc5n1344_3_FASTCARRY
    );
  U_DCT1D_rtlc5n1344_3_CYAND_2939 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1344_3_CYSELG,
      I1 => U_DCT1D_rtlc5n1344_3_CYSELF,
      O => U_DCT1D_rtlc5n1344_3_CYAND
    );
  U_DCT1D_rtlc5n1344_3_CYMUXFAST_2940 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_3_CYMUXG2,
      IB => U_DCT1D_rtlc5n1344_3_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1344_3_CYAND,
      O => U_DCT1D_rtlc5n1344_3_CYMUXFAST
    );
  U_DCT1D_rtlc5n1344_3_CYMUXG2_2941 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_3_CY0G,
      IB => U_DCT1D_rtlc5n1344_3_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1344_3_CYSELG,
      O => U_DCT1D_rtlc5n1344_3_CYMUXG2
    );
  U_DCT1D_rtlc5n1344_3_CY0G_2942 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(4),
      O => U_DCT1D_rtlc5n1344_3_CY0G
    );
  U_DCT1D_rtlc5n1344_3_CYSELG_2943 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z111,
      O => U_DCT1D_rtlc5n1344_3_CYSELG
    );
  U_DCT1D_rtlc5n1344_5_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_5_XORF,
      O => U_DCT1D_rtlc5n1344(5)
    );
  U_DCT1D_rtlc5n1344_5_XORF_2944 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1344_5_CYINIT,
      I1 => U_DCT1D_nx59700z108,
      O => U_DCT1D_rtlc5n1344_5_XORF
    );
  U_DCT1D_rtlc5n1344_5_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_5_CY0F,
      IB => U_DCT1D_rtlc5n1344_5_CYINIT,
      SEL => U_DCT1D_rtlc5n1344_5_CYSELF,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63471_O
    );
  U_DCT1D_rtlc5n1344_5_CYMUXF2_2945 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_5_CY0F,
      IB => U_DCT1D_rtlc5n1344_5_CY0F,
      SEL => U_DCT1D_rtlc5n1344_5_CYSELF,
      O => U_DCT1D_rtlc5n1344_5_CYMUXF2
    );
  U_DCT1D_rtlc5n1344_5_CYINIT_2946 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63474_O,
      O => U_DCT1D_rtlc5n1344_5_CYINIT
    );
  U_DCT1D_rtlc5n1344_5_CY0F_2947 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(5),
      O => U_DCT1D_rtlc5n1344_5_CY0F
    );
  U_DCT1D_rtlc5n1344_5_CYSELF_2948 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z108,
      O => U_DCT1D_rtlc5n1344_5_CYSELF
    );
  U_DCT1D_rtlc5n1344_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_5_XORG,
      O => U_DCT1D_rtlc5n1344(6)
    );
  U_DCT1D_rtlc5n1344_5_XORG_2949 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_491_add_20_ix59700z63471_O,
      I1 => U_DCT1D_nx59700z105,
      O => U_DCT1D_rtlc5n1344_5_XORG
    );
  U_DCT1D_rtlc5n1344_5_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_5_CYMUXFAST,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63467_O
    );
  U_DCT1D_rtlc5n1344_5_FASTCARRY_2950 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63474_O,
      O => U_DCT1D_rtlc5n1344_5_FASTCARRY
    );
  U_DCT1D_rtlc5n1344_5_CYAND_2951 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1344_5_CYSELG,
      I1 => U_DCT1D_rtlc5n1344_5_CYSELF,
      O => U_DCT1D_rtlc5n1344_5_CYAND
    );
  U_DCT1D_rtlc5n1344_5_CYMUXFAST_2952 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_5_CYMUXG2,
      IB => U_DCT1D_rtlc5n1344_5_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1344_5_CYAND,
      O => U_DCT1D_rtlc5n1344_5_CYMUXFAST
    );
  U_DCT1D_rtlc5n1344_5_CYMUXG2_2953 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_5_CY0G,
      IB => U_DCT1D_rtlc5n1344_5_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1344_5_CYSELG,
      O => U_DCT1D_rtlc5n1344_5_CYMUXG2
    );
  U_DCT1D_rtlc5n1344_5_CY0G_2954 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(6),
      O => U_DCT1D_rtlc5n1344_5_CY0G
    );
  U_DCT1D_rtlc5n1344_5_CYSELG_2955 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z105,
      O => U_DCT1D_rtlc5n1344_5_CYSELG
    );
  U_DCT1D_rtlc5n1344_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_7_XORF,
      O => U_DCT1D_rtlc5n1344(7)
    );
  U_DCT1D_rtlc5n1344_7_XORF_2956 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1344_7_CYINIT,
      I1 => U_DCT1D_nx59700z102,
      O => U_DCT1D_rtlc5n1344_7_XORF
    );
  U_DCT1D_rtlc5n1344_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_7_CY0F,
      IB => U_DCT1D_rtlc5n1344_7_CYINIT,
      SEL => U_DCT1D_rtlc5n1344_7_CYSELF,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63463_O
    );
  U_DCT1D_rtlc5n1344_7_CYMUXF2_2957 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_7_CY0F,
      IB => U_DCT1D_rtlc5n1344_7_CY0F,
      SEL => U_DCT1D_rtlc5n1344_7_CYSELF,
      O => U_DCT1D_rtlc5n1344_7_CYMUXF2
    );
  U_DCT1D_rtlc5n1344_7_CYINIT_2958 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63467_O,
      O => U_DCT1D_rtlc5n1344_7_CYINIT
    );
  U_DCT1D_rtlc5n1344_7_CY0F_2959 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(7),
      O => U_DCT1D_rtlc5n1344_7_CY0F
    );
  U_DCT1D_rtlc5n1344_7_CYSELF_2960 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z102,
      O => U_DCT1D_rtlc5n1344_7_CYSELF
    );
  U_DCT1D_rtlc5n1344_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_7_XORG,
      O => U_DCT1D_rtlc5n1344(8)
    );
  U_DCT1D_rtlc5n1344_7_XORG_2961 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_491_add_20_ix59700z63463_O,
      I1 => U_DCT1D_nx59700z99,
      O => U_DCT1D_rtlc5n1344_7_XORG
    );
  U_DCT1D_rtlc5n1344_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_7_CYMUXFAST,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63460_O
    );
  U_DCT1D_rtlc5n1344_7_FASTCARRY_2962 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63467_O,
      O => U_DCT1D_rtlc5n1344_7_FASTCARRY
    );
  U_DCT1D_rtlc5n1344_7_CYAND_2963 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1344_7_CYSELG,
      I1 => U_DCT1D_rtlc5n1344_7_CYSELF,
      O => U_DCT1D_rtlc5n1344_7_CYAND
    );
  U_DCT1D_rtlc5n1344_7_CYMUXFAST_2964 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_7_CYMUXG2,
      IB => U_DCT1D_rtlc5n1344_7_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1344_7_CYAND,
      O => U_DCT1D_rtlc5n1344_7_CYMUXFAST
    );
  U_DCT1D_rtlc5n1344_7_CYMUXG2_2965 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_7_CY0G,
      IB => U_DCT1D_rtlc5n1344_7_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1344_7_CYSELG,
      O => U_DCT1D_rtlc5n1344_7_CYMUXG2
    );
  U_DCT1D_rtlc5n1344_7_CY0G_2966 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(8),
      O => U_DCT1D_rtlc5n1344_7_CY0G
    );
  U_DCT1D_rtlc5n1344_7_CYSELG_2967 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z99,
      O => U_DCT1D_rtlc5n1344_7_CYSELG
    );
  U_DCT1D_rtlc5n1344_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_9_XORF,
      O => U_DCT1D_rtlc5n1344(9)
    );
  U_DCT1D_rtlc5n1344_9_XORF_2968 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1344_9_CYINIT,
      I1 => U_DCT1D_nx59700z96,
      O => U_DCT1D_rtlc5n1344_9_XORF
    );
  U_DCT1D_rtlc5n1344_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_9_CY0F,
      IB => U_DCT1D_rtlc5n1344_9_CYINIT,
      SEL => U_DCT1D_rtlc5n1344_9_CYSELF,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63456_O
    );
  U_DCT1D_rtlc5n1344_9_CYMUXF2_2969 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_9_CY0F,
      IB => U_DCT1D_rtlc5n1344_9_CY0F,
      SEL => U_DCT1D_rtlc5n1344_9_CYSELF,
      O => U_DCT1D_rtlc5n1344_9_CYMUXF2
    );
  U_DCT1D_rtlc5n1344_9_CYINIT_2970 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63460_O,
      O => U_DCT1D_rtlc5n1344_9_CYINIT
    );
  U_DCT1D_rtlc5n1344_9_CY0F_2971 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(9),
      O => U_DCT1D_rtlc5n1344_9_CY0F
    );
  U_DCT1D_rtlc5n1344_9_CYSELF_2972 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z96,
      O => U_DCT1D_rtlc5n1344_9_CYSELF
    );
  U_DCT1D_rtlc5n1344_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_9_XORG,
      O => U_DCT1D_rtlc5n1344(10)
    );
  U_DCT1D_rtlc5n1344_9_XORG_2973 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_491_add_20_ix59700z63456_O,
      I1 => U_DCT1D_nx59700z93,
      O => U_DCT1D_rtlc5n1344_9_XORG
    );
  U_DCT1D_rtlc5n1344_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_9_CYMUXFAST,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63453_O
    );
  U_DCT1D_rtlc5n1344_9_FASTCARRY_2974 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63460_O,
      O => U_DCT1D_rtlc5n1344_9_FASTCARRY
    );
  U_DCT1D_rtlc5n1344_9_CYAND_2975 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1344_9_CYSELG,
      I1 => U_DCT1D_rtlc5n1344_9_CYSELF,
      O => U_DCT1D_rtlc5n1344_9_CYAND
    );
  U_DCT1D_rtlc5n1344_9_CYMUXFAST_2976 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_9_CYMUXG2,
      IB => U_DCT1D_rtlc5n1344_9_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1344_9_CYAND,
      O => U_DCT1D_rtlc5n1344_9_CYMUXFAST
    );
  U_DCT1D_rtlc5n1344_9_CYMUXG2_2977 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_9_CY0G,
      IB => U_DCT1D_rtlc5n1344_9_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1344_9_CYSELG,
      O => U_DCT1D_rtlc5n1344_9_CYMUXG2
    );
  U_DCT1D_rtlc5n1344_9_CY0G_2978 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(10),
      O => U_DCT1D_rtlc5n1344_9_CY0G
    );
  U_DCT1D_rtlc5n1344_9_CYSELG_2979 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z93,
      O => U_DCT1D_rtlc5n1344_9_CYSELG
    );
  U_DCT1D_rtlc5n1344_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_11_XORF,
      O => U_DCT1D_rtlc5n1344(11)
    );
  U_DCT1D_rtlc5n1344_11_XORF_2980 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1344_11_CYINIT,
      I1 => U_DCT1D_nx59700z90,
      O => U_DCT1D_rtlc5n1344_11_XORF
    );
  U_DCT1D_rtlc5n1344_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_11_CY0F,
      IB => U_DCT1D_rtlc5n1344_11_CYINIT,
      SEL => U_DCT1D_rtlc5n1344_11_CYSELF,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63449_O
    );
  U_DCT1D_rtlc5n1344_11_CYMUXF2_2981 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_11_CY0F,
      IB => U_DCT1D_rtlc5n1344_11_CY0F,
      SEL => U_DCT1D_rtlc5n1344_11_CYSELF,
      O => U_DCT1D_rtlc5n1344_11_CYMUXF2
    );
  U_DCT1D_rtlc5n1344_11_CYINIT_2982 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63453_O,
      O => U_DCT1D_rtlc5n1344_11_CYINIT
    );
  U_DCT1D_rtlc5n1344_11_CY0F_2983 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(11),
      O => U_DCT1D_rtlc5n1344_11_CY0F
    );
  U_DCT1D_rtlc5n1344_11_CYSELF_2984 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z90,
      O => U_DCT1D_rtlc5n1344_11_CYSELF
    );
  U_DCT1D_rtlc5n1344_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_11_XORG,
      O => U_DCT1D_rtlc5n1344(12)
    );
  U_DCT1D_rtlc5n1344_11_XORG_2985 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_491_add_20_ix59700z63449_O,
      I1 => U_DCT1D_nx59700z87,
      O => U_DCT1D_rtlc5n1344_11_XORG
    );
  U_DCT1D_rtlc5n1344_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_11_CYMUXFAST,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63446_O
    );
  U_DCT1D_rtlc5n1344_11_FASTCARRY_2986 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63453_O,
      O => U_DCT1D_rtlc5n1344_11_FASTCARRY
    );
  U_DCT1D_rtlc5n1344_11_CYAND_2987 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1344_11_CYSELG,
      I1 => U_DCT1D_rtlc5n1344_11_CYSELF,
      O => U_DCT1D_rtlc5n1344_11_CYAND
    );
  U_DCT1D_rtlc5n1344_11_CYMUXFAST_2988 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_11_CYMUXG2,
      IB => U_DCT1D_rtlc5n1344_11_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1344_11_CYAND,
      O => U_DCT1D_rtlc5n1344_11_CYMUXFAST
    );
  U_DCT1D_rtlc5n1344_11_CYMUXG2_2989 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_11_CY0G,
      IB => U_DCT1D_rtlc5n1344_11_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1344_11_CYSELG,
      O => U_DCT1D_rtlc5n1344_11_CYMUXG2
    );
  U_DCT1D_rtlc5n1344_11_CY0G_2990 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(12),
      O => U_DCT1D_rtlc5n1344_11_CY0G
    );
  U_DCT1D_rtlc5n1344_11_CYSELG_2991 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z87,
      O => U_DCT1D_rtlc5n1344_11_CYSELG
    );
  U_DCT1D_rtlc5n1344_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_13_XORF,
      O => U_DCT1D_rtlc5n1344(13)
    );
  U_DCT1D_rtlc5n1344_13_XORF_2992 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1344_13_CYINIT,
      I1 => U_DCT1D_nx59700z84,
      O => U_DCT1D_rtlc5n1344_13_XORF
    );
  U_DCT1D_rtlc5n1344_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_13_CY0F,
      IB => U_DCT1D_rtlc5n1344_13_CYINIT,
      SEL => U_DCT1D_rtlc5n1344_13_CYSELF,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63442_O
    );
  U_DCT1D_rtlc5n1344_13_CYMUXF2_2993 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_13_CY0F,
      IB => U_DCT1D_rtlc5n1344_13_CY0F,
      SEL => U_DCT1D_rtlc5n1344_13_CYSELF,
      O => U_DCT1D_rtlc5n1344_13_CYMUXF2
    );
  U_DCT1D_rtlc5n1344_13_CYINIT_2994 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63446_O,
      O => U_DCT1D_rtlc5n1344_13_CYINIT
    );
  U_DCT1D_rtlc5n1344_13_CY0F_2995 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(13),
      O => U_DCT1D_rtlc5n1344_13_CY0F
    );
  U_DCT1D_rtlc5n1344_13_CYSELF_2996 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z84,
      O => U_DCT1D_rtlc5n1344_13_CYSELF
    );
  U_DCT1D_rtlc5n1344_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_13_XORG,
      O => U_DCT1D_rtlc5n1344(14)
    );
  U_DCT1D_rtlc5n1344_13_XORG_2997 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_491_add_20_ix59700z63442_O,
      I1 => U_DCT1D_nx59700z81,
      O => U_DCT1D_rtlc5n1344_13_XORG
    );
  U_DCT1D_rtlc5n1344_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_13_CYMUXFAST,
      O => U_DCT1D_rtlc_491_add_20_ix59700z63439_O
    );
  U_DCT1D_rtlc5n1344_13_FASTCARRY_2998 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63446_O,
      O => U_DCT1D_rtlc5n1344_13_FASTCARRY
    );
  U_DCT1D_rtlc5n1344_13_CYAND_2999 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1344_13_CYSELG,
      I1 => U_DCT1D_rtlc5n1344_13_CYSELF,
      O => U_DCT1D_rtlc5n1344_13_CYAND
    );
  U_DCT1D_rtlc5n1344_13_CYMUXFAST_3000 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_13_CYMUXG2,
      IB => U_DCT1D_rtlc5n1344_13_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1344_13_CYAND,
      O => U_DCT1D_rtlc5n1344_13_CYMUXFAST
    );
  U_DCT1D_rtlc5n1344_13_CYMUXG2_3001 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1344_13_CY0G,
      IB => U_DCT1D_rtlc5n1344_13_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1344_13_CYSELG,
      O => U_DCT1D_rtlc5n1344_13_CYMUXG2
    );
  U_DCT1D_rtlc5n1344_13_CY0G_3002 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s(13),
      O => U_DCT1D_rtlc5n1344_13_CY0G
    );
  U_DCT1D_rtlc5n1344_13_CYSELG_3003 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z81,
      O => U_DCT1D_rtlc5n1344_13_CYSELG
    );
  U_DCT1D_nx59700z79_rt_3004 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z79,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z79_rt
    );
  U_DCT1D_rtlc5n1344_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344_15_XORF,
      O => U_DCT1D_rtlc5n1344(15)
    );
  U_DCT1D_rtlc5n1344_15_XORF_3005 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1344_15_CYINIT,
      I1 => U_DCT1D_nx59700z79_rt,
      O => U_DCT1D_rtlc5n1344_15_XORF
    );
  U_DCT1D_rtlc5n1344_15_CYINIT_3006 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_491_add_20_ix59700z63439_O,
      O => U_DCT1D_rtlc5n1344_15_CYINIT
    );
  U_DCT2D_rtlc5n1481_3_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_3_XORF,
      O => U_DCT2D_rtlc5n1481(3)
    );
  U_DCT2D_rtlc5n1481_3_XORF_3007 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1481_3_CYINIT,
      I1 => U_DCT2D_nx65206z162,
      O => U_DCT2D_rtlc5n1481_3_XORF
    );
  U_DCT2D_rtlc5n1481_3_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_3_CY0F,
      IB => U_DCT2D_rtlc5n1481_3_CYINIT,
      SEL => U_DCT2D_rtlc5n1481_3_CYSELF,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63535_O
    );
  U_DCT2D_rtlc5n1481_3_CYINIT_3008 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_3_BXINVNOT,
      O => U_DCT2D_rtlc5n1481_3_CYINIT
    );
  U_DCT2D_rtlc5n1481_3_CY0F_3009 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(1),
      O => U_DCT2D_rtlc5n1481_3_CY0F
    );
  U_DCT2D_rtlc5n1481_3_CYSELF_3010 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z162,
      O => U_DCT2D_rtlc5n1481_3_CYSELF
    );
  U_DCT2D_rtlc5n1481_3_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_30,
      O => U_DCT2D_rtlc5n1481_3_BXINVNOT
    );
  U_DCT2D_rtlc5n1481_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_3_XORG,
      O => U_DCT2D_rtlc5n1481(4)
    );
  U_DCT2D_rtlc5n1481_3_XORG_3011 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_333_add_55_ix65206z63535_O,
      I1 => U_DCT2D_nx65206z159,
      O => U_DCT2D_rtlc5n1481_3_XORG
    );
  U_DCT2D_rtlc5n1481_3_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_3_CYMUXG,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63531_O
    );
  U_DCT2D_rtlc5n1481_3_CYMUXG_3012 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_3_CY0G,
      IB => U_DCT2D_rtlc_333_add_55_ix65206z63535_O,
      SEL => U_DCT2D_rtlc5n1481_3_CYSELG,
      O => U_DCT2D_rtlc5n1481_3_CYMUXG
    );
  U_DCT2D_rtlc5n1481_3_CY0G_3013 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(2),
      O => U_DCT2D_rtlc5n1481_3_CY0G
    );
  U_DCT2D_rtlc5n1481_3_CYSELG_3014 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z159,
      O => U_DCT2D_rtlc5n1481_3_CYSELG
    );
  U_DCT1D_reg_databuf_reg_2_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_2_6_DXMUX,
      CE => U_DCT1D_databuf_reg_2_6_CEINV,
      CLK => U_DCT1D_databuf_reg_2_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_2_6_FFX_RST,
      O => U_DCT1D_databuf_reg_2_Q(6)
    );
  U_DCT1D_databuf_reg_2_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_2_6_FFX_RST
    );
  U_DCT2D_rtlc5n1481_5_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_5_XORF,
      O => U_DCT2D_rtlc5n1481(5)
    );
  U_DCT2D_rtlc5n1481_5_XORF_3015 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1481_5_CYINIT,
      I1 => U_DCT2D_nx65206z156,
      O => U_DCT2D_rtlc5n1481_5_XORF
    );
  U_DCT2D_rtlc5n1481_5_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_5_CY0F,
      IB => U_DCT2D_rtlc5n1481_5_CYINIT,
      SEL => U_DCT2D_rtlc5n1481_5_CYSELF,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63528_O
    );
  U_DCT2D_rtlc5n1481_5_CYMUXF2_3016 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_5_CY0F,
      IB => U_DCT2D_rtlc5n1481_5_CY0F,
      SEL => U_DCT2D_rtlc5n1481_5_CYSELF,
      O => U_DCT2D_rtlc5n1481_5_CYMUXF2
    );
  U_DCT2D_rtlc5n1481_5_CYINIT_3017 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63531_O,
      O => U_DCT2D_rtlc5n1481_5_CYINIT
    );
  U_DCT2D_rtlc5n1481_5_CY0F_3018 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(3),
      O => U_DCT2D_rtlc5n1481_5_CY0F
    );
  U_DCT2D_rtlc5n1481_5_CYSELF_3019 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z156,
      O => U_DCT2D_rtlc5n1481_5_CYSELF
    );
  U_DCT2D_rtlc5n1481_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_5_XORG,
      O => U_DCT2D_rtlc5n1481(6)
    );
  U_DCT2D_rtlc5n1481_5_XORG_3020 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_333_add_55_ix65206z63528_O,
      I1 => U_DCT2D_nx65206z153,
      O => U_DCT2D_rtlc5n1481_5_XORG
    );
  U_DCT2D_rtlc5n1481_5_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_5_CYMUXFAST,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63524_O
    );
  U_DCT2D_rtlc5n1481_5_FASTCARRY_3021 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63531_O,
      O => U_DCT2D_rtlc5n1481_5_FASTCARRY
    );
  U_DCT2D_rtlc5n1481_5_CYAND_3022 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1481_5_CYSELG,
      I1 => U_DCT2D_rtlc5n1481_5_CYSELF,
      O => U_DCT2D_rtlc5n1481_5_CYAND
    );
  U_DCT2D_rtlc5n1481_5_CYMUXFAST_3023 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_5_CYMUXG2,
      IB => U_DCT2D_rtlc5n1481_5_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1481_5_CYAND,
      O => U_DCT2D_rtlc5n1481_5_CYMUXFAST
    );
  U_DCT2D_rtlc5n1481_5_CYMUXG2_3024 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_5_CY0G,
      IB => U_DCT2D_rtlc5n1481_5_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1481_5_CYSELG,
      O => U_DCT2D_rtlc5n1481_5_CYMUXG2
    );
  U_DCT2D_rtlc5n1481_5_CY0G_3025 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(4),
      O => U_DCT2D_rtlc5n1481_5_CY0G
    );
  U_DCT2D_rtlc5n1481_5_CYSELG_3026 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z153,
      O => U_DCT2D_rtlc5n1481_5_CYSELG
    );
  U_DCT2D_rtlc5n1481_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_7_XORF,
      O => U_DCT2D_rtlc5n1481(7)
    );
  U_DCT2D_rtlc5n1481_7_XORF_3027 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1481_7_CYINIT,
      I1 => U_DCT2D_nx65206z150,
      O => U_DCT2D_rtlc5n1481_7_XORF
    );
  U_DCT2D_rtlc5n1481_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_7_CY0F,
      IB => U_DCT2D_rtlc5n1481_7_CYINIT,
      SEL => U_DCT2D_rtlc5n1481_7_CYSELF,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63521_O
    );
  U_DCT2D_rtlc5n1481_7_CYMUXF2_3028 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_7_CY0F,
      IB => U_DCT2D_rtlc5n1481_7_CY0F,
      SEL => U_DCT2D_rtlc5n1481_7_CYSELF,
      O => U_DCT2D_rtlc5n1481_7_CYMUXF2
    );
  U_DCT2D_rtlc5n1481_7_CYINIT_3029 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63524_O,
      O => U_DCT2D_rtlc5n1481_7_CYINIT
    );
  U_DCT2D_rtlc5n1481_7_CY0F_3030 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(5),
      O => U_DCT2D_rtlc5n1481_7_CY0F
    );
  U_DCT2D_rtlc5n1481_7_CYSELF_3031 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z150,
      O => U_DCT2D_rtlc5n1481_7_CYSELF
    );
  U_DCT2D_rtlc5n1481_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_7_XORG,
      O => U_DCT2D_rtlc5n1481(8)
    );
  U_DCT2D_rtlc5n1481_7_XORG_3032 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_333_add_55_ix65206z63521_O,
      I1 => U_DCT2D_nx65206z147,
      O => U_DCT2D_rtlc5n1481_7_XORG
    );
  U_DCT2D_rtlc5n1481_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_7_CYMUXFAST,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63517_O
    );
  U_DCT2D_rtlc5n1481_7_FASTCARRY_3033 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63524_O,
      O => U_DCT2D_rtlc5n1481_7_FASTCARRY
    );
  U_DCT2D_rtlc5n1481_7_CYAND_3034 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1481_7_CYSELG,
      I1 => U_DCT2D_rtlc5n1481_7_CYSELF,
      O => U_DCT2D_rtlc5n1481_7_CYAND
    );
  U_DCT2D_rtlc5n1481_7_CYMUXFAST_3035 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_7_CYMUXG2,
      IB => U_DCT2D_rtlc5n1481_7_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1481_7_CYAND,
      O => U_DCT2D_rtlc5n1481_7_CYMUXFAST
    );
  U_DCT2D_rtlc5n1481_7_CYMUXG2_3036 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_7_CY0G,
      IB => U_DCT2D_rtlc5n1481_7_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1481_7_CYSELG,
      O => U_DCT2D_rtlc5n1481_7_CYMUXG2
    );
  U_DCT2D_rtlc5n1481_7_CY0G_3037 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(6),
      O => U_DCT2D_rtlc5n1481_7_CY0G
    );
  U_DCT2D_rtlc5n1481_7_CYSELG_3038 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z147,
      O => U_DCT2D_rtlc5n1481_7_CYSELG
    );
  U_DCT2D_rtlc5n1481_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_9_XORF,
      O => U_DCT2D_rtlc5n1481(9)
    );
  U_DCT2D_rtlc5n1481_9_XORF_3039 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1481_9_CYINIT,
      I1 => U_DCT2D_nx65206z144,
      O => U_DCT2D_rtlc5n1481_9_XORF
    );
  U_DCT2D_rtlc5n1481_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_9_CY0F,
      IB => U_DCT2D_rtlc5n1481_9_CYINIT,
      SEL => U_DCT2D_rtlc5n1481_9_CYSELF,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63514_O
    );
  U_DCT2D_rtlc5n1481_9_CYMUXF2_3040 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_9_CY0F,
      IB => U_DCT2D_rtlc5n1481_9_CY0F,
      SEL => U_DCT2D_rtlc5n1481_9_CYSELF,
      O => U_DCT2D_rtlc5n1481_9_CYMUXF2
    );
  U_DCT2D_rtlc5n1481_9_CYINIT_3041 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63517_O,
      O => U_DCT2D_rtlc5n1481_9_CYINIT
    );
  U_DCT2D_rtlc5n1481_9_CY0F_3042 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(7),
      O => U_DCT2D_rtlc5n1481_9_CY0F
    );
  U_DCT2D_rtlc5n1481_9_CYSELF_3043 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z144,
      O => U_DCT2D_rtlc5n1481_9_CYSELF
    );
  U_DCT2D_rtlc5n1481_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_9_XORG,
      O => U_DCT2D_rtlc5n1481(10)
    );
  U_DCT2D_rtlc5n1481_9_XORG_3044 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_333_add_55_ix65206z63514_O,
      I1 => U_DCT2D_nx65206z141,
      O => U_DCT2D_rtlc5n1481_9_XORG
    );
  U_DCT2D_rtlc5n1481_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_9_CYMUXFAST,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63510_O
    );
  U_DCT2D_rtlc5n1481_9_FASTCARRY_3045 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63517_O,
      O => U_DCT2D_rtlc5n1481_9_FASTCARRY
    );
  U_DCT2D_rtlc5n1481_9_CYAND_3046 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1481_9_CYSELG,
      I1 => U_DCT2D_rtlc5n1481_9_CYSELF,
      O => U_DCT2D_rtlc5n1481_9_CYAND
    );
  U_DCT2D_rtlc5n1481_9_CYMUXFAST_3047 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_9_CYMUXG2,
      IB => U_DCT2D_rtlc5n1481_9_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1481_9_CYAND,
      O => U_DCT2D_rtlc5n1481_9_CYMUXFAST
    );
  U_DCT2D_rtlc5n1481_9_CYMUXG2_3048 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_9_CY0G,
      IB => U_DCT2D_rtlc5n1481_9_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1481_9_CYSELG,
      O => U_DCT2D_rtlc5n1481_9_CYMUXG2
    );
  U_DCT2D_rtlc5n1481_9_CY0G_3049 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(8),
      O => U_DCT2D_rtlc5n1481_9_CY0G
    );
  U_DCT2D_rtlc5n1481_9_CYSELG_3050 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z141,
      O => U_DCT2D_rtlc5n1481_9_CYSELG
    );
  U_DCT2D_rtlc5n1481_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_11_XORF,
      O => U_DCT2D_rtlc5n1481(11)
    );
  U_DCT2D_rtlc5n1481_11_XORF_3051 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1481_11_CYINIT,
      I1 => U_DCT2D_nx65206z138,
      O => U_DCT2D_rtlc5n1481_11_XORF
    );
  U_DCT2D_rtlc5n1481_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_11_CY0F,
      IB => U_DCT2D_rtlc5n1481_11_CYINIT,
      SEL => U_DCT2D_rtlc5n1481_11_CYSELF,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63506_O
    );
  U_DCT2D_rtlc5n1481_11_CYMUXF2_3052 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_11_CY0F,
      IB => U_DCT2D_rtlc5n1481_11_CY0F,
      SEL => U_DCT2D_rtlc5n1481_11_CYSELF,
      O => U_DCT2D_rtlc5n1481_11_CYMUXF2
    );
  U_DCT2D_rtlc5n1481_11_CYINIT_3053 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63510_O,
      O => U_DCT2D_rtlc5n1481_11_CYINIT
    );
  U_DCT2D_rtlc5n1481_11_CY0F_3054 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(9),
      O => U_DCT2D_rtlc5n1481_11_CY0F
    );
  U_DCT2D_rtlc5n1481_11_CYSELF_3055 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z138,
      O => U_DCT2D_rtlc5n1481_11_CYSELF
    );
  U_DCT2D_rtlc5n1481_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_11_XORG,
      O => U_DCT2D_rtlc5n1481(12)
    );
  U_DCT2D_rtlc5n1481_11_XORG_3056 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_333_add_55_ix65206z63506_O,
      I1 => U_DCT2D_nx65206z135,
      O => U_DCT2D_rtlc5n1481_11_XORG
    );
  U_DCT2D_rtlc5n1481_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_11_CYMUXFAST,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63503_O
    );
  U_DCT2D_rtlc5n1481_11_FASTCARRY_3057 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63510_O,
      O => U_DCT2D_rtlc5n1481_11_FASTCARRY
    );
  U_DCT2D_rtlc5n1481_11_CYAND_3058 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1481_11_CYSELG,
      I1 => U_DCT2D_rtlc5n1481_11_CYSELF,
      O => U_DCT2D_rtlc5n1481_11_CYAND
    );
  U_DCT2D_rtlc5n1481_11_CYMUXFAST_3059 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_11_CYMUXG2,
      IB => U_DCT2D_rtlc5n1481_11_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1481_11_CYAND,
      O => U_DCT2D_rtlc5n1481_11_CYMUXFAST
    );
  U_DCT2D_rtlc5n1481_11_CYMUXG2_3060 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_11_CY0G,
      IB => U_DCT2D_rtlc5n1481_11_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1481_11_CYSELG,
      O => U_DCT2D_rtlc5n1481_11_CYMUXG2
    );
  U_DCT2D_rtlc5n1481_11_CY0G_3061 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(10),
      O => U_DCT2D_rtlc5n1481_11_CY0G
    );
  U_DCT2D_rtlc5n1481_11_CYSELG_3062 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z135,
      O => U_DCT2D_rtlc5n1481_11_CYSELG
    );
  U_DCT2D_rtlc5n1481_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_13_XORF,
      O => U_DCT2D_rtlc5n1481(13)
    );
  U_DCT2D_rtlc5n1481_13_XORF_3063 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1481_13_CYINIT,
      I1 => U_DCT2D_nx65206z132,
      O => U_DCT2D_rtlc5n1481_13_XORF
    );
  U_DCT2D_rtlc5n1481_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_13_CY0F,
      IB => U_DCT2D_rtlc5n1481_13_CYINIT,
      SEL => U_DCT2D_rtlc5n1481_13_CYSELF,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63499_O
    );
  U_DCT2D_rtlc5n1481_13_CYMUXF2_3064 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_13_CY0F,
      IB => U_DCT2D_rtlc5n1481_13_CY0F,
      SEL => U_DCT2D_rtlc5n1481_13_CYSELF,
      O => U_DCT2D_rtlc5n1481_13_CYMUXF2
    );
  U_DCT2D_rtlc5n1481_13_CYINIT_3065 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63503_O,
      O => U_DCT2D_rtlc5n1481_13_CYINIT
    );
  U_DCT2D_rtlc5n1481_13_CY0F_3066 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(11),
      O => U_DCT2D_rtlc5n1481_13_CY0F
    );
  U_DCT2D_rtlc5n1481_13_CYSELF_3067 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z132,
      O => U_DCT2D_rtlc5n1481_13_CYSELF
    );
  U_DCT2D_rtlc5n1481_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_13_XORG,
      O => U_DCT2D_rtlc5n1481(14)
    );
  U_DCT2D_rtlc5n1481_13_XORG_3068 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_333_add_55_ix65206z63499_O,
      I1 => U_DCT2D_nx65206z129,
      O => U_DCT2D_rtlc5n1481_13_XORG
    );
  U_DCT2D_rtlc5n1481_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_13_CYMUXFAST,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63496_O
    );
  U_DCT2D_rtlc5n1481_13_FASTCARRY_3069 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63503_O,
      O => U_DCT2D_rtlc5n1481_13_FASTCARRY
    );
  U_DCT2D_rtlc5n1481_13_CYAND_3070 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1481_13_CYSELG,
      I1 => U_DCT2D_rtlc5n1481_13_CYSELF,
      O => U_DCT2D_rtlc5n1481_13_CYAND
    );
  U_DCT2D_rtlc5n1481_13_CYMUXFAST_3071 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_13_CYMUXG2,
      IB => U_DCT2D_rtlc5n1481_13_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1481_13_CYAND,
      O => U_DCT2D_rtlc5n1481_13_CYMUXFAST
    );
  U_DCT2D_rtlc5n1481_13_CYMUXG2_3072 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_13_CY0G,
      IB => U_DCT2D_rtlc5n1481_13_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1481_13_CYSELG,
      O => U_DCT2D_rtlc5n1481_13_CYMUXG2
    );
  U_DCT2D_rtlc5n1481_13_CY0G_3073 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(12),
      O => U_DCT2D_rtlc5n1481_13_CY0G
    );
  U_DCT2D_rtlc5n1481_13_CYSELG_3074 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z129,
      O => U_DCT2D_rtlc5n1481_13_CYSELG
    );
  U_DCT2D_rtlc5n1481_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_15_XORF,
      O => U_DCT2D_rtlc5n1481(15)
    );
  U_DCT2D_rtlc5n1481_15_XORF_3075 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1481_15_CYINIT,
      I1 => U_DCT2D_nx65206z126,
      O => U_DCT2D_rtlc5n1481_15_XORF
    );
  U_DCT2D_rtlc5n1481_15_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_15_CY0F,
      IB => U_DCT2D_rtlc5n1481_15_CYINIT,
      SEL => U_DCT2D_rtlc5n1481_15_CYSELF,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63492_O
    );
  U_DCT2D_rtlc5n1481_15_CYMUXF2_3076 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_15_CY0F,
      IB => U_DCT2D_rtlc5n1481_15_CY0F,
      SEL => U_DCT2D_rtlc5n1481_15_CYSELF,
      O => U_DCT2D_rtlc5n1481_15_CYMUXF2
    );
  U_DCT2D_rtlc5n1481_15_CYINIT_3077 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63496_O,
      O => U_DCT2D_rtlc5n1481_15_CYINIT
    );
  U_DCT2D_rtlc5n1481_15_CY0F_3078 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(13),
      O => U_DCT2D_rtlc5n1481_15_CY0F
    );
  U_DCT2D_rtlc5n1481_15_CYSELF_3079 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z126,
      O => U_DCT2D_rtlc5n1481_15_CYSELF
    );
  U_DCT2D_rtlc5n1481_15_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_15_XORG,
      O => U_DCT2D_rtlc5n1481(16)
    );
  U_DCT2D_rtlc5n1481_15_XORG_3080 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_333_add_55_ix65206z63492_O,
      I1 => U_DCT2D_nx65206z123,
      O => U_DCT2D_rtlc5n1481_15_XORG
    );
  U_DCT2D_rtlc5n1481_15_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_15_CYMUXFAST,
      O => U_DCT2D_rtlc_333_add_55_ix65206z63489_O
    );
  U_DCT2D_rtlc5n1481_15_FASTCARRY_3081 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63496_O,
      O => U_DCT2D_rtlc5n1481_15_FASTCARRY
    );
  U_DCT2D_rtlc5n1481_15_CYAND_3082 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1481_15_CYSELG,
      I1 => U_DCT2D_rtlc5n1481_15_CYSELF,
      O => U_DCT2D_rtlc5n1481_15_CYAND
    );
  U_DCT2D_rtlc5n1481_15_CYMUXFAST_3083 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_15_CYMUXG2,
      IB => U_DCT2D_rtlc5n1481_15_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1481_15_CYAND,
      O => U_DCT2D_rtlc5n1481_15_CYMUXFAST
    );
  U_DCT2D_rtlc5n1481_15_CYMUXG2_3084 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1481_15_CY0G,
      IB => U_DCT2D_rtlc5n1481_15_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1481_15_CYSELG,
      O => U_DCT2D_rtlc5n1481_15_CYMUXG2
    );
  U_DCT2D_rtlc5n1481_15_CY0G_3085 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s(13),
      O => U_DCT2D_rtlc5n1481_15_CY0G
    );
  U_DCT2D_rtlc5n1481_15_CYSELG_3086 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z123,
      O => U_DCT2D_rtlc5n1481_15_CYSELG
    );
  U_DCT2D_nx65206z121_rt_3087 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_nx65206z121,
      O => U_DCT2D_nx65206z121_rt
    );
  U_DCT2D_rtlc5n1481_17_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1481_17_XORF,
      O => U_DCT2D_rtlc5n1481(17)
    );
  U_DCT2D_rtlc5n1481_17_XORF_3088 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1481_17_CYINIT,
      I1 => U_DCT2D_nx65206z121_rt,
      O => U_DCT2D_rtlc5n1481_17_XORF
    );
  U_DCT2D_rtlc5n1481_17_CYINIT_3089 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_333_add_55_ix65206z63489_O,
      O => U_DCT2D_rtlc5n1481_17_CYINIT
    );
  U_DCT2D_rtlc5n1498_8_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_8_XORF,
      O => U_DCT2D_rtlc5n1498(8)
    );
  U_DCT2D_rtlc5n1498_8_XORF_3090 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1498_8_CYINIT,
      I1 => U_DCT2D_nx65206z411,
      O => U_DCT2D_rtlc5n1498_8_XORF
    );
  U_DCT2D_rtlc5n1498_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_8_CY0F,
      IB => U_DCT2D_rtlc5n1498_8_CYINIT,
      SEL => U_DCT2D_rtlc5n1498_8_CYSELF,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63910_O
    );
  U_DCT2D_rtlc5n1498_8_CYINIT_3091 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_8_BXINVNOT,
      O => U_DCT2D_rtlc5n1498_8_CYINIT
    );
  U_DCT2D_rtlc5n1498_8_CY0F_3092 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(8),
      O => U_DCT2D_rtlc5n1498_8_CY0F
    );
  U_DCT2D_rtlc5n1498_8_CYSELF_3093 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z411,
      O => U_DCT2D_rtlc5n1498_8_CYSELF
    );
  U_DCT2D_rtlc5n1498_8_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_6,
      O => U_DCT2D_rtlc5n1498_8_BXINVNOT
    );
  U_DCT2D_rtlc5n1498_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_8_XORG,
      O => U_DCT2D_rtlc5n1498(9)
    );
  U_DCT2D_rtlc5n1498_8_XORG_3094 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_399_add_69_ix65206z63910_O,
      I1 => U_DCT2D_nx65206z408,
      O => U_DCT2D_rtlc5n1498_8_XORG
    );
  U_DCT2D_rtlc5n1498_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_8_CYMUXG,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63904_O
    );
  U_DCT2D_rtlc5n1498_8_CYMUXG_3095 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_8_CY0G,
      IB => U_DCT2D_rtlc_399_add_69_ix65206z63910_O,
      SEL => U_DCT2D_rtlc5n1498_8_CYSELG,
      O => U_DCT2D_rtlc5n1498_8_CYMUXG
    );
  U_DCT2D_rtlc5n1498_8_CY0G_3096 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(9),
      O => U_DCT2D_rtlc5n1498_8_CY0G
    );
  U_DCT2D_rtlc5n1498_8_CYSELG_3097 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z408,
      O => U_DCT2D_rtlc5n1498_8_CYSELG
    );
  U_DCT2D_rtlc5n1498_10_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_10_XORF,
      O => U_DCT2D_rtlc5n1498(10)
    );
  U_DCT2D_rtlc5n1498_10_XORF_3098 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1498_10_CYINIT,
      I1 => U_DCT2D_nx65206z405,
      O => U_DCT2D_rtlc5n1498_10_XORF
    );
  U_DCT2D_rtlc5n1498_10_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_10_CY0F,
      IB => U_DCT2D_rtlc5n1498_10_CYINIT,
      SEL => U_DCT2D_rtlc5n1498_10_CYSELF,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63898_O
    );
  U_DCT2D_rtlc5n1498_10_CYMUXF2_3099 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_10_CY0F,
      IB => U_DCT2D_rtlc5n1498_10_CY0F,
      SEL => U_DCT2D_rtlc5n1498_10_CYSELF,
      O => U_DCT2D_rtlc5n1498_10_CYMUXF2
    );
  U_DCT2D_rtlc5n1498_10_CYINIT_3100 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63904_O,
      O => U_DCT2D_rtlc5n1498_10_CYINIT
    );
  U_DCT2D_rtlc5n1498_10_CY0F_3101 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(10),
      O => U_DCT2D_rtlc5n1498_10_CY0F
    );
  U_DCT2D_rtlc5n1498_10_CYSELF_3102 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z405,
      O => U_DCT2D_rtlc5n1498_10_CYSELF
    );
  U_DCT2D_rtlc5n1498_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_10_XORG,
      O => U_DCT2D_rtlc5n1498(11)
    );
  U_DCT2D_rtlc5n1498_10_XORG_3103 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_399_add_69_ix65206z63898_O,
      I1 => U_DCT2D_nx65206z402,
      O => U_DCT2D_rtlc5n1498_10_XORG
    );
  U_DCT2D_rtlc5n1498_10_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_10_CYMUXFAST,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63892_O
    );
  U_DCT2D_rtlc5n1498_10_FASTCARRY_3104 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63904_O,
      O => U_DCT2D_rtlc5n1498_10_FASTCARRY
    );
  U_DCT2D_rtlc5n1498_10_CYAND_3105 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1498_10_CYSELG,
      I1 => U_DCT2D_rtlc5n1498_10_CYSELF,
      O => U_DCT2D_rtlc5n1498_10_CYAND
    );
  U_DCT2D_rtlc5n1498_10_CYMUXFAST_3106 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_10_CYMUXG2,
      IB => U_DCT2D_rtlc5n1498_10_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1498_10_CYAND,
      O => U_DCT2D_rtlc5n1498_10_CYMUXFAST
    );
  U_DCT2D_rtlc5n1498_10_CYMUXG2_3107 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_10_CY0G,
      IB => U_DCT2D_rtlc5n1498_10_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1498_10_CYSELG,
      O => U_DCT2D_rtlc5n1498_10_CYMUXG2
    );
  U_DCT2D_rtlc5n1498_10_CY0G_3108 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(11),
      O => U_DCT2D_rtlc5n1498_10_CY0G
    );
  U_DCT2D_rtlc5n1498_10_CYSELG_3109 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z402,
      O => U_DCT2D_rtlc5n1498_10_CYSELG
    );
  U_DCT2D_rtlc5n1498_12_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_12_XORF,
      O => U_DCT2D_rtlc5n1498(12)
    );
  U_DCT2D_rtlc5n1498_12_XORF_3110 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1498_12_CYINIT,
      I1 => U_DCT2D_nx65206z399,
      O => U_DCT2D_rtlc5n1498_12_XORF
    );
  U_DCT2D_rtlc5n1498_12_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_12_CY0F,
      IB => U_DCT2D_rtlc5n1498_12_CYINIT,
      SEL => U_DCT2D_rtlc5n1498_12_CYSELF,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63886_O
    );
  U_DCT2D_rtlc5n1498_12_CYMUXF2_3111 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_12_CY0F,
      IB => U_DCT2D_rtlc5n1498_12_CY0F,
      SEL => U_DCT2D_rtlc5n1498_12_CYSELF,
      O => U_DCT2D_rtlc5n1498_12_CYMUXF2
    );
  U_DCT2D_rtlc5n1498_12_CYINIT_3112 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63892_O,
      O => U_DCT2D_rtlc5n1498_12_CYINIT
    );
  U_DCT2D_rtlc5n1498_12_CY0F_3113 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(12),
      O => U_DCT2D_rtlc5n1498_12_CY0F
    );
  U_DCT2D_rtlc5n1498_12_CYSELF_3114 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z399,
      O => U_DCT2D_rtlc5n1498_12_CYSELF
    );
  U_DCT2D_rtlc5n1498_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_12_XORG,
      O => U_DCT2D_rtlc5n1498(13)
    );
  U_DCT2D_rtlc5n1498_12_XORG_3115 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_399_add_69_ix65206z63886_O,
      I1 => U_DCT2D_nx65206z396,
      O => U_DCT2D_rtlc5n1498_12_XORG
    );
  U_DCT2D_rtlc5n1498_12_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_12_CYMUXFAST,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63880_O
    );
  U_DCT2D_rtlc5n1498_12_FASTCARRY_3116 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63892_O,
      O => U_DCT2D_rtlc5n1498_12_FASTCARRY
    );
  U_DCT2D_rtlc5n1498_12_CYAND_3117 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1498_12_CYSELG,
      I1 => U_DCT2D_rtlc5n1498_12_CYSELF,
      O => U_DCT2D_rtlc5n1498_12_CYAND
    );
  U_DCT2D_rtlc5n1498_12_CYMUXFAST_3118 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_12_CYMUXG2,
      IB => U_DCT2D_rtlc5n1498_12_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1498_12_CYAND,
      O => U_DCT2D_rtlc5n1498_12_CYMUXFAST
    );
  U_DCT2D_rtlc5n1498_12_CYMUXG2_3119 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_12_CY0G,
      IB => U_DCT2D_rtlc5n1498_12_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1498_12_CYSELG,
      O => U_DCT2D_rtlc5n1498_12_CYMUXG2
    );
  U_DCT2D_rtlc5n1498_12_CY0G_3120 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(13),
      O => U_DCT2D_rtlc5n1498_12_CY0G
    );
  U_DCT2D_rtlc5n1498_12_CYSELG_3121 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z396,
      O => U_DCT2D_rtlc5n1498_12_CYSELG
    );
  U_DCT2D_rtlc5n1498_14_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_14_XORF,
      O => U_DCT2D_rtlc5n1498(14)
    );
  U_DCT2D_rtlc5n1498_14_XORF_3122 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1498_14_CYINIT,
      I1 => U_DCT2D_nx65206z393,
      O => U_DCT2D_rtlc5n1498_14_XORF
    );
  U_DCT2D_rtlc5n1498_14_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_14_CY0F,
      IB => U_DCT2D_rtlc5n1498_14_CYINIT,
      SEL => U_DCT2D_rtlc5n1498_14_CYSELF,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63874_O
    );
  U_DCT2D_rtlc5n1498_14_CYMUXF2_3123 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_14_CY0F,
      IB => U_DCT2D_rtlc5n1498_14_CY0F,
      SEL => U_DCT2D_rtlc5n1498_14_CYSELF,
      O => U_DCT2D_rtlc5n1498_14_CYMUXF2
    );
  U_DCT2D_rtlc5n1498_14_CYINIT_3124 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63880_O,
      O => U_DCT2D_rtlc5n1498_14_CYINIT
    );
  U_DCT2D_rtlc5n1498_14_CY0F_3125 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(14),
      O => U_DCT2D_rtlc5n1498_14_CY0F
    );
  U_DCT2D_rtlc5n1498_14_CYSELF_3126 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z393,
      O => U_DCT2D_rtlc5n1498_14_CYSELF
    );
  U_DCT2D_rtlc5n1498_14_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_14_XORG,
      O => U_DCT2D_rtlc5n1498(15)
    );
  U_DCT2D_rtlc5n1498_14_XORG_3127 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_399_add_69_ix65206z63874_O,
      I1 => U_DCT2D_nx65206z390,
      O => U_DCT2D_rtlc5n1498_14_XORG
    );
  U_DCT2D_rtlc5n1498_14_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_14_CYMUXFAST,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63868_O
    );
  U_DCT2D_rtlc5n1498_14_FASTCARRY_3128 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63880_O,
      O => U_DCT2D_rtlc5n1498_14_FASTCARRY
    );
  U_DCT2D_rtlc5n1498_14_CYAND_3129 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1498_14_CYSELG,
      I1 => U_DCT2D_rtlc5n1498_14_CYSELF,
      O => U_DCT2D_rtlc5n1498_14_CYAND
    );
  U_DCT2D_rtlc5n1498_14_CYMUXFAST_3130 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_14_CYMUXG2,
      IB => U_DCT2D_rtlc5n1498_14_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1498_14_CYAND,
      O => U_DCT2D_rtlc5n1498_14_CYMUXFAST
    );
  U_DCT2D_rtlc5n1498_14_CYMUXG2_3131 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_14_CY0G,
      IB => U_DCT2D_rtlc5n1498_14_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1498_14_CYSELG,
      O => U_DCT2D_rtlc5n1498_14_CYMUXG2
    );
  U_DCT2D_rtlc5n1498_14_CY0G_3132 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(15),
      O => U_DCT2D_rtlc5n1498_14_CY0G
    );
  U_DCT2D_rtlc5n1498_14_CYSELG_3133 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z390,
      O => U_DCT2D_rtlc5n1498_14_CYSELG
    );
  U_DCT2D_rtlc5n1498_16_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_16_XORF,
      O => U_DCT2D_rtlc5n1498(16)
    );
  U_DCT2D_rtlc5n1498_16_XORF_3134 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1498_16_CYINIT,
      I1 => U_DCT2D_nx65206z387,
      O => U_DCT2D_rtlc5n1498_16_XORF
    );
  U_DCT2D_rtlc5n1498_16_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_16_CY0F,
      IB => U_DCT2D_rtlc5n1498_16_CYINIT,
      SEL => U_DCT2D_rtlc5n1498_16_CYSELF,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63862_O
    );
  U_DCT2D_rtlc5n1498_16_CYMUXF2_3135 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_16_CY0F,
      IB => U_DCT2D_rtlc5n1498_16_CY0F,
      SEL => U_DCT2D_rtlc5n1498_16_CYSELF,
      O => U_DCT2D_rtlc5n1498_16_CYMUXF2
    );
  U_DCT2D_rtlc5n1498_16_CYINIT_3136 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63868_O,
      O => U_DCT2D_rtlc5n1498_16_CYINIT
    );
  U_DCT2D_rtlc5n1498_16_CY0F_3137 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(16),
      O => U_DCT2D_rtlc5n1498_16_CY0F
    );
  U_DCT2D_rtlc5n1498_16_CYSELF_3138 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z387,
      O => U_DCT2D_rtlc5n1498_16_CYSELF
    );
  U_DCT2D_rtlc5n1498_16_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_16_XORG,
      O => U_DCT2D_rtlc5n1498(17)
    );
  U_DCT2D_rtlc5n1498_16_XORG_3139 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_399_add_69_ix65206z63862_O,
      I1 => U_DCT2D_nx65206z384,
      O => U_DCT2D_rtlc5n1498_16_XORG
    );
  U_DCT2D_rtlc5n1498_16_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_16_CYMUXFAST,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63856_O
    );
  U_DCT2D_rtlc5n1498_16_FASTCARRY_3140 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63868_O,
      O => U_DCT2D_rtlc5n1498_16_FASTCARRY
    );
  U_DCT2D_rtlc5n1498_16_CYAND_3141 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1498_16_CYSELG,
      I1 => U_DCT2D_rtlc5n1498_16_CYSELF,
      O => U_DCT2D_rtlc5n1498_16_CYAND
    );
  U_DCT2D_rtlc5n1498_16_CYMUXFAST_3142 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_16_CYMUXG2,
      IB => U_DCT2D_rtlc5n1498_16_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1498_16_CYAND,
      O => U_DCT2D_rtlc5n1498_16_CYMUXFAST
    );
  U_DCT2D_rtlc5n1498_16_CYMUXG2_3143 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_16_CY0G,
      IB => U_DCT2D_rtlc5n1498_16_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1498_16_CYSELG,
      O => U_DCT2D_rtlc5n1498_16_CYMUXG2
    );
  U_DCT2D_rtlc5n1498_16_CY0G_3144 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(17),
      O => U_DCT2D_rtlc5n1498_16_CY0G
    );
  U_DCT2D_rtlc5n1498_16_CYSELG_3145 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z384,
      O => U_DCT2D_rtlc5n1498_16_CYSELG
    );
  U_DCT2D_rtlc5n1498_18_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_18_XORF,
      O => U_DCT2D_rtlc5n1498(18)
    );
  U_DCT2D_rtlc5n1498_18_XORF_3146 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1498_18_CYINIT,
      I1 => U_DCT2D_nx65206z381,
      O => U_DCT2D_rtlc5n1498_18_XORF
    );
  U_DCT2D_rtlc5n1498_18_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_18_CY0F,
      IB => U_DCT2D_rtlc5n1498_18_CYINIT,
      SEL => U_DCT2D_rtlc5n1498_18_CYSELF,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63851_O
    );
  U_DCT2D_rtlc5n1498_18_CYMUXF2_3147 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_18_CY0F,
      IB => U_DCT2D_rtlc5n1498_18_CY0F,
      SEL => U_DCT2D_rtlc5n1498_18_CYSELF,
      O => U_DCT2D_rtlc5n1498_18_CYMUXF2
    );
  U_DCT2D_rtlc5n1498_18_CYINIT_3148 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63856_O,
      O => U_DCT2D_rtlc5n1498_18_CYINIT
    );
  U_DCT2D_rtlc5n1498_18_CY0F_3149 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(18),
      O => U_DCT2D_rtlc5n1498_18_CY0F
    );
  U_DCT2D_rtlc5n1498_18_CYSELF_3150 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z381,
      O => U_DCT2D_rtlc5n1498_18_CYSELF
    );
  U_DCT2D_rtlc5n1498_18_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_18_XORG,
      O => U_DCT2D_rtlc5n1498(19)
    );
  U_DCT2D_rtlc5n1498_18_XORG_3151 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_399_add_69_ix65206z63851_O,
      I1 => U_DCT2D_nx65206z378,
      O => U_DCT2D_rtlc5n1498_18_XORG
    );
  U_DCT2D_rtlc5n1498_18_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_18_CYMUXFAST,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63847_O
    );
  U_DCT2D_rtlc5n1498_18_FASTCARRY_3152 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63856_O,
      O => U_DCT2D_rtlc5n1498_18_FASTCARRY
    );
  U_DCT2D_rtlc5n1498_18_CYAND_3153 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1498_18_CYSELG,
      I1 => U_DCT2D_rtlc5n1498_18_CYSELF,
      O => U_DCT2D_rtlc5n1498_18_CYAND
    );
  U_DCT2D_rtlc5n1498_18_CYMUXFAST_3154 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_18_CYMUXG2,
      IB => U_DCT2D_rtlc5n1498_18_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1498_18_CYAND,
      O => U_DCT2D_rtlc5n1498_18_CYMUXFAST
    );
  U_DCT2D_rtlc5n1498_18_CYMUXG2_3155 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_18_CY0G,
      IB => U_DCT2D_rtlc5n1498_18_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1498_18_CYSELG,
      O => U_DCT2D_rtlc5n1498_18_CYMUXG2
    );
  U_DCT2D_rtlc5n1498_18_CY0G_3156 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(19),
      O => U_DCT2D_rtlc5n1498_18_CY0G
    );
  U_DCT2D_rtlc5n1498_18_CYSELG_3157 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z378,
      O => U_DCT2D_rtlc5n1498_18_CYSELG
    );
  U_DCT2D_rtlc5n1498_20_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_20_XORF,
      O => U_DCT2D_rtlc5n1498(20)
    );
  U_DCT2D_rtlc5n1498_20_XORF_3158 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1498_20_CYINIT,
      I1 => U_DCT2D_nx65206z375,
      O => U_DCT2D_rtlc5n1498_20_XORF
    );
  U_DCT2D_rtlc5n1498_20_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_20_CY0F,
      IB => U_DCT2D_rtlc5n1498_20_CYINIT,
      SEL => U_DCT2D_rtlc5n1498_20_CYSELF,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63843_O
    );
  U_DCT2D_rtlc5n1498_20_CYMUXF2_3159 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_20_CY0F,
      IB => U_DCT2D_rtlc5n1498_20_CY0F,
      SEL => U_DCT2D_rtlc5n1498_20_CYSELF,
      O => U_DCT2D_rtlc5n1498_20_CYMUXF2
    );
  U_DCT2D_rtlc5n1498_20_CYINIT_3160 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63847_O,
      O => U_DCT2D_rtlc5n1498_20_CYINIT
    );
  U_DCT2D_rtlc5n1498_20_CY0F_3161 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(19),
      O => U_DCT2D_rtlc5n1498_20_CY0F
    );
  U_DCT2D_rtlc5n1498_20_CYSELF_3162 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z375,
      O => U_DCT2D_rtlc5n1498_20_CYSELF
    );
  U_DCT2D_rtlc5n1498_20_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_20_XORG,
      O => U_DCT2D_rtlc5n1498(21)
    );
  U_DCT2D_rtlc5n1498_20_XORG_3163 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_399_add_69_ix65206z63843_O,
      I1 => U_DCT2D_nx65206z372,
      O => U_DCT2D_rtlc5n1498_20_XORG
    );
  U_DCT2D_rtlc5n1498_20_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_20_CYMUXFAST,
      O => U_DCT2D_rtlc_399_add_69_ix65206z63839_O
    );
  U_DCT2D_rtlc5n1498_20_FASTCARRY_3164 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63847_O,
      O => U_DCT2D_rtlc5n1498_20_FASTCARRY
    );
  U_DCT2D_rtlc5n1498_20_CYAND_3165 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1498_20_CYSELG,
      I1 => U_DCT2D_rtlc5n1498_20_CYSELF,
      O => U_DCT2D_rtlc5n1498_20_CYAND
    );
  U_DCT2D_rtlc5n1498_20_CYMUXFAST_3166 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_20_CYMUXG2,
      IB => U_DCT2D_rtlc5n1498_20_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1498_20_CYAND,
      O => U_DCT2D_rtlc5n1498_20_CYMUXFAST
    );
  U_DCT2D_rtlc5n1498_20_CYMUXG2_3167 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1498_20_CY0G,
      IB => U_DCT2D_rtlc5n1498_20_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1498_20_CYSELG,
      O => U_DCT2D_rtlc5n1498_20_CYMUXG2
    );
  U_DCT2D_rtlc5n1498_20_CY0G_3168 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1494(19),
      O => U_DCT2D_rtlc5n1498_20_CY0G
    );
  U_DCT2D_rtlc5n1498_20_CYSELG_3169 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z372,
      O => U_DCT2D_rtlc5n1498_20_CYSELG
    );
  U_DCT2D_rtlc5n1498_22_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1498_22_XORF,
      O => U_DCT2D_rtlc5n1498(22)
    );
  U_DCT2D_rtlc5n1498_22_XORF_3170 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1498_22_CYINIT,
      I1 => U_DCT2D_nx65206z296_rt,
      O => U_DCT2D_rtlc5n1498_22_XORF
    );
  U_DCT2D_rtlc5n1498_22_CYINIT_3171 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_399_add_69_ix65206z63839_O,
      O => U_DCT2D_rtlc5n1498_22_CYINIT
    );
  U_DCT1D_rtlc5n1354_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_4_CY0F,
      IB => U_DCT1D_rtlc5n1354_4_CYINIT,
      SEL => U_DCT1D_rtlc5n1354_4_CYSELF,
      O => U_DCT1D_rtlc_510_add_27_ix59700z63433_O
    );
  U_DCT1D_rtlc5n1354_4_CYINIT_3172 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_4_BXINVNOT,
      O => U_DCT1D_rtlc5n1354_4_CYINIT
    );
  U_DCT1D_rtlc5n1354_4_CY0F_3173 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s(3),
      O => U_DCT1D_rtlc5n1354_4_CY0F
    );
  U_DCT1D_rtlc5n1354_4_CYSELF_3174 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z77,
      O => U_DCT1D_rtlc5n1354_4_CYSELF
    );
  U_DCT1D_rtlc5n1354_4_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_20,
      O => U_DCT1D_rtlc5n1354_4_BXINVNOT
    );
  U_DCT1D_rtlc5n1354_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_4_XORG,
      O => U_DCT1D_rtlc5n1354(4)
    );
  U_DCT1D_rtlc5n1354_4_XORG_3175 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_510_add_27_ix59700z63433_O,
      I1 => U_DCT1D_nx59700z74,
      O => U_DCT1D_rtlc5n1354_4_XORG
    );
  U_DCT1D_rtlc5n1354_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_4_CYMUXG,
      O => U_DCT1D_rtlc_510_add_27_ix59700z63429_O
    );
  U_DCT1D_rtlc5n1354_4_CYMUXG_3176 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_4_CY0G,
      IB => U_DCT1D_rtlc_510_add_27_ix59700z63433_O,
      SEL => U_DCT1D_rtlc5n1354_4_CYSELG,
      O => U_DCT1D_rtlc5n1354_4_CYMUXG
    );
  U_DCT1D_rtlc5n1354_4_CY0G_3177 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s(4),
      O => U_DCT1D_rtlc5n1354_4_CY0G
    );
  U_DCT1D_rtlc5n1354_4_CYSELG_3178 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z74,
      O => U_DCT1D_rtlc5n1354_4_CYSELG
    );
  U_DCT1D_rtlc5n1354_5_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_5_XORF,
      O => U_DCT1D_rtlc5n1354(5)
    );
  U_DCT1D_rtlc5n1354_5_XORF_3179 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1354_5_CYINIT,
      I1 => U_DCT1D_nx59700z71,
      O => U_DCT1D_rtlc5n1354_5_XORF
    );
  U_DCT1D_rtlc5n1354_5_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_5_CY0F,
      IB => U_DCT1D_rtlc5n1354_5_CYINIT,
      SEL => U_DCT1D_rtlc5n1354_5_CYSELF,
      O => U_DCT1D_rtlc_510_add_27_ix59700z63426_O
    );
  U_DCT1D_rtlc5n1354_5_CYMUXF2_3180 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_5_CY0F,
      IB => U_DCT1D_rtlc5n1354_5_CY0F,
      SEL => U_DCT1D_rtlc5n1354_5_CYSELF,
      O => U_DCT1D_rtlc5n1354_5_CYMUXF2
    );
  U_DCT1D_rtlc5n1354_5_CYINIT_3181 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_510_add_27_ix59700z63429_O,
      O => U_DCT1D_rtlc5n1354_5_CYINIT
    );
  U_DCT1D_rtlc5n1354_5_CY0F_3182 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s(5),
      O => U_DCT1D_rtlc5n1354_5_CY0F
    );
  U_DCT1D_rtlc5n1354_5_CYSELF_3183 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z71,
      O => U_DCT1D_rtlc5n1354_5_CYSELF
    );
  U_DCT1D_rtlc5n1354_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_5_XORG,
      O => U_DCT1D_rtlc5n1354(6)
    );
  U_DCT1D_rtlc5n1354_5_XORG_3184 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_510_add_27_ix59700z63426_O,
      I1 => U_DCT1D_nx59700z68,
      O => U_DCT1D_rtlc5n1354_5_XORG
    );
  U_DCT1D_rtlc5n1354_5_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_5_CYMUXFAST,
      O => U_DCT1D_rtlc_510_add_27_ix59700z63422_O
    );
  U_DCT1D_rtlc5n1354_5_FASTCARRY_3185 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_510_add_27_ix59700z63429_O,
      O => U_DCT1D_rtlc5n1354_5_FASTCARRY
    );
  U_DCT1D_rtlc5n1354_5_CYAND_3186 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1354_5_CYSELG,
      I1 => U_DCT1D_rtlc5n1354_5_CYSELF,
      O => U_DCT1D_rtlc5n1354_5_CYAND
    );
  U_DCT1D_rtlc5n1354_5_CYMUXFAST_3187 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_5_CYMUXG2,
      IB => U_DCT1D_rtlc5n1354_5_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1354_5_CYAND,
      O => U_DCT1D_rtlc5n1354_5_CYMUXFAST
    );
  U_DCT1D_rtlc5n1354_5_CYMUXG2_3188 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_5_CY0G,
      IB => U_DCT1D_rtlc5n1354_5_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1354_5_CYSELG,
      O => U_DCT1D_rtlc5n1354_5_CYMUXG2
    );
  U_DCT1D_rtlc5n1354_5_CY0G_3189 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s(6),
      O => U_DCT1D_rtlc5n1354_5_CY0G
    );
  U_DCT1D_rtlc5n1354_5_CYSELG_3190 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z68,
      O => U_DCT1D_rtlc5n1354_5_CYSELG
    );
  U_DCT1D_rtlc5n1354_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_7_XORF,
      O => U_DCT1D_rtlc5n1354(7)
    );
  U_DCT1D_rtlc5n1354_7_XORF_3191 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1354_7_CYINIT,
      I1 => U_DCT1D_nx59700z65,
      O => U_DCT1D_rtlc5n1354_7_XORF
    );
  U_DCT1D_rtlc5n1354_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_7_CY0F,
      IB => U_DCT1D_rtlc5n1354_7_CYINIT,
      SEL => U_DCT1D_rtlc5n1354_7_CYSELF,
      O => U_DCT1D_rtlc_510_add_27_ix59700z63419_O
    );
  U_DCT1D_rtlc5n1354_7_CYMUXF2_3192 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_7_CY0F,
      IB => U_DCT1D_rtlc5n1354_7_CY0F,
      SEL => U_DCT1D_rtlc5n1354_7_CYSELF,
      O => U_DCT1D_rtlc5n1354_7_CYMUXF2
    );
  U_DCT1D_rtlc5n1354_7_CYINIT_3193 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_510_add_27_ix59700z63422_O,
      O => U_DCT1D_rtlc5n1354_7_CYINIT
    );
  U_DCT1D_rtlc5n1354_7_CY0F_3194 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s(7),
      O => U_DCT1D_rtlc5n1354_7_CY0F
    );
  U_DCT1D_rtlc5n1354_7_CYSELF_3195 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z65,
      O => U_DCT1D_rtlc5n1354_7_CYSELF
    );
  U_DCT1D_rtlc5n1354_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_7_XORG,
      O => U_DCT1D_rtlc5n1354(8)
    );
  U_DCT1D_rtlc5n1354_7_XORG_3196 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_510_add_27_ix59700z63419_O,
      I1 => U_DCT1D_nx59700z62,
      O => U_DCT1D_rtlc5n1354_7_XORG
    );
  U_DCT1D_rtlc5n1354_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_7_CYMUXFAST,
      O => U_DCT1D_rtlc_510_add_27_ix59700z63415_O
    );
  U_DCT1D_rtlc5n1354_7_FASTCARRY_3197 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_510_add_27_ix59700z63422_O,
      O => U_DCT1D_rtlc5n1354_7_FASTCARRY
    );
  U_DCT1D_rtlc5n1354_7_CYAND_3198 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1354_7_CYSELG,
      I1 => U_DCT1D_rtlc5n1354_7_CYSELF,
      O => U_DCT1D_rtlc5n1354_7_CYAND
    );
  U_DCT1D_rtlc5n1354_7_CYMUXFAST_3199 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_7_CYMUXG2,
      IB => U_DCT1D_rtlc5n1354_7_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1354_7_CYAND,
      O => U_DCT1D_rtlc5n1354_7_CYMUXFAST
    );
  U_DCT1D_rtlc5n1354_7_CYMUXG2_3200 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_7_CY0G,
      IB => U_DCT1D_rtlc5n1354_7_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1354_7_CYSELG,
      O => U_DCT1D_rtlc5n1354_7_CYMUXG2
    );
  U_DCT1D_rtlc5n1354_7_CY0G_3201 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s(8),
      O => U_DCT1D_rtlc5n1354_7_CY0G
    );
  U_DCT1D_rtlc5n1354_7_CYSELG_3202 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z62,
      O => U_DCT1D_rtlc5n1354_7_CYSELG
    );
  U_DCT1D_rtlc5n1354_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_9_XORF,
      O => U_DCT1D_rtlc5n1354(9)
    );
  U_DCT1D_rtlc5n1354_9_XORF_3203 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1354_9_CYINIT,
      I1 => U_DCT1D_nx59700z59,
      O => U_DCT1D_rtlc5n1354_9_XORF
    );
  U_DCT1D_rtlc5n1354_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_9_CY0F,
      IB => U_DCT1D_rtlc5n1354_9_CYINIT,
      SEL => U_DCT1D_rtlc5n1354_9_CYSELF,
      O => U_DCT1D_rtlc_510_add_27_ix59700z63412_O
    );
  U_DCT1D_rtlc5n1354_9_CYMUXF2_3204 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_9_CY0F,
      IB => U_DCT1D_rtlc5n1354_9_CY0F,
      SEL => U_DCT1D_rtlc5n1354_9_CYSELF,
      O => U_DCT1D_rtlc5n1354_9_CYMUXF2
    );
  U_DCT1D_rtlc5n1354_9_CYINIT_3205 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_510_add_27_ix59700z63415_O,
      O => U_DCT1D_rtlc5n1354_9_CYINIT
    );
  U_DCT1D_rtlc5n1354_9_CY0F_3206 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s(9),
      O => U_DCT1D_rtlc5n1354_9_CY0F
    );
  U_DCT1D_rtlc5n1354_9_CYSELF_3207 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z59,
      O => U_DCT1D_rtlc5n1354_9_CYSELF
    );
  U_DCT1D_rtlc5n1354_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_9_XORG,
      O => U_DCT1D_rtlc5n1354(10)
    );
  U_DCT1D_rtlc5n1354_9_XORG_3208 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_510_add_27_ix59700z63412_O,
      I1 => U_DCT1D_nx59700z56,
      O => U_DCT1D_rtlc5n1354_9_XORG
    );
  U_DCT1D_rtlc5n1354_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_9_CYMUXFAST,
      O => U_DCT1D_rtlc_510_add_27_ix59700z63408_O
    );
  U_DCT1D_rtlc5n1354_9_FASTCARRY_3209 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_510_add_27_ix59700z63415_O,
      O => U_DCT1D_rtlc5n1354_9_FASTCARRY
    );
  U_DCT1D_rtlc5n1354_9_CYAND_3210 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1354_9_CYSELG,
      I1 => U_DCT1D_rtlc5n1354_9_CYSELF,
      O => U_DCT1D_rtlc5n1354_9_CYAND
    );
  U_DCT1D_rtlc5n1354_9_CYMUXFAST_3211 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_9_CYMUXG2,
      IB => U_DCT1D_rtlc5n1354_9_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1354_9_CYAND,
      O => U_DCT1D_rtlc5n1354_9_CYMUXFAST
    );
  U_DCT1D_rtlc5n1354_9_CYMUXG2_3212 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_9_CY0G,
      IB => U_DCT1D_rtlc5n1354_9_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1354_9_CYSELG,
      O => U_DCT1D_rtlc5n1354_9_CYMUXG2
    );
  U_DCT1D_rtlc5n1354_9_CY0G_3213 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s(10),
      O => U_DCT1D_rtlc5n1354_9_CY0G
    );
  U_DCT1D_rtlc5n1354_9_CYSELG_3214 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z56,
      O => U_DCT1D_rtlc5n1354_9_CYSELG
    );
  U_DCT1D_rtlc5n1354_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_11_XORF,
      O => U_DCT1D_rtlc5n1354(11)
    );
  U_DCT1D_rtlc5n1354_11_XORF_3215 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1354_11_CYINIT,
      I1 => U_DCT1D_nx59700z53,
      O => U_DCT1D_rtlc5n1354_11_XORF
    );
  U_DCT1D_rtlc5n1354_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_11_CY0F,
      IB => U_DCT1D_rtlc5n1354_11_CYINIT,
      SEL => U_DCT1D_rtlc5n1354_11_CYSELF,
      O => U_DCT1D_rtlc_510_add_27_ix59700z63405_O
    );
  U_DCT1D_rtlc5n1354_11_CYMUXF2_3216 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_11_CY0F,
      IB => U_DCT1D_rtlc5n1354_11_CY0F,
      SEL => U_DCT1D_rtlc5n1354_11_CYSELF,
      O => U_DCT1D_rtlc5n1354_11_CYMUXF2
    );
  U_DCT1D_rtlc5n1354_11_CYINIT_3217 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_510_add_27_ix59700z63408_O,
      O => U_DCT1D_rtlc5n1354_11_CYINIT
    );
  U_DCT1D_rtlc5n1354_11_CY0F_3218 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s(11),
      O => U_DCT1D_rtlc5n1354_11_CY0F
    );
  U_DCT1D_rtlc5n1354_11_CYSELF_3219 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z53,
      O => U_DCT1D_rtlc5n1354_11_CYSELF
    );
  U_DCT1D_rtlc5n1354_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_11_XORG,
      O => U_DCT1D_rtlc5n1354(12)
    );
  U_DCT1D_rtlc5n1354_11_XORG_3220 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_510_add_27_ix59700z63405_O,
      I1 => U_DCT1D_nx59700z50,
      O => U_DCT1D_rtlc5n1354_11_XORG
    );
  U_DCT1D_rtlc5n1354_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_11_CYMUXFAST,
      O => U_DCT1D_rtlc_510_add_27_ix59700z63401_O
    );
  U_DCT1D_rtlc5n1354_11_FASTCARRY_3221 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_510_add_27_ix59700z63408_O,
      O => U_DCT1D_rtlc5n1354_11_FASTCARRY
    );
  U_DCT1D_rtlc5n1354_11_CYAND_3222 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1354_11_CYSELG,
      I1 => U_DCT1D_rtlc5n1354_11_CYSELF,
      O => U_DCT1D_rtlc5n1354_11_CYAND
    );
  U_DCT1D_rtlc5n1354_11_CYMUXFAST_3223 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_11_CYMUXG2,
      IB => U_DCT1D_rtlc5n1354_11_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1354_11_CYAND,
      O => U_DCT1D_rtlc5n1354_11_CYMUXFAST
    );
  U_DCT1D_rtlc5n1354_11_CYMUXG2_3224 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_11_CY0G,
      IB => U_DCT1D_rtlc5n1354_11_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1354_11_CYSELG,
      O => U_DCT1D_rtlc5n1354_11_CYMUXG2
    );
  U_DCT1D_rtlc5n1354_11_CY0G_3225 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s(12),
      O => U_DCT1D_rtlc5n1354_11_CY0G
    );
  U_DCT1D_rtlc5n1354_11_CYSELG_3226 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z50,
      O => U_DCT1D_rtlc5n1354_11_CYSELG
    );
  U_DCT1D_rtlc5n1354_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_13_XORF,
      O => U_DCT1D_rtlc5n1354(13)
    );
  U_DCT1D_rtlc5n1354_13_XORF_3227 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1354_13_CYINIT,
      I1 => U_DCT1D_nx59700z47,
      O => U_DCT1D_rtlc5n1354_13_XORF
    );
  U_DCT1D_rtlc5n1354_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_13_CY0F,
      IB => U_DCT1D_rtlc5n1354_13_CYINIT,
      SEL => U_DCT1D_rtlc5n1354_13_CYSELF,
      O => U_DCT1D_rtlc_510_add_27_ix59700z63398_O
    );
  U_DCT1D_rtlc5n1354_13_CYMUXF2_3228 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_13_CY0F,
      IB => U_DCT1D_rtlc5n1354_13_CY0F,
      SEL => U_DCT1D_rtlc5n1354_13_CYSELF,
      O => U_DCT1D_rtlc5n1354_13_CYMUXF2
    );
  U_DCT1D_rtlc5n1354_13_CYINIT_3229 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_510_add_27_ix59700z63401_O,
      O => U_DCT1D_rtlc5n1354_13_CYINIT
    );
  U_DCT1D_rtlc5n1354_13_CY0F_3230 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s(13),
      O => U_DCT1D_rtlc5n1354_13_CY0F
    );
  U_DCT1D_rtlc5n1354_13_CYSELF_3231 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z47,
      O => U_DCT1D_rtlc5n1354_13_CYSELF
    );
  U_DCT1D_rtlc5n1354_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_13_XORG,
      O => U_DCT1D_rtlc5n1354(14)
    );
  U_DCT1D_rtlc5n1354_13_XORG_3232 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_510_add_27_ix59700z63398_O,
      I1 => U_DCT1D_nx59700z44,
      O => U_DCT1D_rtlc5n1354_13_XORG
    );
  U_DCT1D_rtlc5n1354_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_13_CYMUXFAST,
      O => U_DCT1D_rtlc_510_add_27_ix59700z63392_O
    );
  U_DCT1D_rtlc5n1354_13_FASTCARRY_3233 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_510_add_27_ix59700z63401_O,
      O => U_DCT1D_rtlc5n1354_13_FASTCARRY
    );
  U_DCT1D_rtlc5n1354_13_CYAND_3234 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1354_13_CYSELG,
      I1 => U_DCT1D_rtlc5n1354_13_CYSELF,
      O => U_DCT1D_rtlc5n1354_13_CYAND
    );
  U_DCT1D_rtlc5n1354_13_CYMUXFAST_3235 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_13_CYMUXG2,
      IB => U_DCT1D_rtlc5n1354_13_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1354_13_CYAND,
      O => U_DCT1D_rtlc5n1354_13_CYMUXFAST
    );
  U_DCT1D_rtlc5n1354_13_CYMUXG2_3236 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1354_13_CY0G,
      IB => U_DCT1D_rtlc5n1354_13_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1354_13_CYSELG,
      O => U_DCT1D_rtlc5n1354_13_CYMUXG2
    );
  U_DCT1D_rtlc5n1354_13_CY0G_3237 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s(13),
      O => U_DCT1D_rtlc5n1354_13_CY0G
    );
  U_DCT1D_rtlc5n1354_13_CYSELG_3238 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z44,
      O => U_DCT1D_rtlc5n1354_13_CYSELG
    );
  U_DCT1D_nx59700z42_rt_3239 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z42,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z42_rt
    );
  U_DCT1D_rtlc5n1354_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1354_15_XORF,
      O => U_DCT1D_rtlc5n1354(15)
    );
  U_DCT1D_rtlc5n1354_15_XORF_3240 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1354_15_CYINIT,
      I1 => U_DCT1D_nx59700z42_rt,
      O => U_DCT1D_rtlc5n1354_15_XORF
    );
  U_DCT1D_rtlc5n1354_15_CYINIT_3241 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_510_add_27_ix59700z63392_O,
      O => U_DCT1D_rtlc5n1354_15_CYINIT
    );
  U_DCT1D_nx59700z493_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z493_XORF,
      O => U_DCT1D_nx59700z493
    );
  U_DCT1D_nx59700z493_XORF_3242 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z493_CYINIT,
      I1 => U_DCT1D_nx59700z493_F,
      O => U_DCT1D_nx59700z493_XORF
    );
  U_DCT1D_nx59700z493_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z493_CY0F,
      IB => U_DCT1D_nx59700z493_CYINIT,
      SEL => U_DCT1D_nx59700z493_CYSELF,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63689_O
    );
  U_DCT1D_nx59700z493_CYINIT_3243 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z493_BXINVNOT,
      O => U_DCT1D_nx59700z493_CYINIT
    );
  U_DCT1D_nx59700z493_CY0F_3244 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z251,
      O => U_DCT1D_nx59700z493_CY0F
    );
  U_DCT1D_nx59700z493_CYSELF_3245 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z493_F,
      O => U_DCT1D_nx59700z493_CYSELF
    );
  U_DCT1D_nx59700z493_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_13,
      O => U_DCT1D_nx59700z493_BXINVNOT
    );
  U_DCT1D_nx59700z493_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z493_XORG,
      O => U_DCT1D_nx59700z490
    );
  U_DCT1D_nx59700z493_XORG_3246 : X_XOR2
    port map (
      I0 => U_DCT1D_ix773_modgen_add_291_ix59700z63689_O,
      I1 => U_DCT1D_nx59700z247,
      O => U_DCT1D_nx59700z493_XORG
    );
  U_DCT1D_nx59700z493_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z493_CYMUXG,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63683_O
    );
  U_DCT1D_nx59700z493_CYMUXG_3247 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z493_CY0G,
      IB => U_DCT1D_ix773_modgen_add_291_ix59700z63689_O,
      SEL => U_DCT1D_nx59700z493_CYSELG,
      O => U_DCT1D_nx59700z493_CYMUXG
    );
  U_DCT1D_nx59700z493_CY0G_3248 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z248,
      O => U_DCT1D_nx59700z493_CY0G
    );
  U_DCT1D_nx59700z493_CYSELG_3249 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z247,
      O => U_DCT1D_nx59700z493_CYSELG
    );
  U_DCT1D_reg_databuf_reg_2_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_2_8_DXMUX,
      CE => U_DCT1D_databuf_reg_2_8_CEINV,
      CLK => U_DCT1D_databuf_reg_2_8_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_2_8_FFX_RST,
      O => U_DCT1D_databuf_reg_2_Q(8)
    );
  U_DCT1D_databuf_reg_2_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_2_8_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_2_8_FFX_RST
    );
  U_DCT1D_databuf_reg_2_8_FFX_RSTAND_3250 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_2_8_FFX_RSTAND
    );
  U_DCT1D_nx59700z487_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z487_XORF,
      O => U_DCT1D_nx59700z487
    );
  U_DCT1D_nx59700z487_XORF_3251 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z487_CYINIT,
      I1 => U_DCT1D_nx59700z244,
      O => U_DCT1D_nx59700z487_XORF
    );
  U_DCT1D_nx59700z487_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z487_CY0F,
      IB => U_DCT1D_nx59700z487_CYINIT,
      SEL => U_DCT1D_nx59700z487_CYSELF,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63677_O
    );
  U_DCT1D_nx59700z487_CYMUXF2_3252 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z487_CY0F,
      IB => U_DCT1D_nx59700z487_CY0F,
      SEL => U_DCT1D_nx59700z487_CYSELF,
      O => U_DCT1D_nx59700z487_CYMUXF2
    );
  U_DCT1D_nx59700z487_CYINIT_3253 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63683_O,
      O => U_DCT1D_nx59700z487_CYINIT
    );
  U_DCT1D_nx59700z487_CY0F_3254 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z245,
      O => U_DCT1D_nx59700z487_CY0F
    );
  U_DCT1D_nx59700z487_CYSELF_3255 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z244,
      O => U_DCT1D_nx59700z487_CYSELF
    );
  U_DCT1D_nx59700z487_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z487_XORG,
      O => U_DCT1D_nx59700z484
    );
  U_DCT1D_nx59700z487_XORG_3256 : X_XOR2
    port map (
      I0 => U_DCT1D_ix773_modgen_add_291_ix59700z63677_O,
      I1 => U_DCT1D_nx59700z241,
      O => U_DCT1D_nx59700z487_XORG
    );
  U_DCT1D_nx59700z487_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z487_CYMUXFAST,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63671_O
    );
  U_DCT1D_nx59700z487_FASTCARRY_3257 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63683_O,
      O => U_DCT1D_nx59700z487_FASTCARRY
    );
  U_DCT1D_nx59700z487_CYAND_3258 : X_AND2
    port map (
      I0 => U_DCT1D_nx59700z487_CYSELG,
      I1 => U_DCT1D_nx59700z487_CYSELF,
      O => U_DCT1D_nx59700z487_CYAND
    );
  U_DCT1D_nx59700z487_CYMUXFAST_3259 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z487_CYMUXG2,
      IB => U_DCT1D_nx59700z487_FASTCARRY,
      SEL => U_DCT1D_nx59700z487_CYAND,
      O => U_DCT1D_nx59700z487_CYMUXFAST
    );
  U_DCT1D_nx59700z487_CYMUXG2_3260 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z487_CY0G,
      IB => U_DCT1D_nx59700z487_CYMUXF2,
      SEL => U_DCT1D_nx59700z487_CYSELG,
      O => U_DCT1D_nx59700z487_CYMUXG2
    );
  U_DCT1D_nx59700z487_CY0G_3261 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z242,
      O => U_DCT1D_nx59700z487_CY0G
    );
  U_DCT1D_nx59700z487_CYSELG_3262 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z241,
      O => U_DCT1D_nx59700z487_CYSELG
    );
  U_DCT1D_nx59700z480_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z480_XORF,
      O => U_DCT1D_nx59700z480
    );
  U_DCT1D_nx59700z480_XORF_3263 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z480_CYINIT,
      I1 => U_DCT1D_nx59700z238,
      O => U_DCT1D_nx59700z480_XORF
    );
  U_DCT1D_nx59700z480_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z480_CY0F,
      IB => U_DCT1D_nx59700z480_CYINIT,
      SEL => U_DCT1D_nx59700z480_CYSELF,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63665_O
    );
  U_DCT1D_nx59700z480_CYMUXF2_3264 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z480_CY0F,
      IB => U_DCT1D_nx59700z480_CY0F,
      SEL => U_DCT1D_nx59700z480_CYSELF,
      O => U_DCT1D_nx59700z480_CYMUXF2
    );
  U_DCT1D_nx59700z480_CYINIT_3265 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63671_O,
      O => U_DCT1D_nx59700z480_CYINIT
    );
  U_DCT1D_nx59700z480_CY0F_3266 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z239,
      O => U_DCT1D_nx59700z480_CY0F
    );
  U_DCT1D_nx59700z480_CYSELF_3267 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z238,
      O => U_DCT1D_nx59700z480_CYSELF
    );
  U_DCT1D_nx59700z480_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z480_XORG,
      O => U_DCT1D_nx59700z476
    );
  U_DCT1D_nx59700z480_XORG_3268 : X_XOR2
    port map (
      I0 => U_DCT1D_ix773_modgen_add_291_ix59700z63665_O,
      I1 => U_DCT1D_nx59700z235,
      O => U_DCT1D_nx59700z480_XORG
    );
  U_DCT1D_nx59700z480_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z480_CYMUXFAST,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63659_O
    );
  U_DCT1D_nx59700z480_FASTCARRY_3269 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63671_O,
      O => U_DCT1D_nx59700z480_FASTCARRY
    );
  U_DCT1D_nx59700z480_CYAND_3270 : X_AND2
    port map (
      I0 => U_DCT1D_nx59700z480_CYSELG,
      I1 => U_DCT1D_nx59700z480_CYSELF,
      O => U_DCT1D_nx59700z480_CYAND
    );
  U_DCT1D_nx59700z480_CYMUXFAST_3271 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z480_CYMUXG2,
      IB => U_DCT1D_nx59700z480_FASTCARRY,
      SEL => U_DCT1D_nx59700z480_CYAND,
      O => U_DCT1D_nx59700z480_CYMUXFAST
    );
  U_DCT1D_nx59700z480_CYMUXG2_3272 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z480_CY0G,
      IB => U_DCT1D_nx59700z480_CYMUXF2,
      SEL => U_DCT1D_nx59700z480_CYSELG,
      O => U_DCT1D_nx59700z480_CYMUXG2
    );
  U_DCT1D_nx59700z480_CY0G_3273 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z236,
      O => U_DCT1D_nx59700z480_CY0G
    );
  U_DCT1D_nx59700z480_CYSELG_3274 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z235,
      O => U_DCT1D_nx59700z480_CYSELG
    );
  U_DCT1D_nx59700z472_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z472_XORF,
      O => U_DCT1D_nx59700z472
    );
  U_DCT1D_nx59700z472_XORF_3275 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z472_CYINIT,
      I1 => U_DCT1D_nx59700z232,
      O => U_DCT1D_nx59700z472_XORF
    );
  U_DCT1D_nx59700z472_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z472_CY0F,
      IB => U_DCT1D_nx59700z472_CYINIT,
      SEL => U_DCT1D_nx59700z472_CYSELF,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63653_O
    );
  U_DCT1D_nx59700z472_CYMUXF2_3276 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z472_CY0F,
      IB => U_DCT1D_nx59700z472_CY0F,
      SEL => U_DCT1D_nx59700z472_CYSELF,
      O => U_DCT1D_nx59700z472_CYMUXF2
    );
  U_DCT1D_nx59700z472_CYINIT_3277 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63659_O,
      O => U_DCT1D_nx59700z472_CYINIT
    );
  U_DCT1D_nx59700z472_CY0F_3278 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z233,
      O => U_DCT1D_nx59700z472_CY0F
    );
  U_DCT1D_nx59700z472_CYSELF_3279 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z232,
      O => U_DCT1D_nx59700z472_CYSELF
    );
  U_DCT1D_nx59700z472_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z472_XORG,
      O => U_DCT1D_nx59700z468
    );
  U_DCT1D_nx59700z472_XORG_3280 : X_XOR2
    port map (
      I0 => U_DCT1D_ix773_modgen_add_291_ix59700z63653_O,
      I1 => U_DCT1D_nx59700z229,
      O => U_DCT1D_nx59700z472_XORG
    );
  U_DCT1D_nx59700z472_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z472_CYMUXFAST,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63647_O
    );
  U_DCT1D_nx59700z472_FASTCARRY_3281 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63659_O,
      O => U_DCT1D_nx59700z472_FASTCARRY
    );
  U_DCT1D_nx59700z472_CYAND_3282 : X_AND2
    port map (
      I0 => U_DCT1D_nx59700z472_CYSELG,
      I1 => U_DCT1D_nx59700z472_CYSELF,
      O => U_DCT1D_nx59700z472_CYAND
    );
  U_DCT1D_nx59700z472_CYMUXFAST_3283 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z472_CYMUXG2,
      IB => U_DCT1D_nx59700z472_FASTCARRY,
      SEL => U_DCT1D_nx59700z472_CYAND,
      O => U_DCT1D_nx59700z472_CYMUXFAST
    );
  U_DCT1D_nx59700z472_CYMUXG2_3284 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z472_CY0G,
      IB => U_DCT1D_nx59700z472_CYMUXF2,
      SEL => U_DCT1D_nx59700z472_CYSELG,
      O => U_DCT1D_nx59700z472_CYMUXG2
    );
  U_DCT1D_nx59700z472_CY0G_3285 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z230,
      O => U_DCT1D_nx59700z472_CY0G
    );
  U_DCT1D_nx59700z472_CYSELG_3286 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z229,
      O => U_DCT1D_nx59700z472_CYSELG
    );
  U_DCT1D_nx59700z464_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z464_XORF,
      O => U_DCT1D_nx59700z464
    );
  U_DCT1D_nx59700z464_XORF_3287 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z464_CYINIT,
      I1 => U_DCT1D_nx59700z226,
      O => U_DCT1D_nx59700z464_XORF
    );
  U_DCT1D_nx59700z464_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z464_CY0F,
      IB => U_DCT1D_nx59700z464_CYINIT,
      SEL => U_DCT1D_nx59700z464_CYSELF,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63641_O
    );
  U_DCT1D_nx59700z464_CYMUXF2_3288 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z464_CY0F,
      IB => U_DCT1D_nx59700z464_CY0F,
      SEL => U_DCT1D_nx59700z464_CYSELF,
      O => U_DCT1D_nx59700z464_CYMUXF2
    );
  U_DCT1D_nx59700z464_CYINIT_3289 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63647_O,
      O => U_DCT1D_nx59700z464_CYINIT
    );
  U_DCT1D_nx59700z464_CY0F_3290 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z227,
      O => U_DCT1D_nx59700z464_CY0F
    );
  U_DCT1D_nx59700z464_CYSELF_3291 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z226,
      O => U_DCT1D_nx59700z464_CYSELF
    );
  U_DCT1D_nx59700z464_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z464_XORG,
      O => U_DCT1D_nx59700z460
    );
  U_DCT1D_nx59700z464_XORG_3292 : X_XOR2
    port map (
      I0 => U_DCT1D_ix773_modgen_add_291_ix59700z63641_O,
      I1 => U_DCT1D_nx59700z223,
      O => U_DCT1D_nx59700z464_XORG
    );
  U_DCT1D_nx59700z464_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z464_CYMUXFAST,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63635_O
    );
  U_DCT1D_nx59700z464_FASTCARRY_3293 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63647_O,
      O => U_DCT1D_nx59700z464_FASTCARRY
    );
  U_DCT1D_nx59700z464_CYAND_3294 : X_AND2
    port map (
      I0 => U_DCT1D_nx59700z464_CYSELG,
      I1 => U_DCT1D_nx59700z464_CYSELF,
      O => U_DCT1D_nx59700z464_CYAND
    );
  U_DCT1D_nx59700z464_CYMUXFAST_3295 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z464_CYMUXG2,
      IB => U_DCT1D_nx59700z464_FASTCARRY,
      SEL => U_DCT1D_nx59700z464_CYAND,
      O => U_DCT1D_nx59700z464_CYMUXFAST
    );
  U_DCT1D_nx59700z464_CYMUXG2_3296 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z464_CY0G,
      IB => U_DCT1D_nx59700z464_CYMUXF2,
      SEL => U_DCT1D_nx59700z464_CYSELG,
      O => U_DCT1D_nx59700z464_CYMUXG2
    );
  U_DCT1D_nx59700z464_CY0G_3297 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z224,
      O => U_DCT1D_nx59700z464_CY0G
    );
  U_DCT1D_nx59700z464_CYSELG_3298 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z223,
      O => U_DCT1D_nx59700z464_CYSELG
    );
  U_DCT1D_nx59700z456_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z456_XORF,
      O => U_DCT1D_nx59700z456
    );
  U_DCT1D_nx59700z456_XORF_3299 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z456_CYINIT,
      I1 => U_DCT1D_nx59700z220,
      O => U_DCT1D_nx59700z456_XORF
    );
  U_DCT1D_nx59700z456_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z456_CY0F,
      IB => U_DCT1D_nx59700z456_CYINIT,
      SEL => U_DCT1D_nx59700z456_CYSELF,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63629_O
    );
  U_DCT1D_nx59700z456_CYMUXF2_3300 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z456_CY0F,
      IB => U_DCT1D_nx59700z456_CY0F,
      SEL => U_DCT1D_nx59700z456_CYSELF,
      O => U_DCT1D_nx59700z456_CYMUXF2
    );
  U_DCT1D_nx59700z456_CYINIT_3301 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63635_O,
      O => U_DCT1D_nx59700z456_CYINIT
    );
  U_DCT1D_nx59700z456_CY0F_3302 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z221,
      O => U_DCT1D_nx59700z456_CY0F
    );
  U_DCT1D_nx59700z456_CYSELF_3303 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z220,
      O => U_DCT1D_nx59700z456_CYSELF
    );
  U_DCT1D_nx59700z456_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z456_XORG,
      O => U_DCT1D_nx59700z452
    );
  U_DCT1D_nx59700z456_XORG_3304 : X_XOR2
    port map (
      I0 => U_DCT1D_ix773_modgen_add_291_ix59700z63629_O,
      I1 => U_DCT1D_nx59700z217,
      O => U_DCT1D_nx59700z456_XORG
    );
  U_DCT1D_nx59700z456_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z456_CYMUXFAST,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63624_O
    );
  U_DCT1D_nx59700z456_FASTCARRY_3305 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63635_O,
      O => U_DCT1D_nx59700z456_FASTCARRY
    );
  U_DCT1D_nx59700z456_CYAND_3306 : X_AND2
    port map (
      I0 => U_DCT1D_nx59700z456_CYSELG,
      I1 => U_DCT1D_nx59700z456_CYSELF,
      O => U_DCT1D_nx59700z456_CYAND
    );
  U_DCT1D_nx59700z456_CYMUXFAST_3307 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z456_CYMUXG2,
      IB => U_DCT1D_nx59700z456_FASTCARRY,
      SEL => U_DCT1D_nx59700z456_CYAND,
      O => U_DCT1D_nx59700z456_CYMUXFAST
    );
  U_DCT1D_nx59700z456_CYMUXG2_3308 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z456_CY0G,
      IB => U_DCT1D_nx59700z456_CYMUXF2,
      SEL => U_DCT1D_nx59700z456_CYSELG,
      O => U_DCT1D_nx59700z456_CYMUXG2
    );
  U_DCT1D_nx59700z456_CY0G_3309 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z218,
      O => U_DCT1D_nx59700z456_CY0G
    );
  U_DCT1D_nx59700z456_CYSELG_3310 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z217,
      O => U_DCT1D_nx59700z456_CYSELG
    );
  U_DCT1D_nx59700z448_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z448_XORF,
      O => U_DCT1D_nx59700z448
    );
  U_DCT1D_nx59700z448_XORF_3311 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z448_CYINIT,
      I1 => U_DCT1D_nx59700z214,
      O => U_DCT1D_nx59700z448_XORF
    );
  U_DCT1D_nx59700z448_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z448_CY0F,
      IB => U_DCT1D_nx59700z448_CYINIT,
      SEL => U_DCT1D_nx59700z448_CYSELF,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63619_O
    );
  U_DCT1D_nx59700z448_CYMUXF2_3312 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z448_CY0F,
      IB => U_DCT1D_nx59700z448_CY0F,
      SEL => U_DCT1D_nx59700z448_CYSELF,
      O => U_DCT1D_nx59700z448_CYMUXF2
    );
  U_DCT1D_nx59700z448_CYINIT_3313 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63624_O,
      O => U_DCT1D_nx59700z448_CYINIT
    );
  U_DCT1D_nx59700z448_CY0F_3314 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z215,
      O => U_DCT1D_nx59700z448_CY0F
    );
  U_DCT1D_nx59700z448_CYSELF_3315 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z214,
      O => U_DCT1D_nx59700z448_CYSELF
    );
  U_DCT1D_nx59700z448_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z448_XORG,
      O => U_DCT1D_nx59700z444
    );
  U_DCT1D_nx59700z448_XORG_3316 : X_XOR2
    port map (
      I0 => U_DCT1D_ix773_modgen_add_291_ix59700z63619_O,
      I1 => U_DCT1D_nx59700z211,
      O => U_DCT1D_nx59700z448_XORG
    );
  U_DCT1D_nx59700z448_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z448_CYMUXFAST,
      O => U_DCT1D_ix773_modgen_add_291_ix59700z63615_O
    );
  U_DCT1D_nx59700z448_FASTCARRY_3317 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63624_O,
      O => U_DCT1D_nx59700z448_FASTCARRY
    );
  U_DCT1D_nx59700z448_CYAND_3318 : X_AND2
    port map (
      I0 => U_DCT1D_nx59700z448_CYSELG,
      I1 => U_DCT1D_nx59700z448_CYSELF,
      O => U_DCT1D_nx59700z448_CYAND
    );
  U_DCT1D_nx59700z448_CYMUXFAST_3319 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z448_CYMUXG2,
      IB => U_DCT1D_nx59700z448_FASTCARRY,
      SEL => U_DCT1D_nx59700z448_CYAND,
      O => U_DCT1D_nx59700z448_CYMUXFAST
    );
  U_DCT1D_nx59700z448_CYMUXG2_3320 : X_MUX2
    port map (
      IA => U_DCT1D_nx59700z448_CY0G,
      IB => U_DCT1D_nx59700z448_CYMUXF2,
      SEL => U_DCT1D_nx59700z448_CYSELG,
      O => U_DCT1D_nx59700z448_CYMUXG2
    );
  U_DCT1D_nx59700z448_CY0G_3321 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z212,
      O => U_DCT1D_nx59700z448_CY0G
    );
  U_DCT1D_nx59700z448_CYSELG_3322 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z211,
      O => U_DCT1D_nx59700z448_CYSELG
    );
  U_DCT1D_nx59700z4_rt_3323 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_nx59700z4,
      O => U_DCT1D_nx59700z4_rt
    );
  U_DCT1D_nx59700z3_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z3_XORF,
      O => U_DCT1D_nx59700z3
    );
  U_DCT1D_nx59700z3_XORF_3324 : X_XOR2
    port map (
      I0 => U_DCT1D_nx59700z3_CYINIT,
      I1 => U_DCT1D_nx59700z4_rt,
      O => U_DCT1D_nx59700z3_XORF
    );
  U_DCT1D_nx59700z3_CYINIT_3325 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix773_modgen_add_291_ix59700z63615_O,
      O => U_DCT1D_nx59700z3_CYINIT
    );
  U_DCT1D_ix59700z64053_O_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_ix59700z64053_O_CY0F,
      IB => U_DCT1D_ix59700z64053_O_CYINIT,
      SEL => U_DCT1D_ix59700z64053_O_CYSELF,
      O => U_DCT1D_ix59700z64056_O
    );
  U_DCT1D_ix59700z64053_O_CYINIT_3326 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GLOBAL_LOGIC1_21,
      O => U_DCT1D_ix59700z64053_O_CYINIT
    );
  U_DCT1D_ix59700z64053_O_CY0F_3327 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(8),
      O => U_DCT1D_ix59700z64053_O_CY0F
    );
  U_DCT1D_ix59700z64053_O_CYSELF_3328 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z528,
      O => U_DCT1D_ix59700z64053_O_CYSELF
    );
  U_DCT1D_ix59700z64053_O_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z64053_O_CYMUXG,
      O => U_DCT1D_ix59700z64053_O
    );
  U_DCT1D_ix59700z64053_O_CYMUXG_3329 : X_MUX2
    port map (
      IA => U_DCT1D_ix59700z64053_O_CY0G,
      IB => U_DCT1D_ix59700z64056_O,
      SEL => U_DCT1D_ix59700z64053_O_CYSELG,
      O => U_DCT1D_ix59700z64053_O_CYMUXG
    );
  U_DCT1D_ix59700z64053_O_CY0G_3330 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(9),
      O => U_DCT1D_ix59700z64053_O_CY0G
    );
  U_DCT1D_ix59700z64053_O_CYSELG_3331 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z526,
      O => U_DCT1D_ix59700z64053_O_CYSELG
    );
  U_DCT1D_ix59700z64047_O_CYMUXF2_3332 : X_MUX2
    port map (
      IA => U_DCT1D_ix59700z64047_O_CY0F,
      IB => U_DCT1D_ix59700z64047_O_CY0F,
      SEL => U_DCT1D_ix59700z64047_O_CYSELF,
      O => U_DCT1D_ix59700z64047_O_CYMUXF2
    );
  U_DCT1D_ix59700z64047_O_CY0F_3333 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(10),
      O => U_DCT1D_ix59700z64047_O_CY0F
    );
  U_DCT1D_ix59700z64047_O_CYSELF_3334 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z524,
      O => U_DCT1D_ix59700z64047_O_CYSELF
    );
  U_DCT1D_ix59700z64047_O_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z64047_O_CYMUXFAST,
      O => U_DCT1D_ix59700z64047_O
    );
  U_DCT1D_ix59700z64047_O_FASTCARRY_3335 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z64053_O,
      O => U_DCT1D_ix59700z64047_O_FASTCARRY
    );
  U_DCT1D_ix59700z64047_O_CYAND_3336 : X_AND2
    port map (
      I0 => U_DCT1D_ix59700z64047_O_CYSELG,
      I1 => U_DCT1D_ix59700z64047_O_CYSELF,
      O => U_DCT1D_ix59700z64047_O_CYAND
    );
  U_DCT1D_ix59700z64047_O_CYMUXFAST_3337 : X_MUX2
    port map (
      IA => U_DCT1D_ix59700z64047_O_CYMUXG2,
      IB => U_DCT1D_ix59700z64047_O_FASTCARRY,
      SEL => U_DCT1D_ix59700z64047_O_CYAND,
      O => U_DCT1D_ix59700z64047_O_CYMUXFAST
    );
  U_DCT1D_ix59700z64047_O_CYMUXG2_3338 : X_MUX2
    port map (
      IA => U_DCT1D_ix59700z64047_O_CY0G,
      IB => U_DCT1D_ix59700z64047_O_CYMUXF2,
      SEL => U_DCT1D_ix59700z64047_O_CYSELG,
      O => U_DCT1D_ix59700z64047_O_CYMUXG2
    );
  U_DCT1D_ix59700z64047_O_CY0G_3339 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(11),
      O => U_DCT1D_ix59700z64047_O_CY0G
    );
  U_DCT1D_ix59700z64047_O_CYSELG_3340 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z522,
      O => U_DCT1D_ix59700z64047_O_CYSELG
    );
  ramdatai_s_0_DXMUX_3341 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_0_FXMUX,
      O => ramdatai_s_0_DXMUX
    );
  ramdatai_s_0_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_0_FXMUX,
      O => U_DCT1D_rtlc5n2660
    );
  ramdatai_s_0_FXMUX_3342 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_0_XORF,
      O => ramdatai_s_0_FXMUX
    );
  ramdatai_s_0_XORF_3343 : X_XOR2
    port map (
      I0 => ramdatai_s_0_CYINIT,
      I1 => U_DCT1D_nx59700z519,
      O => ramdatai_s_0_XORF
    );
  ramdatai_s_0_CYMUXF : X_MUX2
    port map (
      IA => ramdatai_s_0_CY0F,
      IB => ramdatai_s_0_CYINIT,
      SEL => ramdatai_s_0_CYSELF,
      O => U_DCT1D_ix59700z64042_O
    );
  ramdatai_s_0_CYMUXF2_3344 : X_MUX2
    port map (
      IA => ramdatai_s_0_CY0F,
      IB => ramdatai_s_0_CY0F,
      SEL => ramdatai_s_0_CYSELF,
      O => ramdatai_s_0_CYMUXF2
    );
  ramdatai_s_0_CYINIT_3345 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z64047_O,
      O => ramdatai_s_0_CYINIT
    );
  ramdatai_s_0_CY0F_3346 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(12),
      O => ramdatai_s_0_CY0F
    );
  ramdatai_s_0_CYSELF_3347 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z519,
      O => ramdatai_s_0_CYSELF
    );
  ramdatai_s_0_DYMUX_3348 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_0_GYMUX,
      O => ramdatai_s_0_DYMUX
    );
  ramdatai_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_0_GYMUX,
      O => U_DCT1D_rtlc5n2659
    );
  ramdatai_s_0_GYMUX_3349 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_0_XORG,
      O => ramdatai_s_0_GYMUX
    );
  ramdatai_s_0_XORG_3350 : X_XOR2
    port map (
      I0 => U_DCT1D_ix59700z64042_O,
      I1 => U_DCT1D_nx59700z516,
      O => ramdatai_s_0_XORG
    );
  ramdatai_s_0_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_0_CYMUXFAST,
      O => U_DCT1D_ix59700z64038_O
    );
  ramdatai_s_0_FASTCARRY_3351 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z64047_O,
      O => ramdatai_s_0_FASTCARRY
    );
  ramdatai_s_0_CYAND_3352 : X_AND2
    port map (
      I0 => ramdatai_s_0_CYSELG,
      I1 => ramdatai_s_0_CYSELF,
      O => ramdatai_s_0_CYAND
    );
  ramdatai_s_0_CYMUXFAST_3353 : X_MUX2
    port map (
      IA => ramdatai_s_0_CYMUXG2,
      IB => ramdatai_s_0_FASTCARRY,
      SEL => ramdatai_s_0_CYAND,
      O => ramdatai_s_0_CYMUXFAST
    );
  ramdatai_s_0_CYMUXG2_3354 : X_MUX2
    port map (
      IA => ramdatai_s_0_CY0G,
      IB => ramdatai_s_0_CYMUXF2,
      SEL => ramdatai_s_0_CYSELG,
      O => ramdatai_s_0_CYMUXG2
    );
  ramdatai_s_0_CY0G_3355 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(13),
      O => ramdatai_s_0_CY0G
    );
  ramdatai_s_0_CYSELG_3356 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z516,
      O => ramdatai_s_0_CYSELG
    );
  ramdatai_s_0_SRINV_3357 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramdatai_s_0_SRINV
    );
  ramdatai_s_0_CLKINV_3358 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramdatai_s_0_CLKINV
    );
  ramdatai_s_0_CEINV_3359 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => ramdatai_s_0_CEINV
    );
  ramdatai_s_2_DXMUX_3360 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_2_FXMUX,
      O => ramdatai_s_2_DXMUX
    );
  ramdatai_s_2_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_2_FXMUX,
      O => U_DCT1D_rtlc5n2658
    );
  ramdatai_s_2_FXMUX_3361 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_2_XORF,
      O => ramdatai_s_2_FXMUX
    );
  ramdatai_s_2_XORF_3362 : X_XOR2
    port map (
      I0 => ramdatai_s_2_CYINIT,
      I1 => U_DCT1D_nx59700z513,
      O => ramdatai_s_2_XORF
    );
  ramdatai_s_2_CYMUXF : X_MUX2
    port map (
      IA => ramdatai_s_2_CY0F,
      IB => ramdatai_s_2_CYINIT,
      SEL => ramdatai_s_2_CYSELF,
      O => U_DCT1D_ix59700z64033_O
    );
  ramdatai_s_2_CYMUXF2_3363 : X_MUX2
    port map (
      IA => ramdatai_s_2_CY0F,
      IB => ramdatai_s_2_CY0F,
      SEL => ramdatai_s_2_CYSELF,
      O => ramdatai_s_2_CYMUXF2
    );
  ramdatai_s_2_CYINIT_3364 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z64038_O,
      O => ramdatai_s_2_CYINIT
    );
  ramdatai_s_2_CY0F_3365 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(14),
      O => ramdatai_s_2_CY0F
    );
  ramdatai_s_2_CYSELF_3366 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z513,
      O => ramdatai_s_2_CYSELF
    );
  ramdatai_s_2_DYMUX_3367 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_2_GYMUX,
      O => ramdatai_s_2_DYMUX
    );
  ramdatai_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_2_GYMUX,
      O => U_DCT1D_rtlc5n2657
    );
  ramdatai_s_2_GYMUX_3368 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_2_XORG,
      O => ramdatai_s_2_GYMUX
    );
  ramdatai_s_2_XORG_3369 : X_XOR2
    port map (
      I0 => U_DCT1D_ix59700z64033_O,
      I1 => U_DCT1D_nx59700z510,
      O => ramdatai_s_2_XORG
    );
  ramdatai_s_2_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_2_CYMUXFAST,
      O => U_DCT1D_ix59700z64029_O
    );
  ramdatai_s_2_FASTCARRY_3370 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z64038_O,
      O => ramdatai_s_2_FASTCARRY
    );
  ramdatai_s_2_CYAND_3371 : X_AND2
    port map (
      I0 => ramdatai_s_2_CYSELG,
      I1 => ramdatai_s_2_CYSELF,
      O => ramdatai_s_2_CYAND
    );
  ramdatai_s_2_CYMUXFAST_3372 : X_MUX2
    port map (
      IA => ramdatai_s_2_CYMUXG2,
      IB => ramdatai_s_2_FASTCARRY,
      SEL => ramdatai_s_2_CYAND,
      O => ramdatai_s_2_CYMUXFAST
    );
  ramdatai_s_2_CYMUXG2_3373 : X_MUX2
    port map (
      IA => ramdatai_s_2_CY0G,
      IB => ramdatai_s_2_CYMUXF2,
      SEL => ramdatai_s_2_CYSELG,
      O => ramdatai_s_2_CYMUXG2
    );
  ramdatai_s_2_CY0G_3374 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(15),
      O => ramdatai_s_2_CY0G
    );
  ramdatai_s_2_CYSELG_3375 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z510,
      O => ramdatai_s_2_CYSELG
    );
  ramdatai_s_2_SRINV_3376 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramdatai_s_2_SRINV
    );
  ramdatai_s_2_CLKINV_3377 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramdatai_s_2_CLKINV
    );
  ramdatai_s_2_CEINV_3378 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => ramdatai_s_2_CEINV
    );
  ramdatai_s_4_DXMUX_3379 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_4_FXMUX,
      O => ramdatai_s_4_DXMUX
    );
  ramdatai_s_4_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_4_FXMUX,
      O => U_DCT1D_rtlc5n2656
    );
  ramdatai_s_4_FXMUX_3380 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_4_XORF,
      O => ramdatai_s_4_FXMUX
    );
  ramdatai_s_4_XORF_3381 : X_XOR2
    port map (
      I0 => ramdatai_s_4_CYINIT,
      I1 => U_DCT1D_nx59700z507,
      O => ramdatai_s_4_XORF
    );
  ramdatai_s_4_CYMUXF : X_MUX2
    port map (
      IA => ramdatai_s_4_CY0F,
      IB => ramdatai_s_4_CYINIT,
      SEL => ramdatai_s_4_CYSELF,
      O => U_DCT1D_ix59700z64025_O
    );
  ramdatai_s_4_CYMUXF2_3382 : X_MUX2
    port map (
      IA => ramdatai_s_4_CY0F,
      IB => ramdatai_s_4_CY0F,
      SEL => ramdatai_s_4_CYSELF,
      O => ramdatai_s_4_CYMUXF2
    );
  ramdatai_s_4_CYINIT_3383 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z64029_O,
      O => ramdatai_s_4_CYINIT
    );
  ramdatai_s_4_CY0F_3384 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(16),
      O => ramdatai_s_4_CY0F
    );
  ramdatai_s_4_CYSELF_3385 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z507,
      O => ramdatai_s_4_CYSELF
    );
  ramdatai_s_4_DYMUX_3386 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_4_GYMUX,
      O => ramdatai_s_4_DYMUX
    );
  ramdatai_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_4_GYMUX,
      O => U_DCT1D_rtlc5n2655
    );
  ramdatai_s_4_GYMUX_3387 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_4_XORG,
      O => ramdatai_s_4_GYMUX
    );
  ramdatai_s_4_XORG_3388 : X_XOR2
    port map (
      I0 => U_DCT1D_ix59700z64025_O,
      I1 => U_DCT1D_nx59700z504,
      O => ramdatai_s_4_XORG
    );
  ramdatai_s_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_4_CYMUXFAST,
      O => U_DCT1D_ix59700z64020_O
    );
  ramdatai_s_4_FASTCARRY_3389 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z64029_O,
      O => ramdatai_s_4_FASTCARRY
    );
  ramdatai_s_4_CYAND_3390 : X_AND2
    port map (
      I0 => ramdatai_s_4_CYSELG,
      I1 => ramdatai_s_4_CYSELF,
      O => ramdatai_s_4_CYAND
    );
  ramdatai_s_4_CYMUXFAST_3391 : X_MUX2
    port map (
      IA => ramdatai_s_4_CYMUXG2,
      IB => ramdatai_s_4_FASTCARRY,
      SEL => ramdatai_s_4_CYAND,
      O => ramdatai_s_4_CYMUXFAST
    );
  ramdatai_s_4_CYMUXG2_3392 : X_MUX2
    port map (
      IA => ramdatai_s_4_CY0G,
      IB => ramdatai_s_4_CYMUXF2,
      SEL => ramdatai_s_4_CYSELG,
      O => ramdatai_s_4_CYMUXG2
    );
  ramdatai_s_4_CY0G_3393 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(17),
      O => ramdatai_s_4_CY0G
    );
  ramdatai_s_4_CYSELG_3394 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z504,
      O => ramdatai_s_4_CYSELG
    );
  ramdatai_s_4_SRINV_3395 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramdatai_s_4_SRINV
    );
  ramdatai_s_4_CLKINV_3396 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramdatai_s_4_CLKINV
    );
  ramdatai_s_4_CEINV_3397 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => ramdatai_s_4_CEINV
    );
  ramdatai_s_6_DXMUX_3398 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_6_FXMUX,
      O => ramdatai_s_6_DXMUX
    );
  ramdatai_s_6_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_6_FXMUX,
      O => U_DCT1D_rtlc5n2654
    );
  ramdatai_s_6_FXMUX_3399 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_6_XORF,
      O => ramdatai_s_6_FXMUX
    );
  ramdatai_s_6_XORF_3400 : X_XOR2
    port map (
      I0 => ramdatai_s_6_CYINIT,
      I1 => U_DCT1D_nx59700z501,
      O => ramdatai_s_6_XORF
    );
  ramdatai_s_6_CYMUXF : X_MUX2
    port map (
      IA => ramdatai_s_6_CY0F,
      IB => ramdatai_s_6_CYINIT,
      SEL => ramdatai_s_6_CYSELF,
      O => U_DCT1D_ix59700z64016_O
    );
  ramdatai_s_6_CYMUXF2_3401 : X_MUX2
    port map (
      IA => ramdatai_s_6_CY0F,
      IB => ramdatai_s_6_CY0F,
      SEL => ramdatai_s_6_CYSELF,
      O => ramdatai_s_6_CYMUXF2
    );
  ramdatai_s_6_CYINIT_3402 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z64020_O,
      O => ramdatai_s_6_CYINIT
    );
  ramdatai_s_6_CY0F_3403 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(18),
      O => ramdatai_s_6_CY0F
    );
  ramdatai_s_6_CYSELF_3404 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z501,
      O => ramdatai_s_6_CYSELF
    );
  ramdatai_s_6_DYMUX_3405 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_6_GYMUX,
      O => ramdatai_s_6_DYMUX
    );
  ramdatai_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_6_GYMUX,
      O => U_DCT1D_rtlc5n2653
    );
  ramdatai_s_6_GYMUX_3406 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_6_XORG,
      O => ramdatai_s_6_GYMUX
    );
  ramdatai_s_6_XORG_3407 : X_XOR2
    port map (
      I0 => U_DCT1D_ix59700z64016_O,
      I1 => U_DCT1D_nx59700z498,
      O => ramdatai_s_6_XORG
    );
  ramdatai_s_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_6_CYMUXFAST,
      O => U_DCT1D_ix59700z64012_O
    );
  ramdatai_s_6_FASTCARRY_3408 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z64020_O,
      O => ramdatai_s_6_FASTCARRY
    );
  ramdatai_s_6_CYAND_3409 : X_AND2
    port map (
      I0 => ramdatai_s_6_CYSELG,
      I1 => ramdatai_s_6_CYSELF,
      O => ramdatai_s_6_CYAND
    );
  ramdatai_s_6_CYMUXFAST_3410 : X_MUX2
    port map (
      IA => ramdatai_s_6_CYMUXG2,
      IB => ramdatai_s_6_FASTCARRY,
      SEL => ramdatai_s_6_CYAND,
      O => ramdatai_s_6_CYMUXFAST
    );
  ramdatai_s_6_CYMUXG2_3411 : X_MUX2
    port map (
      IA => ramdatai_s_6_CY0G,
      IB => ramdatai_s_6_CYMUXF2,
      SEL => ramdatai_s_6_CYSELG,
      O => ramdatai_s_6_CYMUXG2
    );
  ramdatai_s_6_CY0G_3412 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(19),
      O => ramdatai_s_6_CY0G
    );
  ramdatai_s_6_CYSELG_3413 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z498,
      O => ramdatai_s_6_CYSELG
    );
  ramdatai_s_6_SRINV_3414 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramdatai_s_6_SRINV
    );
  ramdatai_s_6_CLKINV_3415 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramdatai_s_6_CLKINV
    );
  ramdatai_s_6_CEINV_3416 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => ramdatai_s_6_CEINV
    );
  U_DCT1D_nx59700z1_rt_3417 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z1_rt
    );
  ramdatai_s_8_DXMUX_3418 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_8_FXMUX,
      O => ramdatai_s_8_DXMUX
    );
  ramdatai_s_8_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_8_FXMUX,
      O => U_DCT1D_rtlc5n2652
    );
  ramdatai_s_8_FXMUX_3419 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_8_XORF,
      O => ramdatai_s_8_FXMUX
    );
  ramdatai_s_8_XORF_3420 : X_XOR2
    port map (
      I0 => ramdatai_s_8_CYINIT,
      I1 => U_DCT1D_nx59700z495,
      O => ramdatai_s_8_XORF
    );
  ramdatai_s_8_CYMUXF : X_MUX2
    port map (
      IA => ramdatai_s_8_CY0F,
      IB => ramdatai_s_8_CYINIT,
      SEL => ramdatai_s_8_CYSELF,
      O => U_DCT1D_ix59700z64007_O
    );
  ramdatai_s_8_CYINIT_3421 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z64012_O,
      O => ramdatai_s_8_CYINIT
    );
  ramdatai_s_8_CY0F_3422 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1350(20),
      O => ramdatai_s_8_CY0F
    );
  ramdatai_s_8_CYSELF_3423 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z495,
      O => ramdatai_s_8_CYSELF
    );
  ramdatai_s_8_DYMUX_3424 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_8_GYMUX,
      O => ramdatai_s_8_DYMUX
    );
  ramdatai_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_8_GYMUX,
      O => U_DCT1D_rtlc5n2651
    );
  ramdatai_s_8_GYMUX_3425 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_s_8_XORG,
      O => ramdatai_s_8_GYMUX
    );
  ramdatai_s_8_XORG_3426 : X_XOR2
    port map (
      I0 => U_DCT1D_ix59700z64007_O,
      I1 => U_DCT1D_nx59700z1_rt,
      O => ramdatai_s_8_XORG
    );
  ramdatai_s_8_SRINV_3427 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramdatai_s_8_SRINV
    );
  ramdatai_s_8_CLKINV_3428 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramdatai_s_8_CLKINV
    );
  ramdatai_s_8_CEINV_3429 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => ramdatai_s_8_CEINV
    );
  U_DCT1D_ix59700z31689 : X_LUT4
    generic map(
      INIT => X"74B8"
    )
    port map (
      ADR0 => romodatao7_s(1),
      ADR1 => U_DCT1D_state_reg(0),
      ADR2 => romedatao6_s(2),
      ADR3 => romodatao6_s(2),
      O => U_DCT1D_nx59700z371
    );
  U_DCT1D_rtlc5n1347_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_7_XORF,
      O => U_DCT1D_rtlc5n1347(7)
    );
  U_DCT1D_rtlc5n1347_7_XORF_3430 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1347_7_CYINIT,
      I1 => U_DCT1D_nx59700z374,
      O => U_DCT1D_rtlc5n1347_7_XORF
    );
  U_DCT1D_rtlc5n1347_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_7_CY0F,
      IB => U_DCT1D_rtlc5n1347_7_CYINIT,
      SEL => U_DCT1D_rtlc5n1347_7_CYSELF,
      O => U_DCT1D_ix59700z63837_O
    );
  U_DCT1D_rtlc5n1347_7_CYINIT_3431 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_7_BXINVNOT,
      O => U_DCT1D_rtlc5n1347_7_CYINIT
    );
  U_DCT1D_rtlc5n1347_7_CY0F_3432 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z375,
      O => U_DCT1D_rtlc5n1347_7_CY0F
    );
  U_DCT1D_rtlc5n1347_7_FAND : X_AND2
    port map (
      I0 => romodatao6_s(1),
      I1 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z375
    );
  U_DCT1D_rtlc5n1347_7_CYSELF_3433 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z374,
      O => U_DCT1D_rtlc5n1347_7_CYSELF
    );
  U_DCT1D_rtlc5n1347_7_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_10,
      O => U_DCT1D_rtlc5n1347_7_BXINVNOT
    );
  U_DCT1D_rtlc5n1347_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_7_XORG,
      O => U_DCT1D_rtlc5n1347(8)
    );
  U_DCT1D_rtlc5n1347_7_XORG_3434 : X_XOR2
    port map (
      I0 => U_DCT1D_ix59700z63837_O,
      I1 => U_DCT1D_nx59700z371,
      O => U_DCT1D_rtlc5n1347_7_XORG
    );
  U_DCT1D_rtlc5n1347_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_7_CYMUXG,
      O => U_DCT1D_ix59700z63834_O
    );
  U_DCT1D_rtlc5n1347_7_CYMUXG_3435 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_7_CY0G,
      IB => U_DCT1D_ix59700z63837_O,
      SEL => U_DCT1D_rtlc5n1347_7_CYSELG,
      O => U_DCT1D_rtlc5n1347_7_CYMUXG
    );
  U_DCT1D_rtlc5n1347_7_CY0G_3436 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z372,
      O => U_DCT1D_rtlc5n1347_7_CY0G
    );
  U_DCT1D_rtlc5n1347_7_GAND : X_AND2
    port map (
      I0 => U_DCT1D_state_reg(0),
      I1 => romodatao7_s(1),
      O => U_DCT1D_nx59700z372
    );
  U_DCT1D_rtlc5n1347_7_CYSELG_3437 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z371,
      O => U_DCT1D_rtlc5n1347_7_CYSELG
    );
  U_DCT2D_ix60819z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_5_1_Q,
      ADR1 => U_DCT2D_latchbuf_reg_2_1_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx60819z1
    );
  U_DCT1D_ix59700z23985 : X_LUT4
    generic map(
      INIT => X"3C66"
    )
    port map (
      ADR0 => romedatao7_s(3),
      ADR1 => U_DCT1D_nx59700z366,
      ADR2 => romodatao7_s(3),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z365
    );
  U_DCT1D_rtlc5n1347_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_9_XORF,
      O => U_DCT1D_rtlc5n1347(9)
    );
  U_DCT1D_rtlc5n1347_9_XORF_3438 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1347_9_CYINIT,
      I1 => U_DCT1D_nx59700z368,
      O => U_DCT1D_rtlc5n1347_9_XORF
    );
  U_DCT1D_rtlc5n1347_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_9_CY0F,
      IB => U_DCT1D_rtlc5n1347_9_CYINIT,
      SEL => U_DCT1D_rtlc5n1347_9_CYSELF,
      O => U_DCT1D_ix59700z63831_O
    );
  U_DCT1D_rtlc5n1347_9_CYMUXF2_3439 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_9_CY0F,
      IB => U_DCT1D_rtlc5n1347_9_CY0F,
      SEL => U_DCT1D_rtlc5n1347_9_CYSELF,
      O => U_DCT1D_rtlc5n1347_9_CYMUXF2
    );
  U_DCT1D_rtlc5n1347_9_CYINIT_3440 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63834_O,
      O => U_DCT1D_rtlc5n1347_9_CYINIT
    );
  U_DCT1D_rtlc5n1347_9_CY0F_3441 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z369,
      O => U_DCT1D_rtlc5n1347_9_CY0F
    );
  U_DCT1D_rtlc5n1347_9_CYSELF_3442 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z368,
      O => U_DCT1D_rtlc5n1347_9_CYSELF
    );
  U_DCT1D_rtlc5n1347_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_9_XORG,
      O => U_DCT1D_rtlc5n1347(10)
    );
  U_DCT1D_rtlc5n1347_9_XORG_3443 : X_XOR2
    port map (
      I0 => U_DCT1D_ix59700z63831_O,
      I1 => U_DCT1D_nx59700z365,
      O => U_DCT1D_rtlc5n1347_9_XORG
    );
  U_DCT1D_rtlc5n1347_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_9_CYMUXFAST,
      O => U_DCT1D_ix59700z63828_O
    );
  U_DCT1D_rtlc5n1347_9_FASTCARRY_3444 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63834_O,
      O => U_DCT1D_rtlc5n1347_9_FASTCARRY
    );
  U_DCT1D_rtlc5n1347_9_CYAND_3445 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1347_9_CYSELG,
      I1 => U_DCT1D_rtlc5n1347_9_CYSELF,
      O => U_DCT1D_rtlc5n1347_9_CYAND
    );
  U_DCT1D_rtlc5n1347_9_CYMUXFAST_3446 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_9_CYMUXG2,
      IB => U_DCT1D_rtlc5n1347_9_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1347_9_CYAND,
      O => U_DCT1D_rtlc5n1347_9_CYMUXFAST
    );
  U_DCT1D_rtlc5n1347_9_CYMUXG2_3447 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_9_CY0G,
      IB => U_DCT1D_rtlc5n1347_9_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1347_9_CYSELG,
      O => U_DCT1D_rtlc5n1347_9_CYMUXG2
    );
  U_DCT1D_rtlc5n1347_9_CY0G_3448 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z366,
      O => U_DCT1D_rtlc5n1347_9_CY0G
    );
  U_DCT1D_rtlc5n1347_9_CYSELG_3449 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z365,
      O => U_DCT1D_rtlc5n1347_9_CYSELG
    );
  U_DCT1D_ix59700z23979 : X_LUT4
    generic map(
      INIT => X"36C6"
    )
    port map (
      ADR0 => romedatao7_s(5),
      ADR1 => U_DCT1D_nx59700z360,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => romodatao7_s(5),
      O => U_DCT1D_nx59700z359
    );
  U_DCT1D_rtlc5n1347_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_11_XORF,
      O => U_DCT1D_rtlc5n1347(11)
    );
  U_DCT1D_rtlc5n1347_11_XORF_3450 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1347_11_CYINIT,
      I1 => U_DCT1D_nx59700z362,
      O => U_DCT1D_rtlc5n1347_11_XORF
    );
  U_DCT1D_rtlc5n1347_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_11_CY0F,
      IB => U_DCT1D_rtlc5n1347_11_CYINIT,
      SEL => U_DCT1D_rtlc5n1347_11_CYSELF,
      O => U_DCT1D_ix59700z63825_O
    );
  U_DCT1D_rtlc5n1347_11_CYMUXF2_3451 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_11_CY0F,
      IB => U_DCT1D_rtlc5n1347_11_CY0F,
      SEL => U_DCT1D_rtlc5n1347_11_CYSELF,
      O => U_DCT1D_rtlc5n1347_11_CYMUXF2
    );
  U_DCT1D_rtlc5n1347_11_CYINIT_3452 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63828_O,
      O => U_DCT1D_rtlc5n1347_11_CYINIT
    );
  U_DCT1D_rtlc5n1347_11_CY0F_3453 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z363,
      O => U_DCT1D_rtlc5n1347_11_CY0F
    );
  U_DCT1D_rtlc5n1347_11_CYSELF_3454 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z362,
      O => U_DCT1D_rtlc5n1347_11_CYSELF
    );
  U_DCT1D_rtlc5n1347_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_11_XORG,
      O => U_DCT1D_rtlc5n1347(12)
    );
  U_DCT1D_rtlc5n1347_11_XORG_3455 : X_XOR2
    port map (
      I0 => U_DCT1D_ix59700z63825_O,
      I1 => U_DCT1D_nx59700z359,
      O => U_DCT1D_rtlc5n1347_11_XORG
    );
  U_DCT1D_rtlc5n1347_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_11_CYMUXFAST,
      O => U_DCT1D_ix59700z63822_O
    );
  U_DCT1D_rtlc5n1347_11_FASTCARRY_3456 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63828_O,
      O => U_DCT1D_rtlc5n1347_11_FASTCARRY
    );
  U_DCT1D_rtlc5n1347_11_CYAND_3457 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1347_11_CYSELG,
      I1 => U_DCT1D_rtlc5n1347_11_CYSELF,
      O => U_DCT1D_rtlc5n1347_11_CYAND
    );
  U_DCT1D_rtlc5n1347_11_CYMUXFAST_3458 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_11_CYMUXG2,
      IB => U_DCT1D_rtlc5n1347_11_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1347_11_CYAND,
      O => U_DCT1D_rtlc5n1347_11_CYMUXFAST
    );
  U_DCT1D_rtlc5n1347_11_CYMUXG2_3459 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_11_CY0G,
      IB => U_DCT1D_rtlc5n1347_11_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1347_11_CYSELG,
      O => U_DCT1D_rtlc5n1347_11_CYMUXG2
    );
  U_DCT1D_rtlc5n1347_11_CY0G_3460 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z360,
      O => U_DCT1D_rtlc5n1347_11_CY0G
    );
  U_DCT1D_rtlc5n1347_11_CYSELG_3461 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z359,
      O => U_DCT1D_rtlc5n1347_11_CYSELG
    );
  U_DCT1D_ix59700z23973 : X_LUT4
    generic map(
      INIT => X"56A6"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z354,
      ADR1 => romedatao7_s(7),
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => romodatao7_s(7),
      O => U_DCT1D_nx59700z353
    );
  U_DCT1D_rtlc5n1347_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_13_XORF,
      O => U_DCT1D_rtlc5n1347(13)
    );
  U_DCT1D_rtlc5n1347_13_XORF_3462 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1347_13_CYINIT,
      I1 => U_DCT1D_nx59700z356,
      O => U_DCT1D_rtlc5n1347_13_XORF
    );
  U_DCT1D_rtlc5n1347_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_13_CY0F,
      IB => U_DCT1D_rtlc5n1347_13_CYINIT,
      SEL => U_DCT1D_rtlc5n1347_13_CYSELF,
      O => U_DCT1D_ix59700z63819_O
    );
  U_DCT1D_rtlc5n1347_13_CYMUXF2_3463 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_13_CY0F,
      IB => U_DCT1D_rtlc5n1347_13_CY0F,
      SEL => U_DCT1D_rtlc5n1347_13_CYSELF,
      O => U_DCT1D_rtlc5n1347_13_CYMUXF2
    );
  U_DCT1D_rtlc5n1347_13_CYINIT_3464 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63822_O,
      O => U_DCT1D_rtlc5n1347_13_CYINIT
    );
  U_DCT1D_rtlc5n1347_13_CY0F_3465 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z357,
      O => U_DCT1D_rtlc5n1347_13_CY0F
    );
  U_DCT1D_rtlc5n1347_13_CYSELF_3466 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z356,
      O => U_DCT1D_rtlc5n1347_13_CYSELF
    );
  U_DCT1D_rtlc5n1347_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_13_XORG,
      O => U_DCT1D_rtlc5n1347(14)
    );
  U_DCT1D_rtlc5n1347_13_XORG_3467 : X_XOR2
    port map (
      I0 => U_DCT1D_ix59700z63819_O,
      I1 => U_DCT1D_nx59700z353,
      O => U_DCT1D_rtlc5n1347_13_XORG
    );
  U_DCT1D_rtlc5n1347_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_13_CYMUXFAST,
      O => U_DCT1D_ix59700z63816_O
    );
  U_DCT1D_rtlc5n1347_13_FASTCARRY_3468 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63822_O,
      O => U_DCT1D_rtlc5n1347_13_FASTCARRY
    );
  U_DCT1D_rtlc5n1347_13_CYAND_3469 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1347_13_CYSELG,
      I1 => U_DCT1D_rtlc5n1347_13_CYSELF,
      O => U_DCT1D_rtlc5n1347_13_CYAND
    );
  U_DCT1D_rtlc5n1347_13_CYMUXFAST_3470 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_13_CYMUXG2,
      IB => U_DCT1D_rtlc5n1347_13_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1347_13_CYAND,
      O => U_DCT1D_rtlc5n1347_13_CYMUXFAST
    );
  U_DCT1D_rtlc5n1347_13_CYMUXG2_3471 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_13_CY0G,
      IB => U_DCT1D_rtlc5n1347_13_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1347_13_CYSELG,
      O => U_DCT1D_rtlc5n1347_13_CYMUXG2
    );
  U_DCT1D_rtlc5n1347_13_CY0G_3472 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z354,
      O => U_DCT1D_rtlc5n1347_13_CY0G
    );
  U_DCT1D_rtlc5n1347_13_CYSELG_3473 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z353,
      O => U_DCT1D_rtlc5n1347_13_CYSELG
    );
  U_DCT1D_ix59700z23967 : X_LUT4
    generic map(
      INIT => X"56A6"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z348,
      ADR1 => romedatao7_s(9),
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => romodatao7_s(9),
      O => U_DCT1D_nx59700z347
    );
  U_DCT1D_rtlc5n1347_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_15_XORF,
      O => U_DCT1D_rtlc5n1347(15)
    );
  U_DCT1D_rtlc5n1347_15_XORF_3474 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1347_15_CYINIT,
      I1 => U_DCT1D_nx59700z350,
      O => U_DCT1D_rtlc5n1347_15_XORF
    );
  U_DCT1D_rtlc5n1347_15_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_15_CY0F,
      IB => U_DCT1D_rtlc5n1347_15_CYINIT,
      SEL => U_DCT1D_rtlc5n1347_15_CYSELF,
      O => U_DCT1D_ix59700z63813_O
    );
  U_DCT1D_rtlc5n1347_15_CYMUXF2_3475 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_15_CY0F,
      IB => U_DCT1D_rtlc5n1347_15_CY0F,
      SEL => U_DCT1D_rtlc5n1347_15_CYSELF,
      O => U_DCT1D_rtlc5n1347_15_CYMUXF2
    );
  U_DCT1D_rtlc5n1347_15_CYINIT_3476 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63816_O,
      O => U_DCT1D_rtlc5n1347_15_CYINIT
    );
  U_DCT1D_rtlc5n1347_15_CY0F_3477 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z351,
      O => U_DCT1D_rtlc5n1347_15_CY0F
    );
  U_DCT1D_rtlc5n1347_15_CYSELF_3478 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z350,
      O => U_DCT1D_rtlc5n1347_15_CYSELF
    );
  U_DCT1D_rtlc5n1347_15_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_15_XORG,
      O => U_DCT1D_rtlc5n1347(16)
    );
  U_DCT1D_rtlc5n1347_15_XORG_3479 : X_XOR2
    port map (
      I0 => U_DCT1D_ix59700z63813_O,
      I1 => U_DCT1D_nx59700z347,
      O => U_DCT1D_rtlc5n1347_15_XORG
    );
  U_DCT1D_rtlc5n1347_15_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_15_CYMUXFAST,
      O => U_DCT1D_ix59700z63810_O
    );
  U_DCT1D_rtlc5n1347_15_FASTCARRY_3480 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63816_O,
      O => U_DCT1D_rtlc5n1347_15_FASTCARRY
    );
  U_DCT1D_rtlc5n1347_15_CYAND_3481 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1347_15_CYSELG,
      I1 => U_DCT1D_rtlc5n1347_15_CYSELF,
      O => U_DCT1D_rtlc5n1347_15_CYAND
    );
  U_DCT1D_rtlc5n1347_15_CYMUXFAST_3482 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_15_CYMUXG2,
      IB => U_DCT1D_rtlc5n1347_15_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1347_15_CYAND,
      O => U_DCT1D_rtlc5n1347_15_CYMUXFAST
    );
  U_DCT1D_rtlc5n1347_15_CYMUXG2_3483 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_15_CY0G,
      IB => U_DCT1D_rtlc5n1347_15_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1347_15_CYSELG,
      O => U_DCT1D_rtlc5n1347_15_CYMUXG2
    );
  U_DCT1D_rtlc5n1347_15_CY0G_3484 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z348,
      O => U_DCT1D_rtlc5n1347_15_CY0G
    );
  U_DCT1D_rtlc5n1347_15_CYSELG_3485 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z347,
      O => U_DCT1D_rtlc5n1347_15_CYSELG
    );
  U_DCT1D_ix59700z23961 : X_LUT4
    generic map(
      INIT => X"56A6"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z342,
      ADR1 => romedatao7_s(11),
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => romodatao7_s(11),
      O => U_DCT1D_nx59700z341
    );
  U_DCT1D_rtlc5n1347_17_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_17_XORF,
      O => U_DCT1D_rtlc5n1347(17)
    );
  U_DCT1D_rtlc5n1347_17_XORF_3486 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1347_17_CYINIT,
      I1 => U_DCT1D_nx59700z344,
      O => U_DCT1D_rtlc5n1347_17_XORF
    );
  U_DCT1D_rtlc5n1347_17_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_17_CY0F,
      IB => U_DCT1D_rtlc5n1347_17_CYINIT,
      SEL => U_DCT1D_rtlc5n1347_17_CYSELF,
      O => U_DCT1D_ix59700z63807_O
    );
  U_DCT1D_rtlc5n1347_17_CYMUXF2_3487 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_17_CY0F,
      IB => U_DCT1D_rtlc5n1347_17_CY0F,
      SEL => U_DCT1D_rtlc5n1347_17_CYSELF,
      O => U_DCT1D_rtlc5n1347_17_CYMUXF2
    );
  U_DCT1D_rtlc5n1347_17_CYINIT_3488 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63810_O,
      O => U_DCT1D_rtlc5n1347_17_CYINIT
    );
  U_DCT1D_rtlc5n1347_17_CY0F_3489 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z345,
      O => U_DCT1D_rtlc5n1347_17_CY0F
    );
  U_DCT1D_rtlc5n1347_17_CYSELF_3490 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z344,
      O => U_DCT1D_rtlc5n1347_17_CYSELF
    );
  U_DCT1D_rtlc5n1347_17_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_17_XORG,
      O => U_DCT1D_rtlc5n1347(18)
    );
  U_DCT1D_rtlc5n1347_17_XORG_3491 : X_XOR2
    port map (
      I0 => U_DCT1D_ix59700z63807_O,
      I1 => U_DCT1D_nx59700z341,
      O => U_DCT1D_rtlc5n1347_17_XORG
    );
  U_DCT1D_rtlc5n1347_17_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_17_CYMUXFAST,
      O => U_DCT1D_ix59700z63804_O
    );
  U_DCT1D_rtlc5n1347_17_FASTCARRY_3492 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63810_O,
      O => U_DCT1D_rtlc5n1347_17_FASTCARRY
    );
  U_DCT1D_rtlc5n1347_17_CYAND_3493 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1347_17_CYSELG,
      I1 => U_DCT1D_rtlc5n1347_17_CYSELF,
      O => U_DCT1D_rtlc5n1347_17_CYAND
    );
  U_DCT1D_rtlc5n1347_17_CYMUXFAST_3494 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_17_CYMUXG2,
      IB => U_DCT1D_rtlc5n1347_17_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1347_17_CYAND,
      O => U_DCT1D_rtlc5n1347_17_CYMUXFAST
    );
  U_DCT1D_rtlc5n1347_17_CYMUXG2_3495 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_17_CY0G,
      IB => U_DCT1D_rtlc5n1347_17_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1347_17_CYSELG,
      O => U_DCT1D_rtlc5n1347_17_CYMUXG2
    );
  U_DCT1D_rtlc5n1347_17_CY0G_3496 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z342,
      O => U_DCT1D_rtlc5n1347_17_CY0G
    );
  U_DCT1D_rtlc5n1347_17_CYSELG_3497 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z341,
      O => U_DCT1D_rtlc5n1347_17_CYSELG
    );
  U_DCT1D_ix59700z23957 : X_LUT4
    generic map(
      INIT => X"3C66"
    )
    port map (
      ADR0 => romedatao7_s(13),
      ADR1 => U_DCT1D_nx59700z335,
      ADR2 => romodatao7_s(13),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z337
    );
  U_DCT1D_rtlc5n1347_19_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_19_XORF,
      O => U_DCT1D_rtlc5n1347(19)
    );
  U_DCT1D_rtlc5n1347_19_XORF_3498 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1347_19_CYINIT,
      I1 => U_DCT1D_nx59700z339,
      O => U_DCT1D_rtlc5n1347_19_XORF
    );
  U_DCT1D_rtlc5n1347_19_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_19_CY0F,
      IB => U_DCT1D_rtlc5n1347_19_CYINIT,
      SEL => U_DCT1D_rtlc5n1347_19_CYSELF,
      O => U_DCT1D_ix59700z63802_O
    );
  U_DCT1D_rtlc5n1347_19_CYMUXF2_3499 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_19_CY0F,
      IB => U_DCT1D_rtlc5n1347_19_CY0F,
      SEL => U_DCT1D_rtlc5n1347_19_CYSELF,
      O => U_DCT1D_rtlc5n1347_19_CYMUXF2
    );
  U_DCT1D_rtlc5n1347_19_CYINIT_3500 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63804_O,
      O => U_DCT1D_rtlc5n1347_19_CYINIT
    );
  U_DCT1D_rtlc5n1347_19_CY0F_3501 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z335,
      O => U_DCT1D_rtlc5n1347_19_CY0F
    );
  U_DCT1D_rtlc5n1347_19_CYSELF_3502 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z339,
      O => U_DCT1D_rtlc5n1347_19_CYSELF
    );
  U_DCT1D_rtlc5n1347_19_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_19_XORG,
      O => U_DCT1D_rtlc5n1347(20)
    );
  U_DCT1D_rtlc5n1347_19_XORG_3503 : X_XOR2
    port map (
      I0 => U_DCT1D_ix59700z63802_O,
      I1 => U_DCT1D_nx59700z337,
      O => U_DCT1D_rtlc5n1347_19_XORG
    );
  U_DCT1D_rtlc5n1347_19_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_19_CYMUXFAST,
      O => U_DCT1D_ix59700z63800_O
    );
  U_DCT1D_rtlc5n1347_19_FASTCARRY_3504 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63804_O,
      O => U_DCT1D_rtlc5n1347_19_FASTCARRY
    );
  U_DCT1D_rtlc5n1347_19_CYAND_3505 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1347_19_CYSELG,
      I1 => U_DCT1D_rtlc5n1347_19_CYSELF,
      O => U_DCT1D_rtlc5n1347_19_CYAND
    );
  U_DCT1D_rtlc5n1347_19_CYMUXFAST_3506 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_19_CYMUXG2,
      IB => U_DCT1D_rtlc5n1347_19_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1347_19_CYAND,
      O => U_DCT1D_rtlc5n1347_19_CYMUXFAST
    );
  U_DCT1D_rtlc5n1347_19_CYMUXG2_3507 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1347_19_CY0G,
      IB => U_DCT1D_rtlc5n1347_19_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1347_19_CYSELG,
      O => U_DCT1D_rtlc5n1347_19_CYMUXG2
    );
  U_DCT1D_rtlc5n1347_19_CY0G_3508 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z335,
      O => U_DCT1D_rtlc5n1347_19_CY0G
    );
  U_DCT1D_rtlc5n1347_19_CYSELG_3509 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z337,
      O => U_DCT1D_rtlc5n1347_19_CYSELG
    );
  U_DCT1D_nx59700z334_rt_3510 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_nx59700z334,
      O => U_DCT1D_nx59700z334_rt
    );
  U_DCT1D_rtlc5n1347_21_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1347_21_XORF,
      O => U_DCT1D_rtlc5n1347(21)
    );
  U_DCT1D_rtlc5n1347_21_XORF_3511 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1347_21_CYINIT,
      I1 => U_DCT1D_nx59700z334_rt,
      O => U_DCT1D_rtlc5n1347_21_XORF
    );
  U_DCT1D_rtlc5n1347_21_CYINIT_3512 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ix59700z63800_O,
      O => U_DCT1D_rtlc5n1347_21_CYINIT
    );
  U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CY0F,
      IB => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYINIT,
      SEL => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYSELF,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63612_O
    );
  U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYINIT_3513 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_BXINVNOT,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYINIT
    );
  U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CY0F_3514 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(2),
      O => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CY0F
    );
  U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYSELF_3515 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z209,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYSELF
    );
  U_DCT1D_rtlc_496_add_22_ix59700z63608_O_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_0,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_BXINVNOT
    );
  U_DCT1D_rtlc_496_add_22_ix59700z63608_O_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYMUXG,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63608_O
    );
  U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYMUXG_3516 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CY0G,
      IB => U_DCT1D_rtlc_496_add_22_ix59700z63612_O,
      SEL => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYSELG,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYMUXG
    );
  U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CY0G_3517 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(3),
      O => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CY0G
    );
  U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYSELG_3518 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z207,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63608_O_CYSELG
    );
  U_DCT1D_rtlc5n1348_4_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_4_XORF,
      O => U_DCT1D_rtlc5n1348(4)
    );
  U_DCT1D_rtlc5n1348_4_XORF_3519 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1348_4_CYINIT,
      I1 => U_DCT1D_nx59700z204,
      O => U_DCT1D_rtlc5n1348_4_XORF
    );
  U_DCT1D_rtlc5n1348_4_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_4_CY0F,
      IB => U_DCT1D_rtlc5n1348_4_CYINIT,
      SEL => U_DCT1D_rtlc5n1348_4_CYSELF,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63603_O
    );
  U_DCT1D_rtlc5n1348_4_CYMUXF2_3520 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_4_CY0F,
      IB => U_DCT1D_rtlc5n1348_4_CY0F,
      SEL => U_DCT1D_rtlc5n1348_4_CYSELF,
      O => U_DCT1D_rtlc5n1348_4_CYMUXF2
    );
  U_DCT1D_rtlc5n1348_4_CYINIT_3521 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63608_O,
      O => U_DCT1D_rtlc5n1348_4_CYINIT
    );
  U_DCT1D_rtlc5n1348_4_CY0F_3522 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(4),
      O => U_DCT1D_rtlc5n1348_4_CY0F
    );
  U_DCT1D_rtlc5n1348_4_CYSELF_3523 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z204,
      O => U_DCT1D_rtlc5n1348_4_CYSELF
    );
  U_DCT1D_rtlc5n1348_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_4_XORG,
      O => U_DCT1D_rtlc5n1348(5)
    );
  U_DCT1D_rtlc5n1348_4_XORG_3524 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_496_add_22_ix59700z63603_O,
      I1 => U_DCT1D_nx59700z201,
      O => U_DCT1D_rtlc5n1348_4_XORG
    );
  U_DCT1D_rtlc5n1348_4_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_4_CYMUXFAST,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63597_O
    );
  U_DCT1D_rtlc5n1348_4_FASTCARRY_3525 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63608_O,
      O => U_DCT1D_rtlc5n1348_4_FASTCARRY
    );
  U_DCT1D_rtlc5n1348_4_CYAND_3526 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1348_4_CYSELG,
      I1 => U_DCT1D_rtlc5n1348_4_CYSELF,
      O => U_DCT1D_rtlc5n1348_4_CYAND
    );
  U_DCT1D_rtlc5n1348_4_CYMUXFAST_3527 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_4_CYMUXG2,
      IB => U_DCT1D_rtlc5n1348_4_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1348_4_CYAND,
      O => U_DCT1D_rtlc5n1348_4_CYMUXFAST
    );
  U_DCT1D_rtlc5n1348_4_CYMUXG2_3528 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_4_CY0G,
      IB => U_DCT1D_rtlc5n1348_4_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1348_4_CYSELG,
      O => U_DCT1D_rtlc5n1348_4_CYMUXG2
    );
  U_DCT1D_rtlc5n1348_4_CY0G_3529 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(5),
      O => U_DCT1D_rtlc5n1348_4_CY0G
    );
  U_DCT1D_rtlc5n1348_4_CYSELG_3530 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z201,
      O => U_DCT1D_rtlc5n1348_4_CYSELG
    );
  U_DCT1D_rtlc5n1348_6_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_6_XORF,
      O => U_DCT1D_rtlc5n1348(6)
    );
  U_DCT1D_rtlc5n1348_6_XORF_3531 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1348_6_CYINIT,
      I1 => U_DCT1D_nx59700z198,
      O => U_DCT1D_rtlc5n1348_6_XORF
    );
  U_DCT1D_rtlc5n1348_6_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_6_CY0F,
      IB => U_DCT1D_rtlc5n1348_6_CYINIT,
      SEL => U_DCT1D_rtlc5n1348_6_CYSELF,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63592_O
    );
  U_DCT1D_rtlc5n1348_6_CYMUXF2_3532 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_6_CY0F,
      IB => U_DCT1D_rtlc5n1348_6_CY0F,
      SEL => U_DCT1D_rtlc5n1348_6_CYSELF,
      O => U_DCT1D_rtlc5n1348_6_CYMUXF2
    );
  U_DCT1D_rtlc5n1348_6_CYINIT_3533 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63597_O,
      O => U_DCT1D_rtlc5n1348_6_CYINIT
    );
  U_DCT1D_rtlc5n1348_6_CY0F_3534 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(6),
      O => U_DCT1D_rtlc5n1348_6_CY0F
    );
  U_DCT1D_rtlc5n1348_6_CYSELF_3535 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z198,
      O => U_DCT1D_rtlc5n1348_6_CYSELF
    );
  U_DCT1D_rtlc5n1348_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_6_XORG,
      O => U_DCT1D_rtlc5n1348(7)
    );
  U_DCT1D_rtlc5n1348_6_XORG_3536 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_496_add_22_ix59700z63592_O,
      I1 => U_DCT1D_nx59700z195,
      O => U_DCT1D_rtlc5n1348_6_XORG
    );
  U_DCT1D_rtlc5n1348_6_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_6_CYMUXFAST,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63587_O
    );
  U_DCT1D_rtlc5n1348_6_FASTCARRY_3537 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63597_O,
      O => U_DCT1D_rtlc5n1348_6_FASTCARRY
    );
  U_DCT1D_rtlc5n1348_6_CYAND_3538 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1348_6_CYSELG,
      I1 => U_DCT1D_rtlc5n1348_6_CYSELF,
      O => U_DCT1D_rtlc5n1348_6_CYAND
    );
  U_DCT1D_rtlc5n1348_6_CYMUXFAST_3539 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_6_CYMUXG2,
      IB => U_DCT1D_rtlc5n1348_6_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1348_6_CYAND,
      O => U_DCT1D_rtlc5n1348_6_CYMUXFAST
    );
  U_DCT1D_rtlc5n1348_6_CYMUXG2_3540 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_6_CY0G,
      IB => U_DCT1D_rtlc5n1348_6_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1348_6_CYSELG,
      O => U_DCT1D_rtlc5n1348_6_CYMUXG2
    );
  U_DCT1D_rtlc5n1348_6_CY0G_3541 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(7),
      O => U_DCT1D_rtlc5n1348_6_CY0G
    );
  U_DCT1D_rtlc5n1348_6_CYSELG_3542 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z195,
      O => U_DCT1D_rtlc5n1348_6_CYSELG
    );
  U_DCT1D_rtlc5n1348_8_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_8_XORF,
      O => U_DCT1D_rtlc5n1348(8)
    );
  U_DCT1D_rtlc5n1348_8_XORF_3543 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1348_8_CYINIT,
      I1 => U_DCT1D_nx59700z192,
      O => U_DCT1D_rtlc5n1348_8_XORF
    );
  U_DCT1D_rtlc5n1348_8_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_8_CY0F,
      IB => U_DCT1D_rtlc5n1348_8_CYINIT,
      SEL => U_DCT1D_rtlc5n1348_8_CYSELF,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63582_O
    );
  U_DCT1D_rtlc5n1348_8_CYMUXF2_3544 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_8_CY0F,
      IB => U_DCT1D_rtlc5n1348_8_CY0F,
      SEL => U_DCT1D_rtlc5n1348_8_CYSELF,
      O => U_DCT1D_rtlc5n1348_8_CYMUXF2
    );
  U_DCT1D_rtlc5n1348_8_CYINIT_3545 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63587_O,
      O => U_DCT1D_rtlc5n1348_8_CYINIT
    );
  U_DCT1D_rtlc5n1348_8_CY0F_3546 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(8),
      O => U_DCT1D_rtlc5n1348_8_CY0F
    );
  U_DCT1D_rtlc5n1348_8_CYSELF_3547 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z192,
      O => U_DCT1D_rtlc5n1348_8_CYSELF
    );
  U_DCT1D_rtlc5n1348_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_8_XORG,
      O => U_DCT1D_rtlc5n1348(9)
    );
  U_DCT1D_rtlc5n1348_8_XORG_3548 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_496_add_22_ix59700z63582_O,
      I1 => U_DCT1D_nx59700z189,
      O => U_DCT1D_rtlc5n1348_8_XORG
    );
  U_DCT1D_rtlc5n1348_8_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_8_CYMUXFAST,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63577_O
    );
  U_DCT1D_rtlc5n1348_8_FASTCARRY_3549 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63587_O,
      O => U_DCT1D_rtlc5n1348_8_FASTCARRY
    );
  U_DCT1D_rtlc5n1348_8_CYAND_3550 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1348_8_CYSELG,
      I1 => U_DCT1D_rtlc5n1348_8_CYSELF,
      O => U_DCT1D_rtlc5n1348_8_CYAND
    );
  U_DCT1D_rtlc5n1348_8_CYMUXFAST_3551 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_8_CYMUXG2,
      IB => U_DCT1D_rtlc5n1348_8_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1348_8_CYAND,
      O => U_DCT1D_rtlc5n1348_8_CYMUXFAST
    );
  U_DCT1D_rtlc5n1348_8_CYMUXG2_3552 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_8_CY0G,
      IB => U_DCT1D_rtlc5n1348_8_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1348_8_CYSELG,
      O => U_DCT1D_rtlc5n1348_8_CYMUXG2
    );
  U_DCT1D_rtlc5n1348_8_CY0G_3553 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(9),
      O => U_DCT1D_rtlc5n1348_8_CY0G
    );
  U_DCT1D_rtlc5n1348_8_CYSELG_3554 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z189,
      O => U_DCT1D_rtlc5n1348_8_CYSELG
    );
  U_DCT1D_rtlc5n1348_10_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_10_XORF,
      O => U_DCT1D_rtlc5n1348(10)
    );
  U_DCT1D_rtlc5n1348_10_XORF_3555 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1348_10_CYINIT,
      I1 => U_DCT1D_nx59700z186,
      O => U_DCT1D_rtlc5n1348_10_XORF
    );
  U_DCT1D_rtlc5n1348_10_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_10_CY0F,
      IB => U_DCT1D_rtlc5n1348_10_CYINIT,
      SEL => U_DCT1D_rtlc5n1348_10_CYSELF,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63572_O
    );
  U_DCT1D_rtlc5n1348_10_CYMUXF2_3556 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_10_CY0F,
      IB => U_DCT1D_rtlc5n1348_10_CY0F,
      SEL => U_DCT1D_rtlc5n1348_10_CYSELF,
      O => U_DCT1D_rtlc5n1348_10_CYMUXF2
    );
  U_DCT1D_rtlc5n1348_10_CYINIT_3557 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63577_O,
      O => U_DCT1D_rtlc5n1348_10_CYINIT
    );
  U_DCT1D_rtlc5n1348_10_CY0F_3558 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(10),
      O => U_DCT1D_rtlc5n1348_10_CY0F
    );
  U_DCT1D_rtlc5n1348_10_CYSELF_3559 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z186,
      O => U_DCT1D_rtlc5n1348_10_CYSELF
    );
  U_DCT1D_rtlc5n1348_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_10_XORG,
      O => U_DCT1D_rtlc5n1348(11)
    );
  U_DCT1D_rtlc5n1348_10_XORG_3560 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_496_add_22_ix59700z63572_O,
      I1 => U_DCT1D_nx59700z183,
      O => U_DCT1D_rtlc5n1348_10_XORG
    );
  U_DCT1D_rtlc5n1348_10_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_10_CYMUXFAST,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63567_O
    );
  U_DCT1D_rtlc5n1348_10_FASTCARRY_3561 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63577_O,
      O => U_DCT1D_rtlc5n1348_10_FASTCARRY
    );
  U_DCT1D_rtlc5n1348_10_CYAND_3562 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1348_10_CYSELG,
      I1 => U_DCT1D_rtlc5n1348_10_CYSELF,
      O => U_DCT1D_rtlc5n1348_10_CYAND
    );
  U_DCT1D_rtlc5n1348_10_CYMUXFAST_3563 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_10_CYMUXG2,
      IB => U_DCT1D_rtlc5n1348_10_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1348_10_CYAND,
      O => U_DCT1D_rtlc5n1348_10_CYMUXFAST
    );
  U_DCT1D_rtlc5n1348_10_CYMUXG2_3564 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_10_CY0G,
      IB => U_DCT1D_rtlc5n1348_10_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1348_10_CYSELG,
      O => U_DCT1D_rtlc5n1348_10_CYMUXG2
    );
  U_DCT1D_rtlc5n1348_10_CY0G_3565 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(11),
      O => U_DCT1D_rtlc5n1348_10_CY0G
    );
  U_DCT1D_rtlc5n1348_10_CYSELG_3566 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z183,
      O => U_DCT1D_rtlc5n1348_10_CYSELG
    );
  U_DCT1D_rtlc5n1348_12_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_12_XORF,
      O => U_DCT1D_rtlc5n1348(12)
    );
  U_DCT1D_rtlc5n1348_12_XORF_3567 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1348_12_CYINIT,
      I1 => U_DCT1D_nx59700z180,
      O => U_DCT1D_rtlc5n1348_12_XORF
    );
  U_DCT1D_rtlc5n1348_12_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_12_CY0F,
      IB => U_DCT1D_rtlc5n1348_12_CYINIT,
      SEL => U_DCT1D_rtlc5n1348_12_CYSELF,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63561_O
    );
  U_DCT1D_rtlc5n1348_12_CYMUXF2_3568 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_12_CY0F,
      IB => U_DCT1D_rtlc5n1348_12_CY0F,
      SEL => U_DCT1D_rtlc5n1348_12_CYSELF,
      O => U_DCT1D_rtlc5n1348_12_CYMUXF2
    );
  U_DCT1D_rtlc5n1348_12_CYINIT_3569 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63567_O,
      O => U_DCT1D_rtlc5n1348_12_CYINIT
    );
  U_DCT1D_rtlc5n1348_12_CY0F_3570 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(12),
      O => U_DCT1D_rtlc5n1348_12_CY0F
    );
  U_DCT1D_rtlc5n1348_12_CYSELF_3571 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z180,
      O => U_DCT1D_rtlc5n1348_12_CYSELF
    );
  U_DCT1D_rtlc5n1348_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_12_XORG,
      O => U_DCT1D_rtlc5n1348(13)
    );
  U_DCT1D_rtlc5n1348_12_XORG_3572 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_496_add_22_ix59700z63561_O,
      I1 => U_DCT1D_nx59700z177,
      O => U_DCT1D_rtlc5n1348_12_XORG
    );
  U_DCT1D_rtlc5n1348_12_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_12_CYMUXFAST,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63556_O
    );
  U_DCT1D_rtlc5n1348_12_FASTCARRY_3573 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63567_O,
      O => U_DCT1D_rtlc5n1348_12_FASTCARRY
    );
  U_DCT1D_rtlc5n1348_12_CYAND_3574 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1348_12_CYSELG,
      I1 => U_DCT1D_rtlc5n1348_12_CYSELF,
      O => U_DCT1D_rtlc5n1348_12_CYAND
    );
  U_DCT1D_rtlc5n1348_12_CYMUXFAST_3575 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_12_CYMUXG2,
      IB => U_DCT1D_rtlc5n1348_12_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1348_12_CYAND,
      O => U_DCT1D_rtlc5n1348_12_CYMUXFAST
    );
  U_DCT1D_rtlc5n1348_12_CYMUXG2_3576 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_12_CY0G,
      IB => U_DCT1D_rtlc5n1348_12_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1348_12_CYSELG,
      O => U_DCT1D_rtlc5n1348_12_CYMUXG2
    );
  U_DCT1D_rtlc5n1348_12_CY0G_3577 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(13),
      O => U_DCT1D_rtlc5n1348_12_CY0G
    );
  U_DCT1D_rtlc5n1348_12_CYSELG_3578 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z177,
      O => U_DCT1D_rtlc5n1348_12_CYSELG
    );
  U_DCT1D_rtlc5n1348_14_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_14_XORF,
      O => U_DCT1D_rtlc5n1348(14)
    );
  U_DCT1D_rtlc5n1348_14_XORF_3579 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1348_14_CYINIT,
      I1 => U_DCT1D_nx59700z174,
      O => U_DCT1D_rtlc5n1348_14_XORF
    );
  U_DCT1D_rtlc5n1348_14_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_14_CY0F,
      IB => U_DCT1D_rtlc5n1348_14_CYINIT,
      SEL => U_DCT1D_rtlc5n1348_14_CYSELF,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63551_O
    );
  U_DCT1D_rtlc5n1348_14_CYMUXF2_3580 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_14_CY0F,
      IB => U_DCT1D_rtlc5n1348_14_CY0F,
      SEL => U_DCT1D_rtlc5n1348_14_CYSELF,
      O => U_DCT1D_rtlc5n1348_14_CYMUXF2
    );
  U_DCT1D_rtlc5n1348_14_CYINIT_3581 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63556_O,
      O => U_DCT1D_rtlc5n1348_14_CYINIT
    );
  U_DCT1D_rtlc5n1348_14_CY0F_3582 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(14),
      O => U_DCT1D_rtlc5n1348_14_CY0F
    );
  U_DCT1D_rtlc5n1348_14_CYSELF_3583 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z174,
      O => U_DCT1D_rtlc5n1348_14_CYSELF
    );
  U_DCT1D_rtlc5n1348_14_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_14_XORG,
      O => U_DCT1D_rtlc5n1348(15)
    );
  U_DCT1D_rtlc5n1348_14_XORG_3584 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_496_add_22_ix59700z63551_O,
      I1 => U_DCT1D_nx59700z171,
      O => U_DCT1D_rtlc5n1348_14_XORG
    );
  U_DCT1D_rtlc5n1348_14_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_14_CYMUXFAST,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63546_O
    );
  U_DCT1D_rtlc5n1348_14_FASTCARRY_3585 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63556_O,
      O => U_DCT1D_rtlc5n1348_14_FASTCARRY
    );
  U_DCT1D_rtlc5n1348_14_CYAND_3586 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1348_14_CYSELG,
      I1 => U_DCT1D_rtlc5n1348_14_CYSELF,
      O => U_DCT1D_rtlc5n1348_14_CYAND
    );
  U_DCT1D_rtlc5n1348_14_CYMUXFAST_3587 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_14_CYMUXG2,
      IB => U_DCT1D_rtlc5n1348_14_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1348_14_CYAND,
      O => U_DCT1D_rtlc5n1348_14_CYMUXFAST
    );
  U_DCT1D_rtlc5n1348_14_CYMUXG2_3588 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_14_CY0G,
      IB => U_DCT1D_rtlc5n1348_14_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1348_14_CYSELG,
      O => U_DCT1D_rtlc5n1348_14_CYMUXG2
    );
  U_DCT1D_rtlc5n1348_14_CY0G_3589 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(15),
      O => U_DCT1D_rtlc5n1348_14_CY0G
    );
  U_DCT1D_rtlc5n1348_14_CYSELG_3590 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z171,
      O => U_DCT1D_rtlc5n1348_14_CYSELG
    );
  U_DCT1D_rtlc5n1348_16_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_16_XORF,
      O => U_DCT1D_rtlc5n1348(16)
    );
  U_DCT1D_rtlc5n1348_16_XORF_3591 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1348_16_CYINIT,
      I1 => U_DCT1D_nx59700z168,
      O => U_DCT1D_rtlc5n1348_16_XORF
    );
  U_DCT1D_rtlc5n1348_16_CYMUXF : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_16_CY0F,
      IB => U_DCT1D_rtlc5n1348_16_CYINIT,
      SEL => U_DCT1D_rtlc5n1348_16_CYSELF,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63542_O
    );
  U_DCT1D_rtlc5n1348_16_CYMUXF2_3592 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_16_CY0F,
      IB => U_DCT1D_rtlc5n1348_16_CY0F,
      SEL => U_DCT1D_rtlc5n1348_16_CYSELF,
      O => U_DCT1D_rtlc5n1348_16_CYMUXF2
    );
  U_DCT1D_rtlc5n1348_16_CYINIT_3593 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63546_O,
      O => U_DCT1D_rtlc5n1348_16_CYINIT
    );
  U_DCT1D_rtlc5n1348_16_CY0F_3594 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(15),
      O => U_DCT1D_rtlc5n1348_16_CY0F
    );
  U_DCT1D_rtlc5n1348_16_CYSELF_3595 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z168,
      O => U_DCT1D_rtlc5n1348_16_CYSELF
    );
  U_DCT1D_rtlc5n1348_16_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_16_XORG,
      O => U_DCT1D_rtlc5n1348(17)
    );
  U_DCT1D_rtlc5n1348_16_XORG_3596 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc_496_add_22_ix59700z63542_O,
      I1 => U_DCT1D_nx59700z165,
      O => U_DCT1D_rtlc5n1348_16_XORG
    );
  U_DCT1D_rtlc5n1348_16_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_16_CYMUXFAST,
      O => U_DCT1D_rtlc_496_add_22_ix59700z63538_O
    );
  U_DCT1D_rtlc5n1348_16_FASTCARRY_3597 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63546_O,
      O => U_DCT1D_rtlc5n1348_16_FASTCARRY
    );
  U_DCT1D_rtlc5n1348_16_CYAND_3598 : X_AND2
    port map (
      I0 => U_DCT1D_rtlc5n1348_16_CYSELG,
      I1 => U_DCT1D_rtlc5n1348_16_CYSELF,
      O => U_DCT1D_rtlc5n1348_16_CYAND
    );
  U_DCT1D_rtlc5n1348_16_CYMUXFAST_3599 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_16_CYMUXG2,
      IB => U_DCT1D_rtlc5n1348_16_FASTCARRY,
      SEL => U_DCT1D_rtlc5n1348_16_CYAND,
      O => U_DCT1D_rtlc5n1348_16_CYMUXFAST
    );
  U_DCT1D_rtlc5n1348_16_CYMUXG2_3600 : X_MUX2
    port map (
      IA => U_DCT1D_rtlc5n1348_16_CY0G,
      IB => U_DCT1D_rtlc5n1348_16_CYMUXF2,
      SEL => U_DCT1D_rtlc5n1348_16_CYSELG,
      O => U_DCT1D_rtlc5n1348_16_CYMUXG2
    );
  U_DCT1D_rtlc5n1348_16_CY0G_3601 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1344(15),
      O => U_DCT1D_rtlc5n1348_16_CY0G
    );
  U_DCT1D_rtlc5n1348_16_CYSELG_3602 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z165,
      O => U_DCT1D_rtlc5n1348_16_CYSELG
    );
  U_DCT1D_rtlc5n1348_18_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1348_18_XORF,
      O => U_DCT1D_rtlc5n1348(18)
    );
  U_DCT1D_rtlc5n1348_18_XORF_3603 : X_XOR2
    port map (
      I0 => U_DCT1D_rtlc5n1348_18_CYINIT,
      I1 => U_DCT1D_nx59700z78_rt,
      O => U_DCT1D_rtlc5n1348_18_XORF
    );
  U_DCT1D_rtlc5n1348_18_CYINIT_3604 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc_496_add_22_ix59700z63538_O,
      O => U_DCT1D_rtlc5n1348_18_CYINIT
    );
  U_DCT2D_rtlc5n1482_5_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_5_XORF,
      O => U_DCT2D_rtlc5n1482(5)
    );
  U_DCT2D_rtlc5n1482_5_XORF_3605 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1482_5_CYINIT,
      I1 => U_DCT2D_nx65206z454,
      O => U_DCT2D_rtlc5n1482_5_XORF
    );
  U_DCT2D_rtlc5n1482_5_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_5_CY0F,
      IB => U_DCT2D_rtlc5n1482_5_CYINIT,
      SEL => U_DCT2D_rtlc5n1482_5_CYSELF,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63963_O
    );
  U_DCT2D_rtlc5n1482_5_CYINIT_3606 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_5_BXINVNOT,
      O => U_DCT2D_rtlc5n1482_5_CYINIT
    );
  U_DCT2D_rtlc5n1482_5_CY0F_3607 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(1),
      O => U_DCT2D_rtlc5n1482_5_CY0F
    );
  U_DCT2D_rtlc5n1482_5_CYSELF_3608 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z454,
      O => U_DCT2D_rtlc5n1482_5_CYSELF
    );
  U_DCT2D_rtlc5n1482_5_BXINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_24,
      O => U_DCT2D_rtlc5n1482_5_BXINVNOT
    );
  U_DCT2D_rtlc5n1482_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_5_XORG,
      O => U_DCT2D_rtlc5n1482(6)
    );
  U_DCT2D_rtlc5n1482_5_XORG_3609 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_338_add_57_ix65206z63963_O,
      I1 => U_DCT2D_nx65206z451,
      O => U_DCT2D_rtlc5n1482_5_XORG
    );
  U_DCT2D_rtlc5n1482_5_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_5_CYMUXG,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63959_O
    );
  U_DCT2D_rtlc5n1482_5_CYMUXG_3610 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_5_CY0G,
      IB => U_DCT2D_rtlc_338_add_57_ix65206z63963_O,
      SEL => U_DCT2D_rtlc5n1482_5_CYSELG,
      O => U_DCT2D_rtlc5n1482_5_CYMUXG
    );
  U_DCT2D_rtlc5n1482_5_CY0G_3611 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(2),
      O => U_DCT2D_rtlc5n1482_5_CY0G
    );
  U_DCT2D_rtlc5n1482_5_CYSELG_3612 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z451,
      O => U_DCT2D_rtlc5n1482_5_CYSELG
    );
  U_DCT2D_rtlc5n1482_7_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_7_XORF,
      O => U_DCT2D_rtlc5n1482(7)
    );
  U_DCT2D_rtlc5n1482_7_XORF_3613 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1482_7_CYINIT,
      I1 => U_DCT2D_nx65206z448,
      O => U_DCT2D_rtlc5n1482_7_XORF
    );
  U_DCT2D_rtlc5n1482_7_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_7_CY0F,
      IB => U_DCT2D_rtlc5n1482_7_CYINIT,
      SEL => U_DCT2D_rtlc5n1482_7_CYSELF,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63956_O
    );
  U_DCT2D_rtlc5n1482_7_CYMUXF2_3614 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_7_CY0F,
      IB => U_DCT2D_rtlc5n1482_7_CY0F,
      SEL => U_DCT2D_rtlc5n1482_7_CYSELF,
      O => U_DCT2D_rtlc5n1482_7_CYMUXF2
    );
  U_DCT2D_rtlc5n1482_7_CYINIT_3615 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63959_O,
      O => U_DCT2D_rtlc5n1482_7_CYINIT
    );
  U_DCT2D_rtlc5n1482_7_CY0F_3616 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(3),
      O => U_DCT2D_rtlc5n1482_7_CY0F
    );
  U_DCT2D_rtlc5n1482_7_CYSELF_3617 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z448,
      O => U_DCT2D_rtlc5n1482_7_CYSELF
    );
  U_DCT2D_rtlc5n1482_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_7_XORG,
      O => U_DCT2D_rtlc5n1482(8)
    );
  U_DCT2D_rtlc5n1482_7_XORG_3618 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_338_add_57_ix65206z63956_O,
      I1 => U_DCT2D_nx65206z445,
      O => U_DCT2D_rtlc5n1482_7_XORG
    );
  U_DCT2D_rtlc5n1482_7_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_7_CYMUXFAST,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63952_O
    );
  U_DCT2D_rtlc5n1482_7_FASTCARRY_3619 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63959_O,
      O => U_DCT2D_rtlc5n1482_7_FASTCARRY
    );
  U_DCT2D_rtlc5n1482_7_CYAND_3620 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1482_7_CYSELG,
      I1 => U_DCT2D_rtlc5n1482_7_CYSELF,
      O => U_DCT2D_rtlc5n1482_7_CYAND
    );
  U_DCT2D_rtlc5n1482_7_CYMUXFAST_3621 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_7_CYMUXG2,
      IB => U_DCT2D_rtlc5n1482_7_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1482_7_CYAND,
      O => U_DCT2D_rtlc5n1482_7_CYMUXFAST
    );
  U_DCT2D_rtlc5n1482_7_CYMUXG2_3622 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_7_CY0G,
      IB => U_DCT2D_rtlc5n1482_7_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1482_7_CYSELG,
      O => U_DCT2D_rtlc5n1482_7_CYMUXG2
    );
  U_DCT2D_rtlc5n1482_7_CY0G_3623 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(4),
      O => U_DCT2D_rtlc5n1482_7_CY0G
    );
  U_DCT2D_rtlc5n1482_7_CYSELG_3624 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z445,
      O => U_DCT2D_rtlc5n1482_7_CYSELG
    );
  U_DCT2D_rtlc5n1482_9_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_9_XORF,
      O => U_DCT2D_rtlc5n1482(9)
    );
  U_DCT2D_rtlc5n1482_9_XORF_3625 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1482_9_CYINIT,
      I1 => U_DCT2D_nx65206z442,
      O => U_DCT2D_rtlc5n1482_9_XORF
    );
  U_DCT2D_rtlc5n1482_9_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_9_CY0F,
      IB => U_DCT2D_rtlc5n1482_9_CYINIT,
      SEL => U_DCT2D_rtlc5n1482_9_CYSELF,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63949_O
    );
  U_DCT2D_rtlc5n1482_9_CYMUXF2_3626 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_9_CY0F,
      IB => U_DCT2D_rtlc5n1482_9_CY0F,
      SEL => U_DCT2D_rtlc5n1482_9_CYSELF,
      O => U_DCT2D_rtlc5n1482_9_CYMUXF2
    );
  U_DCT2D_rtlc5n1482_9_CYINIT_3627 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63952_O,
      O => U_DCT2D_rtlc5n1482_9_CYINIT
    );
  U_DCT2D_rtlc5n1482_9_CY0F_3628 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(5),
      O => U_DCT2D_rtlc5n1482_9_CY0F
    );
  U_DCT2D_rtlc5n1482_9_CYSELF_3629 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z442,
      O => U_DCT2D_rtlc5n1482_9_CYSELF
    );
  U_DCT2D_rtlc5n1482_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_9_XORG,
      O => U_DCT2D_rtlc5n1482(10)
    );
  U_DCT2D_rtlc5n1482_9_XORG_3630 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_338_add_57_ix65206z63949_O,
      I1 => U_DCT2D_nx65206z439,
      O => U_DCT2D_rtlc5n1482_9_XORG
    );
  U_DCT2D_rtlc5n1482_9_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_9_CYMUXFAST,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63945_O
    );
  U_DCT2D_rtlc5n1482_9_FASTCARRY_3631 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63952_O,
      O => U_DCT2D_rtlc5n1482_9_FASTCARRY
    );
  U_DCT2D_rtlc5n1482_9_CYAND_3632 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1482_9_CYSELG,
      I1 => U_DCT2D_rtlc5n1482_9_CYSELF,
      O => U_DCT2D_rtlc5n1482_9_CYAND
    );
  U_DCT2D_rtlc5n1482_9_CYMUXFAST_3633 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_9_CYMUXG2,
      IB => U_DCT2D_rtlc5n1482_9_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1482_9_CYAND,
      O => U_DCT2D_rtlc5n1482_9_CYMUXFAST
    );
  U_DCT2D_rtlc5n1482_9_CYMUXG2_3634 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_9_CY0G,
      IB => U_DCT2D_rtlc5n1482_9_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1482_9_CYSELG,
      O => U_DCT2D_rtlc5n1482_9_CYMUXG2
    );
  U_DCT2D_rtlc5n1482_9_CY0G_3635 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(6),
      O => U_DCT2D_rtlc5n1482_9_CY0G
    );
  U_DCT2D_rtlc5n1482_9_CYSELG_3636 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z439,
      O => U_DCT2D_rtlc5n1482_9_CYSELG
    );
  U_DCT2D_rtlc5n1482_11_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_11_XORF,
      O => U_DCT2D_rtlc5n1482(11)
    );
  U_DCT2D_rtlc5n1482_11_XORF_3637 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1482_11_CYINIT,
      I1 => U_DCT2D_nx65206z436,
      O => U_DCT2D_rtlc5n1482_11_XORF
    );
  U_DCT2D_rtlc5n1482_11_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_11_CY0F,
      IB => U_DCT2D_rtlc5n1482_11_CYINIT,
      SEL => U_DCT2D_rtlc5n1482_11_CYSELF,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63942_O
    );
  U_DCT2D_rtlc5n1482_11_CYMUXF2_3638 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_11_CY0F,
      IB => U_DCT2D_rtlc5n1482_11_CY0F,
      SEL => U_DCT2D_rtlc5n1482_11_CYSELF,
      O => U_DCT2D_rtlc5n1482_11_CYMUXF2
    );
  U_DCT2D_rtlc5n1482_11_CYINIT_3639 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63945_O,
      O => U_DCT2D_rtlc5n1482_11_CYINIT
    );
  U_DCT2D_rtlc5n1482_11_CY0F_3640 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(7),
      O => U_DCT2D_rtlc5n1482_11_CY0F
    );
  U_DCT2D_rtlc5n1482_11_CYSELF_3641 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z436,
      O => U_DCT2D_rtlc5n1482_11_CYSELF
    );
  U_DCT2D_rtlc5n1482_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_11_XORG,
      O => U_DCT2D_rtlc5n1482(12)
    );
  U_DCT2D_rtlc5n1482_11_XORG_3642 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_338_add_57_ix65206z63942_O,
      I1 => U_DCT2D_nx65206z433,
      O => U_DCT2D_rtlc5n1482_11_XORG
    );
  U_DCT2D_rtlc5n1482_11_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_11_CYMUXFAST,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63938_O
    );
  U_DCT2D_rtlc5n1482_11_FASTCARRY_3643 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63945_O,
      O => U_DCT2D_rtlc5n1482_11_FASTCARRY
    );
  U_DCT2D_rtlc5n1482_11_CYAND_3644 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1482_11_CYSELG,
      I1 => U_DCT2D_rtlc5n1482_11_CYSELF,
      O => U_DCT2D_rtlc5n1482_11_CYAND
    );
  U_DCT2D_rtlc5n1482_11_CYMUXFAST_3645 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_11_CYMUXG2,
      IB => U_DCT2D_rtlc5n1482_11_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1482_11_CYAND,
      O => U_DCT2D_rtlc5n1482_11_CYMUXFAST
    );
  U_DCT2D_rtlc5n1482_11_CYMUXG2_3646 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_11_CY0G,
      IB => U_DCT2D_rtlc5n1482_11_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1482_11_CYSELG,
      O => U_DCT2D_rtlc5n1482_11_CYMUXG2
    );
  U_DCT2D_rtlc5n1482_11_CY0G_3647 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(8),
      O => U_DCT2D_rtlc5n1482_11_CY0G
    );
  U_DCT2D_rtlc5n1482_11_CYSELG_3648 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z433,
      O => U_DCT2D_rtlc5n1482_11_CYSELG
    );
  U_DCT2D_reg_databuf_reg_2_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_2_0_DYMUX,
      CE => U_DCT2D_databuf_reg_2_0_CEINV,
      CLK => U_DCT2D_databuf_reg_2_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_2_0_FFY_RST,
      O => U_DCT2D_databuf_reg_2_Q(1)
    );
  U_DCT2D_databuf_reg_2_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_2_0_FFY_RST
    );
  U_DCT2D_rtlc5n1482_13_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_13_XORF,
      O => U_DCT2D_rtlc5n1482(13)
    );
  U_DCT2D_rtlc5n1482_13_XORF_3649 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1482_13_CYINIT,
      I1 => U_DCT2D_nx65206z430,
      O => U_DCT2D_rtlc5n1482_13_XORF
    );
  U_DCT2D_rtlc5n1482_13_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_13_CY0F,
      IB => U_DCT2D_rtlc5n1482_13_CYINIT,
      SEL => U_DCT2D_rtlc5n1482_13_CYSELF,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63935_O
    );
  U_DCT2D_rtlc5n1482_13_CYMUXF2_3650 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_13_CY0F,
      IB => U_DCT2D_rtlc5n1482_13_CY0F,
      SEL => U_DCT2D_rtlc5n1482_13_CYSELF,
      O => U_DCT2D_rtlc5n1482_13_CYMUXF2
    );
  U_DCT2D_rtlc5n1482_13_CYINIT_3651 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63938_O,
      O => U_DCT2D_rtlc5n1482_13_CYINIT
    );
  U_DCT2D_rtlc5n1482_13_CY0F_3652 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(9),
      O => U_DCT2D_rtlc5n1482_13_CY0F
    );
  U_DCT2D_rtlc5n1482_13_CYSELF_3653 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z430,
      O => U_DCT2D_rtlc5n1482_13_CYSELF
    );
  U_DCT2D_rtlc5n1482_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_13_XORG,
      O => U_DCT2D_rtlc5n1482(14)
    );
  U_DCT2D_rtlc5n1482_13_XORG_3654 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_338_add_57_ix65206z63935_O,
      I1 => U_DCT2D_nx65206z427,
      O => U_DCT2D_rtlc5n1482_13_XORG
    );
  U_DCT2D_rtlc5n1482_13_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_13_CYMUXFAST,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63931_O
    );
  U_DCT2D_rtlc5n1482_13_FASTCARRY_3655 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63938_O,
      O => U_DCT2D_rtlc5n1482_13_FASTCARRY
    );
  U_DCT2D_rtlc5n1482_13_CYAND_3656 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1482_13_CYSELG,
      I1 => U_DCT2D_rtlc5n1482_13_CYSELF,
      O => U_DCT2D_rtlc5n1482_13_CYAND
    );
  U_DCT2D_rtlc5n1482_13_CYMUXFAST_3657 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_13_CYMUXG2,
      IB => U_DCT2D_rtlc5n1482_13_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1482_13_CYAND,
      O => U_DCT2D_rtlc5n1482_13_CYMUXFAST
    );
  U_DCT2D_rtlc5n1482_13_CYMUXG2_3658 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_13_CY0G,
      IB => U_DCT2D_rtlc5n1482_13_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1482_13_CYSELG,
      O => U_DCT2D_rtlc5n1482_13_CYMUXG2
    );
  U_DCT2D_rtlc5n1482_13_CY0G_3659 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(10),
      O => U_DCT2D_rtlc5n1482_13_CY0G
    );
  U_DCT2D_rtlc5n1482_13_CYSELG_3660 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z427,
      O => U_DCT2D_rtlc5n1482_13_CYSELG
    );
  U_DCT2D_rtlc5n1482_15_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_15_XORF,
      O => U_DCT2D_rtlc5n1482(15)
    );
  U_DCT2D_rtlc5n1482_15_XORF_3661 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1482_15_CYINIT,
      I1 => U_DCT2D_nx65206z424,
      O => U_DCT2D_rtlc5n1482_15_XORF
    );
  U_DCT2D_rtlc5n1482_15_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_15_CY0F,
      IB => U_DCT2D_rtlc5n1482_15_CYINIT,
      SEL => U_DCT2D_rtlc5n1482_15_CYSELF,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63928_O
    );
  U_DCT2D_rtlc5n1482_15_CYMUXF2_3662 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_15_CY0F,
      IB => U_DCT2D_rtlc5n1482_15_CY0F,
      SEL => U_DCT2D_rtlc5n1482_15_CYSELF,
      O => U_DCT2D_rtlc5n1482_15_CYMUXF2
    );
  U_DCT2D_rtlc5n1482_15_CYINIT_3663 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63931_O,
      O => U_DCT2D_rtlc5n1482_15_CYINIT
    );
  U_DCT2D_rtlc5n1482_15_CY0F_3664 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(11),
      O => U_DCT2D_rtlc5n1482_15_CY0F
    );
  U_DCT2D_rtlc5n1482_15_CYSELF_3665 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z424,
      O => U_DCT2D_rtlc5n1482_15_CYSELF
    );
  U_DCT2D_rtlc5n1482_15_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_15_XORG,
      O => U_DCT2D_rtlc5n1482(16)
    );
  U_DCT2D_rtlc5n1482_15_XORG_3666 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_338_add_57_ix65206z63928_O,
      I1 => U_DCT2D_nx65206z421,
      O => U_DCT2D_rtlc5n1482_15_XORG
    );
  U_DCT2D_rtlc5n1482_15_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_15_CYMUXFAST,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63924_O
    );
  U_DCT2D_rtlc5n1482_15_FASTCARRY_3667 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63931_O,
      O => U_DCT2D_rtlc5n1482_15_FASTCARRY
    );
  U_DCT2D_rtlc5n1482_15_CYAND_3668 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1482_15_CYSELG,
      I1 => U_DCT2D_rtlc5n1482_15_CYSELF,
      O => U_DCT2D_rtlc5n1482_15_CYAND
    );
  U_DCT2D_rtlc5n1482_15_CYMUXFAST_3669 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_15_CYMUXG2,
      IB => U_DCT2D_rtlc5n1482_15_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1482_15_CYAND,
      O => U_DCT2D_rtlc5n1482_15_CYMUXFAST
    );
  U_DCT2D_rtlc5n1482_15_CYMUXG2_3670 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_15_CY0G,
      IB => U_DCT2D_rtlc5n1482_15_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1482_15_CYSELG,
      O => U_DCT2D_rtlc5n1482_15_CYMUXG2
    );
  U_DCT2D_rtlc5n1482_15_CY0G_3671 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(12),
      O => U_DCT2D_rtlc5n1482_15_CY0G
    );
  U_DCT2D_rtlc5n1482_15_CYSELG_3672 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z421,
      O => U_DCT2D_rtlc5n1482_15_CYSELG
    );
  U_DCT2D_rtlc5n1482_17_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_17_XORF,
      O => U_DCT2D_rtlc5n1482(17)
    );
  U_DCT2D_rtlc5n1482_17_XORF_3673 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1482_17_CYINIT,
      I1 => U_DCT2D_nx65206z418,
      O => U_DCT2D_rtlc5n1482_17_XORF
    );
  U_DCT2D_rtlc5n1482_17_CYMUXF : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_17_CY0F,
      IB => U_DCT2D_rtlc5n1482_17_CYINIT,
      SEL => U_DCT2D_rtlc5n1482_17_CYSELF,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63921_O
    );
  U_DCT2D_rtlc5n1482_17_CYMUXF2_3674 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_17_CY0F,
      IB => U_DCT2D_rtlc5n1482_17_CY0F,
      SEL => U_DCT2D_rtlc5n1482_17_CYSELF,
      O => U_DCT2D_rtlc5n1482_17_CYMUXF2
    );
  U_DCT2D_rtlc5n1482_17_CYINIT_3675 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63924_O,
      O => U_DCT2D_rtlc5n1482_17_CYINIT
    );
  U_DCT2D_rtlc5n1482_17_CY0F_3676 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(13),
      O => U_DCT2D_rtlc5n1482_17_CY0F
    );
  U_DCT2D_rtlc5n1482_17_CYSELF_3677 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z418,
      O => U_DCT2D_rtlc5n1482_17_CYSELF
    );
  U_DCT2D_rtlc5n1482_17_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_17_XORG,
      O => U_DCT2D_rtlc5n1482(18)
    );
  U_DCT2D_rtlc5n1482_17_XORG_3678 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc_338_add_57_ix65206z63921_O,
      I1 => U_DCT2D_nx65206z415,
      O => U_DCT2D_rtlc5n1482_17_XORG
    );
  U_DCT2D_rtlc5n1482_17_COUTUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_17_CYMUXFAST,
      O => U_DCT2D_rtlc_338_add_57_ix65206z63917_O
    );
  U_DCT2D_rtlc5n1482_17_FASTCARRY_3679 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63924_O,
      O => U_DCT2D_rtlc5n1482_17_FASTCARRY
    );
  U_DCT2D_rtlc5n1482_17_CYAND_3680 : X_AND2
    port map (
      I0 => U_DCT2D_rtlc5n1482_17_CYSELG,
      I1 => U_DCT2D_rtlc5n1482_17_CYSELF,
      O => U_DCT2D_rtlc5n1482_17_CYAND
    );
  U_DCT2D_rtlc5n1482_17_CYMUXFAST_3681 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_17_CYMUXG2,
      IB => U_DCT2D_rtlc5n1482_17_FASTCARRY,
      SEL => U_DCT2D_rtlc5n1482_17_CYAND,
      O => U_DCT2D_rtlc5n1482_17_CYMUXFAST
    );
  U_DCT2D_rtlc5n1482_17_CYMUXG2_3682 : X_MUX2
    port map (
      IA => U_DCT2D_rtlc5n1482_17_CY0G,
      IB => U_DCT2D_rtlc5n1482_17_CYMUXF2,
      SEL => U_DCT2D_rtlc5n1482_17_CYSELG,
      O => U_DCT2D_rtlc5n1482_17_CYMUXG2
    );
  U_DCT2D_rtlc5n1482_17_CY0G_3683 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s(13),
      O => U_DCT2D_rtlc5n1482_17_CY0G
    );
  U_DCT2D_rtlc5n1482_17_CYSELG_3684 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z415,
      O => U_DCT2D_rtlc5n1482_17_CYSELG
    );
  U_DCT2D_nx65206z413_rt_3685 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_nx65206z413,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z413_rt
    );
  U_DCT2D_rtlc5n1482_19_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1482_19_XORF,
      O => U_DCT2D_rtlc5n1482(19)
    );
  U_DCT2D_rtlc5n1482_19_XORF_3686 : X_XOR2
    port map (
      I0 => U_DCT2D_rtlc5n1482_19_CYINIT,
      I1 => U_DCT2D_nx65206z413_rt,
      O => U_DCT2D_rtlc5n1482_19_XORF
    );
  U_DCT2D_rtlc5n1482_19_CYINIT_3687 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc_338_add_57_ix65206z63917_O,
      O => U_DCT2D_rtlc5n1482_19_CYINIT
    );
  nx53675z1410_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1410_F5MUX,
      O => nx53675z1410
    );
  nx53675z1410_F5MUX_3688 : X_MUX2
    port map (
      IA => nx53675z1411,
      IB => nx53675z1412,
      SEL => nx53675z1410_BXINV,
      O => nx53675z1410_F5MUX
    );
  nx53675z1410_BXINV_3689 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1410_BXINV
    );
  rome2datao5_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_12_F5MUX,
      O => nx53675z333
    );
  rome2datao5_s_12_F5MUX_3690 : X_MUX2
    port map (
      IA => nx53675z334,
      IB => nx53675z335,
      SEL => rome2datao5_s_12_BXINV,
      O => rome2datao5_s_12_F5MUX
    );
  rome2datao5_s_12_BXINV_3691 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao5_s_12_BXINV
    );
  rome2datao5_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_12_F6MUX,
      O => rome2datao5_s(12)
    );
  rome2datao5_s_12_F6MUX_3692 : X_MUX2
    port map (
      IA => nx53675z330,
      IB => nx53675z333,
      SEL => rome2datao5_s_12_BYINV,
      O => rome2datao5_s_12_F6MUX
    );
  rome2datao5_s_12_BYINV_3693 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao5_s_12_BYINV
    );
  nx53675z330_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z330_F5MUX,
      O => nx53675z330
    );
  nx53675z330_F5MUX_3694 : X_MUX2
    port map (
      IA => nx53675z331,
      IB => nx53675z332,
      SEL => nx53675z330_BXINV,
      O => nx53675z330_F5MUX
    );
  nx53675z330_BXINV_3695 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z330_BXINV
    );
  rome2datao5_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_11_F5MUX,
      O => nx53675z339
    );
  rome2datao5_s_11_F5MUX_3696 : X_MUX2
    port map (
      IA => nx53675z340,
      IB => nx53675z341,
      SEL => rome2datao5_s_11_BXINV,
      O => rome2datao5_s_11_F5MUX
    );
  rome2datao5_s_11_BXINV_3697 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao5_s_11_BXINV
    );
  rome2datao5_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_11_F6MUX,
      O => rome2datao5_s(11)
    );
  rome2datao5_s_11_F6MUX_3698 : X_MUX2
    port map (
      IA => nx53675z336,
      IB => nx53675z339,
      SEL => rome2datao5_s_11_BYINV,
      O => rome2datao5_s_11_F6MUX
    );
  rome2datao5_s_11_BYINV_3699 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao5_s_11_BYINV
    );
  nx53675z336_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z336_F5MUX,
      O => nx53675z336
    );
  nx53675z336_F5MUX_3700 : X_MUX2
    port map (
      IA => nx53675z337,
      IB => nx53675z338,
      SEL => nx53675z336_BXINV,
      O => nx53675z336_F5MUX
    );
  nx53675z336_BXINV_3701 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z336_BXINV
    );
  rome2datao5_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_10_F5MUX,
      O => nx53675z345
    );
  rome2datao5_s_10_F5MUX_3702 : X_MUX2
    port map (
      IA => nx53675z346,
      IB => nx53675z347,
      SEL => rome2datao5_s_10_BXINV,
      O => rome2datao5_s_10_F5MUX
    );
  rome2datao5_s_10_BXINV_3703 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao5_s_10_BXINV
    );
  rome2datao5_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_10_F6MUX,
      O => rome2datao5_s(10)
    );
  rome2datao5_s_10_F6MUX_3704 : X_MUX2
    port map (
      IA => nx53675z342,
      IB => nx53675z345,
      SEL => rome2datao5_s_10_BYINV,
      O => rome2datao5_s_10_F6MUX
    );
  rome2datao5_s_10_BYINV_3705 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao5_s_10_BYINV
    );
  nx53675z342_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z342_F5MUX,
      O => nx53675z342
    );
  nx53675z342_F5MUX_3706 : X_MUX2
    port map (
      IA => nx53675z343,
      IB => nx53675z344,
      SEL => nx53675z342_BXINV,
      O => nx53675z342_F5MUX
    );
  nx53675z342_BXINV_3707 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z342_BXINV
    );
  rome2datao5_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_9_F5MUX,
      O => nx53675z351
    );
  rome2datao5_s_9_F5MUX_3708 : X_MUX2
    port map (
      IA => nx53675z352,
      IB => nx53675z353,
      SEL => rome2datao5_s_9_BXINV,
      O => rome2datao5_s_9_F5MUX
    );
  rome2datao5_s_9_BXINV_3709 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao5_s_9_BXINV
    );
  rome2datao5_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_9_F6MUX,
      O => rome2datao5_s(9)
    );
  rome2datao5_s_9_F6MUX_3710 : X_MUX2
    port map (
      IA => nx53675z348,
      IB => nx53675z351,
      SEL => rome2datao5_s_9_BYINV,
      O => rome2datao5_s_9_F6MUX
    );
  rome2datao5_s_9_BYINV_3711 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao5_s_9_BYINV
    );
  nx53675z348_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z348_F5MUX,
      O => nx53675z348
    );
  nx53675z348_F5MUX_3712 : X_MUX2
    port map (
      IA => nx53675z349,
      IB => nx53675z350,
      SEL => nx53675z348_BXINV,
      O => nx53675z348_F5MUX
    );
  nx53675z348_BXINV_3713 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z348_BXINV
    );
  U_DCT2D_reg_databuf_reg_2_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_2_10_DXMUX,
      CE => U_DCT2D_databuf_reg_2_10_CEINV,
      CLK => U_DCT2D_databuf_reg_2_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_2_10_FFX_RST,
      O => U_DCT2D_databuf_reg_2_Q(10)
    );
  U_DCT2D_databuf_reg_2_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_10_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_2_10_FFX_RST
    );
  U_DCT2D_databuf_reg_2_10_FFX_RSTAND_3714 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_2_10_FFX_RSTAND
    );
  rome2datao5_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_3_F5MUX,
      O => nx53675z386
    );
  rome2datao5_s_3_F5MUX_3715 : X_MUX2
    port map (
      IA => nx53675z387,
      IB => nx53675z388,
      SEL => rome2datao5_s_3_BXINV,
      O => rome2datao5_s_3_F5MUX
    );
  rome2datao5_s_3_BXINV_3716 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao5_s_3_BXINV
    );
  rome2datao5_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_3_F6MUX,
      O => rome2datao5_s(3)
    );
  rome2datao5_s_3_F6MUX_3717 : X_MUX2
    port map (
      IA => nx53675z384,
      IB => nx53675z386,
      SEL => rome2datao5_s_3_BYINV,
      O => rome2datao5_s_3_F6MUX
    );
  rome2datao5_s_3_BYINV_3718 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao5_s_3_BYINV
    );
  nx53675z384_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z384_F5MUX,
      O => nx53675z384
    );
  nx53675z384_F5MUX_3719 : X_MUX2
    port map (
      IA => U2_ROME5_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx53675z385,
      SEL => nx53675z384_BXINV,
      O => nx53675z384_F5MUX
    );
  nx53675z384_BXINV_3720 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z384_BXINV
    );
  rome2datao5_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_2_F5MUX,
      O => U2_ROME5_modgen_rom_ix2_nx_ro64_32_l
    );
  rome2datao5_s_2_F5MUX_3721 : X_MUX2
    port map (
      IA => rome2datao5_s_2_G,
      IB => nx53675z389,
      SEL => rome2datao5_s_2_BXINV,
      O => rome2datao5_s_2_F5MUX
    );
  rome2datao5_s_2_BXINV_3722 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao5_s_2_BXINV
    );
  rome2datao5_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_2_F6MUX,
      O => rome2datao5_s(2)
    );
  rome2datao5_s_2_F6MUX_3723 : X_MUX2
    port map (
      IA => U2_ROME5_modgen_rom_ix2_nx_ro64_32_u,
      IB => U2_ROME5_modgen_rom_ix2_nx_ro64_32_l,
      SEL => rome2datao5_s_2_BYINV,
      O => rome2datao5_s_2_F6MUX
    );
  rome2datao5_s_2_BYINV_3724 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao5_s_2_BYINV
    );
  U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U2_ROME5_modgen_rom_ix2_nx_ro64_32_u
    );
  U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_F5MUX_3725 : X_MUX2
    port map (
      IA => U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U2_ROME5_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_BXINV_3726 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  romo2datao8_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_13_F5MUX,
      O => nx53675z1347
    );
  romo2datao8_s_13_F5MUX_3727 : X_MUX2
    port map (
      IA => nx53675z1348,
      IB => nx53675z1349,
      SEL => romo2datao8_s_13_BXINV,
      O => romo2datao8_s_13_F5MUX
    );
  romo2datao8_s_13_BXINV_3728 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_13_BXINV
    );
  romo2datao8_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_13_F6MUX,
      O => romo2datao8_s(13)
    );
  romo2datao8_s_13_F6MUX_3729 : X_MUX2
    port map (
      IA => nx53675z1345,
      IB => nx53675z1347,
      SEL => romo2datao8_s_13_BYINV,
      O => romo2datao8_s_13_F6MUX
    );
  romo2datao8_s_13_BYINV_3730 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_13_BYINV
    );
  nx53675z1345_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1345_F5MUX,
      O => nx53675z1345
    );
  nx53675z1345_F5MUX_3731 : X_MUX2
    port map (
      IA => nx53675z1345_G,
      IB => nx53675z1346,
      SEL => nx53675z1345_BXINV,
      O => nx53675z1345_F5MUX
    );
  nx53675z1345_BXINV_3732 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1345_BXINV
    );
  romo2datao8_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_1_F5MUX,
      O => nx53675z1419
    );
  romo2datao8_s_1_F5MUX_3733 : X_MUX2
    port map (
      IA => nx53675z1420,
      IB => nx53675z1421,
      SEL => romo2datao8_s_1_BXINV,
      O => romo2datao8_s_1_F5MUX
    );
  romo2datao8_s_1_BXINV_3734 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_1_BXINV
    );
  romo2datao8_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_1_F6MUX,
      O => romo2datao8_s(1)
    );
  romo2datao8_s_1_F6MUX_3735 : X_MUX2
    port map (
      IA => nx53675z1416,
      IB => nx53675z1419,
      SEL => romo2datao8_s_1_BYINV,
      O => romo2datao8_s_1_F6MUX
    );
  romo2datao8_s_1_BYINV_3736 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_1_BYINV
    );
  nx53675z1416_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1416_F5MUX,
      O => nx53675z1416
    );
  nx53675z1416_F5MUX_3737 : X_MUX2
    port map (
      IA => nx53675z1417,
      IB => nx53675z1418,
      SEL => nx53675z1416_BXINV,
      O => nx53675z1416_F5MUX
    );
  nx53675z1416_BXINV_3738 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1416_BXINV
    );
  rome2datao7_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_12_F5MUX,
      O => nx53675z463
    );
  rome2datao7_s_12_F5MUX_3739 : X_MUX2
    port map (
      IA => nx53675z464,
      IB => nx53675z465,
      SEL => rome2datao7_s_12_BXINV,
      O => rome2datao7_s_12_F5MUX
    );
  rome2datao7_s_12_BXINV_3740 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao7_s_12_BXINV
    );
  rome2datao7_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_12_F6MUX,
      O => rome2datao7_s(12)
    );
  rome2datao7_s_12_F6MUX_3741 : X_MUX2
    port map (
      IA => nx53675z460,
      IB => nx53675z463,
      SEL => rome2datao7_s_12_BYINV,
      O => rome2datao7_s_12_F6MUX
    );
  rome2datao7_s_12_BYINV_3742 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao7_s_12_BYINV
    );
  ix53675z61491 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => rome2addro7_s(0),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z461
    );
  nx53675z460_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z460_F5MUX,
      O => nx53675z460
    );
  nx53675z460_F5MUX_3743 : X_MUX2
    port map (
      IA => nx53675z461,
      IB => nx53675z462,
      SEL => nx53675z460_BXINV,
      O => nx53675z460_F5MUX
    );
  nx53675z460_BXINV_3744 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z460_BXINV
    );
  rome2datao7_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_11_F5MUX,
      O => nx53675z469
    );
  rome2datao7_s_11_F5MUX_3745 : X_MUX2
    port map (
      IA => nx53675z470,
      IB => nx53675z471,
      SEL => rome2datao7_s_11_BXINV,
      O => rome2datao7_s_11_F5MUX
    );
  rome2datao7_s_11_BXINV_3746 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao7_s_11_BXINV
    );
  rome2datao7_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_11_F6MUX,
      O => rome2datao7_s(11)
    );
  rome2datao7_s_11_F6MUX_3747 : X_MUX2
    port map (
      IA => nx53675z466,
      IB => nx53675z469,
      SEL => rome2datao7_s_11_BYINV,
      O => rome2datao7_s_11_F6MUX
    );
  rome2datao7_s_11_BYINV_3748 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao7_s_11_BYINV
    );
  nx53675z466_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z466_F5MUX,
      O => nx53675z466
    );
  nx53675z466_F5MUX_3749 : X_MUX2
    port map (
      IA => nx53675z467,
      IB => nx53675z468,
      SEL => nx53675z466_BXINV,
      O => nx53675z466_F5MUX
    );
  nx53675z466_BXINV_3750 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z466_BXINV
    );
  rome2datao7_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_3_F5MUX,
      O => nx53675z516
    );
  rome2datao7_s_3_F5MUX_3751 : X_MUX2
    port map (
      IA => nx53675z517,
      IB => nx53675z518,
      SEL => rome2datao7_s_3_BXINV,
      O => rome2datao7_s_3_F5MUX
    );
  rome2datao7_s_3_BXINV_3752 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao7_s_3_BXINV
    );
  rome2datao7_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_3_F6MUX,
      O => rome2datao7_s(3)
    );
  rome2datao7_s_3_F6MUX_3753 : X_MUX2
    port map (
      IA => nx53675z514,
      IB => nx53675z516,
      SEL => rome2datao7_s_3_BYINV,
      O => rome2datao7_s_3_F6MUX
    );
  rome2datao7_s_3_BYINV_3754 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao7_s_3_BYINV
    );
  nx53675z514_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z514_F5MUX,
      O => nx53675z514
    );
  nx53675z514_F5MUX_3755 : X_MUX2
    port map (
      IA => U2_ROME7_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx53675z515,
      SEL => nx53675z514_BXINV,
      O => nx53675z514_F5MUX
    );
  nx53675z514_BXINV_3756 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z514_BXINV
    );
  rome2datao7_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_2_F5MUX,
      O => U2_ROME7_modgen_rom_ix2_nx_ro64_32_l
    );
  rome2datao7_s_2_F5MUX_3757 : X_MUX2
    port map (
      IA => rome2datao7_s_2_G,
      IB => nx53675z519,
      SEL => rome2datao7_s_2_BXINV,
      O => rome2datao7_s_2_F5MUX
    );
  rome2datao7_s_2_BXINV_3758 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao7_s_2_BXINV
    );
  rome2datao7_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_2_F6MUX,
      O => rome2datao7_s(2)
    );
  rome2datao7_s_2_F6MUX_3759 : X_MUX2
    port map (
      IA => U2_ROME7_modgen_rom_ix2_nx_ro64_32_u,
      IB => U2_ROME7_modgen_rom_ix2_nx_ro64_32_l,
      SEL => rome2datao7_s_2_BYINV,
      O => rome2datao7_s_2_F6MUX
    );
  rome2datao7_s_2_BYINV_3760 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao7_s_2_BYINV
    );
  U_DCT2D_ix50549z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_0_1_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_7_1_Q,
      O => U_DCT2D_nx50549z1
    );
  U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U2_ROME7_modgen_rom_ix2_nx_ro64_32_u
    );
  U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_F5MUX_3761 : X_MUX2
    port map (
      IA => U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U2_ROME7_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_BXINV_3762 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  romo2datao9_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_6_F5MUX,
      O => nx53675z1468
    );
  romo2datao9_s_6_F5MUX_3763 : X_MUX2
    port map (
      IA => nx53675z1469,
      IB => nx53675z1470,
      SEL => romo2datao9_s_6_BXINV,
      O => romo2datao9_s_6_F5MUX
    );
  romo2datao9_s_6_BXINV_3764 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_6_BXINV
    );
  romo2datao9_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_6_F6MUX,
      O => romo2datao9_s(6)
    );
  romo2datao9_s_6_F6MUX_3765 : X_MUX2
    port map (
      IA => nx53675z1465,
      IB => nx53675z1468,
      SEL => romo2datao9_s_6_BYINV,
      O => romo2datao9_s_6_F6MUX
    );
  romo2datao9_s_6_BYINV_3766 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_6_BYINV
    );
  nx53675z1465_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1465_F5MUX,
      O => nx53675z1465
    );
  nx53675z1465_F5MUX_3767 : X_MUX2
    port map (
      IA => nx53675z1466,
      IB => nx53675z1467,
      SEL => nx53675z1465_BXINV,
      O => nx53675z1465_F5MUX
    );
  nx53675z1465_BXINV_3768 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1465_BXINV
    );
  romo2datao9_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_5_F5MUX,
      O => nx53675z1474
    );
  romo2datao9_s_5_F5MUX_3769 : X_MUX2
    port map (
      IA => nx53675z1475,
      IB => nx53675z1476,
      SEL => romo2datao9_s_5_BXINV,
      O => romo2datao9_s_5_F5MUX
    );
  romo2datao9_s_5_BXINV_3770 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_5_BXINV
    );
  romo2datao9_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_5_F6MUX,
      O => romo2datao9_s(5)
    );
  romo2datao9_s_5_F6MUX_3771 : X_MUX2
    port map (
      IA => nx53675z1471,
      IB => nx53675z1474,
      SEL => romo2datao9_s_5_BYINV,
      O => romo2datao9_s_5_F6MUX
    );
  romo2datao9_s_5_BYINV_3772 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_5_BYINV
    );
  nx53675z1471_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1471_F5MUX,
      O => nx53675z1471
    );
  nx53675z1471_F5MUX_3773 : X_MUX2
    port map (
      IA => nx53675z1472,
      IB => nx53675z1473,
      SEL => nx53675z1471_BXINV,
      O => nx53675z1471_F5MUX
    );
  nx53675z1471_BXINV_3774 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1471_BXINV
    );
  romo2datao9_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_4_F5MUX,
      O => nx53675z1480
    );
  romo2datao9_s_4_F5MUX_3775 : X_MUX2
    port map (
      IA => nx53675z1481,
      IB => nx53675z1482,
      SEL => romo2datao9_s_4_BXINV,
      O => romo2datao9_s_4_F5MUX
    );
  romo2datao9_s_4_BXINV_3776 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_4_BXINV
    );
  romo2datao9_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_4_F6MUX,
      O => romo2datao9_s(4)
    );
  romo2datao9_s_4_F6MUX_3777 : X_MUX2
    port map (
      IA => nx53675z1477,
      IB => nx53675z1480,
      SEL => romo2datao9_s_4_BYINV,
      O => romo2datao9_s_4_F6MUX
    );
  romo2datao9_s_4_BYINV_3778 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_4_BYINV
    );
  nx53675z1477_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1477_F5MUX,
      O => nx53675z1477
    );
  nx53675z1477_F5MUX_3779 : X_MUX2
    port map (
      IA => nx53675z1478,
      IB => nx53675z1479,
      SEL => nx53675z1477_BXINV,
      O => nx53675z1477_F5MUX
    );
  nx53675z1477_BXINV_3780 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1477_BXINV
    );
  romo2datao9_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_3_F5MUX,
      O => nx53675z1486
    );
  romo2datao9_s_3_F5MUX_3781 : X_MUX2
    port map (
      IA => nx53675z1487,
      IB => nx53675z1488,
      SEL => romo2datao9_s_3_BXINV,
      O => romo2datao9_s_3_F5MUX
    );
  romo2datao9_s_3_BXINV_3782 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_3_BXINV
    );
  romo2datao9_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_3_F6MUX,
      O => romo2datao9_s(3)
    );
  romo2datao9_s_3_F6MUX_3783 : X_MUX2
    port map (
      IA => nx53675z1483,
      IB => nx53675z1486,
      SEL => romo2datao9_s_3_BYINV,
      O => romo2datao9_s_3_F6MUX
    );
  romo2datao9_s_3_BYINV_3784 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_3_BYINV
    );
  nx53675z1483_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1483_F5MUX,
      O => nx53675z1483
    );
  nx53675z1483_F5MUX_3785 : X_MUX2
    port map (
      IA => nx53675z1484,
      IB => nx53675z1485,
      SEL => nx53675z1483_BXINV,
      O => nx53675z1483_F5MUX
    );
  nx53675z1483_BXINV_3786 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1483_BXINV
    );
  romo2datao8_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_0_F5MUX,
      O => U2_ROMO8_modgen_rom_ix0_nx_ro64_32_l
    );
  romo2datao8_s_0_F5MUX_3787 : X_MUX2
    port map (
      IA => nx53675z1422,
      IB => nx53675z1423,
      SEL => romo2datao8_s_0_BXINV,
      O => romo2datao8_s_0_F5MUX
    );
  romo2datao8_s_0_BXINV_3788 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_0_BXINV
    );
  romo2datao8_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_0_F6MUX,
      O => romo2datao8_s(0)
    );
  romo2datao8_s_0_F6MUX_3789 : X_MUX2
    port map (
      IA => U2_ROMO8_modgen_rom_ix0_nx_ro64_32_u,
      IB => U2_ROMO8_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romo2datao8_s_0_BYINV,
      O => romo2datao8_s_0_F6MUX
    );
  romo2datao8_s_0_BYINV_3790 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_0_BYINV
    );
  U2_ROMO8_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROMO8_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U2_ROMO8_modgen_rom_ix0_nx_ro64_32_u
    );
  U2_ROMO8_modgen_rom_ix0_nx_ro64_32_u_F5MUX_3791 : X_MUX2
    port map (
      IA => U2_ROMO8_modgen_rom_ix0_nx_rm64_16_u,
      IB => U2_ROMO8_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U2_ROMO8_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U2_ROMO8_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U2_ROMO8_modgen_rom_ix0_nx_ro64_32_u_BXINV_3792 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => U2_ROMO8_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romo2datao4_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_4_F5MUX,
      O => nx53675z1085
    );
  romo2datao4_s_4_F5MUX_3793 : X_MUX2
    port map (
      IA => nx53675z1086,
      IB => nx53675z1087,
      SEL => romo2datao4_s_4_BXINV,
      O => romo2datao4_s_4_F5MUX
    );
  romo2datao4_s_4_BXINV_3794 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_4_BXINV
    );
  romo2datao4_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_4_F6MUX,
      O => romo2datao4_s(4)
    );
  romo2datao4_s_4_F6MUX_3795 : X_MUX2
    port map (
      IA => nx53675z1082,
      IB => nx53675z1085,
      SEL => romo2datao4_s_4_BYINV,
      O => romo2datao4_s_4_F6MUX
    );
  romo2datao4_s_4_BYINV_3796 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_4_BYINV
    );
  nx53675z1082_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1082_F5MUX,
      O => nx53675z1082
    );
  nx53675z1082_F5MUX_3797 : X_MUX2
    port map (
      IA => nx53675z1083,
      IB => nx53675z1084,
      SEL => nx53675z1082_BXINV,
      O => nx53675z1082_F5MUX
    );
  nx53675z1082_BXINV_3798 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1082_BXINV
    );
  rome2datao4_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_9_F5MUX,
      O => nx53675z286
    );
  rome2datao4_s_9_F5MUX_3799 : X_MUX2
    port map (
      IA => nx53675z287,
      IB => nx53675z288,
      SEL => rome2datao4_s_9_BXINV,
      O => rome2datao4_s_9_F5MUX
    );
  rome2datao4_s_9_BXINV_3800 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao4_s_9_BXINV
    );
  rome2datao4_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_9_F6MUX,
      O => rome2datao4_s(9)
    );
  rome2datao4_s_9_F6MUX_3801 : X_MUX2
    port map (
      IA => nx53675z283,
      IB => nx53675z286,
      SEL => rome2datao4_s_9_BYINV,
      O => rome2datao4_s_9_F6MUX
    );
  rome2datao4_s_9_BYINV_3802 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao4_s_9_BYINV
    );
  nx53675z283_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z283_F5MUX,
      O => nx53675z283
    );
  nx53675z283_F5MUX_3803 : X_MUX2
    port map (
      IA => nx53675z284,
      IB => nx53675z285,
      SEL => nx53675z283_BXINV,
      O => nx53675z283_F5MUX
    );
  nx53675z283_BXINV_3804 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z283_BXINV
    );
  rome2datao4_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_8_F5MUX,
      O => nx53675z292
    );
  rome2datao4_s_8_F5MUX_3805 : X_MUX2
    port map (
      IA => nx53675z293,
      IB => nx53675z294,
      SEL => rome2datao4_s_8_BXINV,
      O => rome2datao4_s_8_F5MUX
    );
  rome2datao4_s_8_BXINV_3806 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao4_s_8_BXINV
    );
  rome2datao4_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_8_F6MUX,
      O => rome2datao4_s(8)
    );
  rome2datao4_s_8_F6MUX_3807 : X_MUX2
    port map (
      IA => nx53675z289,
      IB => nx53675z292,
      SEL => rome2datao4_s_8_BYINV,
      O => rome2datao4_s_8_F6MUX
    );
  rome2datao4_s_8_BYINV_3808 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao4_s_8_BYINV
    );
  nx53675z289_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z289_F5MUX,
      O => nx53675z289
    );
  nx53675z289_F5MUX_3809 : X_MUX2
    port map (
      IA => nx53675z290,
      IB => nx53675z291,
      SEL => nx53675z289_BXINV,
      O => nx53675z289_F5MUX
    );
  nx53675z289_BXINV_3810 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z289_BXINV
    );
  rome2datao4_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_7_F5MUX,
      O => nx53675z298
    );
  rome2datao4_s_7_F5MUX_3811 : X_MUX2
    port map (
      IA => nx53675z299,
      IB => nx53675z300,
      SEL => rome2datao4_s_7_BXINV,
      O => rome2datao4_s_7_F5MUX
    );
  rome2datao4_s_7_BXINV_3812 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao4_s_7_BXINV
    );
  rome2datao4_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_7_F6MUX,
      O => rome2datao4_s(7)
    );
  rome2datao4_s_7_F6MUX_3813 : X_MUX2
    port map (
      IA => nx53675z295,
      IB => nx53675z298,
      SEL => rome2datao4_s_7_BYINV,
      O => rome2datao4_s_7_F6MUX
    );
  rome2datao4_s_7_BYINV_3814 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao4_s_7_BYINV
    );
  nx53675z295_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z295_F5MUX,
      O => nx53675z295
    );
  nx53675z295_F5MUX_3815 : X_MUX2
    port map (
      IA => nx53675z296,
      IB => nx53675z297,
      SEL => nx53675z295_BXINV,
      O => nx53675z295_F5MUX
    );
  nx53675z295_BXINV_3816 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z295_BXINV
    );
  rome2datao3_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_11_F5MUX,
      O => nx53675z209
    );
  rome2datao3_s_11_F5MUX_3817 : X_MUX2
    port map (
      IA => nx53675z210,
      IB => nx53675z211,
      SEL => rome2datao3_s_11_BXINV,
      O => rome2datao3_s_11_F5MUX
    );
  rome2datao3_s_11_BXINV_3818 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao3_s_11_BXINV
    );
  rome2datao3_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_11_F6MUX,
      O => rome2datao3_s(11)
    );
  rome2datao3_s_11_F6MUX_3819 : X_MUX2
    port map (
      IA => nx53675z206,
      IB => nx53675z209,
      SEL => rome2datao3_s_11_BYINV,
      O => rome2datao3_s_11_F6MUX
    );
  rome2datao3_s_11_BYINV_3820 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao3_s_11_BYINV
    );
  U_DCT2D_reg_databuf_reg_4_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_4_0_DYMUX,
      CE => U_DCT2D_databuf_reg_4_0_CEINV,
      CLK => U_DCT2D_databuf_reg_4_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_4_0_FFY_RST,
      O => U_DCT2D_databuf_reg_4_Q(1)
    );
  U_DCT2D_databuf_reg_4_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_4_0_FFY_RST
    );
  nx53675z206_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z206_F5MUX,
      O => nx53675z206
    );
  nx53675z206_F5MUX_3821 : X_MUX2
    port map (
      IA => nx53675z207,
      IB => nx53675z208,
      SEL => nx53675z206_BXINV,
      O => nx53675z206_F5MUX
    );
  nx53675z206_BXINV_3822 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z206_BXINV
    );
  rome2datao0_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_10_F5MUX,
      O => nx53675z21
    );
  rome2datao0_s_10_F5MUX_3823 : X_MUX2
    port map (
      IA => nx53675z22,
      IB => nx53675z23,
      SEL => rome2datao0_s_10_BXINV,
      O => rome2datao0_s_10_F5MUX
    );
  rome2datao0_s_10_BXINV_3824 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao0_s_10_BXINV
    );
  rome2datao0_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_10_F6MUX,
      O => rome2datao0_s(10)
    );
  rome2datao0_s_10_F6MUX_3825 : X_MUX2
    port map (
      IA => nx53675z18,
      IB => nx53675z21,
      SEL => rome2datao0_s_10_BYINV,
      O => rome2datao0_s_10_F6MUX
    );
  rome2datao0_s_10_BYINV_3826 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao0_s_10_BYINV
    );
  ix53675z34386 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => rome2addro0_s(1),
      ADR1 => rome2addro0_s(0),
      ADR2 => rome2addro0_s(3),
      ADR3 => rome2addro0_s(2),
      O => nx53675z19
    );
  nx53675z18_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z18_F5MUX,
      O => nx53675z18
    );
  nx53675z18_F5MUX_3827 : X_MUX2
    port map (
      IA => nx53675z19,
      IB => nx53675z20,
      SEL => nx53675z18_BXINV,
      O => nx53675z18_F5MUX
    );
  nx53675z18_BXINV_3828 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z18_BXINV
    );
  rome2datao0_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_9_F5MUX,
      O => nx53675z27
    );
  rome2datao0_s_9_F5MUX_3829 : X_MUX2
    port map (
      IA => nx53675z28,
      IB => nx53675z29,
      SEL => rome2datao0_s_9_BXINV,
      O => rome2datao0_s_9_F5MUX
    );
  rome2datao0_s_9_BXINV_3830 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao0_s_9_BXINV
    );
  rome2datao0_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_9_F6MUX,
      O => rome2datao0_s(9)
    );
  rome2datao0_s_9_F6MUX_3831 : X_MUX2
    port map (
      IA => nx53675z24,
      IB => nx53675z27,
      SEL => rome2datao0_s_9_BYINV,
      O => rome2datao0_s_9_F6MUX
    );
  rome2datao0_s_9_BYINV_3832 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao0_s_9_BYINV
    );
  nx53675z24_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z24_F5MUX,
      O => nx53675z24
    );
  nx53675z24_F5MUX_3833 : X_MUX2
    port map (
      IA => nx53675z25,
      IB => nx53675z26,
      SEL => nx53675z24_BXINV,
      O => nx53675z24_F5MUX
    );
  nx53675z24_BXINV_3834 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z24_BXINV
    );
  rome2datao9_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_13_F5MUX,
      O => nx53675z587
    );
  rome2datao9_s_13_F5MUX_3835 : X_MUX2
    port map (
      IA => nx53675z588,
      IB => nx53675z589,
      SEL => rome2datao9_s_13_BXINV,
      O => rome2datao9_s_13_F5MUX
    );
  rome2datao9_s_13_BXINV_3836 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao9_s_13_BXINV
    );
  rome2datao9_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_13_F6MUX,
      O => rome2datao9_s(13)
    );
  rome2datao9_s_13_F6MUX_3837 : X_MUX2
    port map (
      IA => nx53675z585,
      IB => nx53675z587,
      SEL => rome2datao9_s_13_BYINV,
      O => rome2datao9_s_13_F6MUX
    );
  rome2datao9_s_13_BYINV_3838 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao9_s_13_BYINV
    );
  nx53675z585_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z585_F5MUX,
      O => nx53675z585
    );
  nx53675z585_F5MUX_3839 : X_MUX2
    port map (
      IA => nx53675z585_G,
      IB => nx53675z586,
      SEL => nx53675z585_BXINV,
      O => nx53675z585_F5MUX
    );
  nx53675z585_BXINV_3840 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z585_BXINV
    );
  rome2datao8_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_2_F5MUX,
      O => U2_ROME8_modgen_rom_ix2_nx_ro64_32_l
    );
  rome2datao8_s_2_F5MUX_3841 : X_MUX2
    port map (
      IA => rome2datao8_s_2_G,
      IB => nx53675z584,
      SEL => rome2datao8_s_2_BXINV,
      O => rome2datao8_s_2_F5MUX
    );
  rome2datao8_s_2_BXINV_3842 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao8_s_2_BXINV
    );
  rome2datao8_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_2_F6MUX,
      O => rome2datao8_s(2)
    );
  rome2datao8_s_2_F6MUX_3843 : X_MUX2
    port map (
      IA => U2_ROME8_modgen_rom_ix2_nx_ro64_32_u,
      IB => U2_ROME8_modgen_rom_ix2_nx_ro64_32_l,
      SEL => rome2datao8_s_2_BYINV,
      O => rome2datao8_s_2_F6MUX
    );
  rome2datao8_s_2_BYINV_3844 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao8_s_2_BYINV
    );
  U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U2_ROME8_modgen_rom_ix2_nx_ro64_32_u
    );
  U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_F5MUX_3845 : X_MUX2
    port map (
      IA => U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U2_ROME8_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_BXINV_3846 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  rome2datao10_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_12_F5MUX,
      O => nx53675z658
    );
  rome2datao10_s_12_F5MUX_3847 : X_MUX2
    port map (
      IA => nx53675z659,
      IB => nx53675z660,
      SEL => rome2datao10_s_12_BXINV,
      O => rome2datao10_s_12_F5MUX
    );
  rome2datao10_s_12_BXINV_3848 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao10_s_12_BXINV
    );
  rome2datao10_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_12_F6MUX,
      O => rome2datao10_s(12)
    );
  rome2datao10_s_12_F6MUX_3849 : X_MUX2
    port map (
      IA => nx53675z655,
      IB => nx53675z658,
      SEL => rome2datao10_s_12_BYINV,
      O => rome2datao10_s_12_F6MUX
    );
  rome2datao10_s_12_BYINV_3850 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao10_s_12_BYINV
    );
  ix53675z61770 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(0),
      ADR3 => rome2addro10_s(3),
      O => nx53675z656
    );
  nx53675z655_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z655_F5MUX,
      O => nx53675z655
    );
  nx53675z655_F5MUX_3851 : X_MUX2
    port map (
      IA => nx53675z656,
      IB => nx53675z657,
      SEL => nx53675z655_BXINV,
      O => nx53675z655_F5MUX
    );
  nx53675z655_BXINV_3852 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z655_BXINV
    );
  rome2datao10_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_11_F5MUX,
      O => nx53675z664
    );
  rome2datao10_s_11_F5MUX_3853 : X_MUX2
    port map (
      IA => nx53675z665,
      IB => nx53675z666,
      SEL => rome2datao10_s_11_BXINV,
      O => rome2datao10_s_11_F5MUX
    );
  rome2datao10_s_11_BXINV_3854 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao10_s_11_BXINV
    );
  rome2datao10_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_11_F6MUX,
      O => rome2datao10_s(11)
    );
  rome2datao10_s_11_F6MUX_3855 : X_MUX2
    port map (
      IA => nx53675z661,
      IB => nx53675z664,
      SEL => rome2datao10_s_11_BYINV,
      O => rome2datao10_s_11_F6MUX
    );
  rome2datao10_s_11_BYINV_3856 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao10_s_11_BYINV
    );
  U_DCT2D_ix59822z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_2_0_Q,
      ADR1 => U_DCT2D_latchbuf_reg_5_0_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx59822z1
    );
  nx53675z661_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z661_F5MUX,
      O => nx53675z661
    );
  nx53675z661_F5MUX_3857 : X_MUX2
    port map (
      IA => nx53675z662,
      IB => nx53675z663,
      SEL => nx53675z661_BXINV,
      O => nx53675z661_F5MUX
    );
  nx53675z661_BXINV_3858 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z661_BXINV
    );
  rome2datao2_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_8_F5MUX,
      O => nx53675z162
    );
  rome2datao2_s_8_F5MUX_3859 : X_MUX2
    port map (
      IA => nx53675z163,
      IB => nx53675z164,
      SEL => rome2datao2_s_8_BXINV,
      O => rome2datao2_s_8_F5MUX
    );
  rome2datao2_s_8_BXINV_3860 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao2_s_8_BXINV
    );
  rome2datao2_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_8_F6MUX,
      O => rome2datao2_s(8)
    );
  rome2datao2_s_8_F6MUX_3861 : X_MUX2
    port map (
      IA => nx53675z159,
      IB => nx53675z162,
      SEL => rome2datao2_s_8_BYINV,
      O => rome2datao2_s_8_F6MUX
    );
  rome2datao2_s_8_BYINV_3862 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao2_s_8_BYINV
    );
  ix53675z7552 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => rome2addro2_s(0),
      ADR1 => rome2addro2_s(1),
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(3),
      O => nx53675z160
    );
  nx53675z159_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z159_F5MUX,
      O => nx53675z159
    );
  nx53675z159_F5MUX_3863 : X_MUX2
    port map (
      IA => nx53675z160,
      IB => nx53675z161,
      SEL => nx53675z159_BXINV,
      O => nx53675z159_F5MUX
    );
  nx53675z159_BXINV_3864 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z159_BXINV
    );
  rome2datao1_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_8_F5MUX,
      O => nx53675z97
    );
  rome2datao1_s_8_F5MUX_3865 : X_MUX2
    port map (
      IA => nx53675z98,
      IB => nx53675z99,
      SEL => rome2datao1_s_8_BXINV,
      O => rome2datao1_s_8_F5MUX
    );
  rome2datao1_s_8_BXINV_3866 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao1_s_8_BXINV
    );
  rome2datao1_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_8_F6MUX,
      O => rome2datao1_s(8)
    );
  rome2datao1_s_8_F6MUX_3867 : X_MUX2
    port map (
      IA => nx53675z94,
      IB => nx53675z97,
      SEL => rome2datao1_s_8_BYINV,
      O => rome2datao1_s_8_F6MUX
    );
  rome2datao1_s_8_BYINV_3868 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao1_s_8_BYINV
    );
  ix53675z7458 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(3),
      O => nx53675z95
    );
  nx53675z94_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z94_F5MUX,
      O => nx53675z94
    );
  nx53675z94_F5MUX_3869 : X_MUX2
    port map (
      IA => nx53675z95,
      IB => nx53675z96,
      SEL => nx53675z94_BXINV,
      O => nx53675z94_F5MUX
    );
  nx53675z94_BXINV_3870 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z94_BXINV
    );
  rome2datao1_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_7_F5MUX,
      O => nx53675z103
    );
  rome2datao1_s_7_F5MUX_3871 : X_MUX2
    port map (
      IA => nx53675z104,
      IB => nx53675z105,
      SEL => rome2datao1_s_7_BXINV,
      O => rome2datao1_s_7_F5MUX
    );
  rome2datao1_s_7_BXINV_3872 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao1_s_7_BXINV
    );
  rome2datao1_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_7_F6MUX,
      O => rome2datao1_s(7)
    );
  rome2datao1_s_7_F6MUX_3873 : X_MUX2
    port map (
      IA => nx53675z100,
      IB => nx53675z103,
      SEL => rome2datao1_s_7_BYINV,
      O => rome2datao1_s_7_F6MUX
    );
  rome2datao1_s_7_BYINV_3874 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao1_s_7_BYINV
    );
  nx53675z100_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z100_F5MUX,
      O => nx53675z100
    );
  nx53675z100_F5MUX_3875 : X_MUX2
    port map (
      IA => nx53675z101,
      IB => nx53675z102,
      SEL => nx53675z100_BXINV,
      O => nx53675z100_F5MUX
    );
  nx53675z100_BXINV_3876 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z100_BXINV
    );
  rome2datao1_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_6_F5MUX,
      O => nx53675z109
    );
  rome2datao1_s_6_F5MUX_3877 : X_MUX2
    port map (
      IA => nx53675z110,
      IB => nx53675z111,
      SEL => rome2datao1_s_6_BXINV,
      O => rome2datao1_s_6_F5MUX
    );
  rome2datao1_s_6_BXINV_3878 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao1_s_6_BXINV
    );
  rome2datao1_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_6_F6MUX,
      O => rome2datao1_s(6)
    );
  rome2datao1_s_6_F6MUX_3879 : X_MUX2
    port map (
      IA => nx53675z106,
      IB => nx53675z109,
      SEL => rome2datao1_s_6_BYINV,
      O => rome2datao1_s_6_F6MUX
    );
  rome2datao1_s_6_BYINV_3880 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao1_s_6_BYINV
    );
  nx53675z106_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z106_F5MUX,
      O => nx53675z106
    );
  nx53675z106_F5MUX_3881 : X_MUX2
    port map (
      IA => nx53675z107,
      IB => nx53675z108,
      SEL => nx53675z106_BXINV,
      O => nx53675z106_F5MUX
    );
  nx53675z106_BXINV_3882 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z106_BXINV
    );
  rome2datao1_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_5_F5MUX,
      O => nx53675z115
    );
  rome2datao1_s_5_F5MUX_3883 : X_MUX2
    port map (
      IA => nx53675z116,
      IB => nx53675z117,
      SEL => rome2datao1_s_5_BXINV,
      O => rome2datao1_s_5_F5MUX
    );
  rome2datao1_s_5_BXINV_3884 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao1_s_5_BXINV
    );
  rome2datao1_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_5_F6MUX,
      O => rome2datao1_s(5)
    );
  rome2datao1_s_5_F6MUX_3885 : X_MUX2
    port map (
      IA => nx53675z112,
      IB => nx53675z115,
      SEL => rome2datao1_s_5_BYINV,
      O => rome2datao1_s_5_F6MUX
    );
  rome2datao1_s_5_BYINV_3886 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao1_s_5_BYINV
    );
  nx53675z112_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z112_F5MUX,
      O => nx53675z112
    );
  nx53675z112_F5MUX_3887 : X_MUX2
    port map (
      IA => nx53675z113,
      IB => nx53675z114,
      SEL => nx53675z112_BXINV,
      O => nx53675z112_F5MUX
    );
  nx53675z112_BXINV_3888 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z112_BXINV
    );
  rome2datao0_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_8_F5MUX,
      O => nx53675z33
    );
  rome2datao0_s_8_F5MUX_3889 : X_MUX2
    port map (
      IA => nx53675z34,
      IB => nx53675z35,
      SEL => rome2datao0_s_8_BXINV,
      O => rome2datao0_s_8_F5MUX
    );
  rome2datao0_s_8_BXINV_3890 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao0_s_8_BXINV
    );
  rome2datao0_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_8_F6MUX,
      O => rome2datao0_s(8)
    );
  rome2datao0_s_8_F6MUX_3891 : X_MUX2
    port map (
      IA => nx53675z30,
      IB => nx53675z33,
      SEL => rome2datao0_s_8_BYINV,
      O => rome2datao0_s_8_F6MUX
    );
  rome2datao0_s_8_BYINV_3892 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao0_s_8_BYINV
    );
  nx53675z30_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z30_F5MUX,
      O => nx53675z30
    );
  nx53675z30_F5MUX_3893 : X_MUX2
    port map (
      IA => nx53675z31,
      IB => nx53675z32,
      SEL => nx53675z30_BXINV,
      O => nx53675z30_F5MUX
    );
  nx53675z30_BXINV_3894 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z30_BXINV
    );
  rome2datao0_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_7_F5MUX,
      O => nx53675z39
    );
  rome2datao0_s_7_F5MUX_3895 : X_MUX2
    port map (
      IA => nx53675z40,
      IB => nx53675z41,
      SEL => rome2datao0_s_7_BXINV,
      O => rome2datao0_s_7_F5MUX
    );
  rome2datao0_s_7_BXINV_3896 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao0_s_7_BXINV
    );
  rome2datao0_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_7_F6MUX,
      O => rome2datao0_s(7)
    );
  rome2datao0_s_7_F6MUX_3897 : X_MUX2
    port map (
      IA => nx53675z36,
      IB => nx53675z39,
      SEL => rome2datao0_s_7_BYINV,
      O => rome2datao0_s_7_F6MUX
    );
  rome2datao0_s_7_BYINV_3898 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao0_s_7_BYINV
    );
  nx53675z36_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z36_F5MUX,
      O => nx53675z36
    );
  nx53675z36_F5MUX_3899 : X_MUX2
    port map (
      IA => nx53675z37,
      IB => nx53675z38,
      SEL => nx53675z36_BXINV,
      O => nx53675z36_F5MUX
    );
  nx53675z36_BXINV_3900 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z36_BXINV
    );
  rome2datao0_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_6_F5MUX,
      O => nx53675z45
    );
  rome2datao0_s_6_F5MUX_3901 : X_MUX2
    port map (
      IA => nx53675z46,
      IB => nx53675z47,
      SEL => rome2datao0_s_6_BXINV,
      O => rome2datao0_s_6_F5MUX
    );
  rome2datao0_s_6_BXINV_3902 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao0_s_6_BXINV
    );
  rome2datao0_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_6_F6MUX,
      O => rome2datao0_s(6)
    );
  rome2datao0_s_6_F6MUX_3903 : X_MUX2
    port map (
      IA => nx53675z42,
      IB => nx53675z45,
      SEL => rome2datao0_s_6_BYINV,
      O => rome2datao0_s_6_F6MUX
    );
  rome2datao0_s_6_BYINV_3904 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao0_s_6_BYINV
    );
  nx53675z42_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z42_F5MUX,
      O => nx53675z42
    );
  nx53675z42_F5MUX_3905 : X_MUX2
    port map (
      IA => nx53675z43,
      IB => nx53675z44,
      SEL => nx53675z42_BXINV,
      O => nx53675z42_F5MUX
    );
  nx53675z42_BXINV_3906 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z42_BXINV
    );
  rome2datao0_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_5_F5MUX,
      O => nx53675z51
    );
  rome2datao0_s_5_F5MUX_3907 : X_MUX2
    port map (
      IA => nx53675z52,
      IB => nx53675z53,
      SEL => rome2datao0_s_5_BXINV,
      O => rome2datao0_s_5_F5MUX
    );
  rome2datao0_s_5_BXINV_3908 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao0_s_5_BXINV
    );
  rome2datao0_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_5_F6MUX,
      O => rome2datao0_s(5)
    );
  rome2datao0_s_5_F6MUX_3909 : X_MUX2
    port map (
      IA => nx53675z48,
      IB => nx53675z51,
      SEL => rome2datao0_s_5_BYINV,
      O => rome2datao0_s_5_F6MUX
    );
  rome2datao0_s_5_BYINV_3910 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao0_s_5_BYINV
    );
  U_DCT2D_reg_databuf_reg_2_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_2_0_DXMUX,
      CE => U_DCT2D_databuf_reg_2_0_CEINV,
      CLK => U_DCT2D_databuf_reg_2_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_2_0_FFX_RST,
      O => U_DCT2D_databuf_reg_2_Q(0)
    );
  U_DCT2D_databuf_reg_2_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_2_0_FFX_RST
    );
  nx53675z48_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z48_F5MUX,
      O => nx53675z48
    );
  nx53675z48_F5MUX_3911 : X_MUX2
    port map (
      IA => nx53675z49,
      IB => nx53675z50,
      SEL => nx53675z48_BXINV,
      O => nx53675z48_F5MUX
    );
  nx53675z48_BXINV_3912 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z48_BXINV
    );
  rome2datao0_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_4_F5MUX,
      O => nx53675z57
    );
  rome2datao0_s_4_F5MUX_3913 : X_MUX2
    port map (
      IA => nx53675z58,
      IB => nx53675z59,
      SEL => rome2datao0_s_4_BXINV,
      O => rome2datao0_s_4_F5MUX
    );
  rome2datao0_s_4_BXINV_3914 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao0_s_4_BXINV
    );
  rome2datao0_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_4_F6MUX,
      O => rome2datao0_s(4)
    );
  rome2datao0_s_4_F6MUX_3915 : X_MUX2
    port map (
      IA => nx53675z54,
      IB => nx53675z57,
      SEL => rome2datao0_s_4_BYINV,
      O => rome2datao0_s_4_F6MUX
    );
  rome2datao0_s_4_BYINV_3916 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao0_s_4_BYINV
    );
  nx53675z54_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z54_F5MUX,
      O => nx53675z54
    );
  nx53675z54_F5MUX_3917 : X_MUX2
    port map (
      IA => nx53675z55,
      IB => nx53675z56,
      SEL => nx53675z54_BXINV,
      O => nx53675z54_F5MUX
    );
  nx53675z54_BXINV_3918 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z54_BXINV
    );
  U_DCT2D_ix62813z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_2_3_Q,
      ADR1 => U_DCT2D_latchbuf_reg_5_3_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx62813z1
    );
  rome2datao9_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_12_F5MUX,
      O => nx53675z593
    );
  rome2datao9_s_12_F5MUX_3919 : X_MUX2
    port map (
      IA => nx53675z594,
      IB => nx53675z595,
      SEL => rome2datao9_s_12_BXINV,
      O => rome2datao9_s_12_F5MUX
    );
  rome2datao9_s_12_BXINV_3920 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao9_s_12_BXINV
    );
  rome2datao9_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_12_F6MUX,
      O => rome2datao9_s(12)
    );
  rome2datao9_s_12_F6MUX_3921 : X_MUX2
    port map (
      IA => nx53675z590,
      IB => nx53675z593,
      SEL => rome2datao9_s_12_BYINV,
      O => rome2datao9_s_12_F6MUX
    );
  rome2datao9_s_12_BYINV_3922 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao9_s_12_BYINV
    );
  nx53675z590_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z590_F5MUX,
      O => nx53675z590
    );
  nx53675z590_F5MUX_3923 : X_MUX2
    port map (
      IA => nx53675z591,
      IB => nx53675z592,
      SEL => nx53675z590_BXINV,
      O => nx53675z590_F5MUX
    );
  nx53675z590_BXINV_3924 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z590_BXINV
    );
  rome2datao9_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_11_F5MUX,
      O => nx53675z599
    );
  rome2datao9_s_11_F5MUX_3925 : X_MUX2
    port map (
      IA => nx53675z600,
      IB => nx53675z601,
      SEL => rome2datao9_s_11_BXINV,
      O => rome2datao9_s_11_F5MUX
    );
  rome2datao9_s_11_BXINV_3926 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao9_s_11_BXINV
    );
  rome2datao9_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_11_F6MUX,
      O => rome2datao9_s(11)
    );
  rome2datao9_s_11_F6MUX_3927 : X_MUX2
    port map (
      IA => nx53675z596,
      IB => nx53675z599,
      SEL => rome2datao9_s_11_BYINV,
      O => rome2datao9_s_11_F6MUX
    );
  rome2datao9_s_11_BYINV_3928 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao9_s_11_BYINV
    );
  nx53675z596_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z596_F5MUX,
      O => nx53675z596
    );
  nx53675z596_F5MUX_3929 : X_MUX2
    port map (
      IA => nx53675z597,
      IB => nx53675z598,
      SEL => nx53675z596_BXINV,
      O => nx53675z596_F5MUX
    );
  nx53675z596_BXINV_3930 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z596_BXINV
    );
  rome2datao9_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_10_F5MUX,
      O => nx53675z605
    );
  rome2datao9_s_10_F5MUX_3931 : X_MUX2
    port map (
      IA => nx53675z606,
      IB => nx53675z607,
      SEL => rome2datao9_s_10_BXINV,
      O => rome2datao9_s_10_F5MUX
    );
  rome2datao9_s_10_BXINV_3932 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao9_s_10_BXINV
    );
  rome2datao9_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_10_F6MUX,
      O => rome2datao9_s(10)
    );
  rome2datao9_s_10_F6MUX_3933 : X_MUX2
    port map (
      IA => nx53675z602,
      IB => nx53675z605,
      SEL => rome2datao9_s_10_BYINV,
      O => rome2datao9_s_10_F6MUX
    );
  rome2datao9_s_10_BYINV_3934 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao9_s_10_BYINV
    );
  nx53675z602_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z602_F5MUX,
      O => nx53675z602
    );
  nx53675z602_F5MUX_3935 : X_MUX2
    port map (
      IA => nx53675z603,
      IB => nx53675z604,
      SEL => nx53675z602_BXINV,
      O => nx53675z602_F5MUX
    );
  nx53675z602_BXINV_3936 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z602_BXINV
    );
  rome2datao9_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_9_F5MUX,
      O => nx53675z611
    );
  rome2datao9_s_9_F5MUX_3937 : X_MUX2
    port map (
      IA => nx53675z612,
      IB => nx53675z613,
      SEL => rome2datao9_s_9_BXINV,
      O => rome2datao9_s_9_F5MUX
    );
  rome2datao9_s_9_BXINV_3938 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao9_s_9_BXINV
    );
  rome2datao9_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_9_F6MUX,
      O => rome2datao9_s(9)
    );
  rome2datao9_s_9_F6MUX_3939 : X_MUX2
    port map (
      IA => nx53675z608,
      IB => nx53675z611,
      SEL => rome2datao9_s_9_BYINV,
      O => rome2datao9_s_9_F6MUX
    );
  rome2datao9_s_9_BYINV_3940 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao9_s_9_BYINV
    );
  nx53675z608_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z608_F5MUX,
      O => nx53675z608
    );
  nx53675z608_F5MUX_3941 : X_MUX2
    port map (
      IA => nx53675z609,
      IB => nx53675z610,
      SEL => nx53675z608_BXINV,
      O => nx53675z608_F5MUX
    );
  nx53675z608_BXINV_3942 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z608_BXINV
    );
  rome2datao9_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_8_F5MUX,
      O => nx53675z617
    );
  rome2datao9_s_8_F5MUX_3943 : X_MUX2
    port map (
      IA => nx53675z618,
      IB => nx53675z619,
      SEL => rome2datao9_s_8_BXINV,
      O => rome2datao9_s_8_F5MUX
    );
  rome2datao9_s_8_BXINV_3944 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao9_s_8_BXINV
    );
  rome2datao9_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_8_F6MUX,
      O => rome2datao9_s(8)
    );
  rome2datao9_s_8_F6MUX_3945 : X_MUX2
    port map (
      IA => nx53675z614,
      IB => nx53675z617,
      SEL => rome2datao9_s_8_BYINV,
      O => rome2datao9_s_8_F6MUX
    );
  rome2datao9_s_8_BYINV_3946 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao9_s_8_BYINV
    );
  nx53675z614_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z614_F5MUX,
      O => nx53675z614
    );
  nx53675z614_F5MUX_3947 : X_MUX2
    port map (
      IA => nx53675z615,
      IB => nx53675z616,
      SEL => nx53675z614_BXINV,
      O => nx53675z614_F5MUX
    );
  nx53675z614_BXINV_3948 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z614_BXINV
    );
  romo2datao1_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_13_F5MUX,
      O => nx53675z794
    );
  romo2datao1_s_13_F5MUX_3949 : X_MUX2
    port map (
      IA => nx53675z795,
      IB => nx53675z796,
      SEL => romo2datao1_s_13_BXINV,
      O => romo2datao1_s_13_F5MUX
    );
  romo2datao1_s_13_BXINV_3950 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_13_BXINV
    );
  romo2datao1_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_13_F6MUX,
      O => romo2datao1_s(13)
    );
  romo2datao1_s_13_F6MUX_3951 : X_MUX2
    port map (
      IA => nx53675z792,
      IB => nx53675z794,
      SEL => romo2datao1_s_13_BYINV,
      O => romo2datao1_s_13_F6MUX
    );
  romo2datao1_s_13_BYINV_3952 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_13_BYINV
    );
  nx53675z792_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z792_F5MUX,
      O => nx53675z792
    );
  nx53675z792_F5MUX_3953 : X_MUX2
    port map (
      IA => nx53675z792_G,
      IB => nx53675z793,
      SEL => nx53675z792_BXINV,
      O => nx53675z792_F5MUX
    );
  nx53675z792_BXINV_3954 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z792_BXINV
    );
  romo2datao0_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_12_F5MUX,
      O => nx53675z723
    );
  romo2datao0_s_12_F5MUX_3955 : X_MUX2
    port map (
      IA => nx53675z724,
      IB => nx53675z725,
      SEL => romo2datao0_s_12_BXINV,
      O => romo2datao0_s_12_F5MUX
    );
  romo2datao0_s_12_BXINV_3956 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_12_BXINV
    );
  romo2datao0_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_12_F6MUX,
      O => romo2datao0_s(12)
    );
  romo2datao0_s_12_F6MUX_3957 : X_MUX2
    port map (
      IA => nx53675z720,
      IB => nx53675z723,
      SEL => romo2datao0_s_12_BYINV,
      O => romo2datao0_s_12_F6MUX
    );
  romo2datao0_s_12_BYINV_3958 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_12_BYINV
    );
  ix53675z59687 : X_LUT4
    generic map(
      INIT => X"8880"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(3),
      ADR2 => romo2addro0_s(1),
      ADR3 => romo2addro0_s(0),
      O => nx53675z721
    );
  nx53675z720_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z720_F5MUX,
      O => nx53675z720
    );
  nx53675z720_F5MUX_3959 : X_MUX2
    port map (
      IA => nx53675z721,
      IB => nx53675z722,
      SEL => nx53675z720_BXINV,
      O => nx53675z720_F5MUX
    );
  nx53675z720_BXINV_3960 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z720_BXINV
    );
  romo2datao0_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_11_F5MUX,
      O => nx53675z729
    );
  romo2datao0_s_11_F5MUX_3961 : X_MUX2
    port map (
      IA => nx53675z730,
      IB => nx53675z731,
      SEL => romo2datao0_s_11_BXINV,
      O => romo2datao0_s_11_F5MUX
    );
  romo2datao0_s_11_BXINV_3962 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_11_BXINV
    );
  romo2datao0_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_11_F6MUX,
      O => romo2datao0_s(11)
    );
  romo2datao0_s_11_F6MUX_3963 : X_MUX2
    port map (
      IA => nx53675z726,
      IB => nx53675z729,
      SEL => romo2datao0_s_11_BYINV,
      O => romo2datao0_s_11_F6MUX
    );
  romo2datao0_s_11_BYINV_3964 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_11_BYINV
    );
  nx53675z726_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z726_F5MUX,
      O => nx53675z726
    );
  nx53675z726_F5MUX_3965 : X_MUX2
    port map (
      IA => nx53675z727,
      IB => nx53675z728,
      SEL => nx53675z726_BXINV,
      O => nx53675z726_F5MUX
    );
  nx53675z726_BXINV_3966 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z726_BXINV
    );
  romo2datao0_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_10_F5MUX,
      O => nx53675z735
    );
  romo2datao0_s_10_F5MUX_3967 : X_MUX2
    port map (
      IA => nx53675z736,
      IB => nx53675z737,
      SEL => romo2datao0_s_10_BXINV,
      O => romo2datao0_s_10_F5MUX
    );
  romo2datao0_s_10_BXINV_3968 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_10_BXINV
    );
  romo2datao0_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_10_F6MUX,
      O => romo2datao0_s(10)
    );
  romo2datao0_s_10_F6MUX_3969 : X_MUX2
    port map (
      IA => nx53675z732,
      IB => nx53675z735,
      SEL => romo2datao0_s_10_BYINV,
      O => romo2datao0_s_10_F6MUX
    );
  romo2datao0_s_10_BYINV_3970 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_10_BYINV
    );
  nx53675z732_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z732_F5MUX,
      O => nx53675z732
    );
  nx53675z732_F5MUX_3971 : X_MUX2
    port map (
      IA => nx53675z733,
      IB => nx53675z734,
      SEL => nx53675z732_BXINV,
      O => nx53675z732_F5MUX
    );
  nx53675z732_BXINV_3972 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z732_BXINV
    );
  romo2datao7_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_9_F5MUX,
      O => nx53675z1292
    );
  romo2datao7_s_9_F5MUX_3973 : X_MUX2
    port map (
      IA => nx53675z1293,
      IB => nx53675z1294,
      SEL => romo2datao7_s_9_BXINV,
      O => romo2datao7_s_9_F5MUX
    );
  romo2datao7_s_9_BXINV_3974 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_9_BXINV
    );
  romo2datao7_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_9_F6MUX,
      O => romo2datao7_s(9)
    );
  romo2datao7_s_9_F6MUX_3975 : X_MUX2
    port map (
      IA => nx53675z1289,
      IB => nx53675z1292,
      SEL => romo2datao7_s_9_BYINV,
      O => romo2datao7_s_9_F6MUX
    );
  romo2datao7_s_9_BYINV_3976 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_9_BYINV
    );
  ix53675z23968 : X_LUT4
    generic map(
      INIT => X"1A0E"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(3),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1290
    );
  nx53675z1289_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1289_F5MUX,
      O => nx53675z1289
    );
  nx53675z1289_F5MUX_3977 : X_MUX2
    port map (
      IA => nx53675z1290,
      IB => nx53675z1291,
      SEL => nx53675z1289_BXINV,
      O => nx53675z1289_F5MUX
    );
  nx53675z1289_BXINV_3978 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1289_BXINV
    );
  romo2datao7_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_8_F5MUX,
      O => nx53675z1298
    );
  romo2datao7_s_8_F5MUX_3979 : X_MUX2
    port map (
      IA => nx53675z1299,
      IB => nx53675z1300,
      SEL => romo2datao7_s_8_BXINV,
      O => romo2datao7_s_8_F5MUX
    );
  romo2datao7_s_8_BXINV_3980 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_8_BXINV
    );
  romo2datao7_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_8_F6MUX,
      O => romo2datao7_s(8)
    );
  romo2datao7_s_8_F6MUX_3981 : X_MUX2
    port map (
      IA => nx53675z1295,
      IB => nx53675z1298,
      SEL => romo2datao7_s_8_BYINV,
      O => romo2datao7_s_8_F6MUX
    );
  romo2datao7_s_8_BYINV_3982 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_8_BYINV
    );
  nx53675z1295_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1295_F5MUX,
      O => nx53675z1295
    );
  nx53675z1295_F5MUX_3983 : X_MUX2
    port map (
      IA => nx53675z1296,
      IB => nx53675z1297,
      SEL => nx53675z1295_BXINV,
      O => nx53675z1295_F5MUX
    );
  nx53675z1295_BXINV_3984 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1295_BXINV
    );
  romo2datao7_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_7_F5MUX,
      O => nx53675z1304
    );
  romo2datao7_s_7_F5MUX_3985 : X_MUX2
    port map (
      IA => nx53675z1305,
      IB => nx53675z1306,
      SEL => romo2datao7_s_7_BXINV,
      O => romo2datao7_s_7_F5MUX
    );
  romo2datao7_s_7_BXINV_3986 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_7_BXINV
    );
  romo2datao7_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_7_F6MUX,
      O => romo2datao7_s(7)
    );
  romo2datao7_s_7_F6MUX_3987 : X_MUX2
    port map (
      IA => nx53675z1301,
      IB => nx53675z1304,
      SEL => romo2datao7_s_7_BYINV,
      O => romo2datao7_s_7_F6MUX
    );
  romo2datao7_s_7_BYINV_3988 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_7_BYINV
    );
  nx53675z1301_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1301_F5MUX,
      O => nx53675z1301
    );
  nx53675z1301_F5MUX_3989 : X_MUX2
    port map (
      IA => nx53675z1302,
      IB => nx53675z1303,
      SEL => nx53675z1301_BXINV,
      O => nx53675z1301_F5MUX
    );
  nx53675z1301_BXINV_3990 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1301_BXINV
    );
  romo2datao7_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_6_F5MUX,
      O => nx53675z1310
    );
  romo2datao7_s_6_F5MUX_3991 : X_MUX2
    port map (
      IA => nx53675z1311,
      IB => nx53675z1312,
      SEL => romo2datao7_s_6_BXINV,
      O => romo2datao7_s_6_F5MUX
    );
  romo2datao7_s_6_BXINV_3992 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_6_BXINV
    );
  romo2datao7_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_6_F6MUX,
      O => romo2datao7_s(6)
    );
  romo2datao7_s_6_F6MUX_3993 : X_MUX2
    port map (
      IA => nx53675z1307,
      IB => nx53675z1310,
      SEL => romo2datao7_s_6_BYINV,
      O => romo2datao7_s_6_F6MUX
    );
  romo2datao7_s_6_BYINV_3994 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_6_BYINV
    );
  nx53675z1307_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1307_F5MUX,
      O => nx53675z1307
    );
  nx53675z1307_F5MUX_3995 : X_MUX2
    port map (
      IA => nx53675z1308,
      IB => nx53675z1309,
      SEL => nx53675z1307_BXINV,
      O => nx53675z1307_F5MUX
    );
  nx53675z1307_BXINV_3996 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1307_BXINV
    );
  romo2datao8_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_11_F5MUX,
      O => nx53675z1359
    );
  romo2datao8_s_11_F5MUX_3997 : X_MUX2
    port map (
      IA => nx53675z1360,
      IB => nx53675z1361,
      SEL => romo2datao8_s_11_BXINV,
      O => romo2datao8_s_11_F5MUX
    );
  romo2datao8_s_11_BXINV_3998 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_11_BXINV
    );
  romo2datao8_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_11_F6MUX,
      O => romo2datao8_s(11)
    );
  romo2datao8_s_11_F6MUX_3999 : X_MUX2
    port map (
      IA => nx53675z1356,
      IB => nx53675z1359,
      SEL => romo2datao8_s_11_BYINV,
      O => romo2datao8_s_11_F6MUX
    );
  romo2datao8_s_11_BYINV_4000 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_11_BYINV
    );
  ix53675z11145 : X_LUT4
    generic map(
      INIT => X"3C68"
    )
    port map (
      ADR0 => romo2addro8_s(0),
      ADR1 => romo2addro8_s(2),
      ADR2 => romo2addro8_s(3),
      ADR3 => romo2addro8_s(1),
      O => nx53675z1357
    );
  nx53675z1356_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1356_F5MUX,
      O => nx53675z1356
    );
  nx53675z1356_F5MUX_4001 : X_MUX2
    port map (
      IA => nx53675z1357,
      IB => nx53675z1358,
      SEL => nx53675z1356_BXINV,
      O => nx53675z1356_F5MUX
    );
  nx53675z1356_BXINV_4002 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1356_BXINV
    );
  romo2datao8_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_10_F5MUX,
      O => nx53675z1365
    );
  romo2datao8_s_10_F5MUX_4003 : X_MUX2
    port map (
      IA => nx53675z1366,
      IB => nx53675z1367,
      SEL => romo2datao8_s_10_BXINV,
      O => romo2datao8_s_10_F5MUX
    );
  romo2datao8_s_10_BXINV_4004 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_10_BXINV
    );
  romo2datao8_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_10_F6MUX,
      O => romo2datao8_s(10)
    );
  romo2datao8_s_10_F6MUX_4005 : X_MUX2
    port map (
      IA => nx53675z1362,
      IB => nx53675z1365,
      SEL => romo2datao8_s_10_BYINV,
      O => romo2datao8_s_10_F6MUX
    );
  romo2datao8_s_10_BYINV_4006 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_10_BYINV
    );
  nx53675z1362_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1362_F5MUX,
      O => nx53675z1362
    );
  nx53675z1362_F5MUX_4007 : X_MUX2
    port map (
      IA => nx53675z1363,
      IB => nx53675z1364,
      SEL => nx53675z1362_BXINV,
      O => nx53675z1362_F5MUX
    );
  nx53675z1362_BXINV_4008 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1362_BXINV
    );
  rome2datao10_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_10_F5MUX,
      O => nx53675z670
    );
  rome2datao10_s_10_F5MUX_4009 : X_MUX2
    port map (
      IA => nx53675z671,
      IB => nx53675z672,
      SEL => rome2datao10_s_10_BXINV,
      O => rome2datao10_s_10_F5MUX
    );
  rome2datao10_s_10_BXINV_4010 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao10_s_10_BXINV
    );
  rome2datao10_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_10_F6MUX,
      O => rome2datao10_s(10)
    );
  rome2datao10_s_10_F6MUX_4011 : X_MUX2
    port map (
      IA => nx53675z667,
      IB => nx53675z670,
      SEL => rome2datao10_s_10_BYINV,
      O => rome2datao10_s_10_F6MUX
    );
  rome2datao10_s_10_BYINV_4012 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao10_s_10_BYINV
    );
  nx53675z667_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z667_F5MUX,
      O => nx53675z667
    );
  nx53675z667_F5MUX_4013 : X_MUX2
    port map (
      IA => nx53675z668,
      IB => nx53675z669,
      SEL => nx53675z667_BXINV,
      O => nx53675z667_F5MUX
    );
  nx53675z667_BXINV_4014 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z667_BXINV
    );
  rome2datao10_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_9_F5MUX,
      O => nx53675z676
    );
  rome2datao10_s_9_F5MUX_4015 : X_MUX2
    port map (
      IA => nx53675z677,
      IB => nx53675z678,
      SEL => rome2datao10_s_9_BXINV,
      O => rome2datao10_s_9_F5MUX
    );
  rome2datao10_s_9_BXINV_4016 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao10_s_9_BXINV
    );
  rome2datao10_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_9_F6MUX,
      O => rome2datao10_s(9)
    );
  rome2datao10_s_9_F6MUX_4017 : X_MUX2
    port map (
      IA => nx53675z673,
      IB => nx53675z676,
      SEL => rome2datao10_s_9_BYINV,
      O => rome2datao10_s_9_F6MUX
    );
  rome2datao10_s_9_BYINV_4018 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao10_s_9_BYINV
    );
  nx53675z673_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z673_F5MUX,
      O => nx53675z673
    );
  nx53675z673_F5MUX_4019 : X_MUX2
    port map (
      IA => nx53675z674,
      IB => nx53675z675,
      SEL => nx53675z673_BXINV,
      O => nx53675z673_F5MUX
    );
  nx53675z673_BXINV_4020 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z673_BXINV
    );
  rome2datao10_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_8_F5MUX,
      O => nx53675z682
    );
  rome2datao10_s_8_F5MUX_4021 : X_MUX2
    port map (
      IA => nx53675z683,
      IB => nx53675z684,
      SEL => rome2datao10_s_8_BXINV,
      O => rome2datao10_s_8_F5MUX
    );
  rome2datao10_s_8_BXINV_4022 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao10_s_8_BXINV
    );
  rome2datao10_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_8_F6MUX,
      O => rome2datao10_s(8)
    );
  rome2datao10_s_8_F6MUX_4023 : X_MUX2
    port map (
      IA => nx53675z679,
      IB => nx53675z682,
      SEL => rome2datao10_s_8_BYINV,
      O => rome2datao10_s_8_F6MUX
    );
  rome2datao10_s_8_BYINV_4024 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao10_s_8_BYINV
    );
  U_DCT2D_reg_databuf_reg_2_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_2_2_DYMUX,
      CE => U_DCT2D_databuf_reg_2_2_CEINV,
      CLK => U_DCT2D_databuf_reg_2_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_2_2_FFY_RST,
      O => U_DCT2D_databuf_reg_2_Q(3)
    );
  U_DCT2D_databuf_reg_2_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_2_2_FFY_RST
    );
  nx53675z679_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z679_F5MUX,
      O => nx53675z679
    );
  nx53675z679_F5MUX_4025 : X_MUX2
    port map (
      IA => nx53675z680,
      IB => nx53675z681,
      SEL => nx53675z679_BXINV,
      O => nx53675z679_F5MUX
    );
  nx53675z679_BXINV_4026 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z679_BXINV
    );
  rome2datao10_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_7_F5MUX,
      O => nx53675z688
    );
  rome2datao10_s_7_F5MUX_4027 : X_MUX2
    port map (
      IA => nx53675z689,
      IB => nx53675z690,
      SEL => rome2datao10_s_7_BXINV,
      O => rome2datao10_s_7_F5MUX
    );
  rome2datao10_s_7_BXINV_4028 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao10_s_7_BXINV
    );
  rome2datao10_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_7_F6MUX,
      O => rome2datao10_s(7)
    );
  rome2datao10_s_7_F6MUX_4029 : X_MUX2
    port map (
      IA => nx53675z685,
      IB => nx53675z688,
      SEL => rome2datao10_s_7_BYINV,
      O => rome2datao10_s_7_F6MUX
    );
  rome2datao10_s_7_BYINV_4030 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao10_s_7_BYINV
    );
  nx53675z685_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z685_F5MUX,
      O => nx53675z685
    );
  nx53675z685_F5MUX_4031 : X_MUX2
    port map (
      IA => nx53675z686,
      IB => nx53675z687,
      SEL => nx53675z685_BXINV,
      O => nx53675z685_F5MUX
    );
  nx53675z685_BXINV_4032 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z685_BXINV
    );
  rome2datao10_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_6_F5MUX,
      O => nx53675z694
    );
  rome2datao10_s_6_F5MUX_4033 : X_MUX2
    port map (
      IA => nx53675z695,
      IB => nx53675z696,
      SEL => rome2datao10_s_6_BXINV,
      O => rome2datao10_s_6_F5MUX
    );
  rome2datao10_s_6_BXINV_4034 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao10_s_6_BXINV
    );
  rome2datao10_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_6_F6MUX,
      O => rome2datao10_s(6)
    );
  rome2datao10_s_6_F6MUX_4035 : X_MUX2
    port map (
      IA => nx53675z691,
      IB => nx53675z694,
      SEL => rome2datao10_s_6_BYINV,
      O => rome2datao10_s_6_F6MUX
    );
  rome2datao10_s_6_BYINV_4036 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao10_s_6_BYINV
    );
  nx53675z691_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z691_F5MUX,
      O => nx53675z691
    );
  nx53675z691_F5MUX_4037 : X_MUX2
    port map (
      IA => nx53675z692,
      IB => nx53675z693,
      SEL => nx53675z691_BXINV,
      O => nx53675z691_F5MUX
    );
  nx53675z691_BXINV_4038 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z691_BXINV
    );
  rome2datao2_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_7_F5MUX,
      O => nx53675z168
    );
  rome2datao2_s_7_F5MUX_4039 : X_MUX2
    port map (
      IA => nx53675z169,
      IB => nx53675z170,
      SEL => rome2datao2_s_7_BXINV,
      O => rome2datao2_s_7_F5MUX
    );
  rome2datao2_s_7_BXINV_4040 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao2_s_7_BXINV
    );
  rome2datao2_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_7_F6MUX,
      O => rome2datao2_s(7)
    );
  rome2datao2_s_7_F6MUX_4041 : X_MUX2
    port map (
      IA => nx53675z165,
      IB => nx53675z168,
      SEL => rome2datao2_s_7_BYINV,
      O => rome2datao2_s_7_F6MUX
    );
  rome2datao2_s_7_BYINV_4042 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao2_s_7_BYINV
    );
  nx53675z165_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z165_F5MUX,
      O => nx53675z165
    );
  nx53675z165_F5MUX_4043 : X_MUX2
    port map (
      IA => nx53675z166,
      IB => nx53675z167,
      SEL => nx53675z165_BXINV,
      O => nx53675z165_F5MUX
    );
  nx53675z165_BXINV_4044 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z165_BXINV
    );
  rome2datao2_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_6_F5MUX,
      O => nx53675z174
    );
  rome2datao2_s_6_F5MUX_4045 : X_MUX2
    port map (
      IA => nx53675z175,
      IB => nx53675z176,
      SEL => rome2datao2_s_6_BXINV,
      O => rome2datao2_s_6_F5MUX
    );
  rome2datao2_s_6_BXINV_4046 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao2_s_6_BXINV
    );
  rome2datao2_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_6_F6MUX,
      O => rome2datao2_s(6)
    );
  rome2datao2_s_6_F6MUX_4047 : X_MUX2
    port map (
      IA => nx53675z171,
      IB => nx53675z174,
      SEL => rome2datao2_s_6_BYINV,
      O => rome2datao2_s_6_F6MUX
    );
  rome2datao2_s_6_BYINV_4048 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao2_s_6_BYINV
    );
  nx53675z171_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z171_F5MUX,
      O => nx53675z171
    );
  nx53675z171_F5MUX_4049 : X_MUX2
    port map (
      IA => nx53675z172,
      IB => nx53675z173,
      SEL => nx53675z171_BXINV,
      O => nx53675z171_F5MUX
    );
  nx53675z171_BXINV_4050 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z171_BXINV
    );
  rome2datao2_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_5_F5MUX,
      O => nx53675z180
    );
  rome2datao2_s_5_F5MUX_4051 : X_MUX2
    port map (
      IA => nx53675z181,
      IB => nx53675z182,
      SEL => rome2datao2_s_5_BXINV,
      O => rome2datao2_s_5_F5MUX
    );
  rome2datao2_s_5_BXINV_4052 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao2_s_5_BXINV
    );
  rome2datao2_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_5_F6MUX,
      O => rome2datao2_s(5)
    );
  rome2datao2_s_5_F6MUX_4053 : X_MUX2
    port map (
      IA => nx53675z177,
      IB => nx53675z180,
      SEL => rome2datao2_s_5_BYINV,
      O => rome2datao2_s_5_F6MUX
    );
  rome2datao2_s_5_BYINV_4054 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao2_s_5_BYINV
    );
  U_DCT2D_ix61816z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_2_2_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_5_2_Q,
      O => U_DCT2D_nx61816z1
    );
  nx53675z177_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z177_F5MUX,
      O => nx53675z177
    );
  nx53675z177_F5MUX_4055 : X_MUX2
    port map (
      IA => nx53675z178,
      IB => nx53675z179,
      SEL => nx53675z177_BXINV,
      O => nx53675z177_F5MUX
    );
  nx53675z177_BXINV_4056 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z177_BXINV
    );
  rome2datao2_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_4_F5MUX,
      O => nx53675z186
    );
  rome2datao2_s_4_F5MUX_4057 : X_MUX2
    port map (
      IA => nx53675z187,
      IB => nx53675z188,
      SEL => rome2datao2_s_4_BXINV,
      O => rome2datao2_s_4_F5MUX
    );
  rome2datao2_s_4_BXINV_4058 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao2_s_4_BXINV
    );
  rome2datao2_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_4_F6MUX,
      O => rome2datao2_s(4)
    );
  rome2datao2_s_4_F6MUX_4059 : X_MUX2
    port map (
      IA => nx53675z183,
      IB => nx53675z186,
      SEL => rome2datao2_s_4_BYINV,
      O => rome2datao2_s_4_F6MUX
    );
  rome2datao2_s_4_BYINV_4060 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao2_s_4_BYINV
    );
  nx53675z183_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z183_F5MUX,
      O => nx53675z183
    );
  nx53675z183_F5MUX_4061 : X_MUX2
    port map (
      IA => nx53675z184,
      IB => nx53675z185,
      SEL => nx53675z183_BXINV,
      O => nx53675z183_F5MUX
    );
  nx53675z183_BXINV_4062 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z183_BXINV
    );
  rome2datao2_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_3_F5MUX,
      O => nx53675z191
    );
  rome2datao2_s_3_F5MUX_4063 : X_MUX2
    port map (
      IA => nx53675z192,
      IB => nx53675z193,
      SEL => rome2datao2_s_3_BXINV,
      O => rome2datao2_s_3_F5MUX
    );
  rome2datao2_s_3_BXINV_4064 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao2_s_3_BXINV
    );
  rome2datao2_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_3_F6MUX,
      O => rome2datao2_s(3)
    );
  rome2datao2_s_3_F6MUX_4065 : X_MUX2
    port map (
      IA => nx53675z189,
      IB => nx53675z191,
      SEL => rome2datao2_s_3_BYINV,
      O => rome2datao2_s_3_F6MUX
    );
  rome2datao2_s_3_BYINV_4066 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao2_s_3_BYINV
    );
  nx53675z189_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z189_F5MUX,
      O => nx53675z189
    );
  nx53675z189_F5MUX_4067 : X_MUX2
    port map (
      IA => U2_ROME2_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx53675z190,
      SEL => nx53675z189_BXINV,
      O => nx53675z189_F5MUX
    );
  nx53675z189_BXINV_4068 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z189_BXINV
    );
  rome2datao2_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_13_F5MUX,
      O => nx53675z132
    );
  rome2datao2_s_13_F5MUX_4069 : X_MUX2
    port map (
      IA => nx53675z133,
      IB => nx53675z134,
      SEL => rome2datao2_s_13_BXINV,
      O => rome2datao2_s_13_F5MUX
    );
  rome2datao2_s_13_BXINV_4070 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao2_s_13_BXINV
    );
  rome2datao2_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_13_F6MUX,
      O => rome2datao2_s(13)
    );
  rome2datao2_s_13_F6MUX_4071 : X_MUX2
    port map (
      IA => nx53675z130,
      IB => nx53675z132,
      SEL => rome2datao2_s_13_BYINV,
      O => rome2datao2_s_13_F6MUX
    );
  rome2datao2_s_13_BYINV_4072 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao2_s_13_BYINV
    );
  nx53675z130_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z130_F5MUX,
      O => nx53675z130
    );
  nx53675z130_F5MUX_4073 : X_MUX2
    port map (
      IA => nx53675z130_G,
      IB => nx53675z131,
      SEL => nx53675z130_BXINV,
      O => nx53675z130_F5MUX
    );
  nx53675z130_BXINV_4074 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z130_BXINV
    );
  rome2datao1_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_12_F5MUX,
      O => nx53675z73
    );
  rome2datao1_s_12_F5MUX_4075 : X_MUX2
    port map (
      IA => nx53675z74,
      IB => nx53675z75,
      SEL => rome2datao1_s_12_BXINV,
      O => rome2datao1_s_12_F5MUX
    );
  rome2datao1_s_12_BXINV_4076 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao1_s_12_BXINV
    );
  rome2datao1_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_12_F6MUX,
      O => rome2datao1_s(12)
    );
  rome2datao1_s_12_F6MUX_4077 : X_MUX2
    port map (
      IA => nx53675z70,
      IB => nx53675z73,
      SEL => rome2datao1_s_12_BYINV,
      O => rome2datao1_s_12_F6MUX
    );
  rome2datao1_s_12_BYINV_4078 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao1_s_12_BYINV
    );
  nx53675z70_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z70_F5MUX,
      O => nx53675z70
    );
  nx53675z70_F5MUX_4079 : X_MUX2
    port map (
      IA => nx53675z71,
      IB => nx53675z72,
      SEL => nx53675z70_BXINV,
      O => nx53675z70_F5MUX
    );
  nx53675z70_BXINV_4080 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z70_BXINV
    );
  romo2datao9_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_13_F5MUX,
      O => nx53675z1426
    );
  romo2datao9_s_13_F5MUX_4081 : X_MUX2
    port map (
      IA => nx53675z1427,
      IB => nx53675z1428,
      SEL => romo2datao9_s_13_BXINV,
      O => romo2datao9_s_13_F5MUX
    );
  romo2datao9_s_13_BXINV_4082 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_13_BXINV
    );
  romo2datao9_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_13_F6MUX,
      O => romo2datao9_s(13)
    );
  romo2datao9_s_13_F6MUX_4083 : X_MUX2
    port map (
      IA => nx53675z1424,
      IB => nx53675z1426,
      SEL => romo2datao9_s_13_BYINV,
      O => romo2datao9_s_13_F6MUX
    );
  romo2datao9_s_13_BYINV_4084 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_13_BYINV
    );
  nx53675z1424_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1424_F5MUX,
      O => nx53675z1424
    );
  nx53675z1424_F5MUX_4085 : X_MUX2
    port map (
      IA => nx53675z1424_G,
      IB => nx53675z1425,
      SEL => nx53675z1424_BXINV,
      O => nx53675z1424_F5MUX
    );
  nx53675z1424_BXINV_4086 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1424_BXINV
    );
  rome2datao10_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_13_F5MUX,
      O => nx53675z652
    );
  rome2datao10_s_13_F5MUX_4087 : X_MUX2
    port map (
      IA => nx53675z653,
      IB => nx53675z654,
      SEL => rome2datao10_s_13_BXINV,
      O => rome2datao10_s_13_F5MUX
    );
  rome2datao10_s_13_BXINV_4088 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao10_s_13_BXINV
    );
  rome2datao10_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_13_F6MUX,
      O => rome2datao10_s(13)
    );
  rome2datao10_s_13_F6MUX_4089 : X_MUX2
    port map (
      IA => nx53675z650,
      IB => nx53675z652,
      SEL => rome2datao10_s_13_BYINV,
      O => rome2datao10_s_13_F6MUX
    );
  rome2datao10_s_13_BYINV_4090 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao10_s_13_BYINV
    );
  nx53675z650_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z650_F5MUX,
      O => nx53675z650
    );
  nx53675z650_F5MUX_4091 : X_MUX2
    port map (
      IA => nx53675z650_G,
      IB => nx53675z651,
      SEL => nx53675z650_BXINV,
      O => nx53675z650_F5MUX
    );
  nx53675z650_BXINV_4092 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z650_BXINV
    );
  rome2datao4_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_6_F5MUX,
      O => nx53675z304
    );
  rome2datao4_s_6_F5MUX_4093 : X_MUX2
    port map (
      IA => nx53675z305,
      IB => nx53675z306,
      SEL => rome2datao4_s_6_BXINV,
      O => rome2datao4_s_6_F5MUX
    );
  rome2datao4_s_6_BXINV_4094 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao4_s_6_BXINV
    );
  rome2datao4_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_6_F6MUX,
      O => rome2datao4_s(6)
    );
  rome2datao4_s_6_F6MUX_4095 : X_MUX2
    port map (
      IA => nx53675z301,
      IB => nx53675z304,
      SEL => rome2datao4_s_6_BYINV,
      O => rome2datao4_s_6_F6MUX
    );
  rome2datao4_s_6_BYINV_4096 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao4_s_6_BYINV
    );
  ix53675z34228 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(1),
      ADR2 => rome2addro4_s(3),
      ADR3 => rome2addro4_s(2),
      O => nx53675z302
    );
  nx53675z301_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z301_F5MUX,
      O => nx53675z301
    );
  nx53675z301_F5MUX_4097 : X_MUX2
    port map (
      IA => nx53675z302,
      IB => nx53675z303,
      SEL => nx53675z301_BXINV,
      O => nx53675z301_F5MUX
    );
  nx53675z301_BXINV_4098 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z301_BXINV
    );
  rome2datao4_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_5_F5MUX,
      O => nx53675z310
    );
  rome2datao4_s_5_F5MUX_4099 : X_MUX2
    port map (
      IA => nx53675z311,
      IB => nx53675z312,
      SEL => rome2datao4_s_5_BXINV,
      O => rome2datao4_s_5_F5MUX
    );
  rome2datao4_s_5_BXINV_4100 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao4_s_5_BXINV
    );
  rome2datao4_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_5_F6MUX,
      O => rome2datao4_s(5)
    );
  rome2datao4_s_5_F6MUX_4101 : X_MUX2
    port map (
      IA => nx53675z307,
      IB => nx53675z310,
      SEL => rome2datao4_s_5_BYINV,
      O => rome2datao4_s_5_F6MUX
    );
  rome2datao4_s_5_BYINV_4102 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao4_s_5_BYINV
    );
  nx53675z307_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z307_F5MUX,
      O => nx53675z307
    );
  nx53675z307_F5MUX_4103 : X_MUX2
    port map (
      IA => nx53675z308,
      IB => nx53675z309,
      SEL => nx53675z307_BXINV,
      O => nx53675z307_F5MUX
    );
  nx53675z307_BXINV_4104 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z307_BXINV
    );
  rome2datao1_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_13_F5MUX,
      O => nx53675z67
    );
  rome2datao1_s_13_F5MUX_4105 : X_MUX2
    port map (
      IA => nx53675z68,
      IB => nx53675z69,
      SEL => rome2datao1_s_13_BXINV,
      O => rome2datao1_s_13_F5MUX
    );
  rome2datao1_s_13_BXINV_4106 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao1_s_13_BXINV
    );
  rome2datao1_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_13_F6MUX,
      O => rome2datao1_s(13)
    );
  rome2datao1_s_13_F6MUX_4107 : X_MUX2
    port map (
      IA => nx53675z65,
      IB => nx53675z67,
      SEL => rome2datao1_s_13_BYINV,
      O => rome2datao1_s_13_F6MUX
    );
  rome2datao1_s_13_BYINV_4108 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao1_s_13_BYINV
    );
  nx53675z65_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z65_F5MUX,
      O => nx53675z65
    );
  nx53675z65_F5MUX_4109 : X_MUX2
    port map (
      IA => nx53675z65_G,
      IB => nx53675z66,
      SEL => nx53675z65_BXINV,
      O => nx53675z65_F5MUX
    );
  nx53675z65_BXINV_4110 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z65_BXINV
    );
  rome2datao1_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_11_F5MUX,
      O => nx53675z79
    );
  rome2datao1_s_11_F5MUX_4111 : X_MUX2
    port map (
      IA => nx53675z80,
      IB => nx53675z81,
      SEL => rome2datao1_s_11_BXINV,
      O => rome2datao1_s_11_F5MUX
    );
  rome2datao1_s_11_BXINV_4112 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao1_s_11_BXINV
    );
  rome2datao1_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_11_F6MUX,
      O => rome2datao1_s(11)
    );
  rome2datao1_s_11_F6MUX_4113 : X_MUX2
    port map (
      IA => nx53675z76,
      IB => nx53675z79,
      SEL => rome2datao1_s_11_BYINV,
      O => rome2datao1_s_11_F6MUX
    );
  rome2datao1_s_11_BYINV_4114 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao1_s_11_BYINV
    );
  U_DCT2D_reg_databuf_reg_2_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_2_2_DXMUX,
      CE => U_DCT2D_databuf_reg_2_2_CEINV,
      CLK => U_DCT2D_databuf_reg_2_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_2_2_FFX_RST,
      O => U_DCT2D_databuf_reg_2_Q(2)
    );
  U_DCT2D_databuf_reg_2_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_2_2_FFX_RST
    );
  nx53675z76_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z76_F5MUX,
      O => nx53675z76
    );
  nx53675z76_F5MUX_4115 : X_MUX2
    port map (
      IA => nx53675z77,
      IB => nx53675z78,
      SEL => nx53675z76_BXINV,
      O => nx53675z76_F5MUX
    );
  nx53675z76_BXINV_4116 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z76_BXINV
    );
  rome2datao1_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_10_F5MUX,
      O => nx53675z85
    );
  rome2datao1_s_10_F5MUX_4117 : X_MUX2
    port map (
      IA => nx53675z86,
      IB => nx53675z87,
      SEL => rome2datao1_s_10_BXINV,
      O => rome2datao1_s_10_F5MUX
    );
  rome2datao1_s_10_BXINV_4118 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao1_s_10_BXINV
    );
  rome2datao1_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_10_F6MUX,
      O => rome2datao1_s(10)
    );
  rome2datao1_s_10_F6MUX_4119 : X_MUX2
    port map (
      IA => nx53675z82,
      IB => nx53675z85,
      SEL => rome2datao1_s_10_BYINV,
      O => rome2datao1_s_10_F6MUX
    );
  rome2datao1_s_10_BYINV_4120 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao1_s_10_BYINV
    );
  nx53675z82_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z82_F5MUX,
      O => nx53675z82
    );
  nx53675z82_F5MUX_4121 : X_MUX2
    port map (
      IA => nx53675z83,
      IB => nx53675z84,
      SEL => nx53675z82_BXINV,
      O => nx53675z82_F5MUX
    );
  nx53675z82_BXINV_4122 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z82_BXINV
    );
  U_DCT2D_ix64807z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_5_5_Q,
      ADR1 => U_DCT2D_latchbuf_reg_2_5_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx64807z1
    );
  rome2datao1_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_4_F5MUX,
      O => nx53675z121
    );
  rome2datao1_s_4_F5MUX_4123 : X_MUX2
    port map (
      IA => nx53675z122,
      IB => nx53675z123,
      SEL => rome2datao1_s_4_BXINV,
      O => rome2datao1_s_4_F5MUX
    );
  rome2datao1_s_4_BXINV_4124 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao1_s_4_BXINV
    );
  rome2datao1_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_4_F6MUX,
      O => rome2datao1_s(4)
    );
  rome2datao1_s_4_F6MUX_4125 : X_MUX2
    port map (
      IA => nx53675z118,
      IB => nx53675z121,
      SEL => rome2datao1_s_4_BYINV,
      O => rome2datao1_s_4_F6MUX
    );
  rome2datao1_s_4_BYINV_4126 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao1_s_4_BYINV
    );
  nx53675z118_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z118_F5MUX,
      O => nx53675z118
    );
  nx53675z118_F5MUX_4127 : X_MUX2
    port map (
      IA => nx53675z119,
      IB => nx53675z120,
      SEL => nx53675z118_BXINV,
      O => nx53675z118_F5MUX
    );
  nx53675z118_BXINV_4128 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z118_BXINV
    );
  rome2datao1_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_3_F5MUX,
      O => nx53675z126
    );
  rome2datao1_s_3_F5MUX_4129 : X_MUX2
    port map (
      IA => nx53675z127,
      IB => nx53675z128,
      SEL => rome2datao1_s_3_BXINV,
      O => rome2datao1_s_3_F5MUX
    );
  rome2datao1_s_3_BXINV_4130 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao1_s_3_BXINV
    );
  rome2datao1_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_3_F6MUX,
      O => rome2datao1_s(3)
    );
  rome2datao1_s_3_F6MUX_4131 : X_MUX2
    port map (
      IA => nx53675z124,
      IB => nx53675z126,
      SEL => rome2datao1_s_3_BYINV,
      O => rome2datao1_s_3_F6MUX
    );
  rome2datao1_s_3_BYINV_4132 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao1_s_3_BYINV
    );
  nx53675z124_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z124_F5MUX,
      O => nx53675z124
    );
  nx53675z124_F5MUX_4133 : X_MUX2
    port map (
      IA => U2_ROME1_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx53675z125,
      SEL => nx53675z124_BXINV,
      O => nx53675z124_F5MUX
    );
  nx53675z124_BXINV_4134 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z124_BXINV
    );
  rome2datao1_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_2_F5MUX,
      O => U2_ROME1_modgen_rom_ix2_nx_ro64_32_l
    );
  rome2datao1_s_2_F5MUX_4135 : X_MUX2
    port map (
      IA => rome2datao1_s_2_G,
      IB => nx53675z129,
      SEL => rome2datao1_s_2_BXINV,
      O => rome2datao1_s_2_F5MUX
    );
  rome2datao1_s_2_BXINV_4136 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao1_s_2_BXINV
    );
  rome2datao1_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_2_F6MUX,
      O => rome2datao1_s(2)
    );
  rome2datao1_s_2_F6MUX_4137 : X_MUX2
    port map (
      IA => U2_ROME1_modgen_rom_ix2_nx_ro64_32_u,
      IB => U2_ROME1_modgen_rom_ix2_nx_ro64_32_l,
      SEL => rome2datao1_s_2_BYINV,
      O => rome2datao1_s_2_F6MUX
    );
  rome2datao1_s_2_BYINV_4138 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao1_s_2_BYINV
    );
  U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U2_ROME1_modgen_rom_ix2_nx_ro64_32_u
    );
  U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_F5MUX_4139 : X_MUX2
    port map (
      IA => U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U2_ROME1_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_BXINV_4140 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  rome2datao0_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_12_F5MUX,
      O => nx53675z9
    );
  rome2datao0_s_12_F5MUX_4141 : X_MUX2
    port map (
      IA => nx53675z10,
      IB => nx53675z11,
      SEL => rome2datao0_s_12_BXINV,
      O => rome2datao0_s_12_F5MUX
    );
  rome2datao0_s_12_BXINV_4142 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao0_s_12_BXINV
    );
  rome2datao0_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_12_F6MUX,
      O => rome2datao0_s(12)
    );
  rome2datao0_s_12_F6MUX_4143 : X_MUX2
    port map (
      IA => nx53675z6,
      IB => nx53675z9,
      SEL => rome2datao0_s_12_BYINV,
      O => rome2datao0_s_12_F6MUX
    );
  rome2datao0_s_12_BYINV_4144 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao0_s_12_BYINV
    );
  nx53675z6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z6_F5MUX,
      O => nx53675z6
    );
  nx53675z6_F5MUX_4145 : X_MUX2
    port map (
      IA => nx53675z7,
      IB => nx53675z8,
      SEL => nx53675z6_BXINV,
      O => nx53675z6_F5MUX
    );
  nx53675z6_BXINV_4146 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z6_BXINV
    );
  rome2datao0_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_11_F5MUX,
      O => nx53675z15
    );
  rome2datao0_s_11_F5MUX_4147 : X_MUX2
    port map (
      IA => nx53675z16,
      IB => nx53675z17,
      SEL => rome2datao0_s_11_BXINV,
      O => rome2datao0_s_11_F5MUX
    );
  rome2datao0_s_11_BXINV_4148 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao0_s_11_BXINV
    );
  rome2datao0_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_11_F6MUX,
      O => rome2datao0_s(11)
    );
  rome2datao0_s_11_F6MUX_4149 : X_MUX2
    port map (
      IA => nx53675z12,
      IB => nx53675z15,
      SEL => rome2datao0_s_11_BYINV,
      O => rome2datao0_s_11_F6MUX
    );
  rome2datao0_s_11_BYINV_4150 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao0_s_11_BYINV
    );
  nx53675z12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z12_F5MUX,
      O => nx53675z12
    );
  nx53675z12_F5MUX_4151 : X_MUX2
    port map (
      IA => nx53675z13,
      IB => nx53675z14,
      SEL => nx53675z12_BXINV,
      O => nx53675z12_F5MUX
    );
  nx53675z12_BXINV_4152 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z12_BXINV
    );
  rome2datao0_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_3_F5MUX,
      O => nx53675z62
    );
  rome2datao0_s_3_F5MUX_4153 : X_MUX2
    port map (
      IA => nx53675z63,
      IB => nx53675z64,
      SEL => rome2datao0_s_3_BXINV,
      O => rome2datao0_s_3_F5MUX
    );
  rome2datao0_s_3_BXINV_4154 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao0_s_3_BXINV
    );
  rome2datao0_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_3_F6MUX,
      O => rome2datao0_s(3)
    );
  rome2datao0_s_3_F6MUX_4155 : X_MUX2
    port map (
      IA => nx53675z60,
      IB => nx53675z62,
      SEL => rome2datao0_s_3_BYINV,
      O => rome2datao0_s_3_F6MUX
    );
  rome2datao0_s_3_BYINV_4156 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao0_s_3_BYINV
    );
  nx53675z60_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z60_F5MUX,
      O => nx53675z60
    );
  nx53675z60_F5MUX_4157 : X_MUX2
    port map (
      IA => U2_ROME0_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx53675z61,
      SEL => nx53675z60_BXINV,
      O => nx53675z60_F5MUX
    );
  nx53675z60_BXINV_4158 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z60_BXINV
    );
  rome2datao9_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_7_F5MUX,
      O => nx53675z623
    );
  rome2datao9_s_7_F5MUX_4159 : X_MUX2
    port map (
      IA => nx53675z624,
      IB => nx53675z625,
      SEL => rome2datao9_s_7_BXINV,
      O => rome2datao9_s_7_F5MUX
    );
  rome2datao9_s_7_BXINV_4160 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao9_s_7_BXINV
    );
  rome2datao9_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_7_F6MUX,
      O => rome2datao9_s(7)
    );
  rome2datao9_s_7_F6MUX_4161 : X_MUX2
    port map (
      IA => nx53675z620,
      IB => nx53675z623,
      SEL => rome2datao9_s_7_BYINV,
      O => rome2datao9_s_7_F6MUX
    );
  rome2datao9_s_7_BYINV_4162 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao9_s_7_BYINV
    );
  nx53675z620_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z620_F5MUX,
      O => nx53675z620
    );
  nx53675z620_F5MUX_4163 : X_MUX2
    port map (
      IA => nx53675z621,
      IB => nx53675z622,
      SEL => nx53675z620_BXINV,
      O => nx53675z620_F5MUX
    );
  nx53675z620_BXINV_4164 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z620_BXINV
    );
  rome2datao9_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_6_F5MUX,
      O => nx53675z629
    );
  rome2datao9_s_6_F5MUX_4165 : X_MUX2
    port map (
      IA => nx53675z630,
      IB => nx53675z631,
      SEL => rome2datao9_s_6_BXINV,
      O => rome2datao9_s_6_F5MUX
    );
  rome2datao9_s_6_BXINV_4166 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao9_s_6_BXINV
    );
  rome2datao9_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_6_F6MUX,
      O => rome2datao9_s(6)
    );
  rome2datao9_s_6_F6MUX_4167 : X_MUX2
    port map (
      IA => nx53675z626,
      IB => nx53675z629,
      SEL => rome2datao9_s_6_BYINV,
      O => rome2datao9_s_6_F6MUX
    );
  rome2datao9_s_6_BYINV_4168 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao9_s_6_BYINV
    );
  nx53675z626_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z626_F5MUX,
      O => nx53675z626
    );
  nx53675z626_F5MUX_4169 : X_MUX2
    port map (
      IA => nx53675z627,
      IB => nx53675z628,
      SEL => nx53675z626_BXINV,
      O => nx53675z626_F5MUX
    );
  nx53675z626_BXINV_4170 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z626_BXINV
    );
  rome2datao9_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_5_F5MUX,
      O => nx53675z635
    );
  rome2datao9_s_5_F5MUX_4171 : X_MUX2
    port map (
      IA => nx53675z636,
      IB => nx53675z637,
      SEL => rome2datao9_s_5_BXINV,
      O => rome2datao9_s_5_F5MUX
    );
  rome2datao9_s_5_BXINV_4172 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao9_s_5_BXINV
    );
  rome2datao9_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_5_F6MUX,
      O => rome2datao9_s(5)
    );
  rome2datao9_s_5_F6MUX_4173 : X_MUX2
    port map (
      IA => nx53675z632,
      IB => nx53675z635,
      SEL => rome2datao9_s_5_BYINV,
      O => rome2datao9_s_5_F6MUX
    );
  rome2datao9_s_5_BYINV_4174 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao9_s_5_BYINV
    );
  nx53675z632_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z632_F5MUX,
      O => nx53675z632
    );
  nx53675z632_F5MUX_4175 : X_MUX2
    port map (
      IA => nx53675z633,
      IB => nx53675z634,
      SEL => nx53675z632_BXINV,
      O => nx53675z632_F5MUX
    );
  nx53675z632_BXINV_4176 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z632_BXINV
    );
  rome2datao9_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_4_F5MUX,
      O => nx53675z641
    );
  rome2datao9_s_4_F5MUX_4177 : X_MUX2
    port map (
      IA => nx53675z642,
      IB => nx53675z643,
      SEL => rome2datao9_s_4_BXINV,
      O => rome2datao9_s_4_F5MUX
    );
  rome2datao9_s_4_BXINV_4178 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao9_s_4_BXINV
    );
  rome2datao9_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_4_F6MUX,
      O => rome2datao9_s(4)
    );
  rome2datao9_s_4_F6MUX_4179 : X_MUX2
    port map (
      IA => nx53675z638,
      IB => nx53675z641,
      SEL => rome2datao9_s_4_BYINV,
      O => rome2datao9_s_4_F6MUX
    );
  rome2datao9_s_4_BYINV_4180 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao9_s_4_BYINV
    );
  nx53675z638_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z638_F5MUX,
      O => nx53675z638
    );
  nx53675z638_F5MUX_4181 : X_MUX2
    port map (
      IA => nx53675z639,
      IB => nx53675z640,
      SEL => nx53675z638_BXINV,
      O => nx53675z638_F5MUX
    );
  nx53675z638_BXINV_4182 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z638_BXINV
    );
  rome2datao9_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_3_F5MUX,
      O => nx53675z646
    );
  rome2datao9_s_3_F5MUX_4183 : X_MUX2
    port map (
      IA => nx53675z647,
      IB => nx53675z648,
      SEL => rome2datao9_s_3_BXINV,
      O => rome2datao9_s_3_F5MUX
    );
  rome2datao9_s_3_BXINV_4184 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao9_s_3_BXINV
    );
  rome2datao9_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_3_F6MUX,
      O => rome2datao9_s(3)
    );
  rome2datao9_s_3_F6MUX_4185 : X_MUX2
    port map (
      IA => nx53675z644,
      IB => nx53675z646,
      SEL => rome2datao9_s_3_BYINV,
      O => rome2datao9_s_3_F6MUX
    );
  rome2datao9_s_3_BYINV_4186 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao9_s_3_BYINV
    );
  nx53675z644_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z644_F5MUX,
      O => nx53675z644
    );
  nx53675z644_F5MUX_4187 : X_MUX2
    port map (
      IA => U2_ROME9_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx53675z645,
      SEL => nx53675z644_BXINV,
      O => nx53675z644_F5MUX
    );
  nx53675z644_BXINV_4188 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z644_BXINV
    );
  rome2datao0_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_13_F5MUX,
      O => nx53675z3
    );
  rome2datao0_s_13_F5MUX_4189 : X_MUX2
    port map (
      IA => nx53675z4,
      IB => nx53675z5,
      SEL => rome2datao0_s_13_BXINV,
      O => rome2datao0_s_13_F5MUX
    );
  rome2datao0_s_13_BXINV_4190 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao0_s_13_BXINV
    );
  rome2datao0_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao0_s_13_F6MUX,
      O => rome2datao0_s(13)
    );
  rome2datao0_s_13_F6MUX_4191 : X_MUX2
    port map (
      IA => nx53675z1,
      IB => nx53675z3,
      SEL => rome2datao0_s_13_BYINV,
      O => rome2datao0_s_13_F6MUX
    );
  rome2datao0_s_13_BYINV_4192 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao0_s_13_BYINV
    );
  nx53675z1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1_F5MUX,
      O => nx53675z1
    );
  nx53675z1_F5MUX_4193 : X_MUX2
    port map (
      IA => nx53675z1_G,
      IB => nx53675z2,
      SEL => nx53675z1_BXINV,
      O => nx53675z1_F5MUX
    );
  nx53675z1_BXINV_4194 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z1_BXINV
    );
  romo2datao2_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_13_F5MUX,
      O => nx53675z873
    );
  romo2datao2_s_13_F5MUX_4195 : X_MUX2
    port map (
      IA => nx53675z874,
      IB => nx53675z875,
      SEL => romo2datao2_s_13_BXINV,
      O => romo2datao2_s_13_F5MUX
    );
  romo2datao2_s_13_BXINV_4196 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_13_BXINV
    );
  romo2datao2_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_13_F6MUX,
      O => romo2datao2_s(13)
    );
  romo2datao2_s_13_F6MUX_4197 : X_MUX2
    port map (
      IA => nx53675z871,
      IB => nx53675z873,
      SEL => romo2datao2_s_13_BYINV,
      O => romo2datao2_s_13_F6MUX
    );
  romo2datao2_s_13_BYINV_4198 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_13_BYINV
    );
  nx53675z871_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z871_F5MUX,
      O => nx53675z871
    );
  nx53675z871_F5MUX_4199 : X_MUX2
    port map (
      IA => nx53675z871_G,
      IB => nx53675z872,
      SEL => nx53675z871_BXINV,
      O => nx53675z871_F5MUX
    );
  nx53675z871_BXINV_4200 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z871_BXINV
    );
  romo2datao2_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_2_F5MUX,
      O => nx53675z939
    );
  romo2datao2_s_2_F5MUX_4201 : X_MUX2
    port map (
      IA => nx53675z940,
      IB => nx53675z941,
      SEL => romo2datao2_s_2_BXINV,
      O => romo2datao2_s_2_F5MUX
    );
  romo2datao2_s_2_BXINV_4202 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_2_BXINV
    );
  romo2datao2_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_2_F6MUX,
      O => romo2datao2_s(2)
    );
  romo2datao2_s_2_F6MUX_4203 : X_MUX2
    port map (
      IA => nx53675z936,
      IB => nx53675z939,
      SEL => romo2datao2_s_2_BYINV,
      O => romo2datao2_s_2_F6MUX
    );
  romo2datao2_s_2_BYINV_4204 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_2_BYINV
    );
  nx53675z936_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z936_F5MUX,
      O => nx53675z936
    );
  nx53675z936_F5MUX_4205 : X_MUX2
    port map (
      IA => nx53675z937,
      IB => nx53675z938,
      SEL => nx53675z936_BXINV,
      O => nx53675z936_F5MUX
    );
  nx53675z936_BXINV_4206 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z936_BXINV
    );
  romo2datao1_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_12_F5MUX,
      O => nx53675z800
    );
  romo2datao1_s_12_F5MUX_4207 : X_MUX2
    port map (
      IA => nx53675z801,
      IB => nx53675z802,
      SEL => romo2datao1_s_12_BXINV,
      O => romo2datao1_s_12_F5MUX
    );
  romo2datao1_s_12_BXINV_4208 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_12_BXINV
    );
  romo2datao1_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_12_F6MUX,
      O => romo2datao1_s(12)
    );
  romo2datao1_s_12_F6MUX_4209 : X_MUX2
    port map (
      IA => nx53675z797,
      IB => nx53675z800,
      SEL => romo2datao1_s_12_BYINV,
      O => romo2datao1_s_12_F6MUX
    );
  romo2datao1_s_12_BYINV_4210 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_12_BYINV
    );
  nx53675z797_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z797_F5MUX,
      O => nx53675z797
    );
  nx53675z797_F5MUX_4211 : X_MUX2
    port map (
      IA => nx53675z798,
      IB => nx53675z799,
      SEL => nx53675z797_BXINV,
      O => nx53675z797_F5MUX
    );
  nx53675z797_BXINV_4212 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z797_BXINV
    );
  romo2datao1_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_11_F5MUX,
      O => nx53675z806
    );
  romo2datao1_s_11_F5MUX_4213 : X_MUX2
    port map (
      IA => nx53675z807,
      IB => nx53675z808,
      SEL => romo2datao1_s_11_BXINV,
      O => romo2datao1_s_11_F5MUX
    );
  romo2datao1_s_11_BXINV_4214 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_11_BXINV
    );
  romo2datao1_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_11_F6MUX,
      O => romo2datao1_s(11)
    );
  romo2datao1_s_11_F6MUX_4215 : X_MUX2
    port map (
      IA => nx53675z803,
      IB => nx53675z806,
      SEL => romo2datao1_s_11_BYINV,
      O => romo2datao1_s_11_F6MUX
    );
  romo2datao1_s_11_BYINV_4216 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_11_BYINV
    );
  nx53675z803_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z803_F5MUX,
      O => nx53675z803
    );
  nx53675z803_F5MUX_4217 : X_MUX2
    port map (
      IA => nx53675z804,
      IB => nx53675z805,
      SEL => nx53675z803_BXINV,
      O => nx53675z803_F5MUX
    );
  nx53675z803_BXINV_4218 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z803_BXINV
    );
  romo2datao1_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_10_F5MUX,
      O => nx53675z812
    );
  romo2datao1_s_10_F5MUX_4219 : X_MUX2
    port map (
      IA => nx53675z813,
      IB => nx53675z814,
      SEL => romo2datao1_s_10_BXINV,
      O => romo2datao1_s_10_F5MUX
    );
  romo2datao1_s_10_BXINV_4220 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_10_BXINV
    );
  romo2datao1_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_10_F6MUX,
      O => romo2datao1_s(10)
    );
  romo2datao1_s_10_F6MUX_4221 : X_MUX2
    port map (
      IA => nx53675z809,
      IB => nx53675z812,
      SEL => romo2datao1_s_10_BYINV,
      O => romo2datao1_s_10_F6MUX
    );
  romo2datao1_s_10_BYINV_4222 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_10_BYINV
    );
  nx53675z809_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z809_F5MUX,
      O => nx53675z809
    );
  nx53675z809_F5MUX_4223 : X_MUX2
    port map (
      IA => nx53675z810,
      IB => nx53675z811,
      SEL => nx53675z809_BXINV,
      O => nx53675z809_F5MUX
    );
  nx53675z809_BXINV_4224 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z809_BXINV
    );
  romo2datao1_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_9_F5MUX,
      O => nx53675z818
    );
  romo2datao1_s_9_F5MUX_4225 : X_MUX2
    port map (
      IA => nx53675z819,
      IB => nx53675z820,
      SEL => romo2datao1_s_9_BXINV,
      O => romo2datao1_s_9_F5MUX
    );
  romo2datao1_s_9_BXINV_4226 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_9_BXINV
    );
  romo2datao1_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_9_F6MUX,
      O => romo2datao1_s(9)
    );
  romo2datao1_s_9_F6MUX_4227 : X_MUX2
    port map (
      IA => nx53675z815,
      IB => nx53675z818,
      SEL => romo2datao1_s_9_BYINV,
      O => romo2datao1_s_9_F6MUX
    );
  romo2datao1_s_9_BYINV_4228 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_9_BYINV
    );
  U_DCT2D_reg_databuf_reg_2_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_2_4_DYMUX,
      CE => U_DCT2D_databuf_reg_2_4_CEINV,
      CLK => U_DCT2D_databuf_reg_2_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_2_4_FFY_RST,
      O => U_DCT2D_databuf_reg_2_Q(5)
    );
  U_DCT2D_databuf_reg_2_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_2_4_FFY_RST
    );
  nx53675z815_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z815_F5MUX,
      O => nx53675z815
    );
  nx53675z815_F5MUX_4229 : X_MUX2
    port map (
      IA => nx53675z816,
      IB => nx53675z817,
      SEL => nx53675z815_BXINV,
      O => nx53675z815_F5MUX
    );
  nx53675z815_BXINV_4230 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z815_BXINV
    );
  romo2datao1_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_8_F5MUX,
      O => nx53675z824
    );
  romo2datao1_s_8_F5MUX_4231 : X_MUX2
    port map (
      IA => nx53675z825,
      IB => nx53675z826,
      SEL => romo2datao1_s_8_BXINV,
      O => romo2datao1_s_8_F5MUX
    );
  romo2datao1_s_8_BXINV_4232 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_8_BXINV
    );
  romo2datao1_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_8_F6MUX,
      O => romo2datao1_s(8)
    );
  romo2datao1_s_8_F6MUX_4233 : X_MUX2
    port map (
      IA => nx53675z821,
      IB => nx53675z824,
      SEL => romo2datao1_s_8_BYINV,
      O => romo2datao1_s_8_F6MUX
    );
  romo2datao1_s_8_BYINV_4234 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_8_BYINV
    );
  nx53675z821_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z821_F5MUX,
      O => nx53675z821
    );
  nx53675z821_F5MUX_4235 : X_MUX2
    port map (
      IA => nx53675z822,
      IB => nx53675z823,
      SEL => nx53675z821_BXINV,
      O => nx53675z821_F5MUX
    );
  nx53675z821_BXINV_4236 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z821_BXINV
    );
  romo2datao1_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_0_F5MUX,
      O => U2_ROMO1_modgen_rom_ix0_nx_ro64_32_l
    );
  romo2datao1_s_0_F5MUX_4237 : X_MUX2
    port map (
      IA => nx53675z869,
      IB => nx53675z870,
      SEL => romo2datao1_s_0_BXINV,
      O => romo2datao1_s_0_F5MUX
    );
  romo2datao1_s_0_BXINV_4238 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_0_BXINV
    );
  romo2datao1_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_0_F6MUX,
      O => romo2datao1_s(0)
    );
  romo2datao1_s_0_F6MUX_4239 : X_MUX2
    port map (
      IA => U2_ROMO1_modgen_rom_ix0_nx_ro64_32_u,
      IB => U2_ROMO1_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romo2datao1_s_0_BYINV,
      O => romo2datao1_s_0_F6MUX
    );
  romo2datao1_s_0_BYINV_4240 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_0_BYINV
    );
  U2_ROMO1_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROMO1_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U2_ROMO1_modgen_rom_ix0_nx_ro64_32_u
    );
  U2_ROMO1_modgen_rom_ix0_nx_ro64_32_u_F5MUX_4241 : X_MUX2
    port map (
      IA => U2_ROMO1_modgen_rom_ix0_nx_rm64_16_u,
      IB => U2_ROMO1_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U2_ROMO1_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U2_ROMO1_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U2_ROMO1_modgen_rom_ix0_nx_ro64_32_u_BXINV_4242 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => U2_ROMO1_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romo2datao0_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_9_F5MUX,
      O => nx53675z741
    );
  romo2datao0_s_9_F5MUX_4243 : X_MUX2
    port map (
      IA => nx53675z742,
      IB => nx53675z743,
      SEL => romo2datao0_s_9_BXINV,
      O => romo2datao0_s_9_F5MUX
    );
  romo2datao0_s_9_BXINV_4244 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_9_BXINV
    );
  romo2datao0_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_9_F6MUX,
      O => romo2datao0_s(9)
    );
  romo2datao0_s_9_F6MUX_4245 : X_MUX2
    port map (
      IA => nx53675z738,
      IB => nx53675z741,
      SEL => romo2datao0_s_9_BYINV,
      O => romo2datao0_s_9_F6MUX
    );
  romo2datao0_s_9_BYINV_4246 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_9_BYINV
    );
  nx53675z738_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z738_F5MUX,
      O => nx53675z738
    );
  nx53675z738_F5MUX_4247 : X_MUX2
    port map (
      IA => nx53675z739,
      IB => nx53675z740,
      SEL => nx53675z738_BXINV,
      O => nx53675z738_F5MUX
    );
  nx53675z738_BXINV_4248 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z738_BXINV
    );
  romo2datao0_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_8_F5MUX,
      O => nx53675z747
    );
  romo2datao0_s_8_F5MUX_4249 : X_MUX2
    port map (
      IA => nx53675z748,
      IB => nx53675z749,
      SEL => romo2datao0_s_8_BXINV,
      O => romo2datao0_s_8_F5MUX
    );
  romo2datao0_s_8_BXINV_4250 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_8_BXINV
    );
  romo2datao0_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_8_F6MUX,
      O => romo2datao0_s(8)
    );
  romo2datao0_s_8_F6MUX_4251 : X_MUX2
    port map (
      IA => nx53675z744,
      IB => nx53675z747,
      SEL => romo2datao0_s_8_BYINV,
      O => romo2datao0_s_8_F6MUX
    );
  romo2datao0_s_8_BYINV_4252 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_8_BYINV
    );
  nx53675z744_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z744_F5MUX,
      O => nx53675z744
    );
  nx53675z744_F5MUX_4253 : X_MUX2
    port map (
      IA => nx53675z745,
      IB => nx53675z746,
      SEL => nx53675z744_BXINV,
      O => nx53675z744_F5MUX
    );
  nx53675z744_BXINV_4254 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z744_BXINV
    );
  romo2datao0_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_7_F5MUX,
      O => nx53675z753
    );
  romo2datao0_s_7_F5MUX_4255 : X_MUX2
    port map (
      IA => nx53675z754,
      IB => nx53675z755,
      SEL => romo2datao0_s_7_BXINV,
      O => romo2datao0_s_7_F5MUX
    );
  romo2datao0_s_7_BXINV_4256 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_7_BXINV
    );
  romo2datao0_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_7_F6MUX,
      O => romo2datao0_s(7)
    );
  romo2datao0_s_7_F6MUX_4257 : X_MUX2
    port map (
      IA => nx53675z750,
      IB => nx53675z753,
      SEL => romo2datao0_s_7_BYINV,
      O => romo2datao0_s_7_F6MUX
    );
  romo2datao0_s_7_BYINV_4258 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_7_BYINV
    );
  U_DCT2D_ix63810z1321 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_2_4_Q,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_5_4_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx63810z1
    );
  nx53675z750_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z750_F5MUX,
      O => nx53675z750
    );
  nx53675z750_F5MUX_4259 : X_MUX2
    port map (
      IA => nx53675z751,
      IB => nx53675z752,
      SEL => nx53675z750_BXINV,
      O => nx53675z750_F5MUX
    );
  nx53675z750_BXINV_4260 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z750_BXINV
    );
  romo2datao0_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_6_F5MUX,
      O => nx53675z759
    );
  romo2datao0_s_6_F5MUX_4261 : X_MUX2
    port map (
      IA => nx53675z760,
      IB => nx53675z761,
      SEL => romo2datao0_s_6_BXINV,
      O => romo2datao0_s_6_F5MUX
    );
  romo2datao0_s_6_BXINV_4262 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_6_BXINV
    );
  romo2datao0_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_6_F6MUX,
      O => romo2datao0_s(6)
    );
  romo2datao0_s_6_F6MUX_4263 : X_MUX2
    port map (
      IA => nx53675z756,
      IB => nx53675z759,
      SEL => romo2datao0_s_6_BYINV,
      O => romo2datao0_s_6_F6MUX
    );
  romo2datao0_s_6_BYINV_4264 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_6_BYINV
    );
  nx53675z756_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z756_F5MUX,
      O => nx53675z756
    );
  nx53675z756_F5MUX_4265 : X_MUX2
    port map (
      IA => nx53675z757,
      IB => nx53675z758,
      SEL => nx53675z756_BXINV,
      O => nx53675z756_F5MUX
    );
  nx53675z756_BXINV_4266 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z756_BXINV
    );
  romo2datao0_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_5_F5MUX,
      O => nx53675z765
    );
  romo2datao0_s_5_F5MUX_4267 : X_MUX2
    port map (
      IA => nx53675z766,
      IB => nx53675z767,
      SEL => romo2datao0_s_5_BXINV,
      O => romo2datao0_s_5_F5MUX
    );
  romo2datao0_s_5_BXINV_4268 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_5_BXINV
    );
  romo2datao0_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_5_F6MUX,
      O => romo2datao0_s(5)
    );
  romo2datao0_s_5_F6MUX_4269 : X_MUX2
    port map (
      IA => nx53675z762,
      IB => nx53675z765,
      SEL => romo2datao0_s_5_BYINV,
      O => romo2datao0_s_5_F6MUX
    );
  romo2datao0_s_5_BYINV_4270 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_5_BYINV
    );
  nx53675z762_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z762_F5MUX,
      O => nx53675z762
    );
  nx53675z762_F5MUX_4271 : X_MUX2
    port map (
      IA => nx53675z763,
      IB => nx53675z764,
      SEL => nx53675z762_BXINV,
      O => nx53675z762_F5MUX
    );
  nx53675z762_BXINV_4272 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z762_BXINV
    );
  rome2datao3_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_12_F5MUX,
      O => nx53675z203
    );
  rome2datao3_s_12_F5MUX_4273 : X_MUX2
    port map (
      IA => nx53675z204,
      IB => nx53675z205,
      SEL => rome2datao3_s_12_BXINV,
      O => rome2datao3_s_12_F5MUX
    );
  rome2datao3_s_12_BXINV_4274 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao3_s_12_BXINV
    );
  rome2datao3_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_12_F6MUX,
      O => rome2datao3_s(12)
    );
  rome2datao3_s_12_F6MUX_4275 : X_MUX2
    port map (
      IA => nx53675z200,
      IB => nx53675z203,
      SEL => rome2datao3_s_12_BYINV,
      O => rome2datao3_s_12_F6MUX
    );
  rome2datao3_s_12_BYINV_4276 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao3_s_12_BYINV
    );
  ix53675z61119 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => rome2addro3_s(0),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(2),
      ADR3 => rome2addro3_s(3),
      O => nx53675z201
    );
  nx53675z200_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z200_F5MUX,
      O => nx53675z200
    );
  nx53675z200_F5MUX_4277 : X_MUX2
    port map (
      IA => nx53675z201,
      IB => nx53675z202,
      SEL => nx53675z200_BXINV,
      O => nx53675z200_F5MUX
    );
  nx53675z200_BXINV_4278 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z200_BXINV
    );
  rome2datao3_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_6_F5MUX,
      O => nx53675z239
    );
  rome2datao3_s_6_F5MUX_4279 : X_MUX2
    port map (
      IA => nx53675z240,
      IB => nx53675z241,
      SEL => rome2datao3_s_6_BXINV,
      O => rome2datao3_s_6_F5MUX
    );
  rome2datao3_s_6_BXINV_4280 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao3_s_6_BXINV
    );
  rome2datao3_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_6_F6MUX,
      O => rome2datao3_s(6)
    );
  rome2datao3_s_6_F6MUX_4281 : X_MUX2
    port map (
      IA => nx53675z236,
      IB => nx53675z239,
      SEL => rome2datao3_s_6_BYINV,
      O => rome2datao3_s_6_F6MUX
    );
  rome2datao3_s_6_BYINV_4282 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao3_s_6_BYINV
    );
  nx53675z236_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z236_F5MUX,
      O => nx53675z236
    );
  nx53675z236_F5MUX_4283 : X_MUX2
    port map (
      IA => nx53675z237,
      IB => nx53675z238,
      SEL => nx53675z236_BXINV,
      O => nx53675z236_F5MUX
    );
  nx53675z236_BXINV_4284 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z236_BXINV
    );
  rome2datao3_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_4_F5MUX,
      O => nx53675z251
    );
  rome2datao3_s_4_F5MUX_4285 : X_MUX2
    port map (
      IA => nx53675z252,
      IB => nx53675z253,
      SEL => rome2datao3_s_4_BXINV,
      O => rome2datao3_s_4_F5MUX
    );
  rome2datao3_s_4_BXINV_4286 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao3_s_4_BXINV
    );
  rome2datao3_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_4_F6MUX,
      O => rome2datao3_s(4)
    );
  rome2datao3_s_4_F6MUX_4287 : X_MUX2
    port map (
      IA => nx53675z248,
      IB => nx53675z251,
      SEL => rome2datao3_s_4_BYINV,
      O => rome2datao3_s_4_F6MUX
    );
  rome2datao3_s_4_BYINV_4288 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao3_s_4_BYINV
    );
  nx53675z248_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z248_F5MUX,
      O => nx53675z248
    );
  nx53675z248_F5MUX_4289 : X_MUX2
    port map (
      IA => nx53675z249,
      IB => nx53675z250,
      SEL => nx53675z248_BXINV,
      O => nx53675z248_F5MUX
    );
  nx53675z248_BXINV_4290 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z248_BXINV
    );
  rome2datao3_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_2_F5MUX,
      O => U2_ROME3_modgen_rom_ix2_nx_ro64_32_l
    );
  rome2datao3_s_2_F5MUX_4291 : X_MUX2
    port map (
      IA => rome2datao3_s_2_G,
      IB => nx53675z259,
      SEL => rome2datao3_s_2_BXINV,
      O => rome2datao3_s_2_F5MUX
    );
  rome2datao3_s_2_BXINV_4292 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao3_s_2_BXINV
    );
  rome2datao3_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_2_F6MUX,
      O => rome2datao3_s(2)
    );
  rome2datao3_s_2_F6MUX_4293 : X_MUX2
    port map (
      IA => U2_ROME3_modgen_rom_ix2_nx_ro64_32_u,
      IB => U2_ROME3_modgen_rom_ix2_nx_ro64_32_l,
      SEL => rome2datao3_s_2_BYINV,
      O => rome2datao3_s_2_F6MUX
    );
  rome2datao3_s_2_BYINV_4294 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao3_s_2_BYINV
    );
  U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U2_ROME3_modgen_rom_ix2_nx_ro64_32_u
    );
  U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_F5MUX_4295 : X_MUX2
    port map (
      IA => U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U2_ROME3_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_BXINV_4296 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  romo2datao3_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_3_F5MUX,
      O => nx53675z1012
    );
  romo2datao3_s_3_F5MUX_4297 : X_MUX2
    port map (
      IA => nx53675z1013,
      IB => nx53675z1014,
      SEL => romo2datao3_s_3_BXINV,
      O => romo2datao3_s_3_F5MUX
    );
  romo2datao3_s_3_BXINV_4298 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_3_BXINV
    );
  romo2datao3_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_3_F6MUX,
      O => romo2datao3_s(3)
    );
  romo2datao3_s_3_F6MUX_4299 : X_MUX2
    port map (
      IA => nx53675z1009,
      IB => nx53675z1012,
      SEL => romo2datao3_s_3_BYINV,
      O => romo2datao3_s_3_F6MUX
    );
  romo2datao3_s_3_BYINV_4300 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_3_BYINV
    );
  ix53675z6773 : X_LUT4
    generic map(
      INIT => X"3388"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => romo2addro3_s(2),
      ADR2 => VCC,
      ADR3 => romo2addro3_s(3),
      O => nx53675z1010
    );
  nx53675z1009_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1009_F5MUX,
      O => nx53675z1009
    );
  nx53675z1009_F5MUX_4301 : X_MUX2
    port map (
      IA => nx53675z1010,
      IB => nx53675z1011,
      SEL => nx53675z1009_BXINV,
      O => nx53675z1009_F5MUX
    );
  nx53675z1009_BXINV_4302 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1009_BXINV
    );
  rome2datao3_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_13_F5MUX,
      O => nx53675z197
    );
  rome2datao3_s_13_F5MUX_4303 : X_MUX2
    port map (
      IA => nx53675z198,
      IB => nx53675z199,
      SEL => rome2datao3_s_13_BXINV,
      O => rome2datao3_s_13_F5MUX
    );
  rome2datao3_s_13_BXINV_4304 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao3_s_13_BXINV
    );
  rome2datao3_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_13_F6MUX,
      O => rome2datao3_s(13)
    );
  rome2datao3_s_13_F6MUX_4305 : X_MUX2
    port map (
      IA => nx53675z195,
      IB => nx53675z197,
      SEL => rome2datao3_s_13_BYINV,
      O => rome2datao3_s_13_F6MUX
    );
  rome2datao3_s_13_BYINV_4306 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao3_s_13_BYINV
    );
  nx53675z195_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z195_F5MUX,
      O => nx53675z195
    );
  nx53675z195_F5MUX_4307 : X_MUX2
    port map (
      IA => nx53675z195_G,
      IB => nx53675z196,
      SEL => nx53675z195_BXINV,
      O => nx53675z195_F5MUX
    );
  nx53675z195_BXINV_4308 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z195_BXINV
    );
  romo2datao8_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_9_F5MUX,
      O => nx53675z1371
    );
  romo2datao8_s_9_F5MUX_4309 : X_MUX2
    port map (
      IA => nx53675z1372,
      IB => nx53675z1373,
      SEL => romo2datao8_s_9_BXINV,
      O => romo2datao8_s_9_F5MUX
    );
  romo2datao8_s_9_BXINV_4310 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_9_BXINV
    );
  romo2datao8_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_9_F6MUX,
      O => romo2datao8_s(9)
    );
  romo2datao8_s_9_F6MUX_4311 : X_MUX2
    port map (
      IA => nx53675z1368,
      IB => nx53675z1371,
      SEL => romo2datao8_s_9_BYINV,
      O => romo2datao8_s_9_F6MUX
    );
  romo2datao8_s_9_BYINV_4312 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_9_BYINV
    );
  nx53675z1368_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1368_F5MUX,
      O => nx53675z1368
    );
  nx53675z1368_F5MUX_4313 : X_MUX2
    port map (
      IA => nx53675z1369,
      IB => nx53675z1370,
      SEL => nx53675z1368_BXINV,
      O => nx53675z1368_F5MUX
    );
  nx53675z1368_BXINV_4314 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1368_BXINV
    );
  romo2datao8_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_8_F5MUX,
      O => nx53675z1377
    );
  romo2datao8_s_8_F5MUX_4315 : X_MUX2
    port map (
      IA => nx53675z1378,
      IB => nx53675z1379,
      SEL => romo2datao8_s_8_BXINV,
      O => romo2datao8_s_8_F5MUX
    );
  romo2datao8_s_8_BXINV_4316 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_8_BXINV
    );
  romo2datao8_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_8_F6MUX,
      O => romo2datao8_s(8)
    );
  romo2datao8_s_8_F6MUX_4317 : X_MUX2
    port map (
      IA => nx53675z1374,
      IB => nx53675z1377,
      SEL => romo2datao8_s_8_BYINV,
      O => romo2datao8_s_8_F6MUX
    );
  romo2datao8_s_8_BYINV_4318 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_8_BYINV
    );
  U_DCT2D_reg_databuf_reg_2_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_2_4_DXMUX,
      CE => U_DCT2D_databuf_reg_2_4_CEINV,
      CLK => U_DCT2D_databuf_reg_2_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_2_4_FFX_RST,
      O => U_DCT2D_databuf_reg_2_Q(4)
    );
  U_DCT2D_databuf_reg_2_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_2_4_FFX_RST
    );
  nx53675z1374_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1374_F5MUX,
      O => nx53675z1374
    );
  nx53675z1374_F5MUX_4319 : X_MUX2
    port map (
      IA => nx53675z1375,
      IB => nx53675z1376,
      SEL => nx53675z1374_BXINV,
      O => nx53675z1374_F5MUX
    );
  nx53675z1374_BXINV_4320 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1374_BXINV
    );
  romo2datao8_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_7_F5MUX,
      O => nx53675z1383
    );
  romo2datao8_s_7_F5MUX_4321 : X_MUX2
    port map (
      IA => nx53675z1384,
      IB => nx53675z1385,
      SEL => romo2datao8_s_7_BXINV,
      O => romo2datao8_s_7_F5MUX
    );
  romo2datao8_s_7_BXINV_4322 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_7_BXINV
    );
  romo2datao8_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_7_F6MUX,
      O => romo2datao8_s(7)
    );
  romo2datao8_s_7_F6MUX_4323 : X_MUX2
    port map (
      IA => nx53675z1380,
      IB => nx53675z1383,
      SEL => romo2datao8_s_7_BYINV,
      O => romo2datao8_s_7_F6MUX
    );
  romo2datao8_s_7_BYINV_4324 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_7_BYINV
    );
  nx53675z1380_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1380_F5MUX,
      O => nx53675z1380
    );
  nx53675z1380_F5MUX_4325 : X_MUX2
    port map (
      IA => nx53675z1381,
      IB => nx53675z1382,
      SEL => nx53675z1380_BXINV,
      O => nx53675z1380_F5MUX
    );
  nx53675z1380_BXINV_4326 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1380_BXINV
    );
  U_DCT2D_ix1265z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_5_7_Q,
      ADR1 => U_DCT2D_latchbuf_reg_2_7_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx1265z1
    );
  romo2datao8_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_6_F5MUX,
      O => nx53675z1389
    );
  romo2datao8_s_6_F5MUX_4327 : X_MUX2
    port map (
      IA => nx53675z1390,
      IB => nx53675z1391,
      SEL => romo2datao8_s_6_BXINV,
      O => romo2datao8_s_6_F5MUX
    );
  romo2datao8_s_6_BXINV_4328 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_6_BXINV
    );
  romo2datao8_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_6_F6MUX,
      O => romo2datao8_s(6)
    );
  romo2datao8_s_6_F6MUX_4329 : X_MUX2
    port map (
      IA => nx53675z1386,
      IB => nx53675z1389,
      SEL => romo2datao8_s_6_BYINV,
      O => romo2datao8_s_6_F6MUX
    );
  romo2datao8_s_6_BYINV_4330 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_6_BYINV
    );
  nx53675z1386_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1386_F5MUX,
      O => nx53675z1386
    );
  nx53675z1386_F5MUX_4331 : X_MUX2
    port map (
      IA => nx53675z1387,
      IB => nx53675z1388,
      SEL => nx53675z1386_BXINV,
      O => nx53675z1386_F5MUX
    );
  nx53675z1386_BXINV_4332 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1386_BXINV
    );
  romo2datao8_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_5_F5MUX,
      O => nx53675z1395
    );
  romo2datao8_s_5_F5MUX_4333 : X_MUX2
    port map (
      IA => nx53675z1396,
      IB => nx53675z1397,
      SEL => romo2datao8_s_5_BXINV,
      O => romo2datao8_s_5_F5MUX
    );
  romo2datao8_s_5_BXINV_4334 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_5_BXINV
    );
  romo2datao8_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_5_F6MUX,
      O => romo2datao8_s(5)
    );
  romo2datao8_s_5_F6MUX_4335 : X_MUX2
    port map (
      IA => nx53675z1392,
      IB => nx53675z1395,
      SEL => romo2datao8_s_5_BYINV,
      O => romo2datao8_s_5_F6MUX
    );
  romo2datao8_s_5_BYINV_4336 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_5_BYINV
    );
  nx53675z1392_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1392_F5MUX,
      O => nx53675z1392
    );
  nx53675z1392_F5MUX_4337 : X_MUX2
    port map (
      IA => nx53675z1393,
      IB => nx53675z1394,
      SEL => nx53675z1392_BXINV,
      O => nx53675z1392_F5MUX
    );
  nx53675z1392_BXINV_4338 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1392_BXINV
    );
  romo2datao7_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_5_F5MUX,
      O => nx53675z1316
    );
  romo2datao7_s_5_F5MUX_4339 : X_MUX2
    port map (
      IA => nx53675z1317,
      IB => nx53675z1318,
      SEL => romo2datao7_s_5_BXINV,
      O => romo2datao7_s_5_F5MUX
    );
  romo2datao7_s_5_BXINV_4340 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_5_BXINV
    );
  romo2datao7_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_5_F6MUX,
      O => romo2datao7_s(5)
    );
  romo2datao7_s_5_F6MUX_4341 : X_MUX2
    port map (
      IA => nx53675z1313,
      IB => nx53675z1316,
      SEL => romo2datao7_s_5_BYINV,
      O => romo2datao7_s_5_F6MUX
    );
  romo2datao7_s_5_BYINV_4342 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_5_BYINV
    );
  nx53675z1313_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1313_F5MUX,
      O => nx53675z1313
    );
  nx53675z1313_F5MUX_4343 : X_MUX2
    port map (
      IA => nx53675z1314,
      IB => nx53675z1315,
      SEL => nx53675z1313_BXINV,
      O => nx53675z1313_F5MUX
    );
  nx53675z1313_BXINV_4344 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1313_BXINV
    );
  romo2datao7_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_4_F5MUX,
      O => nx53675z1322
    );
  romo2datao7_s_4_F5MUX_4345 : X_MUX2
    port map (
      IA => nx53675z1323,
      IB => nx53675z1324,
      SEL => romo2datao7_s_4_BXINV,
      O => romo2datao7_s_4_F5MUX
    );
  romo2datao7_s_4_BXINV_4346 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_4_BXINV
    );
  romo2datao7_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_4_F6MUX,
      O => romo2datao7_s(4)
    );
  romo2datao7_s_4_F6MUX_4347 : X_MUX2
    port map (
      IA => nx53675z1319,
      IB => nx53675z1322,
      SEL => romo2datao7_s_4_BYINV,
      O => romo2datao7_s_4_F6MUX
    );
  romo2datao7_s_4_BYINV_4348 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_4_BYINV
    );
  nx53675z1319_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1319_F5MUX,
      O => nx53675z1319
    );
  nx53675z1319_F5MUX_4349 : X_MUX2
    port map (
      IA => nx53675z1320,
      IB => nx53675z1321,
      SEL => nx53675z1319_BXINV,
      O => nx53675z1319_F5MUX
    );
  nx53675z1319_BXINV_4350 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1319_BXINV
    );
  romo2datao7_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_3_F5MUX,
      O => nx53675z1328
    );
  romo2datao7_s_3_F5MUX_4351 : X_MUX2
    port map (
      IA => nx53675z1329,
      IB => nx53675z1330,
      SEL => romo2datao7_s_3_BXINV,
      O => romo2datao7_s_3_F5MUX
    );
  romo2datao7_s_3_BXINV_4352 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_3_BXINV
    );
  romo2datao7_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_3_F6MUX,
      O => romo2datao7_s(3)
    );
  romo2datao7_s_3_F6MUX_4353 : X_MUX2
    port map (
      IA => nx53675z1325,
      IB => nx53675z1328,
      SEL => romo2datao7_s_3_BYINV,
      O => romo2datao7_s_3_F6MUX
    );
  romo2datao7_s_3_BYINV_4354 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_3_BYINV
    );
  nx53675z1325_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1325_F5MUX,
      O => nx53675z1325
    );
  nx53675z1325_F5MUX_4355 : X_MUX2
    port map (
      IA => nx53675z1326,
      IB => nx53675z1327,
      SEL => nx53675z1325_BXINV,
      O => nx53675z1325_F5MUX
    );
  nx53675z1325_BXINV_4356 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1325_BXINV
    );
  romo2datao7_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_2_F5MUX,
      O => nx53675z1334
    );
  romo2datao7_s_2_F5MUX_4357 : X_MUX2
    port map (
      IA => nx53675z1335,
      IB => nx53675z1336,
      SEL => romo2datao7_s_2_BXINV,
      O => romo2datao7_s_2_F5MUX
    );
  romo2datao7_s_2_BXINV_4358 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_2_BXINV
    );
  romo2datao7_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_2_F6MUX,
      O => romo2datao7_s(2)
    );
  romo2datao7_s_2_F6MUX_4359 : X_MUX2
    port map (
      IA => nx53675z1331,
      IB => nx53675z1334,
      SEL => romo2datao7_s_2_BYINV,
      O => romo2datao7_s_2_F6MUX
    );
  romo2datao7_s_2_BYINV_4360 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_2_BYINV
    );
  nx53675z1331_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1331_F5MUX,
      O => nx53675z1331
    );
  nx53675z1331_F5MUX_4361 : X_MUX2
    port map (
      IA => nx53675z1332,
      IB => nx53675z1333,
      SEL => nx53675z1331_BXINV,
      O => nx53675z1331_F5MUX
    );
  nx53675z1331_BXINV_4362 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1331_BXINV
    );
  romo2datao7_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_1_F5MUX,
      O => nx53675z1340
    );
  romo2datao7_s_1_F5MUX_4363 : X_MUX2
    port map (
      IA => nx53675z1341,
      IB => nx53675z1342,
      SEL => romo2datao7_s_1_BXINV,
      O => romo2datao7_s_1_F5MUX
    );
  romo2datao7_s_1_BXINV_4364 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_1_BXINV
    );
  romo2datao7_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_1_F6MUX,
      O => romo2datao7_s(1)
    );
  romo2datao7_s_1_F6MUX_4365 : X_MUX2
    port map (
      IA => nx53675z1337,
      IB => nx53675z1340,
      SEL => romo2datao7_s_1_BYINV,
      O => romo2datao7_s_1_F6MUX
    );
  romo2datao7_s_1_BYINV_4366 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_1_BYINV
    );
  nx53675z1337_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1337_F5MUX,
      O => nx53675z1337
    );
  nx53675z1337_F5MUX_4367 : X_MUX2
    port map (
      IA => nx53675z1338,
      IB => nx53675z1339,
      SEL => nx53675z1337_BXINV,
      O => nx53675z1337_F5MUX
    );
  nx53675z1337_BXINV_4368 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1337_BXINV
    );
  rome2datao5_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_5_F5MUX,
      O => nx53675z375
    );
  rome2datao5_s_5_F5MUX_4369 : X_MUX2
    port map (
      IA => nx53675z376,
      IB => nx53675z377,
      SEL => rome2datao5_s_5_BXINV,
      O => rome2datao5_s_5_F5MUX
    );
  rome2datao5_s_5_BXINV_4370 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao5_s_5_BXINV
    );
  rome2datao5_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_5_F6MUX,
      O => rome2datao5_s(5)
    );
  rome2datao5_s_5_F6MUX_4371 : X_MUX2
    port map (
      IA => nx53675z372,
      IB => nx53675z375,
      SEL => rome2datao5_s_5_BYINV,
      O => rome2datao5_s_5_F6MUX
    );
  rome2datao5_s_5_BYINV_4372 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao5_s_5_BYINV
    );
  ix53675z61639 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro5_s(1),
      ADR1 => rome2addro5_s(3),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z373
    );
  nx53675z372_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z372_F5MUX,
      O => nx53675z372
    );
  nx53675z372_F5MUX_4373 : X_MUX2
    port map (
      IA => nx53675z373,
      IB => nx53675z374,
      SEL => nx53675z372_BXINV,
      O => nx53675z372_F5MUX
    );
  nx53675z372_BXINV_4374 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z372_BXINV
    );
  rome2datao5_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_4_F5MUX,
      O => nx53675z381
    );
  rome2datao5_s_4_F5MUX_4375 : X_MUX2
    port map (
      IA => nx53675z382,
      IB => nx53675z383,
      SEL => rome2datao5_s_4_BXINV,
      O => rome2datao5_s_4_F5MUX
    );
  rome2datao5_s_4_BXINV_4376 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao5_s_4_BXINV
    );
  rome2datao5_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_4_F6MUX,
      O => rome2datao5_s(4)
    );
  rome2datao5_s_4_F6MUX_4377 : X_MUX2
    port map (
      IA => nx53675z378,
      IB => nx53675z381,
      SEL => rome2datao5_s_4_BYINV,
      O => rome2datao5_s_4_F6MUX
    );
  rome2datao5_s_4_BYINV_4378 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao5_s_4_BYINV
    );
  nx53675z378_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z378_F5MUX,
      O => nx53675z378
    );
  nx53675z378_F5MUX_4379 : X_MUX2
    port map (
      IA => nx53675z379,
      IB => nx53675z380,
      SEL => nx53675z378_BXINV,
      O => nx53675z378_F5MUX
    );
  nx53675z378_BXINV_4380 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z378_BXINV
    );
  romo2datao7_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_0_F5MUX,
      O => U2_ROMO7_modgen_rom_ix0_nx_ro64_32_l
    );
  romo2datao7_s_0_F5MUX_4381 : X_MUX2
    port map (
      IA => nx53675z1343,
      IB => nx53675z1344,
      SEL => romo2datao7_s_0_BXINV,
      O => romo2datao7_s_0_F5MUX
    );
  romo2datao7_s_0_BXINV_4382 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_0_BXINV
    );
  romo2datao7_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_0_F6MUX,
      O => romo2datao7_s(0)
    );
  romo2datao7_s_0_F6MUX_4383 : X_MUX2
    port map (
      IA => U2_ROMO7_modgen_rom_ix0_nx_ro64_32_u,
      IB => U2_ROMO7_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romo2datao7_s_0_BYINV,
      O => romo2datao7_s_0_F6MUX
    );
  romo2datao7_s_0_BYINV_4384 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_0_BYINV
    );
  U2_ROMO7_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROMO7_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U2_ROMO7_modgen_rom_ix0_nx_ro64_32_u
    );
  U2_ROMO7_modgen_rom_ix0_nx_ro64_32_u_F5MUX_4385 : X_MUX2
    port map (
      IA => U2_ROMO7_modgen_rom_ix0_nx_rm64_16_u,
      IB => U2_ROMO7_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U2_ROMO7_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U2_ROMO7_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U2_ROMO7_modgen_rom_ix0_nx_ro64_32_u_BXINV_4386 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => U2_ROMO7_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  rome2datao10_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_5_F5MUX,
      O => nx53675z700
    );
  rome2datao10_s_5_F5MUX_4387 : X_MUX2
    port map (
      IA => nx53675z701,
      IB => nx53675z702,
      SEL => rome2datao10_s_5_BXINV,
      O => rome2datao10_s_5_F5MUX
    );
  rome2datao10_s_5_BXINV_4388 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao10_s_5_BXINV
    );
  rome2datao10_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_5_F6MUX,
      O => rome2datao10_s(5)
    );
  rome2datao10_s_5_F6MUX_4389 : X_MUX2
    port map (
      IA => nx53675z697,
      IB => nx53675z700,
      SEL => rome2datao10_s_5_BYINV,
      O => rome2datao10_s_5_F6MUX
    );
  rome2datao10_s_5_BYINV_4390 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao10_s_5_BYINV
    );
  nx53675z697_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z697_F5MUX,
      O => nx53675z697
    );
  nx53675z697_F5MUX_4391 : X_MUX2
    port map (
      IA => nx53675z698,
      IB => nx53675z699,
      SEL => nx53675z697_BXINV,
      O => nx53675z697_F5MUX
    );
  nx53675z697_BXINV_4392 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z697_BXINV
    );
  rome2datao10_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_4_F5MUX,
      O => nx53675z706
    );
  rome2datao10_s_4_F5MUX_4393 : X_MUX2
    port map (
      IA => nx53675z707,
      IB => nx53675z708,
      SEL => rome2datao10_s_4_BXINV,
      O => rome2datao10_s_4_F5MUX
    );
  rome2datao10_s_4_BXINV_4394 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao10_s_4_BXINV
    );
  rome2datao10_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_4_F6MUX,
      O => rome2datao10_s(4)
    );
  rome2datao10_s_4_F6MUX_4395 : X_MUX2
    port map (
      IA => nx53675z703,
      IB => nx53675z706,
      SEL => rome2datao10_s_4_BYINV,
      O => rome2datao10_s_4_F6MUX
    );
  rome2datao10_s_4_BYINV_4396 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao10_s_4_BYINV
    );
  nx53675z703_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z703_F5MUX,
      O => nx53675z703
    );
  nx53675z703_F5MUX_4397 : X_MUX2
    port map (
      IA => nx53675z704,
      IB => nx53675z705,
      SEL => nx53675z703_BXINV,
      O => nx53675z703_F5MUX
    );
  nx53675z703_BXINV_4398 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z703_BXINV
    );
  rome2datao10_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_3_F5MUX,
      O => nx53675z711
    );
  rome2datao10_s_3_F5MUX_4399 : X_MUX2
    port map (
      IA => nx53675z712,
      IB => nx53675z713,
      SEL => rome2datao10_s_3_BXINV,
      O => rome2datao10_s_3_F5MUX
    );
  rome2datao10_s_3_BXINV_4400 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao10_s_3_BXINV
    );
  rome2datao10_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_3_F6MUX,
      O => rome2datao10_s(3)
    );
  rome2datao10_s_3_F6MUX_4401 : X_MUX2
    port map (
      IA => nx53675z709,
      IB => nx53675z711,
      SEL => rome2datao10_s_3_BYINV,
      O => rome2datao10_s_3_F6MUX
    );
  rome2datao10_s_3_BYINV_4402 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao10_s_3_BYINV
    );
  nx53675z709_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z709_F5MUX,
      O => nx53675z709
    );
  nx53675z709_F5MUX_4403 : X_MUX2
    port map (
      IA => U2_ROME10_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx53675z710,
      SEL => nx53675z709_BXINV,
      O => nx53675z709_F5MUX
    );
  nx53675z709_BXINV_4404 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z709_BXINV
    );
  rome2datao10_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_2_F5MUX,
      O => U2_ROME10_modgen_rom_ix2_nx_ro64_32_l
    );
  rome2datao10_s_2_F5MUX_4405 : X_MUX2
    port map (
      IA => rome2datao10_s_2_G,
      IB => nx53675z714,
      SEL => rome2datao10_s_2_BXINV,
      O => rome2datao10_s_2_F5MUX
    );
  rome2datao10_s_2_BXINV_4406 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao10_s_2_BXINV
    );
  rome2datao10_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao10_s_2_F6MUX,
      O => rome2datao10_s(2)
    );
  rome2datao10_s_2_F6MUX_4407 : X_MUX2
    port map (
      IA => U2_ROME10_modgen_rom_ix2_nx_ro64_32_u,
      IB => U2_ROME10_modgen_rom_ix2_nx_ro64_32_l,
      SEL => rome2datao10_s_2_BYINV,
      O => rome2datao10_s_2_F6MUX
    );
  rome2datao10_s_2_BYINV_4408 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao10_s_2_BYINV
    );
  U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U2_ROME10_modgen_rom_ix2_nx_ro64_32_u
    );
  U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_F5MUX_4409 : X_MUX2
    port map (
      IA => U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U2_ROME10_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_BXINV_4410 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  rome2datao5_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_13_F5MUX,
      O => nx53675z327
    );
  rome2datao5_s_13_F5MUX_4411 : X_MUX2
    port map (
      IA => nx53675z328,
      IB => nx53675z329,
      SEL => rome2datao5_s_13_BXINV,
      O => rome2datao5_s_13_F5MUX
    );
  rome2datao5_s_13_BXINV_4412 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao5_s_13_BXINV
    );
  rome2datao5_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_13_F6MUX,
      O => rome2datao5_s(13)
    );
  rome2datao5_s_13_F6MUX_4413 : X_MUX2
    port map (
      IA => nx53675z325,
      IB => nx53675z327,
      SEL => rome2datao5_s_13_BYINV,
      O => rome2datao5_s_13_F6MUX
    );
  rome2datao5_s_13_BYINV_4414 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao5_s_13_BYINV
    );
  nx53675z325_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z325_F5MUX,
      O => nx53675z325
    );
  nx53675z325_F5MUX_4415 : X_MUX2
    port map (
      IA => nx53675z325_G,
      IB => nx53675z326,
      SEL => nx53675z325_BXINV,
      O => nx53675z325_F5MUX
    );
  nx53675z325_BXINV_4416 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z325_BXINV
    );
  rome2datao2_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_12_F5MUX,
      O => nx53675z138
    );
  rome2datao2_s_12_F5MUX_4417 : X_MUX2
    port map (
      IA => nx53675z139,
      IB => nx53675z140,
      SEL => rome2datao2_s_12_BXINV,
      O => rome2datao2_s_12_F5MUX
    );
  rome2datao2_s_12_BXINV_4418 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao2_s_12_BXINV
    );
  rome2datao2_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_12_F6MUX,
      O => rome2datao2_s(12)
    );
  rome2datao2_s_12_F6MUX_4419 : X_MUX2
    port map (
      IA => nx53675z135,
      IB => nx53675z138,
      SEL => rome2datao2_s_12_BYINV,
      O => rome2datao2_s_12_F6MUX
    );
  rome2datao2_s_12_BYINV_4420 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao2_s_12_BYINV
    );
  nx53675z135_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z135_F5MUX,
      O => nx53675z135
    );
  nx53675z135_F5MUX_4421 : X_MUX2
    port map (
      IA => nx53675z136,
      IB => nx53675z137,
      SEL => nx53675z135_BXINV,
      O => nx53675z135_F5MUX
    );
  nx53675z135_BXINV_4422 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z135_BXINV
    );
  rome2datao2_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_11_F5MUX,
      O => nx53675z144
    );
  rome2datao2_s_11_F5MUX_4423 : X_MUX2
    port map (
      IA => nx53675z145,
      IB => nx53675z146,
      SEL => rome2datao2_s_11_BXINV,
      O => rome2datao2_s_11_F5MUX
    );
  rome2datao2_s_11_BXINV_4424 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao2_s_11_BXINV
    );
  rome2datao2_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_11_F6MUX,
      O => rome2datao2_s(11)
    );
  rome2datao2_s_11_F6MUX_4425 : X_MUX2
    port map (
      IA => nx53675z141,
      IB => nx53675z144,
      SEL => rome2datao2_s_11_BYINV,
      O => rome2datao2_s_11_F6MUX
    );
  rome2datao2_s_11_BYINV_4426 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao2_s_11_BYINV
    );
  nx53675z141_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z141_F5MUX,
      O => nx53675z141
    );
  nx53675z141_F5MUX_4427 : X_MUX2
    port map (
      IA => nx53675z142,
      IB => nx53675z143,
      SEL => nx53675z141_BXINV,
      O => nx53675z141_F5MUX
    );
  nx53675z141_BXINV_4428 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z141_BXINV
    );
  rome2datao2_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_10_F5MUX,
      O => nx53675z150
    );
  rome2datao2_s_10_F5MUX_4429 : X_MUX2
    port map (
      IA => nx53675z151,
      IB => nx53675z152,
      SEL => rome2datao2_s_10_BXINV,
      O => rome2datao2_s_10_F5MUX
    );
  rome2datao2_s_10_BXINV_4430 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao2_s_10_BXINV
    );
  rome2datao2_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_10_F6MUX,
      O => rome2datao2_s(10)
    );
  rome2datao2_s_10_F6MUX_4431 : X_MUX2
    port map (
      IA => nx53675z147,
      IB => nx53675z150,
      SEL => rome2datao2_s_10_BYINV,
      O => rome2datao2_s_10_F6MUX
    );
  rome2datao2_s_10_BYINV_4432 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao2_s_10_BYINV
    );
  U_DCT2D_reg_databuf_reg_2_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_2_6_DYMUX,
      CE => U_DCT2D_databuf_reg_2_6_CEINV,
      CLK => U_DCT2D_databuf_reg_2_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_2_6_FFY_RST,
      O => U_DCT2D_databuf_reg_2_Q(7)
    );
  U_DCT2D_databuf_reg_2_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_2_6_FFY_RST
    );
  nx53675z147_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z147_F5MUX,
      O => nx53675z147
    );
  nx53675z147_F5MUX_4433 : X_MUX2
    port map (
      IA => nx53675z148,
      IB => nx53675z149,
      SEL => nx53675z147_BXINV,
      O => nx53675z147_F5MUX
    );
  nx53675z147_BXINV_4434 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z147_BXINV
    );
  rome2datao2_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_9_F5MUX,
      O => nx53675z156
    );
  rome2datao2_s_9_F5MUX_4435 : X_MUX2
    port map (
      IA => nx53675z157,
      IB => nx53675z158,
      SEL => rome2datao2_s_9_BXINV,
      O => rome2datao2_s_9_F5MUX
    );
  rome2datao2_s_9_BXINV_4436 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao2_s_9_BXINV
    );
  rome2datao2_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_9_F6MUX,
      O => rome2datao2_s(9)
    );
  rome2datao2_s_9_F6MUX_4437 : X_MUX2
    port map (
      IA => nx53675z153,
      IB => nx53675z156,
      SEL => rome2datao2_s_9_BYINV,
      O => rome2datao2_s_9_F6MUX
    );
  rome2datao2_s_9_BYINV_4438 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao2_s_9_BYINV
    );
  nx53675z153_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z153_F5MUX,
      O => nx53675z153
    );
  nx53675z153_F5MUX_4439 : X_MUX2
    port map (
      IA => nx53675z154,
      IB => nx53675z155,
      SEL => nx53675z153_BXINV,
      O => nx53675z153_F5MUX
    );
  nx53675z153_BXINV_4440 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z153_BXINV
    );
  rome2datao2_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_2_F5MUX,
      O => U2_ROME2_modgen_rom_ix2_nx_ro64_32_l
    );
  rome2datao2_s_2_F5MUX_4441 : X_MUX2
    port map (
      IA => rome2datao2_s_2_G,
      IB => nx53675z194,
      SEL => rome2datao2_s_2_BXINV,
      O => rome2datao2_s_2_F5MUX
    );
  rome2datao2_s_2_BXINV_4442 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao2_s_2_BXINV
    );
  rome2datao2_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao2_s_2_F6MUX,
      O => rome2datao2_s(2)
    );
  rome2datao2_s_2_F6MUX_4443 : X_MUX2
    port map (
      IA => U2_ROME2_modgen_rom_ix2_nx_ro64_32_u,
      IB => U2_ROME2_modgen_rom_ix2_nx_ro64_32_l,
      SEL => rome2datao2_s_2_BYINV,
      O => rome2datao2_s_2_F6MUX
    );
  rome2datao2_s_2_BYINV_4444 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao2_s_2_BYINV
    );
  U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U2_ROME2_modgen_rom_ix2_nx_ro64_32_u
    );
  U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_F5MUX_4445 : X_MUX2
    port map (
      IA => U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U2_ROME2_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_BXINV_4446 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  romo2datao9_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_11_F5MUX,
      O => nx53675z1438
    );
  romo2datao9_s_11_F5MUX_4447 : X_MUX2
    port map (
      IA => nx53675z1439,
      IB => nx53675z1440,
      SEL => romo2datao9_s_11_BXINV,
      O => romo2datao9_s_11_F5MUX
    );
  romo2datao9_s_11_BXINV_4448 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_11_BXINV
    );
  romo2datao9_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_11_F6MUX,
      O => romo2datao9_s(11)
    );
  romo2datao9_s_11_F6MUX_4449 : X_MUX2
    port map (
      IA => nx53675z1435,
      IB => nx53675z1438,
      SEL => romo2datao9_s_11_BYINV,
      O => romo2datao9_s_11_F6MUX
    );
  romo2datao9_s_11_BYINV_4450 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_11_BYINV
    );
  nx53675z1435_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1435_F5MUX,
      O => nx53675z1435
    );
  nx53675z1435_F5MUX_4451 : X_MUX2
    port map (
      IA => nx53675z1436,
      IB => nx53675z1437,
      SEL => nx53675z1435_BXINV,
      O => nx53675z1435_F5MUX
    );
  nx53675z1435_BXINV_4452 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1435_BXINV
    );
  romo2datao9_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_10_F5MUX,
      O => nx53675z1444
    );
  romo2datao9_s_10_F5MUX_4453 : X_MUX2
    port map (
      IA => nx53675z1445,
      IB => nx53675z1446,
      SEL => romo2datao9_s_10_BXINV,
      O => romo2datao9_s_10_F5MUX
    );
  romo2datao9_s_10_BXINV_4454 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_10_BXINV
    );
  romo2datao9_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_10_F6MUX,
      O => romo2datao9_s(10)
    );
  romo2datao9_s_10_F6MUX_4455 : X_MUX2
    port map (
      IA => nx53675z1441,
      IB => nx53675z1444,
      SEL => romo2datao9_s_10_BYINV,
      O => romo2datao9_s_10_F6MUX
    );
  romo2datao9_s_10_BYINV_4456 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_10_BYINV
    );
  nx53675z1441_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1441_F5MUX,
      O => nx53675z1441
    );
  nx53675z1441_F5MUX_4457 : X_MUX2
    port map (
      IA => nx53675z1442,
      IB => nx53675z1443,
      SEL => nx53675z1441_BXINV,
      O => nx53675z1441_F5MUX
    );
  nx53675z1441_BXINV_4458 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1441_BXINV
    );
  romo2datao9_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_9_F5MUX,
      O => nx53675z1450
    );
  romo2datao9_s_9_F5MUX_4459 : X_MUX2
    port map (
      IA => nx53675z1451,
      IB => nx53675z1452,
      SEL => romo2datao9_s_9_BXINV,
      O => romo2datao9_s_9_F5MUX
    );
  romo2datao9_s_9_BXINV_4460 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_9_BXINV
    );
  romo2datao9_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_9_F6MUX,
      O => romo2datao9_s(9)
    );
  romo2datao9_s_9_F6MUX_4461 : X_MUX2
    port map (
      IA => nx53675z1447,
      IB => nx53675z1450,
      SEL => romo2datao9_s_9_BYINV,
      O => romo2datao9_s_9_F6MUX
    );
  romo2datao9_s_9_BYINV_4462 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_9_BYINV
    );
  U_DCT2D_ix268z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_2_6_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_5_6_Q,
      O => U_DCT2D_nx268z1
    );
  nx53675z1447_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1447_F5MUX,
      O => nx53675z1447
    );
  nx53675z1447_F5MUX_4463 : X_MUX2
    port map (
      IA => nx53675z1448,
      IB => nx53675z1449,
      SEL => nx53675z1447_BXINV,
      O => nx53675z1447_F5MUX
    );
  nx53675z1447_BXINV_4464 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1447_BXINV
    );
  romo2datao9_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_8_F5MUX,
      O => nx53675z1456
    );
  romo2datao9_s_8_F5MUX_4465 : X_MUX2
    port map (
      IA => nx53675z1457,
      IB => nx53675z1458,
      SEL => romo2datao9_s_8_BXINV,
      O => romo2datao9_s_8_F5MUX
    );
  romo2datao9_s_8_BXINV_4466 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_8_BXINV
    );
  romo2datao9_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_8_F6MUX,
      O => romo2datao9_s(8)
    );
  romo2datao9_s_8_F6MUX_4467 : X_MUX2
    port map (
      IA => nx53675z1453,
      IB => nx53675z1456,
      SEL => romo2datao9_s_8_BYINV,
      O => romo2datao9_s_8_F6MUX
    );
  romo2datao9_s_8_BYINV_4468 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_8_BYINV
    );
  nx53675z1453_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1453_F5MUX,
      O => nx53675z1453
    );
  nx53675z1453_F5MUX_4469 : X_MUX2
    port map (
      IA => nx53675z1454,
      IB => nx53675z1455,
      SEL => nx53675z1453_BXINV,
      O => nx53675z1453_F5MUX
    );
  nx53675z1453_BXINV_4470 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1453_BXINV
    );
  romo2datao9_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_7_F5MUX,
      O => nx53675z1462
    );
  romo2datao9_s_7_F5MUX_4471 : X_MUX2
    port map (
      IA => nx53675z1463,
      IB => nx53675z1464,
      SEL => romo2datao9_s_7_BXINV,
      O => romo2datao9_s_7_F5MUX
    );
  romo2datao9_s_7_BXINV_4472 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_7_BXINV
    );
  romo2datao9_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_7_F6MUX,
      O => romo2datao9_s(7)
    );
  romo2datao9_s_7_F6MUX_4473 : X_MUX2
    port map (
      IA => nx53675z1459,
      IB => nx53675z1462,
      SEL => romo2datao9_s_7_BYINV,
      O => romo2datao9_s_7_F6MUX
    );
  romo2datao9_s_7_BYINV_4474 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_7_BYINV
    );
  nx53675z1459_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1459_F5MUX,
      O => nx53675z1459
    );
  nx53675z1459_F5MUX_4475 : X_MUX2
    port map (
      IA => nx53675z1460,
      IB => nx53675z1461,
      SEL => nx53675z1459_BXINV,
      O => nx53675z1459_F5MUX
    );
  nx53675z1459_BXINV_4476 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1459_BXINV
    );
  rome2datao6_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_13_F5MUX,
      O => nx53675z392
    );
  rome2datao6_s_13_F5MUX_4477 : X_MUX2
    port map (
      IA => nx53675z393,
      IB => nx53675z394,
      SEL => rome2datao6_s_13_BXINV,
      O => rome2datao6_s_13_F5MUX
    );
  rome2datao6_s_13_BXINV_4478 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao6_s_13_BXINV
    );
  rome2datao6_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_13_F6MUX,
      O => rome2datao6_s(13)
    );
  rome2datao6_s_13_F6MUX_4479 : X_MUX2
    port map (
      IA => nx53675z390,
      IB => nx53675z392,
      SEL => rome2datao6_s_13_BYINV,
      O => rome2datao6_s_13_F6MUX
    );
  rome2datao6_s_13_BYINV_4480 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao6_s_13_BYINV
    );
  nx53675z390_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z390_F5MUX,
      O => nx53675z390
    );
  nx53675z390_F5MUX_4481 : X_MUX2
    port map (
      IA => nx53675z390_G,
      IB => nx53675z391,
      SEL => nx53675z390_BXINV,
      O => nx53675z390_F5MUX
    );
  nx53675z390_BXINV_4482 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z390_BXINV
    );
  rome2datao4_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_12_F5MUX,
      O => nx53675z268
    );
  rome2datao4_s_12_F5MUX_4483 : X_MUX2
    port map (
      IA => nx53675z269,
      IB => nx53675z270,
      SEL => rome2datao4_s_12_BXINV,
      O => rome2datao4_s_12_F5MUX
    );
  rome2datao4_s_12_BXINV_4484 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao4_s_12_BXINV
    );
  rome2datao4_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_12_F6MUX,
      O => rome2datao4_s(12)
    );
  rome2datao4_s_12_F6MUX_4485 : X_MUX2
    port map (
      IA => nx53675z265,
      IB => nx53675z268,
      SEL => rome2datao4_s_12_BYINV,
      O => rome2datao4_s_12_F6MUX
    );
  rome2datao4_s_12_BYINV_4486 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao4_s_12_BYINV
    );
  nx53675z265_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z265_F5MUX,
      O => nx53675z265
    );
  nx53675z265_F5MUX_4487 : X_MUX2
    port map (
      IA => nx53675z266,
      IB => nx53675z267,
      SEL => nx53675z265_BXINV,
      O => nx53675z265_F5MUX
    );
  nx53675z265_BXINV_4488 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z265_BXINV
    );
  rome2datao4_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_11_F5MUX,
      O => nx53675z274
    );
  rome2datao4_s_11_F5MUX_4489 : X_MUX2
    port map (
      IA => nx53675z275,
      IB => nx53675z276,
      SEL => rome2datao4_s_11_BXINV,
      O => rome2datao4_s_11_F5MUX
    );
  rome2datao4_s_11_BXINV_4490 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao4_s_11_BXINV
    );
  rome2datao4_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_11_F6MUX,
      O => rome2datao4_s(11)
    );
  rome2datao4_s_11_F6MUX_4491 : X_MUX2
    port map (
      IA => nx53675z271,
      IB => nx53675z274,
      SEL => rome2datao4_s_11_BYINV,
      O => rome2datao4_s_11_F6MUX
    );
  rome2datao4_s_11_BYINV_4492 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao4_s_11_BYINV
    );
  nx53675z271_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z271_F5MUX,
      O => nx53675z271
    );
  nx53675z271_F5MUX_4493 : X_MUX2
    port map (
      IA => nx53675z272,
      IB => nx53675z273,
      SEL => nx53675z271_BXINV,
      O => nx53675z271_F5MUX
    );
  nx53675z271_BXINV_4494 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z271_BXINV
    );
  rome2datao4_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_10_F5MUX,
      O => nx53675z280
    );
  rome2datao4_s_10_F5MUX_4495 : X_MUX2
    port map (
      IA => nx53675z281,
      IB => nx53675z282,
      SEL => rome2datao4_s_10_BXINV,
      O => rome2datao4_s_10_F5MUX
    );
  rome2datao4_s_10_BXINV_4496 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao4_s_10_BXINV
    );
  rome2datao4_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_10_F6MUX,
      O => rome2datao4_s(10)
    );
  rome2datao4_s_10_F6MUX_4497 : X_MUX2
    port map (
      IA => nx53675z277,
      IB => nx53675z280,
      SEL => rome2datao4_s_10_BYINV,
      O => rome2datao4_s_10_F6MUX
    );
  rome2datao4_s_10_BYINV_4498 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao4_s_10_BYINV
    );
  nx53675z277_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z277_F5MUX,
      O => nx53675z277
    );
  nx53675z277_F5MUX_4499 : X_MUX2
    port map (
      IA => nx53675z278,
      IB => nx53675z279,
      SEL => nx53675z277_BXINV,
      O => nx53675z277_F5MUX
    );
  nx53675z277_BXINV_4500 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z277_BXINV
    );
  rome2datao4_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_4_F5MUX,
      O => nx53675z316
    );
  rome2datao4_s_4_F5MUX_4501 : X_MUX2
    port map (
      IA => nx53675z317,
      IB => nx53675z318,
      SEL => rome2datao4_s_4_BXINV,
      O => rome2datao4_s_4_F5MUX
    );
  rome2datao4_s_4_BXINV_4502 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao4_s_4_BXINV
    );
  rome2datao4_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_4_F6MUX,
      O => rome2datao4_s(4)
    );
  rome2datao4_s_4_F6MUX_4503 : X_MUX2
    port map (
      IA => nx53675z313,
      IB => nx53675z316,
      SEL => rome2datao4_s_4_BYINV,
      O => rome2datao4_s_4_F6MUX
    );
  rome2datao4_s_4_BYINV_4504 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao4_s_4_BYINV
    );
  nx53675z313_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z313_F5MUX,
      O => nx53675z313
    );
  nx53675z313_F5MUX_4505 : X_MUX2
    port map (
      IA => nx53675z314,
      IB => nx53675z315,
      SEL => nx53675z313_BXINV,
      O => nx53675z313_F5MUX
    );
  nx53675z313_BXINV_4506 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z313_BXINV
    );
  rome2datao4_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_3_F5MUX,
      O => nx53675z321
    );
  rome2datao4_s_3_F5MUX_4507 : X_MUX2
    port map (
      IA => nx53675z322,
      IB => nx53675z323,
      SEL => rome2datao4_s_3_BXINV,
      O => rome2datao4_s_3_F5MUX
    );
  rome2datao4_s_3_BXINV_4508 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao4_s_3_BXINV
    );
  rome2datao4_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_3_F6MUX,
      O => rome2datao4_s(3)
    );
  rome2datao4_s_3_F6MUX_4509 : X_MUX2
    port map (
      IA => nx53675z319,
      IB => nx53675z321,
      SEL => rome2datao4_s_3_BYINV,
      O => rome2datao4_s_3_F6MUX
    );
  rome2datao4_s_3_BYINV_4510 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao4_s_3_BYINV
    );
  nx53675z319_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z319_F5MUX,
      O => nx53675z319
    );
  nx53675z319_F5MUX_4511 : X_MUX2
    port map (
      IA => U2_ROME4_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx53675z320,
      SEL => nx53675z319_BXINV,
      O => nx53675z319_F5MUX
    );
  nx53675z319_BXINV_4512 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z319_BXINV
    );
  rome2datao4_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_2_F5MUX,
      O => U2_ROME4_modgen_rom_ix2_nx_ro64_32_l
    );
  rome2datao4_s_2_F5MUX_4513 : X_MUX2
    port map (
      IA => rome2datao4_s_2_G,
      IB => nx53675z324,
      SEL => rome2datao4_s_2_BXINV,
      O => rome2datao4_s_2_F5MUX
    );
  rome2datao4_s_2_BXINV_4514 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao4_s_2_BXINV
    );
  rome2datao4_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_2_F6MUX,
      O => rome2datao4_s(2)
    );
  rome2datao4_s_2_F6MUX_4515 : X_MUX2
    port map (
      IA => U2_ROME4_modgen_rom_ix2_nx_ro64_32_u,
      IB => U2_ROME4_modgen_rom_ix2_nx_ro64_32_l,
      SEL => rome2datao4_s_2_BYINV,
      O => rome2datao4_s_2_F6MUX
    );
  rome2datao4_s_2_BYINV_4516 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao4_s_2_BYINV
    );
  U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U2_ROME4_modgen_rom_ix2_nx_ro64_32_u
    );
  U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_F5MUX_4517 : X_MUX2
    port map (
      IA => U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U2_ROME4_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_BXINV_4518 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  rome2datao1_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_9_F5MUX,
      O => nx53675z91
    );
  rome2datao1_s_9_F5MUX_4519 : X_MUX2
    port map (
      IA => nx53675z92,
      IB => nx53675z93,
      SEL => rome2datao1_s_9_BXINV,
      O => rome2datao1_s_9_F5MUX
    );
  rome2datao1_s_9_BXINV_4520 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao1_s_9_BXINV
    );
  rome2datao1_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao1_s_9_F6MUX,
      O => rome2datao1_s(9)
    );
  rome2datao1_s_9_F6MUX_4521 : X_MUX2
    port map (
      IA => nx53675z88,
      IB => nx53675z91,
      SEL => rome2datao1_s_9_BYINV,
      O => rome2datao1_s_9_F6MUX
    );
  rome2datao1_s_9_BYINV_4522 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao1_s_9_BYINV
    );
  U_DCT2D_reg_databuf_reg_2_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_2_6_DXMUX,
      CE => U_DCT2D_databuf_reg_2_6_CEINV,
      CLK => U_DCT2D_databuf_reg_2_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_2_6_FFX_RST,
      O => U_DCT2D_databuf_reg_2_Q(6)
    );
  U_DCT2D_databuf_reg_2_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_2_6_FFX_RST
    );
  nx53675z88_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z88_F5MUX,
      O => nx53675z88
    );
  nx53675z88_F5MUX_4523 : X_MUX2
    port map (
      IA => nx53675z89,
      IB => nx53675z90,
      SEL => nx53675z88_BXINV,
      O => nx53675z88_F5MUX
    );
  nx53675z88_BXINV_4524 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z88_BXINV
    );
  romo2datao10_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_12_F5MUX,
      O => nx53675z1511
    );
  romo2datao10_s_12_F5MUX_4525 : X_MUX2
    port map (
      IA => nx53675z1512,
      IB => nx53675z1513,
      SEL => romo2datao10_s_12_BXINV,
      O => romo2datao10_s_12_F5MUX
    );
  romo2datao10_s_12_BXINV_4526 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_12_BXINV
    );
  romo2datao10_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_12_F6MUX,
      O => romo2datao10_s(12)
    );
  romo2datao10_s_12_F6MUX_4527 : X_MUX2
    port map (
      IA => nx53675z1508,
      IB => nx53675z1511,
      SEL => romo2datao10_s_12_BYINV,
      O => romo2datao10_s_12_F6MUX
    );
  romo2datao10_s_12_BYINV_4528 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_12_BYINV
    );
  ix53675z60805 : X_LUT4
    generic map(
      INIT => X"C080"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1509
    );
  nx53675z1508_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1508_F5MUX,
      O => nx53675z1508
    );
  nx53675z1508_F5MUX_4529 : X_MUX2
    port map (
      IA => nx53675z1509,
      IB => nx53675z1510,
      SEL => nx53675z1508_BXINV,
      O => nx53675z1508_F5MUX
    );
  nx53675z1508_BXINV_4530 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1508_BXINV
    );
  U_DCT2D_ix3259z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_5_10_Q,
      ADR1 => U_DCT2D_latchbuf_reg_2_10_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx3259z1
    );
  romo2datao3_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_12_F5MUX,
      O => nx53675z958
    );
  romo2datao3_s_12_F5MUX_4531 : X_MUX2
    port map (
      IA => nx53675z959,
      IB => nx53675z960,
      SEL => romo2datao3_s_12_BXINV,
      O => romo2datao3_s_12_F5MUX
    );
  romo2datao3_s_12_BXINV_4532 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_12_BXINV
    );
  romo2datao3_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_12_F6MUX,
      O => romo2datao3_s(12)
    );
  romo2datao3_s_12_F6MUX_4533 : X_MUX2
    port map (
      IA => nx53675z955,
      IB => nx53675z958,
      SEL => romo2datao3_s_12_BYINV,
      O => romo2datao3_s_12_F6MUX
    );
  romo2datao3_s_12_BYINV_4534 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_12_BYINV
    );
  nx53675z955_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z955_F5MUX,
      O => nx53675z955
    );
  nx53675z955_F5MUX_4535 : X_MUX2
    port map (
      IA => nx53675z956,
      IB => nx53675z957,
      SEL => nx53675z955_BXINV,
      O => nx53675z955_F5MUX
    );
  nx53675z955_BXINV_4536 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z955_BXINV
    );
  romo2datao3_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_2_F5MUX,
      O => nx53675z1018
    );
  romo2datao3_s_2_F5MUX_4537 : X_MUX2
    port map (
      IA => nx53675z1019,
      IB => nx53675z1020,
      SEL => romo2datao3_s_2_BXINV,
      O => romo2datao3_s_2_F5MUX
    );
  romo2datao3_s_2_BXINV_4538 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_2_BXINV
    );
  romo2datao3_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_2_F6MUX,
      O => romo2datao3_s(2)
    );
  romo2datao3_s_2_F6MUX_4539 : X_MUX2
    port map (
      IA => nx53675z1015,
      IB => nx53675z1018,
      SEL => romo2datao3_s_2_BYINV,
      O => romo2datao3_s_2_F6MUX
    );
  romo2datao3_s_2_BYINV_4540 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_2_BYINV
    );
  nx53675z1015_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1015_F5MUX,
      O => nx53675z1015
    );
  nx53675z1015_F5MUX_4541 : X_MUX2
    port map (
      IA => nx53675z1016,
      IB => nx53675z1017,
      SEL => nx53675z1015_BXINV,
      O => nx53675z1015_F5MUX
    );
  nx53675z1015_BXINV_4542 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1015_BXINV
    );
  romo2datao2_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_12_F5MUX,
      O => nx53675z879
    );
  romo2datao2_s_12_F5MUX_4543 : X_MUX2
    port map (
      IA => nx53675z880,
      IB => nx53675z881,
      SEL => romo2datao2_s_12_BXINV,
      O => romo2datao2_s_12_F5MUX
    );
  romo2datao2_s_12_BXINV_4544 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_12_BXINV
    );
  romo2datao2_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_12_F6MUX,
      O => romo2datao2_s(12)
    );
  romo2datao2_s_12_F6MUX_4545 : X_MUX2
    port map (
      IA => nx53675z876,
      IB => nx53675z879,
      SEL => romo2datao2_s_12_BYINV,
      O => romo2datao2_s_12_F6MUX
    );
  romo2datao2_s_12_BYINV_4546 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_12_BYINV
    );
  nx53675z876_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z876_F5MUX,
      O => nx53675z876
    );
  nx53675z876_F5MUX_4547 : X_MUX2
    port map (
      IA => nx53675z877,
      IB => nx53675z878,
      SEL => nx53675z876_BXINV,
      O => nx53675z876_F5MUX
    );
  nx53675z876_BXINV_4548 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z876_BXINV
    );
  romo2datao2_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_11_F5MUX,
      O => nx53675z885
    );
  romo2datao2_s_11_F5MUX_4549 : X_MUX2
    port map (
      IA => nx53675z886,
      IB => nx53675z887,
      SEL => romo2datao2_s_11_BXINV,
      O => romo2datao2_s_11_F5MUX
    );
  romo2datao2_s_11_BXINV_4550 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_11_BXINV
    );
  romo2datao2_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_11_F6MUX,
      O => romo2datao2_s(11)
    );
  romo2datao2_s_11_F6MUX_4551 : X_MUX2
    port map (
      IA => nx53675z882,
      IB => nx53675z885,
      SEL => romo2datao2_s_11_BYINV,
      O => romo2datao2_s_11_F6MUX
    );
  romo2datao2_s_11_BYINV_4552 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_11_BYINV
    );
  nx53675z882_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z882_F5MUX,
      O => nx53675z882
    );
  nx53675z882_F5MUX_4553 : X_MUX2
    port map (
      IA => nx53675z883,
      IB => nx53675z884,
      SEL => nx53675z882_BXINV,
      O => nx53675z882_F5MUX
    );
  nx53675z882_BXINV_4554 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z882_BXINV
    );
  romo2datao2_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_10_F5MUX,
      O => nx53675z891
    );
  romo2datao2_s_10_F5MUX_4555 : X_MUX2
    port map (
      IA => nx53675z892,
      IB => nx53675z893,
      SEL => romo2datao2_s_10_BXINV,
      O => romo2datao2_s_10_F5MUX
    );
  romo2datao2_s_10_BXINV_4556 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_10_BXINV
    );
  romo2datao2_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_10_F6MUX,
      O => romo2datao2_s(10)
    );
  romo2datao2_s_10_F6MUX_4557 : X_MUX2
    port map (
      IA => nx53675z888,
      IB => nx53675z891,
      SEL => romo2datao2_s_10_BYINV,
      O => romo2datao2_s_10_F6MUX
    );
  romo2datao2_s_10_BYINV_4558 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_10_BYINV
    );
  nx53675z888_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z888_F5MUX,
      O => nx53675z888
    );
  nx53675z888_F5MUX_4559 : X_MUX2
    port map (
      IA => nx53675z889,
      IB => nx53675z890,
      SEL => nx53675z888_BXINV,
      O => nx53675z888_F5MUX
    );
  nx53675z888_BXINV_4560 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z888_BXINV
    );
  romo2datao2_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_9_F5MUX,
      O => nx53675z897
    );
  romo2datao2_s_9_F5MUX_4561 : X_MUX2
    port map (
      IA => nx53675z898,
      IB => nx53675z899,
      SEL => romo2datao2_s_9_BXINV,
      O => romo2datao2_s_9_F5MUX
    );
  romo2datao2_s_9_BXINV_4562 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_9_BXINV
    );
  romo2datao2_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_9_F6MUX,
      O => romo2datao2_s(9)
    );
  romo2datao2_s_9_F6MUX_4563 : X_MUX2
    port map (
      IA => nx53675z894,
      IB => nx53675z897,
      SEL => romo2datao2_s_9_BYINV,
      O => romo2datao2_s_9_F6MUX
    );
  romo2datao2_s_9_BYINV_4564 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_9_BYINV
    );
  nx53675z894_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z894_F5MUX,
      O => nx53675z894
    );
  nx53675z894_F5MUX_4565 : X_MUX2
    port map (
      IA => nx53675z895,
      IB => nx53675z896,
      SEL => nx53675z894_BXINV,
      O => nx53675z894_F5MUX
    );
  nx53675z894_BXINV_4566 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z894_BXINV
    );
  romo2datao2_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_8_F5MUX,
      O => nx53675z903
    );
  romo2datao2_s_8_F5MUX_4567 : X_MUX2
    port map (
      IA => nx53675z904,
      IB => nx53675z905,
      SEL => romo2datao2_s_8_BXINV,
      O => romo2datao2_s_8_F5MUX
    );
  romo2datao2_s_8_BXINV_4568 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_8_BXINV
    );
  romo2datao2_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_8_F6MUX,
      O => romo2datao2_s(8)
    );
  romo2datao2_s_8_F6MUX_4569 : X_MUX2
    port map (
      IA => nx53675z900,
      IB => nx53675z903,
      SEL => romo2datao2_s_8_BYINV,
      O => romo2datao2_s_8_F6MUX
    );
  romo2datao2_s_8_BYINV_4570 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_8_BYINV
    );
  nx53675z900_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z900_F5MUX,
      O => nx53675z900
    );
  nx53675z900_F5MUX_4571 : X_MUX2
    port map (
      IA => nx53675z901,
      IB => nx53675z902,
      SEL => nx53675z900_BXINV,
      O => nx53675z900_F5MUX
    );
  nx53675z900_BXINV_4572 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z900_BXINV
    );
  rome2datao9_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_2_F5MUX,
      O => U2_ROME9_modgen_rom_ix2_nx_ro64_32_l
    );
  rome2datao9_s_2_F5MUX_4573 : X_MUX2
    port map (
      IA => rome2datao9_s_2_G,
      IB => nx53675z649,
      SEL => rome2datao9_s_2_BXINV,
      O => rome2datao9_s_2_F5MUX
    );
  rome2datao9_s_2_BXINV_4574 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao9_s_2_BXINV
    );
  rome2datao9_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao9_s_2_F6MUX,
      O => rome2datao9_s(2)
    );
  rome2datao9_s_2_F6MUX_4575 : X_MUX2
    port map (
      IA => U2_ROME9_modgen_rom_ix2_nx_ro64_32_u,
      IB => U2_ROME9_modgen_rom_ix2_nx_ro64_32_l,
      SEL => rome2datao9_s_2_BYINV,
      O => rome2datao9_s_2_F6MUX
    );
  rome2datao9_s_2_BYINV_4576 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao9_s_2_BYINV
    );
  U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U2_ROME9_modgen_rom_ix2_nx_ro64_32_u
    );
  U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_F5MUX_4577 : X_MUX2
    port map (
      IA => U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U2_ROME9_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_BXINV_4578 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  romo2datao10_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_13_F5MUX,
      O => nx53675z1505
    );
  romo2datao10_s_13_F5MUX_4579 : X_MUX2
    port map (
      IA => nx53675z1506,
      IB => nx53675z1507,
      SEL => romo2datao10_s_13_BXINV,
      O => romo2datao10_s_13_F5MUX
    );
  romo2datao10_s_13_BXINV_4580 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_13_BXINV
    );
  romo2datao10_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_13_F6MUX,
      O => romo2datao10_s(13)
    );
  romo2datao10_s_13_F6MUX_4581 : X_MUX2
    port map (
      IA => nx53675z1503,
      IB => nx53675z1505,
      SEL => romo2datao10_s_13_BYINV,
      O => romo2datao10_s_13_F6MUX
    );
  romo2datao10_s_13_BYINV_4582 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_13_BYINV
    );
  nx53675z1503_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1503_F5MUX,
      O => nx53675z1503
    );
  nx53675z1503_F5MUX_4583 : X_MUX2
    port map (
      IA => nx53675z1503_G,
      IB => nx53675z1504,
      SEL => nx53675z1503_BXINV,
      O => nx53675z1503_F5MUX
    );
  nx53675z1503_BXINV_4584 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1503_BXINV
    );
  romo2datao10_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_10_F5MUX,
      O => nx53675z1523
    );
  romo2datao10_s_10_F5MUX_4585 : X_MUX2
    port map (
      IA => nx53675z1524,
      IB => nx53675z1525,
      SEL => romo2datao10_s_10_BXINV,
      O => romo2datao10_s_10_F5MUX
    );
  romo2datao10_s_10_BXINV_4586 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_10_BXINV
    );
  romo2datao10_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_10_F6MUX,
      O => romo2datao10_s(10)
    );
  romo2datao10_s_10_F6MUX_4587 : X_MUX2
    port map (
      IA => nx53675z1520,
      IB => nx53675z1523,
      SEL => romo2datao10_s_10_BYINV,
      O => romo2datao10_s_10_F6MUX
    );
  romo2datao10_s_10_BYINV_4588 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_10_BYINV
    );
  nx53675z1520_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1520_F5MUX,
      O => nx53675z1520
    );
  nx53675z1520_F5MUX_4589 : X_MUX2
    port map (
      IA => nx53675z1521,
      IB => nx53675z1522,
      SEL => nx53675z1520_BXINV,
      O => nx53675z1520_F5MUX
    );
  nx53675z1520_BXINV_4590 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1520_BXINV
    );
  romo2datao10_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_2_F5MUX,
      O => nx53675z1571
    );
  romo2datao10_s_2_F5MUX_4591 : X_MUX2
    port map (
      IA => nx53675z1572,
      IB => nx53675z1573,
      SEL => romo2datao10_s_2_BXINV,
      O => romo2datao10_s_2_F5MUX
    );
  romo2datao10_s_2_BXINV_4592 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_2_BXINV
    );
  romo2datao10_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_2_F6MUX,
      O => romo2datao10_s(2)
    );
  romo2datao10_s_2_F6MUX_4593 : X_MUX2
    port map (
      IA => nx53675z1568,
      IB => nx53675z1571,
      SEL => romo2datao10_s_2_BYINV,
      O => romo2datao10_s_2_F6MUX
    );
  romo2datao10_s_2_BYINV_4594 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_2_BYINV
    );
  nx53675z1568_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1568_F5MUX,
      O => nx53675z1568
    );
  nx53675z1568_F5MUX_4595 : X_MUX2
    port map (
      IA => nx53675z1569,
      IB => nx53675z1570,
      SEL => nx53675z1568_BXINV,
      O => nx53675z1568_F5MUX
    );
  nx53675z1568_BXINV_4596 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1568_BXINV
    );
  romo2datao10_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_1_F5MUX,
      O => nx53675z1577
    );
  romo2datao10_s_1_F5MUX_4597 : X_MUX2
    port map (
      IA => nx53675z1578,
      IB => nx53675z1579,
      SEL => romo2datao10_s_1_BXINV,
      O => romo2datao10_s_1_F5MUX
    );
  romo2datao10_s_1_BXINV_4598 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_1_BXINV
    );
  romo2datao10_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_1_F6MUX,
      O => romo2datao10_s(1)
    );
  romo2datao10_s_1_F6MUX_4599 : X_MUX2
    port map (
      IA => nx53675z1574,
      IB => nx53675z1577,
      SEL => romo2datao10_s_1_BYINV,
      O => romo2datao10_s_1_F6MUX
    );
  romo2datao10_s_1_BYINV_4600 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_1_BYINV
    );
  nx53675z1574_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1574_F5MUX,
      O => nx53675z1574
    );
  nx53675z1574_F5MUX_4601 : X_MUX2
    port map (
      IA => nx53675z1575,
      IB => nx53675z1576,
      SEL => nx53675z1574_BXINV,
      O => nx53675z1574_F5MUX
    );
  nx53675z1574_BXINV_4602 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1574_BXINV
    );
  romo2datao10_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_0_F5MUX,
      O => U2_ROMO10_modgen_rom_ix0_nx_ro64_32_l
    );
  romo2datao10_s_0_F5MUX_4603 : X_MUX2
    port map (
      IA => nx53675z1580,
      IB => nx53675z1581,
      SEL => romo2datao10_s_0_BXINV,
      O => romo2datao10_s_0_F5MUX
    );
  romo2datao10_s_0_BXINV_4604 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_0_BXINV
    );
  romo2datao10_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_0_F6MUX,
      O => romo2datao10_s(0)
    );
  romo2datao10_s_0_F6MUX_4605 : X_MUX2
    port map (
      IA => U2_ROMO10_modgen_rom_ix0_nx_ro64_32_u,
      IB => U2_ROMO10_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romo2datao10_s_0_BYINV,
      O => romo2datao10_s_0_F6MUX
    );
  romo2datao10_s_0_BYINV_4606 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_0_BYINV
    );
  U2_ROMO10_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROMO10_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U2_ROMO10_modgen_rom_ix0_nx_ro64_32_u
    );
  U2_ROMO10_modgen_rom_ix0_nx_ro64_32_u_F5MUX_4607 : X_MUX2
    port map (
      IA => U2_ROMO10_modgen_rom_ix0_nx_rm64_16_u,
      IB => U2_ROMO10_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U2_ROMO10_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U2_ROMO10_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U2_ROMO10_modgen_rom_ix0_nx_ro64_32_u_BXINV_4608 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => U2_ROMO10_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romo2datao9_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_0_F5MUX,
      O => U2_ROMO9_modgen_rom_ix0_nx_ro64_32_l
    );
  romo2datao9_s_0_F5MUX_4609 : X_MUX2
    port map (
      IA => nx53675z1501,
      IB => nx53675z1502,
      SEL => romo2datao9_s_0_BXINV,
      O => romo2datao9_s_0_F5MUX
    );
  romo2datao9_s_0_BXINV_4610 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_0_BXINV
    );
  romo2datao9_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_0_F6MUX,
      O => romo2datao9_s(0)
    );
  romo2datao9_s_0_F6MUX_4611 : X_MUX2
    port map (
      IA => U2_ROMO9_modgen_rom_ix0_nx_ro64_32_u,
      IB => U2_ROMO9_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romo2datao9_s_0_BYINV,
      O => romo2datao9_s_0_F6MUX
    );
  romo2datao9_s_0_BYINV_4612 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_0_BYINV
    );
  U2_ROMO9_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROMO9_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U2_ROMO9_modgen_rom_ix0_nx_ro64_32_u
    );
  U2_ROMO9_modgen_rom_ix0_nx_ro64_32_u_F5MUX_4613 : X_MUX2
    port map (
      IA => U2_ROMO9_modgen_rom_ix0_nx_rm64_16_u,
      IB => U2_ROMO9_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U2_ROMO9_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U2_ROMO9_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U2_ROMO9_modgen_rom_ix0_nx_ro64_32_u_BXINV_4614 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => U2_ROMO9_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romo2datao4_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_5_F5MUX,
      O => nx53675z1079
    );
  romo2datao4_s_5_F5MUX_4615 : X_MUX2
    port map (
      IA => nx53675z1080,
      IB => nx53675z1081,
      SEL => romo2datao4_s_5_BXINV,
      O => romo2datao4_s_5_F5MUX
    );
  romo2datao4_s_5_BXINV_4616 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_5_BXINV
    );
  romo2datao4_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_5_F6MUX,
      O => romo2datao4_s(5)
    );
  romo2datao4_s_5_F6MUX_4617 : X_MUX2
    port map (
      IA => nx53675z1076,
      IB => nx53675z1079,
      SEL => romo2datao4_s_5_BYINV,
      O => romo2datao4_s_5_F6MUX
    );
  romo2datao4_s_5_BYINV_4618 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_5_BYINV
    );
  ix53675z19914 : X_LUT4
    generic map(
      INIT => X"4964"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1077
    );
  nx53675z1076_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1076_F5MUX,
      O => nx53675z1076
    );
  nx53675z1076_F5MUX_4619 : X_MUX2
    port map (
      IA => nx53675z1077,
      IB => nx53675z1078,
      SEL => nx53675z1076_BXINV,
      O => nx53675z1076_F5MUX
    );
  nx53675z1076_BXINV_4620 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1076_BXINV
    );
  romo2datao3_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_13_F5MUX,
      O => nx53675z952
    );
  romo2datao3_s_13_F5MUX_4621 : X_MUX2
    port map (
      IA => nx53675z953,
      IB => nx53675z954,
      SEL => romo2datao3_s_13_BXINV,
      O => romo2datao3_s_13_F5MUX
    );
  romo2datao3_s_13_BXINV_4622 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_13_BXINV
    );
  romo2datao3_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_13_F6MUX,
      O => romo2datao3_s(13)
    );
  romo2datao3_s_13_F6MUX_4623 : X_MUX2
    port map (
      IA => nx53675z950,
      IB => nx53675z952,
      SEL => romo2datao3_s_13_BYINV,
      O => romo2datao3_s_13_F6MUX
    );
  romo2datao3_s_13_BYINV_4624 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_13_BYINV
    );
  nx53675z950_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z950_F5MUX,
      O => nx53675z950
    );
  nx53675z950_F5MUX_4625 : X_MUX2
    port map (
      IA => nx53675z950_G,
      IB => nx53675z951,
      SEL => nx53675z950_BXINV,
      O => nx53675z950_F5MUX
    );
  nx53675z950_BXINV_4626 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z950_BXINV
    );
  romo2datao2_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_1_F5MUX,
      O => nx53675z945
    );
  romo2datao2_s_1_F5MUX_4627 : X_MUX2
    port map (
      IA => nx53675z946,
      IB => nx53675z947,
      SEL => romo2datao2_s_1_BXINV,
      O => romo2datao2_s_1_F5MUX
    );
  romo2datao2_s_1_BXINV_4628 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_1_BXINV
    );
  romo2datao2_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_1_F6MUX,
      O => romo2datao2_s(1)
    );
  romo2datao2_s_1_F6MUX_4629 : X_MUX2
    port map (
      IA => nx53675z942,
      IB => nx53675z945,
      SEL => romo2datao2_s_1_BYINV,
      O => romo2datao2_s_1_F6MUX
    );
  romo2datao2_s_1_BYINV_4630 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_1_BYINV
    );
  nx53675z942_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z942_F5MUX,
      O => nx53675z942
    );
  nx53675z942_F5MUX_4631 : X_MUX2
    port map (
      IA => nx53675z943,
      IB => nx53675z944,
      SEL => nx53675z942_BXINV,
      O => nx53675z942_F5MUX
    );
  nx53675z942_BXINV_4632 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z942_BXINV
    );
  romo2datao2_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_0_F5MUX,
      O => U2_ROMO2_modgen_rom_ix0_nx_ro64_32_l
    );
  romo2datao2_s_0_F5MUX_4633 : X_MUX2
    port map (
      IA => nx53675z948,
      IB => nx53675z949,
      SEL => romo2datao2_s_0_BXINV,
      O => romo2datao2_s_0_F5MUX
    );
  romo2datao2_s_0_BXINV_4634 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_0_BXINV
    );
  romo2datao2_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_0_F6MUX,
      O => romo2datao2_s(0)
    );
  romo2datao2_s_0_F6MUX_4635 : X_MUX2
    port map (
      IA => U2_ROMO2_modgen_rom_ix0_nx_ro64_32_u,
      IB => U2_ROMO2_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romo2datao2_s_0_BYINV,
      O => romo2datao2_s_0_F6MUX
    );
  romo2datao2_s_0_BYINV_4636 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_0_BYINV
    );
  U_DCT2D_reg_databuf_reg_2_9_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_2_8_DYMUX,
      CE => U_DCT2D_databuf_reg_2_8_CEINV,
      CLK => U_DCT2D_databuf_reg_2_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_2_8_FFY_RST,
      O => U_DCT2D_databuf_reg_2_Q(9)
    );
  U_DCT2D_databuf_reg_2_8_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_2_8_FFY_RST
    );
  U2_ROMO2_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROMO2_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U2_ROMO2_modgen_rom_ix0_nx_ro64_32_u
    );
  U2_ROMO2_modgen_rom_ix0_nx_ro64_32_u_F5MUX_4637 : X_MUX2
    port map (
      IA => U2_ROMO2_modgen_rom_ix0_nx_rm64_16_u,
      IB => U2_ROMO2_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U2_ROMO2_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U2_ROMO2_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U2_ROMO2_modgen_rom_ix0_nx_ro64_32_u_BXINV_4638 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => U2_ROMO2_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romo2datao1_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_7_F5MUX,
      O => nx53675z830
    );
  romo2datao1_s_7_F5MUX_4639 : X_MUX2
    port map (
      IA => nx53675z831,
      IB => nx53675z832,
      SEL => romo2datao1_s_7_BXINV,
      O => romo2datao1_s_7_F5MUX
    );
  romo2datao1_s_7_BXINV_4640 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_7_BXINV
    );
  romo2datao1_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_7_F6MUX,
      O => romo2datao1_s(7)
    );
  romo2datao1_s_7_F6MUX_4641 : X_MUX2
    port map (
      IA => nx53675z827,
      IB => nx53675z830,
      SEL => romo2datao1_s_7_BYINV,
      O => romo2datao1_s_7_F6MUX
    );
  romo2datao1_s_7_BYINV_4642 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_7_BYINV
    );
  nx53675z827_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z827_F5MUX,
      O => nx53675z827
    );
  nx53675z827_F5MUX_4643 : X_MUX2
    port map (
      IA => nx53675z828,
      IB => nx53675z829,
      SEL => nx53675z827_BXINV,
      O => nx53675z827_F5MUX
    );
  nx53675z827_BXINV_4644 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z827_BXINV
    );
  romo2datao1_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_6_F5MUX,
      O => nx53675z836
    );
  romo2datao1_s_6_F5MUX_4645 : X_MUX2
    port map (
      IA => nx53675z837,
      IB => nx53675z838,
      SEL => romo2datao1_s_6_BXINV,
      O => romo2datao1_s_6_F5MUX
    );
  romo2datao1_s_6_BXINV_4646 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_6_BXINV
    );
  romo2datao1_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_6_F6MUX,
      O => romo2datao1_s(6)
    );
  romo2datao1_s_6_F6MUX_4647 : X_MUX2
    port map (
      IA => nx53675z833,
      IB => nx53675z836,
      SEL => romo2datao1_s_6_BYINV,
      O => romo2datao1_s_6_F6MUX
    );
  romo2datao1_s_6_BYINV_4648 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_6_BYINV
    );
  nx53675z833_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z833_F5MUX,
      O => nx53675z833
    );
  nx53675z833_F5MUX_4649 : X_MUX2
    port map (
      IA => nx53675z834,
      IB => nx53675z835,
      SEL => nx53675z833_BXINV,
      O => nx53675z833_F5MUX
    );
  nx53675z833_BXINV_4650 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z833_BXINV
    );
  romo2datao1_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_5_F5MUX,
      O => nx53675z842
    );
  romo2datao1_s_5_F5MUX_4651 : X_MUX2
    port map (
      IA => nx53675z843,
      IB => nx53675z844,
      SEL => romo2datao1_s_5_BXINV,
      O => romo2datao1_s_5_F5MUX
    );
  romo2datao1_s_5_BXINV_4652 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_5_BXINV
    );
  romo2datao1_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_5_F6MUX,
      O => romo2datao1_s(5)
    );
  romo2datao1_s_5_F6MUX_4653 : X_MUX2
    port map (
      IA => nx53675z839,
      IB => nx53675z842,
      SEL => romo2datao1_s_5_BYINV,
      O => romo2datao1_s_5_F6MUX
    );
  romo2datao1_s_5_BYINV_4654 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_5_BYINV
    );
  nx53675z839_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z839_F5MUX,
      O => nx53675z839
    );
  nx53675z839_F5MUX_4655 : X_MUX2
    port map (
      IA => nx53675z840,
      IB => nx53675z841,
      SEL => nx53675z839_BXINV,
      O => nx53675z839_F5MUX
    );
  nx53675z839_BXINV_4656 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z839_BXINV
    );
  romo2datao1_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_4_F5MUX,
      O => nx53675z848
    );
  romo2datao1_s_4_F5MUX_4657 : X_MUX2
    port map (
      IA => nx53675z849,
      IB => nx53675z850,
      SEL => romo2datao1_s_4_BXINV,
      O => romo2datao1_s_4_F5MUX
    );
  romo2datao1_s_4_BXINV_4658 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_4_BXINV
    );
  romo2datao1_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_4_F6MUX,
      O => romo2datao1_s(4)
    );
  romo2datao1_s_4_F6MUX_4659 : X_MUX2
    port map (
      IA => nx53675z845,
      IB => nx53675z848,
      SEL => romo2datao1_s_4_BYINV,
      O => romo2datao1_s_4_F6MUX
    );
  romo2datao1_s_4_BYINV_4660 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_4_BYINV
    );
  nx53675z845_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z845_F5MUX,
      O => nx53675z845
    );
  nx53675z845_F5MUX_4661 : X_MUX2
    port map (
      IA => nx53675z846,
      IB => nx53675z847,
      SEL => nx53675z845_BXINV,
      O => nx53675z845_F5MUX
    );
  nx53675z845_BXINV_4662 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z845_BXINV
    );
  romo2datao1_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_3_F5MUX,
      O => nx53675z854
    );
  romo2datao1_s_3_F5MUX_4663 : X_MUX2
    port map (
      IA => nx53675z855,
      IB => nx53675z856,
      SEL => romo2datao1_s_3_BXINV,
      O => romo2datao1_s_3_F5MUX
    );
  romo2datao1_s_3_BXINV_4664 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_3_BXINV
    );
  romo2datao1_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_3_F6MUX,
      O => romo2datao1_s(3)
    );
  romo2datao1_s_3_F6MUX_4665 : X_MUX2
    port map (
      IA => nx53675z851,
      IB => nx53675z854,
      SEL => romo2datao1_s_3_BYINV,
      O => romo2datao1_s_3_F6MUX
    );
  romo2datao1_s_3_BYINV_4666 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_3_BYINV
    );
  U_DCT2D_ix2262z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_5_8_Q,
      ADR1 => U_DCT2D_latchbuf_reg_2_8_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx2262z1
    );
  nx53675z851_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z851_F5MUX,
      O => nx53675z851
    );
  nx53675z851_F5MUX_4667 : X_MUX2
    port map (
      IA => nx53675z852,
      IB => nx53675z853,
      SEL => nx53675z851_BXINV,
      O => nx53675z851_F5MUX
    );
  nx53675z851_BXINV_4668 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z851_BXINV
    );
  rome2datao6_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_12_F5MUX,
      O => nx53675z398
    );
  rome2datao6_s_12_F5MUX_4669 : X_MUX2
    port map (
      IA => nx53675z399,
      IB => nx53675z400,
      SEL => rome2datao6_s_12_BXINV,
      O => rome2datao6_s_12_F5MUX
    );
  rome2datao6_s_12_BXINV_4670 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao6_s_12_BXINV
    );
  rome2datao6_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_12_F6MUX,
      O => rome2datao6_s(12)
    );
  rome2datao6_s_12_F6MUX_4671 : X_MUX2
    port map (
      IA => nx53675z395,
      IB => nx53675z398,
      SEL => rome2datao6_s_12_BYINV,
      O => rome2datao6_s_12_F6MUX
    );
  rome2datao6_s_12_BYINV_4672 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao6_s_12_BYINV
    );
  nx53675z395_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z395_F5MUX,
      O => nx53675z395
    );
  nx53675z395_F5MUX_4673 : X_MUX2
    port map (
      IA => nx53675z396,
      IB => nx53675z397,
      SEL => nx53675z395_BXINV,
      O => nx53675z395_F5MUX
    );
  nx53675z395_BXINV_4674 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z395_BXINV
    );
  rome2datao6_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_4_F5MUX,
      O => nx53675z446
    );
  rome2datao6_s_4_F5MUX_4675 : X_MUX2
    port map (
      IA => nx53675z447,
      IB => nx53675z448,
      SEL => rome2datao6_s_4_BXINV,
      O => rome2datao6_s_4_F5MUX
    );
  rome2datao6_s_4_BXINV_4676 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao6_s_4_BXINV
    );
  rome2datao6_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_4_F6MUX,
      O => rome2datao6_s(4)
    );
  rome2datao6_s_4_F6MUX_4677 : X_MUX2
    port map (
      IA => nx53675z443,
      IB => nx53675z446,
      SEL => rome2datao6_s_4_BYINV,
      O => rome2datao6_s_4_F6MUX
    );
  rome2datao6_s_4_BYINV_4678 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao6_s_4_BYINV
    );
  nx53675z443_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z443_F5MUX,
      O => nx53675z443
    );
  nx53675z443_F5MUX_4679 : X_MUX2
    port map (
      IA => nx53675z444,
      IB => nx53675z445,
      SEL => nx53675z443_BXINV,
      O => nx53675z443_F5MUX
    );
  nx53675z443_BXINV_4680 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z443_BXINV
    );
  rome2datao6_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_3_F5MUX,
      O => nx53675z451
    );
  rome2datao6_s_3_F5MUX_4681 : X_MUX2
    port map (
      IA => nx53675z452,
      IB => nx53675z453,
      SEL => rome2datao6_s_3_BXINV,
      O => rome2datao6_s_3_F5MUX
    );
  rome2datao6_s_3_BXINV_4682 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao6_s_3_BXINV
    );
  rome2datao6_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_3_F6MUX,
      O => rome2datao6_s(3)
    );
  rome2datao6_s_3_F6MUX_4683 : X_MUX2
    port map (
      IA => nx53675z449,
      IB => nx53675z451,
      SEL => rome2datao6_s_3_BYINV,
      O => rome2datao6_s_3_F6MUX
    );
  rome2datao6_s_3_BYINV_4684 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao6_s_3_BYINV
    );
  nx53675z449_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z449_F5MUX,
      O => nx53675z449
    );
  nx53675z449_F5MUX_4685 : X_MUX2
    port map (
      IA => U2_ROME6_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx53675z450,
      SEL => nx53675z449_BXINV,
      O => nx53675z449_F5MUX
    );
  nx53675z449_BXINV_4686 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z449_BXINV
    );
  rome2datao6_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_2_F5MUX,
      O => U2_ROME6_modgen_rom_ix2_nx_ro64_32_l
    );
  rome2datao6_s_2_F5MUX_4687 : X_MUX2
    port map (
      IA => rome2datao6_s_2_G,
      IB => nx53675z454,
      SEL => rome2datao6_s_2_BXINV,
      O => rome2datao6_s_2_F5MUX
    );
  rome2datao6_s_2_BXINV_4688 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao6_s_2_BXINV
    );
  rome2datao6_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_2_F6MUX,
      O => rome2datao6_s(2)
    );
  rome2datao6_s_2_F6MUX_4689 : X_MUX2
    port map (
      IA => U2_ROME6_modgen_rom_ix2_nx_ro64_32_u,
      IB => U2_ROME6_modgen_rom_ix2_nx_ro64_32_l,
      SEL => rome2datao6_s_2_BYINV,
      O => rome2datao6_s_2_F6MUX
    );
  rome2datao6_s_2_BYINV_4690 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao6_s_2_BYINV
    );
  U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U2_ROME6_modgen_rom_ix2_nx_ro64_32_u
    );
  U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_F5MUX_4691 : X_MUX2
    port map (
      IA => U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U2_ROME6_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_BXINV_4692 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  romo2datao0_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_4_F5MUX,
      O => nx53675z771
    );
  romo2datao0_s_4_F5MUX_4693 : X_MUX2
    port map (
      IA => nx53675z772,
      IB => nx53675z773,
      SEL => romo2datao0_s_4_BXINV,
      O => romo2datao0_s_4_F5MUX
    );
  romo2datao0_s_4_BXINV_4694 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_4_BXINV
    );
  romo2datao0_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_4_F6MUX,
      O => romo2datao0_s(4)
    );
  romo2datao0_s_4_F6MUX_4695 : X_MUX2
    port map (
      IA => nx53675z768,
      IB => nx53675z771,
      SEL => romo2datao0_s_4_BYINV,
      O => romo2datao0_s_4_F6MUX
    );
  romo2datao0_s_4_BYINV_4696 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_4_BYINV
    );
  nx53675z768_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z768_F5MUX,
      O => nx53675z768
    );
  nx53675z768_F5MUX_4697 : X_MUX2
    port map (
      IA => nx53675z769,
      IB => nx53675z770,
      SEL => nx53675z768_BXINV,
      O => nx53675z768_F5MUX
    );
  nx53675z768_BXINV_4698 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z768_BXINV
    );
  romo2datao0_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_3_F5MUX,
      O => nx53675z777
    );
  romo2datao0_s_3_F5MUX_4699 : X_MUX2
    port map (
      IA => nx53675z778,
      IB => nx53675z779,
      SEL => romo2datao0_s_3_BXINV,
      O => romo2datao0_s_3_F5MUX
    );
  romo2datao0_s_3_BXINV_4700 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_3_BXINV
    );
  romo2datao0_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_3_F6MUX,
      O => romo2datao0_s(3)
    );
  romo2datao0_s_3_F6MUX_4701 : X_MUX2
    port map (
      IA => nx53675z774,
      IB => nx53675z777,
      SEL => romo2datao0_s_3_BYINV,
      O => romo2datao0_s_3_F6MUX
    );
  romo2datao0_s_3_BYINV_4702 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_3_BYINV
    );
  nx53675z774_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z774_F5MUX,
      O => nx53675z774
    );
  nx53675z774_F5MUX_4703 : X_MUX2
    port map (
      IA => nx53675z775,
      IB => nx53675z776,
      SEL => nx53675z774_BXINV,
      O => nx53675z774_F5MUX
    );
  nx53675z774_BXINV_4704 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z774_BXINV
    );
  romo2datao0_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_2_F5MUX,
      O => nx53675z783
    );
  romo2datao0_s_2_F5MUX_4705 : X_MUX2
    port map (
      IA => nx53675z784,
      IB => nx53675z785,
      SEL => romo2datao0_s_2_BXINV,
      O => romo2datao0_s_2_F5MUX
    );
  romo2datao0_s_2_BXINV_4706 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_2_BXINV
    );
  romo2datao0_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_2_F6MUX,
      O => romo2datao0_s(2)
    );
  romo2datao0_s_2_F6MUX_4707 : X_MUX2
    port map (
      IA => nx53675z780,
      IB => nx53675z783,
      SEL => romo2datao0_s_2_BYINV,
      O => romo2datao0_s_2_F6MUX
    );
  romo2datao0_s_2_BYINV_4708 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_2_BYINV
    );
  nx53675z780_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z780_F5MUX,
      O => nx53675z780
    );
  nx53675z780_F5MUX_4709 : X_MUX2
    port map (
      IA => nx53675z781,
      IB => nx53675z782,
      SEL => nx53675z780_BXINV,
      O => nx53675z780_F5MUX
    );
  nx53675z780_BXINV_4710 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z780_BXINV
    );
  romo2datao0_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_1_F5MUX,
      O => nx53675z789
    );
  romo2datao0_s_1_F5MUX_4711 : X_MUX2
    port map (
      IA => nx53675z790,
      IB => nx53675z791,
      SEL => romo2datao0_s_1_BXINV,
      O => romo2datao0_s_1_F5MUX
    );
  romo2datao0_s_1_BXINV_4712 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_1_BXINV
    );
  romo2datao0_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_1_F6MUX,
      O => romo2datao0_s(1)
    );
  romo2datao0_s_1_F6MUX_4713 : X_MUX2
    port map (
      IA => nx53675z786,
      IB => nx53675z789,
      SEL => romo2datao0_s_1_BYINV,
      O => romo2datao0_s_1_F6MUX
    );
  romo2datao0_s_1_BYINV_4714 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_1_BYINV
    );
  nx53675z786_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z786_F5MUX,
      O => nx53675z786
    );
  nx53675z786_F5MUX_4715 : X_MUX2
    port map (
      IA => nx53675z787,
      IB => nx53675z788,
      SEL => nx53675z786_BXINV,
      O => nx53675z786_F5MUX
    );
  nx53675z786_BXINV_4716 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z786_BXINV
    );
  rome2datao3_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_10_F5MUX,
      O => nx53675z215
    );
  rome2datao3_s_10_F5MUX_4717 : X_MUX2
    port map (
      IA => nx53675z216,
      IB => nx53675z217,
      SEL => rome2datao3_s_10_BXINV,
      O => rome2datao3_s_10_F5MUX
    );
  rome2datao3_s_10_BXINV_4718 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao3_s_10_BXINV
    );
  rome2datao3_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_10_F6MUX,
      O => rome2datao3_s(10)
    );
  rome2datao3_s_10_F6MUX_4719 : X_MUX2
    port map (
      IA => nx53675z212,
      IB => nx53675z215,
      SEL => rome2datao3_s_10_BYINV,
      O => rome2datao3_s_10_F6MUX
    );
  rome2datao3_s_10_BYINV_4720 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao3_s_10_BYINV
    );
  nx53675z212_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z212_F5MUX,
      O => nx53675z212
    );
  nx53675z212_F5MUX_4721 : X_MUX2
    port map (
      IA => nx53675z213,
      IB => nx53675z214,
      SEL => nx53675z212_BXINV,
      O => nx53675z212_F5MUX
    );
  nx53675z212_BXINV_4722 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z212_BXINV
    );
  rome2datao3_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_8_F5MUX,
      O => nx53675z227
    );
  rome2datao3_s_8_F5MUX_4723 : X_MUX2
    port map (
      IA => nx53675z228,
      IB => nx53675z229,
      SEL => rome2datao3_s_8_BXINV,
      O => rome2datao3_s_8_F5MUX
    );
  rome2datao3_s_8_BXINV_4724 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao3_s_8_BXINV
    );
  rome2datao3_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_8_F6MUX,
      O => rome2datao3_s(8)
    );
  rome2datao3_s_8_F6MUX_4725 : X_MUX2
    port map (
      IA => nx53675z224,
      IB => nx53675z227,
      SEL => rome2datao3_s_8_BYINV,
      O => rome2datao3_s_8_F6MUX
    );
  rome2datao3_s_8_BYINV_4726 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao3_s_8_BYINV
    );
  U_DCT2D_reg_databuf_reg_2_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_2_8_DXMUX,
      CE => U_DCT2D_databuf_reg_2_8_CEINV,
      CLK => U_DCT2D_databuf_reg_2_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_2_8_FFX_RST,
      O => U_DCT2D_databuf_reg_2_Q(8)
    );
  U_DCT2D_databuf_reg_2_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_2_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_2_8_FFX_RST
    );
  nx53675z224_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z224_F5MUX,
      O => nx53675z224
    );
  nx53675z224_F5MUX_4727 : X_MUX2
    port map (
      IA => nx53675z225,
      IB => nx53675z226,
      SEL => nx53675z224_BXINV,
      O => nx53675z224_F5MUX
    );
  nx53675z224_BXINV_4728 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z224_BXINV
    );
  romo2datao4_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_11_F5MUX,
      O => nx53675z1043
    );
  romo2datao4_s_11_F5MUX_4729 : X_MUX2
    port map (
      IA => nx53675z1044,
      IB => nx53675z1045,
      SEL => romo2datao4_s_11_BXINV,
      O => romo2datao4_s_11_F5MUX
    );
  romo2datao4_s_11_BXINV_4730 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_11_BXINV
    );
  romo2datao4_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_11_F6MUX,
      O => romo2datao4_s(11)
    );
  romo2datao4_s_11_F6MUX_4731 : X_MUX2
    port map (
      IA => nx53675z1040,
      IB => nx53675z1043,
      SEL => romo2datao4_s_11_BYINV,
      O => romo2datao4_s_11_F6MUX
    );
  romo2datao4_s_11_BYINV_4732 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_11_BYINV
    );
  nx53675z1040_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1040_F5MUX,
      O => nx53675z1040
    );
  nx53675z1040_F5MUX_4733 : X_MUX2
    port map (
      IA => nx53675z1041,
      IB => nx53675z1042,
      SEL => nx53675z1040_BXINV,
      O => nx53675z1040_F5MUX
    );
  nx53675z1040_BXINV_4734 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1040_BXINV
    );
  romo2datao3_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_1_F5MUX,
      O => nx53675z1024
    );
  romo2datao3_s_1_F5MUX_4735 : X_MUX2
    port map (
      IA => nx53675z1025,
      IB => nx53675z1026,
      SEL => romo2datao3_s_1_BXINV,
      O => romo2datao3_s_1_F5MUX
    );
  romo2datao3_s_1_BXINV_4736 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_1_BXINV
    );
  romo2datao3_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_1_F6MUX,
      O => romo2datao3_s(1)
    );
  romo2datao3_s_1_F6MUX_4737 : X_MUX2
    port map (
      IA => nx53675z1021,
      IB => nx53675z1024,
      SEL => romo2datao3_s_1_BYINV,
      O => romo2datao3_s_1_F6MUX
    );
  romo2datao3_s_1_BYINV_4738 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_1_BYINV
    );
  nx53675z1021_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1021_F5MUX,
      O => nx53675z1021
    );
  nx53675z1021_F5MUX_4739 : X_MUX2
    port map (
      IA => nx53675z1022,
      IB => nx53675z1023,
      SEL => nx53675z1021_BXINV,
      O => nx53675z1021_F5MUX
    );
  nx53675z1021_BXINV_4740 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1021_BXINV
    );
  romo2datao0_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_13_F5MUX,
      O => nx53675z717
    );
  romo2datao0_s_13_F5MUX_4741 : X_MUX2
    port map (
      IA => nx53675z718,
      IB => nx53675z719,
      SEL => romo2datao0_s_13_BXINV,
      O => romo2datao0_s_13_F5MUX
    );
  romo2datao0_s_13_BXINV_4742 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao0_s_13_BXINV
    );
  romo2datao0_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao0_s_13_F6MUX,
      O => romo2datao0_s(13)
    );
  romo2datao0_s_13_F6MUX_4743 : X_MUX2
    port map (
      IA => nx53675z715,
      IB => nx53675z717,
      SEL => romo2datao0_s_13_BYINV,
      O => romo2datao0_s_13_F6MUX
    );
  romo2datao0_s_13_BYINV_4744 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao0_s_13_BYINV
    );
  nx53675z715_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z715_F5MUX,
      O => nx53675z715
    );
  nx53675z715_F5MUX_4745 : X_MUX2
    port map (
      IA => nx53675z715_G,
      IB => nx53675z716,
      SEL => nx53675z715_BXINV,
      O => nx53675z715_F5MUX
    );
  nx53675z715_BXINV_4746 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z715_BXINV
    );
  romo2datao8_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_12_F5MUX,
      O => nx53675z1353
    );
  romo2datao8_s_12_F5MUX_4747 : X_MUX2
    port map (
      IA => nx53675z1354,
      IB => nx53675z1355,
      SEL => romo2datao8_s_12_BXINV,
      O => romo2datao8_s_12_F5MUX
    );
  romo2datao8_s_12_BXINV_4748 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_12_BXINV
    );
  romo2datao8_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_12_F6MUX,
      O => romo2datao8_s(12)
    );
  romo2datao8_s_12_F6MUX_4749 : X_MUX2
    port map (
      IA => nx53675z1350,
      IB => nx53675z1353,
      SEL => romo2datao8_s_12_BYINV,
      O => romo2datao8_s_12_F6MUX
    );
  romo2datao8_s_12_BYINV_4750 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_12_BYINV
    );
  nx53675z1350_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1350_F5MUX,
      O => nx53675z1350
    );
  nx53675z1350_F5MUX_4751 : X_MUX2
    port map (
      IA => nx53675z1351,
      IB => nx53675z1352,
      SEL => nx53675z1350_BXINV,
      O => nx53675z1350_F5MUX
    );
  nx53675z1350_BXINV_4752 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1350_BXINV
    );
  romo2datao8_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_4_F5MUX,
      O => nx53675z1401
    );
  romo2datao8_s_4_F5MUX_4753 : X_MUX2
    port map (
      IA => nx53675z1402,
      IB => nx53675z1403,
      SEL => romo2datao8_s_4_BXINV,
      O => romo2datao8_s_4_F5MUX
    );
  romo2datao8_s_4_BXINV_4754 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_4_BXINV
    );
  romo2datao8_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_4_F6MUX,
      O => romo2datao8_s(4)
    );
  romo2datao8_s_4_F6MUX_4755 : X_MUX2
    port map (
      IA => nx53675z1398,
      IB => nx53675z1401,
      SEL => romo2datao8_s_4_BYINV,
      O => romo2datao8_s_4_F6MUX
    );
  romo2datao8_s_4_BYINV_4756 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_4_BYINV
    );
  nx53675z1398_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1398_F5MUX,
      O => nx53675z1398
    );
  nx53675z1398_F5MUX_4757 : X_MUX2
    port map (
      IA => nx53675z1399,
      IB => nx53675z1400,
      SEL => nx53675z1398_BXINV,
      O => nx53675z1398_F5MUX
    );
  nx53675z1398_BXINV_4758 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1398_BXINV
    );
  romo2datao8_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_3_F5MUX,
      O => nx53675z1407
    );
  romo2datao8_s_3_F5MUX_4759 : X_MUX2
    port map (
      IA => nx53675z1408,
      IB => nx53675z1409,
      SEL => romo2datao8_s_3_BXINV,
      O => romo2datao8_s_3_F5MUX
    );
  romo2datao8_s_3_BXINV_4760 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_3_BXINV
    );
  romo2datao8_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_3_F6MUX,
      O => romo2datao8_s(3)
    );
  romo2datao8_s_3_F6MUX_4761 : X_MUX2
    port map (
      IA => nx53675z1404,
      IB => nx53675z1407,
      SEL => romo2datao8_s_3_BYINV,
      O => romo2datao8_s_3_F6MUX
    );
  romo2datao8_s_3_BYINV_4762 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_3_BYINV
    );
  nx53675z1404_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1404_F5MUX,
      O => nx53675z1404
    );
  nx53675z1404_F5MUX_4763 : X_MUX2
    port map (
      IA => nx53675z1405,
      IB => nx53675z1406,
      SEL => nx53675z1404_BXINV,
      O => nx53675z1404_F5MUX
    );
  nx53675z1404_BXINV_4764 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1404_BXINV
    );
  romo2datao8_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_2_F5MUX,
      O => nx53675z1413
    );
  romo2datao8_s_2_F5MUX_4765 : X_MUX2
    port map (
      IA => nx53675z1414,
      IB => nx53675z1415,
      SEL => romo2datao8_s_2_BXINV,
      O => romo2datao8_s_2_F5MUX
    );
  romo2datao8_s_2_BXINV_4766 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao8_s_2_BXINV
    );
  romo2datao8_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao8_s_2_F6MUX,
      O => romo2datao8_s(2)
    );
  romo2datao8_s_2_F6MUX_4767 : X_MUX2
    port map (
      IA => nx53675z1410,
      IB => nx53675z1413,
      SEL => romo2datao8_s_2_BYINV,
      O => romo2datao8_s_2_F6MUX
    );
  romo2datao8_s_2_BYINV_4768 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao8_s_2_BYINV
    );
  rome2datao3_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_7_F5MUX,
      O => nx53675z233
    );
  rome2datao3_s_7_F5MUX_4769 : X_MUX2
    port map (
      IA => nx53675z234,
      IB => nx53675z235,
      SEL => rome2datao3_s_7_BXINV,
      O => rome2datao3_s_7_F5MUX
    );
  rome2datao3_s_7_BXINV_4770 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao3_s_7_BXINV
    );
  rome2datao3_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_7_F6MUX,
      O => rome2datao3_s(7)
    );
  rome2datao3_s_7_F6MUX_4771 : X_MUX2
    port map (
      IA => nx53675z230,
      IB => nx53675z233,
      SEL => rome2datao3_s_7_BYINV,
      O => rome2datao3_s_7_F6MUX
    );
  rome2datao3_s_7_BYINV_4772 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao3_s_7_BYINV
    );
  nx53675z230_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z230_F5MUX,
      O => nx53675z230
    );
  nx53675z230_F5MUX_4773 : X_MUX2
    port map (
      IA => nx53675z231,
      IB => nx53675z232,
      SEL => nx53675z230_BXINV,
      O => nx53675z230_F5MUX
    );
  nx53675z230_BXINV_4774 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z230_BXINV
    );
  romo2datao9_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_2_F5MUX,
      O => nx53675z1492
    );
  romo2datao9_s_2_F5MUX_4775 : X_MUX2
    port map (
      IA => nx53675z1493,
      IB => nx53675z1494,
      SEL => romo2datao9_s_2_BXINV,
      O => romo2datao9_s_2_F5MUX
    );
  romo2datao9_s_2_BXINV_4776 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_2_BXINV
    );
  romo2datao9_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_2_F6MUX,
      O => romo2datao9_s(2)
    );
  romo2datao9_s_2_F6MUX_4777 : X_MUX2
    port map (
      IA => nx53675z1489,
      IB => nx53675z1492,
      SEL => romo2datao9_s_2_BYINV,
      O => romo2datao9_s_2_F6MUX
    );
  romo2datao9_s_2_BYINV_4778 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_2_BYINV
    );
  nx53675z1489_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1489_F5MUX,
      O => nx53675z1489
    );
  nx53675z1489_F5MUX_4779 : X_MUX2
    port map (
      IA => nx53675z1490,
      IB => nx53675z1491,
      SEL => nx53675z1489_BXINV,
      O => nx53675z1489_F5MUX
    );
  nx53675z1489_BXINV_4780 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1489_BXINV
    );
  romo2datao4_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_12_F5MUX,
      O => nx53675z1037
    );
  romo2datao4_s_12_F5MUX_4781 : X_MUX2
    port map (
      IA => nx53675z1038,
      IB => nx53675z1039,
      SEL => romo2datao4_s_12_BXINV,
      O => romo2datao4_s_12_F5MUX
    );
  romo2datao4_s_12_BXINV_4782 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_12_BXINV
    );
  romo2datao4_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_12_F6MUX,
      O => romo2datao4_s(12)
    );
  romo2datao4_s_12_F6MUX_4783 : X_MUX2
    port map (
      IA => nx53675z1034,
      IB => nx53675z1037,
      SEL => romo2datao4_s_12_BYINV,
      O => romo2datao4_s_12_F6MUX
    );
  romo2datao4_s_12_BYINV_4784 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_12_BYINV
    );
  nx53675z1034_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1034_F5MUX,
      O => nx53675z1034
    );
  nx53675z1034_F5MUX_4785 : X_MUX2
    port map (
      IA => nx53675z1035,
      IB => nx53675z1036,
      SEL => nx53675z1034_BXINV,
      O => nx53675z1034_F5MUX
    );
  nx53675z1034_BXINV_4786 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1034_BXINV
    );
  romo2datao3_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_10_F5MUX,
      O => nx53675z970
    );
  romo2datao3_s_10_F5MUX_4787 : X_MUX2
    port map (
      IA => nx53675z971,
      IB => nx53675z972,
      SEL => romo2datao3_s_10_BXINV,
      O => romo2datao3_s_10_F5MUX
    );
  romo2datao3_s_10_BXINV_4788 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_10_BXINV
    );
  romo2datao3_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_10_F6MUX,
      O => romo2datao3_s(10)
    );
  romo2datao3_s_10_F6MUX_4789 : X_MUX2
    port map (
      IA => nx53675z967,
      IB => nx53675z970,
      SEL => romo2datao3_s_10_BYINV,
      O => romo2datao3_s_10_F6MUX
    );
  romo2datao3_s_10_BYINV_4790 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_10_BYINV
    );
  nx53675z967_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z967_F5MUX,
      O => nx53675z967
    );
  nx53675z967_F5MUX_4791 : X_MUX2
    port map (
      IA => nx53675z968,
      IB => nx53675z969,
      SEL => nx53675z967_BXINV,
      O => nx53675z967_F5MUX
    );
  nx53675z967_BXINV_4792 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z967_BXINV
    );
  romo2datao3_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_8_F5MUX,
      O => nx53675z982
    );
  romo2datao3_s_8_F5MUX_4793 : X_MUX2
    port map (
      IA => nx53675z983,
      IB => nx53675z984,
      SEL => romo2datao3_s_8_BXINV,
      O => romo2datao3_s_8_F5MUX
    );
  romo2datao3_s_8_BXINV_4794 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_8_BXINV
    );
  romo2datao3_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_8_F6MUX,
      O => romo2datao3_s(8)
    );
  romo2datao3_s_8_F6MUX_4795 : X_MUX2
    port map (
      IA => nx53675z979,
      IB => nx53675z982,
      SEL => romo2datao3_s_8_BYINV,
      O => romo2datao3_s_8_F6MUX
    );
  romo2datao3_s_8_BYINV_4796 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_8_BYINV
    );
  nx53675z979_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z979_F5MUX,
      O => nx53675z979
    );
  nx53675z979_F5MUX_4797 : X_MUX2
    port map (
      IA => nx53675z980,
      IB => nx53675z981,
      SEL => nx53675z979_BXINV,
      O => nx53675z979_F5MUX
    );
  nx53675z979_BXINV_4798 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z979_BXINV
    );
  romo2datao3_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_0_F5MUX,
      O => U2_ROMO3_modgen_rom_ix0_nx_ro64_32_l
    );
  romo2datao3_s_0_F5MUX_4799 : X_MUX2
    port map (
      IA => nx53675z1027,
      IB => nx53675z1028,
      SEL => romo2datao3_s_0_BXINV,
      O => romo2datao3_s_0_F5MUX
    );
  romo2datao3_s_0_BXINV_4800 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_0_BXINV
    );
  romo2datao3_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_0_F6MUX,
      O => romo2datao3_s(0)
    );
  romo2datao3_s_0_F6MUX_4801 : X_MUX2
    port map (
      IA => U2_ROMO3_modgen_rom_ix0_nx_ro64_32_u,
      IB => U2_ROMO3_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romo2datao3_s_0_BYINV,
      O => romo2datao3_s_0_F6MUX
    );
  romo2datao3_s_0_BYINV_4802 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_0_BYINV
    );
  U2_ROMO3_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROMO3_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U2_ROMO3_modgen_rom_ix0_nx_ro64_32_u
    );
  U2_ROMO3_modgen_rom_ix0_nx_ro64_32_u_F5MUX_4803 : X_MUX2
    port map (
      IA => U2_ROMO3_modgen_rom_ix0_nx_rm64_16_u,
      IB => U2_ROMO3_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U2_ROMO3_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U2_ROMO3_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U2_ROMO3_modgen_rom_ix0_nx_ro64_32_u_BXINV_4804 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => U2_ROMO3_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romo2datao2_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_7_F5MUX,
      O => nx53675z909
    );
  romo2datao2_s_7_F5MUX_4805 : X_MUX2
    port map (
      IA => nx53675z910,
      IB => nx53675z911,
      SEL => romo2datao2_s_7_BXINV,
      O => romo2datao2_s_7_F5MUX
    );
  romo2datao2_s_7_BXINV_4806 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_7_BXINV
    );
  romo2datao2_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_7_F6MUX,
      O => romo2datao2_s(7)
    );
  romo2datao2_s_7_F6MUX_4807 : X_MUX2
    port map (
      IA => nx53675z906,
      IB => nx53675z909,
      SEL => romo2datao2_s_7_BYINV,
      O => romo2datao2_s_7_F6MUX
    );
  romo2datao2_s_7_BYINV_4808 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_7_BYINV
    );
  nx53675z906_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z906_F5MUX,
      O => nx53675z906
    );
  nx53675z906_F5MUX_4809 : X_MUX2
    port map (
      IA => nx53675z907,
      IB => nx53675z908,
      SEL => nx53675z906_BXINV,
      O => nx53675z906_F5MUX
    );
  nx53675z906_BXINV_4810 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z906_BXINV
    );
  U_DCT2D_ix49552z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_0_0_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_7_0_Q,
      O => U_DCT2D_nx49552z1
    );
  romo2datao2_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_6_F5MUX,
      O => nx53675z915
    );
  romo2datao2_s_6_F5MUX_4811 : X_MUX2
    port map (
      IA => nx53675z916,
      IB => nx53675z917,
      SEL => romo2datao2_s_6_BXINV,
      O => romo2datao2_s_6_F5MUX
    );
  romo2datao2_s_6_BXINV_4812 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_6_BXINV
    );
  romo2datao2_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_6_F6MUX,
      O => romo2datao2_s(6)
    );
  romo2datao2_s_6_F6MUX_4813 : X_MUX2
    port map (
      IA => nx53675z912,
      IB => nx53675z915,
      SEL => romo2datao2_s_6_BYINV,
      O => romo2datao2_s_6_F6MUX
    );
  romo2datao2_s_6_BYINV_4814 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_6_BYINV
    );
  nx53675z912_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z912_F5MUX,
      O => nx53675z912
    );
  nx53675z912_F5MUX_4815 : X_MUX2
    port map (
      IA => nx53675z913,
      IB => nx53675z914,
      SEL => nx53675z912_BXINV,
      O => nx53675z912_F5MUX
    );
  nx53675z912_BXINV_4816 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z912_BXINV
    );
  romo2datao2_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_5_F5MUX,
      O => nx53675z921
    );
  romo2datao2_s_5_F5MUX_4817 : X_MUX2
    port map (
      IA => nx53675z922,
      IB => nx53675z923,
      SEL => romo2datao2_s_5_BXINV,
      O => romo2datao2_s_5_F5MUX
    );
  romo2datao2_s_5_BXINV_4818 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_5_BXINV
    );
  romo2datao2_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_5_F6MUX,
      O => romo2datao2_s(5)
    );
  romo2datao2_s_5_F6MUX_4819 : X_MUX2
    port map (
      IA => nx53675z918,
      IB => nx53675z921,
      SEL => romo2datao2_s_5_BYINV,
      O => romo2datao2_s_5_F6MUX
    );
  romo2datao2_s_5_BYINV_4820 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_5_BYINV
    );
  nx53675z918_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z918_F5MUX,
      O => nx53675z918
    );
  nx53675z918_F5MUX_4821 : X_MUX2
    port map (
      IA => nx53675z919,
      IB => nx53675z920,
      SEL => nx53675z918_BXINV,
      O => nx53675z918_F5MUX
    );
  nx53675z918_BXINV_4822 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z918_BXINV
    );
  romo2datao2_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_4_F5MUX,
      O => nx53675z927
    );
  romo2datao2_s_4_F5MUX_4823 : X_MUX2
    port map (
      IA => nx53675z928,
      IB => nx53675z929,
      SEL => romo2datao2_s_4_BXINV,
      O => romo2datao2_s_4_F5MUX
    );
  romo2datao2_s_4_BXINV_4824 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_4_BXINV
    );
  romo2datao2_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_4_F6MUX,
      O => romo2datao2_s(4)
    );
  romo2datao2_s_4_F6MUX_4825 : X_MUX2
    port map (
      IA => nx53675z924,
      IB => nx53675z927,
      SEL => romo2datao2_s_4_BYINV,
      O => romo2datao2_s_4_F6MUX
    );
  romo2datao2_s_4_BYINV_4826 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_4_BYINV
    );
  nx53675z924_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z924_F5MUX,
      O => nx53675z924
    );
  nx53675z924_F5MUX_4827 : X_MUX2
    port map (
      IA => nx53675z925,
      IB => nx53675z926,
      SEL => nx53675z924_BXINV,
      O => nx53675z924_F5MUX
    );
  nx53675z924_BXINV_4828 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z924_BXINV
    );
  romo2datao10_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_9_F5MUX,
      O => nx53675z1529
    );
  romo2datao10_s_9_F5MUX_4829 : X_MUX2
    port map (
      IA => nx53675z1530,
      IB => nx53675z1531,
      SEL => romo2datao10_s_9_BXINV,
      O => romo2datao10_s_9_F5MUX
    );
  romo2datao10_s_9_BXINV_4830 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_9_BXINV
    );
  romo2datao10_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_9_F6MUX,
      O => romo2datao10_s(9)
    );
  romo2datao10_s_9_F6MUX_4831 : X_MUX2
    port map (
      IA => nx53675z1526,
      IB => nx53675z1529,
      SEL => romo2datao10_s_9_BYINV,
      O => romo2datao10_s_9_F6MUX
    );
  romo2datao10_s_9_BYINV_4832 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_9_BYINV
    );
  nx53675z1526_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1526_F5MUX,
      O => nx53675z1526
    );
  nx53675z1526_F5MUX_4833 : X_MUX2
    port map (
      IA => nx53675z1527,
      IB => nx53675z1528,
      SEL => nx53675z1526_BXINV,
      O => nx53675z1526_F5MUX
    );
  nx53675z1526_BXINV_4834 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1526_BXINV
    );
  romo2datao10_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_8_F5MUX,
      O => nx53675z1535
    );
  romo2datao10_s_8_F5MUX_4835 : X_MUX2
    port map (
      IA => nx53675z1536,
      IB => nx53675z1537,
      SEL => romo2datao10_s_8_BXINV,
      O => romo2datao10_s_8_F5MUX
    );
  romo2datao10_s_8_BXINV_4836 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_8_BXINV
    );
  romo2datao10_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_8_F6MUX,
      O => romo2datao10_s(8)
    );
  romo2datao10_s_8_F6MUX_4837 : X_MUX2
    port map (
      IA => nx53675z1532,
      IB => nx53675z1535,
      SEL => romo2datao10_s_8_BYINV,
      O => romo2datao10_s_8_F6MUX
    );
  romo2datao10_s_8_BYINV_4838 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_8_BYINV
    );
  nx53675z1532_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1532_F5MUX,
      O => nx53675z1532
    );
  nx53675z1532_F5MUX_4839 : X_MUX2
    port map (
      IA => nx53675z1533,
      IB => nx53675z1534,
      SEL => nx53675z1532_BXINV,
      O => nx53675z1532_F5MUX
    );
  nx53675z1532_BXINV_4840 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1532_BXINV
    );
  romo2datao10_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_7_F5MUX,
      O => nx53675z1541
    );
  romo2datao10_s_7_F5MUX_4841 : X_MUX2
    port map (
      IA => nx53675z1542,
      IB => nx53675z1543,
      SEL => romo2datao10_s_7_BXINV,
      O => romo2datao10_s_7_F5MUX
    );
  romo2datao10_s_7_BXINV_4842 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_7_BXINV
    );
  romo2datao10_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_7_F6MUX,
      O => romo2datao10_s(7)
    );
  romo2datao10_s_7_F6MUX_4843 : X_MUX2
    port map (
      IA => nx53675z1538,
      IB => nx53675z1541,
      SEL => romo2datao10_s_7_BYINV,
      O => romo2datao10_s_7_F6MUX
    );
  romo2datao10_s_7_BYINV_4844 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_7_BYINV
    );
  nx53675z1538_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1538_F5MUX,
      O => nx53675z1538
    );
  nx53675z1538_F5MUX_4845 : X_MUX2
    port map (
      IA => nx53675z1539,
      IB => nx53675z1540,
      SEL => nx53675z1538_BXINV,
      O => nx53675z1538_F5MUX
    );
  nx53675z1538_BXINV_4846 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1538_BXINV
    );
  romo2datao10_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_6_F5MUX,
      O => nx53675z1547
    );
  romo2datao10_s_6_F5MUX_4847 : X_MUX2
    port map (
      IA => nx53675z1548,
      IB => nx53675z1549,
      SEL => romo2datao10_s_6_BXINV,
      O => romo2datao10_s_6_F5MUX
    );
  romo2datao10_s_6_BXINV_4848 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_6_BXINV
    );
  romo2datao10_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_6_F6MUX,
      O => romo2datao10_s(6)
    );
  romo2datao10_s_6_F6MUX_4849 : X_MUX2
    port map (
      IA => nx53675z1544,
      IB => nx53675z1547,
      SEL => romo2datao10_s_6_BYINV,
      O => romo2datao10_s_6_F6MUX
    );
  romo2datao10_s_6_BYINV_4850 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_6_BYINV
    );
  nx53675z1544_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1544_F5MUX,
      O => nx53675z1544
    );
  nx53675z1544_F5MUX_4851 : X_MUX2
    port map (
      IA => nx53675z1545,
      IB => nx53675z1546,
      SEL => nx53675z1544_BXINV,
      O => nx53675z1544_F5MUX
    );
  nx53675z1544_BXINV_4852 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1544_BXINV
    );
  romo2datao10_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_5_F5MUX,
      O => nx53675z1553
    );
  romo2datao10_s_5_F5MUX_4853 : X_MUX2
    port map (
      IA => nx53675z1554,
      IB => nx53675z1555,
      SEL => romo2datao10_s_5_BXINV,
      O => romo2datao10_s_5_F5MUX
    );
  romo2datao10_s_5_BXINV_4854 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_5_BXINV
    );
  romo2datao10_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_5_F6MUX,
      O => romo2datao10_s(5)
    );
  romo2datao10_s_5_F6MUX_4855 : X_MUX2
    port map (
      IA => nx53675z1550,
      IB => nx53675z1553,
      SEL => romo2datao10_s_5_BYINV,
      O => romo2datao10_s_5_F6MUX
    );
  romo2datao10_s_5_BYINV_4856 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_5_BYINV
    );
  nx53675z1550_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1550_F5MUX,
      O => nx53675z1550
    );
  nx53675z1550_F5MUX_4857 : X_MUX2
    port map (
      IA => nx53675z1551,
      IB => nx53675z1552,
      SEL => nx53675z1550_BXINV,
      O => nx53675z1550_F5MUX
    );
  nx53675z1550_BXINV_4858 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1550_BXINV
    );
  romo2datao4_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_13_F5MUX,
      O => nx53675z1031
    );
  romo2datao4_s_13_F5MUX_4859 : X_MUX2
    port map (
      IA => nx53675z1032,
      IB => nx53675z1033,
      SEL => romo2datao4_s_13_BXINV,
      O => romo2datao4_s_13_F5MUX
    );
  romo2datao4_s_13_BXINV_4860 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_13_BXINV
    );
  romo2datao4_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_13_F6MUX,
      O => romo2datao4_s(13)
    );
  romo2datao4_s_13_F6MUX_4861 : X_MUX2
    port map (
      IA => nx53675z1029,
      IB => nx53675z1031,
      SEL => romo2datao4_s_13_BYINV,
      O => romo2datao4_s_13_F6MUX
    );
  romo2datao4_s_13_BYINV_4862 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_13_BYINV
    );
  nx53675z1029_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1029_F5MUX,
      O => nx53675z1029
    );
  nx53675z1029_F5MUX_4863 : X_MUX2
    port map (
      IA => nx53675z1029_G,
      IB => nx53675z1030,
      SEL => nx53675z1029_BXINV,
      O => nx53675z1029_F5MUX
    );
  nx53675z1029_BXINV_4864 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1029_BXINV
    );
  U_DCT2D_reg_databuf_reg_4_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_4_0_DXMUX,
      CE => U_DCT2D_databuf_reg_4_0_CEINV,
      CLK => U_DCT2D_databuf_reg_4_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_4_0_FFX_RST,
      O => U_DCT2D_databuf_reg_4_Q(0)
    );
  U_DCT2D_databuf_reg_4_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_4_0_FFX_RST
    );
  romo2datao1_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_2_F5MUX,
      O => nx53675z860
    );
  romo2datao1_s_2_F5MUX_4865 : X_MUX2
    port map (
      IA => nx53675z861,
      IB => nx53675z862,
      SEL => romo2datao1_s_2_BXINV,
      O => romo2datao1_s_2_F5MUX
    );
  romo2datao1_s_2_BXINV_4866 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_2_BXINV
    );
  romo2datao1_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_2_F6MUX,
      O => romo2datao1_s(2)
    );
  romo2datao1_s_2_F6MUX_4867 : X_MUX2
    port map (
      IA => nx53675z857,
      IB => nx53675z860,
      SEL => romo2datao1_s_2_BYINV,
      O => romo2datao1_s_2_F6MUX
    );
  romo2datao1_s_2_BYINV_4868 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_2_BYINV
    );
  nx53675z857_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z857_F5MUX,
      O => nx53675z857
    );
  nx53675z857_F5MUX_4869 : X_MUX2
    port map (
      IA => nx53675z858,
      IB => nx53675z859,
      SEL => nx53675z857_BXINV,
      O => nx53675z857_F5MUX
    );
  nx53675z857_BXINV_4870 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z857_BXINV
    );
  romo2datao1_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_1_F5MUX,
      O => nx53675z866
    );
  romo2datao1_s_1_F5MUX_4871 : X_MUX2
    port map (
      IA => nx53675z867,
      IB => nx53675z868,
      SEL => romo2datao1_s_1_BXINV,
      O => romo2datao1_s_1_F5MUX
    );
  romo2datao1_s_1_BXINV_4872 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao1_s_1_BXINV
    );
  romo2datao1_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao1_s_1_F6MUX,
      O => romo2datao1_s(1)
    );
  romo2datao1_s_1_F6MUX_4873 : X_MUX2
    port map (
      IA => nx53675z863,
      IB => nx53675z866,
      SEL => romo2datao1_s_1_BYINV,
      O => romo2datao1_s_1_F6MUX
    );
  romo2datao1_s_1_BYINV_4874 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao1_s_1_BYINV
    );
  U_DCT2D_ix52543z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_0_3_Q,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_7_3_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx52543z1
    );
  nx53675z863_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z863_F5MUX,
      O => nx53675z863
    );
  nx53675z863_F5MUX_4875 : X_MUX2
    port map (
      IA => nx53675z864,
      IB => nx53675z865,
      SEL => nx53675z863_BXINV,
      O => nx53675z863_F5MUX
    );
  nx53675z863_BXINV_4876 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z863_BXINV
    );
  rome2datao7_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_13_F5MUX,
      O => nx53675z457
    );
  rome2datao7_s_13_F5MUX_4877 : X_MUX2
    port map (
      IA => nx53675z458,
      IB => nx53675z459,
      SEL => rome2datao7_s_13_BXINV,
      O => rome2datao7_s_13_F5MUX
    );
  rome2datao7_s_13_BXINV_4878 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao7_s_13_BXINV
    );
  rome2datao7_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_13_F6MUX,
      O => rome2datao7_s(13)
    );
  rome2datao7_s_13_F6MUX_4879 : X_MUX2
    port map (
      IA => nx53675z455,
      IB => nx53675z457,
      SEL => rome2datao7_s_13_BYINV,
      O => rome2datao7_s_13_F6MUX
    );
  rome2datao7_s_13_BYINV_4880 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao7_s_13_BYINV
    );
  nx53675z455_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z455_F5MUX,
      O => nx53675z455
    );
  nx53675z455_F5MUX_4881 : X_MUX2
    port map (
      IA => nx53675z455_G,
      IB => nx53675z456,
      SEL => nx53675z455_BXINV,
      O => nx53675z455_F5MUX
    );
  nx53675z455_BXINV_4882 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z455_BXINV
    );
  rome2datao6_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_11_F5MUX,
      O => nx53675z404
    );
  rome2datao6_s_11_F5MUX_4883 : X_MUX2
    port map (
      IA => nx53675z405,
      IB => nx53675z406,
      SEL => rome2datao6_s_11_BXINV,
      O => rome2datao6_s_11_F5MUX
    );
  rome2datao6_s_11_BXINV_4884 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao6_s_11_BXINV
    );
  rome2datao6_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_11_F6MUX,
      O => rome2datao6_s(11)
    );
  rome2datao6_s_11_F6MUX_4885 : X_MUX2
    port map (
      IA => nx53675z401,
      IB => nx53675z404,
      SEL => rome2datao6_s_11_BYINV,
      O => rome2datao6_s_11_F6MUX
    );
  rome2datao6_s_11_BYINV_4886 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao6_s_11_BYINV
    );
  nx53675z401_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z401_F5MUX,
      O => nx53675z401
    );
  nx53675z401_F5MUX_4887 : X_MUX2
    port map (
      IA => nx53675z402,
      IB => nx53675z403,
      SEL => nx53675z401_BXINV,
      O => nx53675z401_F5MUX
    );
  nx53675z401_BXINV_4888 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z401_BXINV
    );
  rome2datao6_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_10_F5MUX,
      O => nx53675z410
    );
  rome2datao6_s_10_F5MUX_4889 : X_MUX2
    port map (
      IA => nx53675z411,
      IB => nx53675z412,
      SEL => rome2datao6_s_10_BXINV,
      O => rome2datao6_s_10_F5MUX
    );
  rome2datao6_s_10_BXINV_4890 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao6_s_10_BXINV
    );
  rome2datao6_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_10_F6MUX,
      O => rome2datao6_s(10)
    );
  rome2datao6_s_10_F6MUX_4891 : X_MUX2
    port map (
      IA => nx53675z407,
      IB => nx53675z410,
      SEL => rome2datao6_s_10_BYINV,
      O => rome2datao6_s_10_F6MUX
    );
  rome2datao6_s_10_BYINV_4892 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao6_s_10_BYINV
    );
  nx53675z407_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z407_F5MUX,
      O => nx53675z407
    );
  nx53675z407_F5MUX_4893 : X_MUX2
    port map (
      IA => nx53675z408,
      IB => nx53675z409,
      SEL => nx53675z407_BXINV,
      O => nx53675z407_F5MUX
    );
  nx53675z407_BXINV_4894 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z407_BXINV
    );
  rome2datao6_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_9_F5MUX,
      O => nx53675z416
    );
  rome2datao6_s_9_F5MUX_4895 : X_MUX2
    port map (
      IA => nx53675z417,
      IB => nx53675z418,
      SEL => rome2datao6_s_9_BXINV,
      O => rome2datao6_s_9_F5MUX
    );
  rome2datao6_s_9_BXINV_4896 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao6_s_9_BXINV
    );
  rome2datao6_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_9_F6MUX,
      O => rome2datao6_s(9)
    );
  rome2datao6_s_9_F6MUX_4897 : X_MUX2
    port map (
      IA => nx53675z413,
      IB => nx53675z416,
      SEL => rome2datao6_s_9_BYINV,
      O => rome2datao6_s_9_F6MUX
    );
  rome2datao6_s_9_BYINV_4898 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao6_s_9_BYINV
    );
  nx53675z413_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z413_F5MUX,
      O => nx53675z413
    );
  nx53675z413_F5MUX_4899 : X_MUX2
    port map (
      IA => nx53675z414,
      IB => nx53675z415,
      SEL => nx53675z413_BXINV,
      O => nx53675z413_F5MUX
    );
  nx53675z413_BXINV_4900 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z413_BXINV
    );
  rome2datao6_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_8_F5MUX,
      O => nx53675z422
    );
  rome2datao6_s_8_F5MUX_4901 : X_MUX2
    port map (
      IA => nx53675z423,
      IB => nx53675z424,
      SEL => rome2datao6_s_8_BXINV,
      O => rome2datao6_s_8_F5MUX
    );
  rome2datao6_s_8_BXINV_4902 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao6_s_8_BXINV
    );
  rome2datao6_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_8_F6MUX,
      O => rome2datao6_s(8)
    );
  rome2datao6_s_8_F6MUX_4903 : X_MUX2
    port map (
      IA => nx53675z419,
      IB => nx53675z422,
      SEL => rome2datao6_s_8_BYINV,
      O => rome2datao6_s_8_F6MUX
    );
  rome2datao6_s_8_BYINV_4904 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao6_s_8_BYINV
    );
  nx53675z419_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z419_F5MUX,
      O => nx53675z419
    );
  nx53675z419_F5MUX_4905 : X_MUX2
    port map (
      IA => nx53675z420,
      IB => nx53675z421,
      SEL => nx53675z419_BXINV,
      O => nx53675z419_F5MUX
    );
  nx53675z419_BXINV_4906 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z419_BXINV
    );
  rome2datao6_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_7_F5MUX,
      O => nx53675z428
    );
  rome2datao6_s_7_F5MUX_4907 : X_MUX2
    port map (
      IA => nx53675z429,
      IB => nx53675z430,
      SEL => rome2datao6_s_7_BXINV,
      O => rome2datao6_s_7_F5MUX
    );
  rome2datao6_s_7_BXINV_4908 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao6_s_7_BXINV
    );
  rome2datao6_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_7_F6MUX,
      O => rome2datao6_s(7)
    );
  rome2datao6_s_7_F6MUX_4909 : X_MUX2
    port map (
      IA => nx53675z425,
      IB => nx53675z428,
      SEL => rome2datao6_s_7_BYINV,
      O => rome2datao6_s_7_F6MUX
    );
  rome2datao6_s_7_BYINV_4910 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao6_s_7_BYINV
    );
  nx53675z425_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z425_F5MUX,
      O => nx53675z425
    );
  nx53675z425_F5MUX_4911 : X_MUX2
    port map (
      IA => nx53675z426,
      IB => nx53675z427,
      SEL => nx53675z425_BXINV,
      O => nx53675z425_F5MUX
    );
  nx53675z425_BXINV_4912 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z425_BXINV
    );
  romo2datao4_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_3_F5MUX,
      O => nx53675z1091
    );
  romo2datao4_s_3_F5MUX_4913 : X_MUX2
    port map (
      IA => nx53675z1092,
      IB => nx53675z1093,
      SEL => romo2datao4_s_3_BXINV,
      O => romo2datao4_s_3_F5MUX
    );
  romo2datao4_s_3_BXINV_4914 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_3_BXINV
    );
  romo2datao4_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_3_F6MUX,
      O => romo2datao4_s(3)
    );
  romo2datao4_s_3_F6MUX_4915 : X_MUX2
    port map (
      IA => nx53675z1088,
      IB => nx53675z1091,
      SEL => romo2datao4_s_3_BYINV,
      O => romo2datao4_s_3_F6MUX
    );
  romo2datao4_s_3_BYINV_4916 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_3_BYINV
    );
  nx53675z1088_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1088_F5MUX,
      O => nx53675z1088
    );
  nx53675z1088_F5MUX_4917 : X_MUX2
    port map (
      IA => nx53675z1089,
      IB => nx53675z1090,
      SEL => nx53675z1088_BXINV,
      O => nx53675z1088_F5MUX
    );
  nx53675z1088_BXINV_4918 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1088_BXINV
    );
  romo2datao4_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_1_F5MUX,
      O => nx53675z1103
    );
  romo2datao4_s_1_F5MUX_4919 : X_MUX2
    port map (
      IA => nx53675z1104,
      IB => nx53675z1105,
      SEL => romo2datao4_s_1_BXINV,
      O => romo2datao4_s_1_F5MUX
    );
  romo2datao4_s_1_BXINV_4920 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_1_BXINV
    );
  romo2datao4_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_1_F6MUX,
      O => romo2datao4_s(1)
    );
  romo2datao4_s_1_F6MUX_4921 : X_MUX2
    port map (
      IA => nx53675z1100,
      IB => nx53675z1103,
      SEL => romo2datao4_s_1_BYINV,
      O => romo2datao4_s_1_F6MUX
    );
  romo2datao4_s_1_BYINV_4922 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_1_BYINV
    );
  nx53675z1100_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1100_F5MUX,
      O => nx53675z1100
    );
  nx53675z1100_F5MUX_4923 : X_MUX2
    port map (
      IA => nx53675z1101,
      IB => nx53675z1102,
      SEL => nx53675z1100_BXINV,
      O => nx53675z1100_F5MUX
    );
  nx53675z1100_BXINV_4924 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1100_BXINV
    );
  romo2datao6_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_8_F5MUX,
      O => nx53675z1219
    );
  romo2datao6_s_8_F5MUX_4925 : X_MUX2
    port map (
      IA => nx53675z1220,
      IB => nx53675z1221,
      SEL => romo2datao6_s_8_BXINV,
      O => romo2datao6_s_8_F5MUX
    );
  romo2datao6_s_8_BXINV_4926 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_8_BXINV
    );
  romo2datao6_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_8_F6MUX,
      O => romo2datao6_s(8)
    );
  romo2datao6_s_8_F6MUX_4927 : X_MUX2
    port map (
      IA => nx53675z1216,
      IB => nx53675z1219,
      SEL => romo2datao6_s_8_BYINV,
      O => romo2datao6_s_8_F6MUX
    );
  romo2datao6_s_8_BYINV_4928 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_8_BYINV
    );
  ix53675z5922 : X_LUT4
    generic map(
      INIT => X"0B42"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(2),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1217
    );
  nx53675z1216_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1216_F5MUX,
      O => nx53675z1216
    );
  nx53675z1216_F5MUX_4929 : X_MUX2
    port map (
      IA => nx53675z1217,
      IB => nx53675z1218,
      SEL => nx53675z1216_BXINV,
      O => nx53675z1216_F5MUX
    );
  nx53675z1216_BXINV_4930 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1216_BXINV
    );
  romo2datao6_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_7_F5MUX,
      O => nx53675z1225
    );
  romo2datao6_s_7_F5MUX_4931 : X_MUX2
    port map (
      IA => nx53675z1226,
      IB => nx53675z1227,
      SEL => romo2datao6_s_7_BXINV,
      O => romo2datao6_s_7_F5MUX
    );
  romo2datao6_s_7_BXINV_4932 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_7_BXINV
    );
  romo2datao6_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_7_F6MUX,
      O => romo2datao6_s(7)
    );
  romo2datao6_s_7_F6MUX_4933 : X_MUX2
    port map (
      IA => nx53675z1222,
      IB => nx53675z1225,
      SEL => romo2datao6_s_7_BYINV,
      O => romo2datao6_s_7_F6MUX
    );
  romo2datao6_s_7_BYINV_4934 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_7_BYINV
    );
  nx53675z1222_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1222_F5MUX,
      O => nx53675z1222
    );
  nx53675z1222_F5MUX_4935 : X_MUX2
    port map (
      IA => nx53675z1223,
      IB => nx53675z1224,
      SEL => nx53675z1222_BXINV,
      O => nx53675z1222_F5MUX
    );
  nx53675z1222_BXINV_4936 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1222_BXINV
    );
  romo2datao5_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_13_F5MUX,
      O => nx53675z1110
    );
  romo2datao5_s_13_F5MUX_4937 : X_MUX2
    port map (
      IA => nx53675z1111,
      IB => nx53675z1112,
      SEL => romo2datao5_s_13_BXINV,
      O => romo2datao5_s_13_F5MUX
    );
  romo2datao5_s_13_BXINV_4938 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_13_BXINV
    );
  romo2datao5_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_13_F6MUX,
      O => romo2datao5_s(13)
    );
  romo2datao5_s_13_F6MUX_4939 : X_MUX2
    port map (
      IA => nx53675z1108,
      IB => nx53675z1110,
      SEL => romo2datao5_s_13_BYINV,
      O => romo2datao5_s_13_F6MUX
    );
  romo2datao5_s_13_BYINV_4940 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_13_BYINV
    );
  nx53675z1108_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1108_F5MUX,
      O => nx53675z1108
    );
  nx53675z1108_F5MUX_4941 : X_MUX2
    port map (
      IA => nx53675z1108_G,
      IB => nx53675z1109,
      SEL => nx53675z1108_BXINV,
      O => nx53675z1108_F5MUX
    );
  nx53675z1108_BXINV_4942 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1108_BXINV
    );
  romo2datao5_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_6_F5MUX,
      O => nx53675z1152
    );
  romo2datao5_s_6_F5MUX_4943 : X_MUX2
    port map (
      IA => nx53675z1153,
      IB => nx53675z1154,
      SEL => romo2datao5_s_6_BXINV,
      O => romo2datao5_s_6_F5MUX
    );
  romo2datao5_s_6_BXINV_4944 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_6_BXINV
    );
  romo2datao5_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_6_F6MUX,
      O => romo2datao5_s(6)
    );
  romo2datao5_s_6_F6MUX_4945 : X_MUX2
    port map (
      IA => nx53675z1149,
      IB => nx53675z1152,
      SEL => romo2datao5_s_6_BYINV,
      O => romo2datao5_s_6_F6MUX
    );
  romo2datao5_s_6_BYINV_4946 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_6_BYINV
    );
  nx53675z1149_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1149_F5MUX,
      O => nx53675z1149
    );
  nx53675z1149_F5MUX_4947 : X_MUX2
    port map (
      IA => nx53675z1150,
      IB => nx53675z1151,
      SEL => nx53675z1149_BXINV,
      O => nx53675z1149_F5MUX
    );
  nx53675z1149_BXINV_4948 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1149_BXINV
    );
  romo2datao5_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_5_F5MUX,
      O => nx53675z1158
    );
  romo2datao5_s_5_F5MUX_4949 : X_MUX2
    port map (
      IA => nx53675z1159,
      IB => nx53675z1160,
      SEL => romo2datao5_s_5_BXINV,
      O => romo2datao5_s_5_F5MUX
    );
  romo2datao5_s_5_BXINV_4950 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_5_BXINV
    );
  romo2datao5_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_5_F6MUX,
      O => romo2datao5_s(5)
    );
  romo2datao5_s_5_F6MUX_4951 : X_MUX2
    port map (
      IA => nx53675z1155,
      IB => nx53675z1158,
      SEL => romo2datao5_s_5_BYINV,
      O => romo2datao5_s_5_F6MUX
    );
  romo2datao5_s_5_BYINV_4952 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_5_BYINV
    );
  nx53675z1155_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1155_F5MUX,
      O => nx53675z1155
    );
  nx53675z1155_F5MUX_4953 : X_MUX2
    port map (
      IA => nx53675z1156,
      IB => nx53675z1157,
      SEL => nx53675z1155_BXINV,
      O => nx53675z1155_F5MUX
    );
  nx53675z1155_BXINV_4954 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1155_BXINV
    );
  romo2datao5_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_4_F5MUX,
      O => nx53675z1164
    );
  romo2datao5_s_4_F5MUX_4955 : X_MUX2
    port map (
      IA => nx53675z1165,
      IB => nx53675z1166,
      SEL => romo2datao5_s_4_BXINV,
      O => romo2datao5_s_4_F5MUX
    );
  romo2datao5_s_4_BXINV_4956 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_4_BXINV
    );
  romo2datao5_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_4_F6MUX,
      O => romo2datao5_s(4)
    );
  romo2datao5_s_4_F6MUX_4957 : X_MUX2
    port map (
      IA => nx53675z1161,
      IB => nx53675z1164,
      SEL => romo2datao5_s_4_BYINV,
      O => romo2datao5_s_4_F6MUX
    );
  romo2datao5_s_4_BYINV_4958 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_4_BYINV
    );
  nx53675z1161_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1161_F5MUX,
      O => nx53675z1161
    );
  nx53675z1161_F5MUX_4959 : X_MUX2
    port map (
      IA => nx53675z1162,
      IB => nx53675z1163,
      SEL => nx53675z1161_BXINV,
      O => nx53675z1161_F5MUX
    );
  nx53675z1161_BXINV_4960 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1161_BXINV
    );
  romo2datao5_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_3_F5MUX,
      O => nx53675z1170
    );
  romo2datao5_s_3_F5MUX_4961 : X_MUX2
    port map (
      IA => nx53675z1171,
      IB => nx53675z1172,
      SEL => romo2datao5_s_3_BXINV,
      O => romo2datao5_s_3_F5MUX
    );
  romo2datao5_s_3_BXINV_4962 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_3_BXINV
    );
  romo2datao5_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_3_F6MUX,
      O => romo2datao5_s(3)
    );
  romo2datao5_s_3_F6MUX_4963 : X_MUX2
    port map (
      IA => nx53675z1167,
      IB => nx53675z1170,
      SEL => romo2datao5_s_3_BYINV,
      O => romo2datao5_s_3_F6MUX
    );
  romo2datao5_s_3_BYINV_4964 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_3_BYINV
    );
  nx53675z1167_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1167_F5MUX,
      O => nx53675z1167
    );
  nx53675z1167_F5MUX_4965 : X_MUX2
    port map (
      IA => nx53675z1168,
      IB => nx53675z1169,
      SEL => nx53675z1167_BXINV,
      O => nx53675z1167_F5MUX
    );
  nx53675z1167_BXINV_4966 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1167_BXINV
    );
  romo2datao4_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_0_F5MUX,
      O => U2_ROMO4_modgen_rom_ix0_nx_ro64_32_l
    );
  romo2datao4_s_0_F5MUX_4967 : X_MUX2
    port map (
      IA => nx53675z1106,
      IB => nx53675z1107,
      SEL => romo2datao4_s_0_BXINV,
      O => romo2datao4_s_0_F5MUX
    );
  romo2datao4_s_0_BXINV_4968 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_0_BXINV
    );
  romo2datao4_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_0_F6MUX,
      O => romo2datao4_s(0)
    );
  romo2datao4_s_0_F6MUX_4969 : X_MUX2
    port map (
      IA => U2_ROMO4_modgen_rom_ix0_nx_ro64_32_u,
      IB => U2_ROMO4_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romo2datao4_s_0_BYINV,
      O => romo2datao4_s_0_F6MUX
    );
  romo2datao4_s_0_BYINV_4970 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_0_BYINV
    );
  U2_ROMO4_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROMO4_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U2_ROMO4_modgen_rom_ix0_nx_ro64_32_u
    );
  U2_ROMO4_modgen_rom_ix0_nx_ro64_32_u_F5MUX_4971 : X_MUX2
    port map (
      IA => U2_ROMO4_modgen_rom_ix0_nx_rm64_16_u,
      IB => U2_ROMO4_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U2_ROMO4_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U2_ROMO4_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U2_ROMO4_modgen_rom_ix0_nx_ro64_32_u_BXINV_4972 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => U2_ROMO4_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  rome2datao8_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_12_F5MUX,
      O => nx53675z528
    );
  rome2datao8_s_12_F5MUX_4973 : X_MUX2
    port map (
      IA => nx53675z529,
      IB => nx53675z530,
      SEL => rome2datao8_s_12_BXINV,
      O => rome2datao8_s_12_F5MUX
    );
  rome2datao8_s_12_BXINV_4974 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao8_s_12_BXINV
    );
  rome2datao8_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_12_F6MUX,
      O => rome2datao8_s(12)
    );
  rome2datao8_s_12_F6MUX_4975 : X_MUX2
    port map (
      IA => nx53675z525,
      IB => nx53675z528,
      SEL => rome2datao8_s_12_BYINV,
      O => rome2datao8_s_12_F6MUX
    );
  rome2datao8_s_12_BYINV_4976 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao8_s_12_BYINV
    );
  nx53675z525_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z525_F5MUX,
      O => nx53675z525
    );
  nx53675z525_F5MUX_4977 : X_MUX2
    port map (
      IA => nx53675z526,
      IB => nx53675z527,
      SEL => nx53675z525_BXINV,
      O => nx53675z525_F5MUX
    );
  nx53675z525_BXINV_4978 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z525_BXINV
    );
  U_DCT2D_reg_databuf_reg_4_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_4_2_DYMUX,
      CE => U_DCT2D_databuf_reg_4_2_CEINV,
      CLK => U_DCT2D_databuf_reg_4_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_4_2_FFY_RST,
      O => U_DCT2D_databuf_reg_4_Q(3)
    );
  U_DCT2D_databuf_reg_4_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_4_2_FFY_RST
    );
  rome2datao8_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_11_F5MUX,
      O => nx53675z534
    );
  rome2datao8_s_11_F5MUX_4979 : X_MUX2
    port map (
      IA => nx53675z535,
      IB => nx53675z536,
      SEL => rome2datao8_s_11_BXINV,
      O => rome2datao8_s_11_F5MUX
    );
  rome2datao8_s_11_BXINV_4980 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao8_s_11_BXINV
    );
  rome2datao8_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_11_F6MUX,
      O => rome2datao8_s(11)
    );
  rome2datao8_s_11_F6MUX_4981 : X_MUX2
    port map (
      IA => nx53675z531,
      IB => nx53675z534,
      SEL => rome2datao8_s_11_BYINV,
      O => rome2datao8_s_11_F6MUX
    );
  rome2datao8_s_11_BYINV_4982 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao8_s_11_BYINV
    );
  nx53675z531_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z531_F5MUX,
      O => nx53675z531
    );
  nx53675z531_F5MUX_4983 : X_MUX2
    port map (
      IA => nx53675z532,
      IB => nx53675z533,
      SEL => nx53675z531_BXINV,
      O => nx53675z531_F5MUX
    );
  nx53675z531_BXINV_4984 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z531_BXINV
    );
  rome2datao8_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_10_F5MUX,
      O => nx53675z540
    );
  rome2datao8_s_10_F5MUX_4985 : X_MUX2
    port map (
      IA => nx53675z541,
      IB => nx53675z542,
      SEL => rome2datao8_s_10_BXINV,
      O => rome2datao8_s_10_F5MUX
    );
  rome2datao8_s_10_BXINV_4986 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao8_s_10_BXINV
    );
  rome2datao8_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_10_F6MUX,
      O => rome2datao8_s(10)
    );
  rome2datao8_s_10_F6MUX_4987 : X_MUX2
    port map (
      IA => nx53675z537,
      IB => nx53675z540,
      SEL => rome2datao8_s_10_BYINV,
      O => rome2datao8_s_10_F6MUX
    );
  rome2datao8_s_10_BYINV_4988 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao8_s_10_BYINV
    );
  nx53675z537_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z537_F5MUX,
      O => nx53675z537
    );
  nx53675z537_F5MUX_4989 : X_MUX2
    port map (
      IA => nx53675z538,
      IB => nx53675z539,
      SEL => nx53675z537_BXINV,
      O => nx53675z537_F5MUX
    );
  nx53675z537_BXINV_4990 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z537_BXINV
    );
  rome2datao8_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_9_F5MUX,
      O => nx53675z546
    );
  rome2datao8_s_9_F5MUX_4991 : X_MUX2
    port map (
      IA => nx53675z547,
      IB => nx53675z548,
      SEL => rome2datao8_s_9_BXINV,
      O => rome2datao8_s_9_F5MUX
    );
  rome2datao8_s_9_BXINV_4992 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao8_s_9_BXINV
    );
  rome2datao8_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_9_F6MUX,
      O => rome2datao8_s(9)
    );
  rome2datao8_s_9_F6MUX_4993 : X_MUX2
    port map (
      IA => nx53675z543,
      IB => nx53675z546,
      SEL => rome2datao8_s_9_BYINV,
      O => rome2datao8_s_9_F6MUX
    );
  rome2datao8_s_9_BYINV_4994 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao8_s_9_BYINV
    );
  nx53675z543_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z543_F5MUX,
      O => nx53675z543
    );
  nx53675z543_F5MUX_4995 : X_MUX2
    port map (
      IA => nx53675z544,
      IB => nx53675z545,
      SEL => nx53675z543_BXINV,
      O => nx53675z543_F5MUX
    );
  nx53675z543_BXINV_4996 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z543_BXINV
    );
  rome2datao4_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_13_F5MUX,
      O => nx53675z262
    );
  rome2datao4_s_13_F5MUX_4997 : X_MUX2
    port map (
      IA => nx53675z263,
      IB => nx53675z264,
      SEL => rome2datao4_s_13_BXINV,
      O => rome2datao4_s_13_F5MUX
    );
  rome2datao4_s_13_BXINV_4998 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao4_s_13_BXINV
    );
  rome2datao4_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao4_s_13_F6MUX,
      O => rome2datao4_s(13)
    );
  rome2datao4_s_13_F6MUX_4999 : X_MUX2
    port map (
      IA => nx53675z260,
      IB => nx53675z262,
      SEL => rome2datao4_s_13_BYINV,
      O => rome2datao4_s_13_F6MUX
    );
  rome2datao4_s_13_BYINV_5000 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao4_s_13_BYINV
    );
  nx53675z260_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z260_F5MUX,
      O => nx53675z260
    );
  nx53675z260_F5MUX_5001 : X_MUX2
    port map (
      IA => nx53675z260_G,
      IB => nx53675z261,
      SEL => nx53675z260_BXINV,
      O => nx53675z260_F5MUX
    );
  nx53675z260_BXINV_5002 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z260_BXINV
    );
  rome2datao8_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_13_F5MUX,
      O => nx53675z522
    );
  rome2datao8_s_13_F5MUX_5003 : X_MUX2
    port map (
      IA => nx53675z523,
      IB => nx53675z524,
      SEL => rome2datao8_s_13_BXINV,
      O => rome2datao8_s_13_F5MUX
    );
  rome2datao8_s_13_BXINV_5004 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao8_s_13_BXINV
    );
  rome2datao8_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_13_F6MUX,
      O => rome2datao8_s(13)
    );
  rome2datao8_s_13_F6MUX_5005 : X_MUX2
    port map (
      IA => nx53675z520,
      IB => nx53675z522,
      SEL => rome2datao8_s_13_BYINV,
      O => rome2datao8_s_13_F6MUX
    );
  rome2datao8_s_13_BYINV_5006 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao8_s_13_BYINV
    );
  nx53675z520_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z520_F5MUX,
      O => nx53675z520
    );
  nx53675z520_F5MUX_5007 : X_MUX2
    port map (
      IA => nx53675z520_G,
      IB => nx53675z521,
      SEL => nx53675z520_BXINV,
      O => nx53675z520_F5MUX
    );
  nx53675z520_BXINV_5008 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z520_BXINV
    );
  U_DCT2D_ix51546z1324 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_0_2_Q,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_7_2_Q,
      O => U_DCT2D_nx51546z1
    );
  rome2datao5_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_8_F5MUX,
      O => nx53675z357
    );
  rome2datao5_s_8_F5MUX_5009 : X_MUX2
    port map (
      IA => nx53675z358,
      IB => nx53675z359,
      SEL => rome2datao5_s_8_BXINV,
      O => rome2datao5_s_8_F5MUX
    );
  rome2datao5_s_8_BXINV_5010 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao5_s_8_BXINV
    );
  rome2datao5_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_8_F6MUX,
      O => rome2datao5_s(8)
    );
  rome2datao5_s_8_F6MUX_5011 : X_MUX2
    port map (
      IA => nx53675z354,
      IB => nx53675z357,
      SEL => rome2datao5_s_8_BYINV,
      O => rome2datao5_s_8_F6MUX
    );
  rome2datao5_s_8_BYINV_5012 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao5_s_8_BYINV
    );
  nx53675z354_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z354_F5MUX,
      O => nx53675z354
    );
  nx53675z354_F5MUX_5013 : X_MUX2
    port map (
      IA => nx53675z355,
      IB => nx53675z356,
      SEL => nx53675z354_BXINV,
      O => nx53675z354_F5MUX
    );
  nx53675z354_BXINV_5014 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z354_BXINV
    );
  rome2datao5_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_7_F5MUX,
      O => nx53675z363
    );
  rome2datao5_s_7_F5MUX_5015 : X_MUX2
    port map (
      IA => nx53675z364,
      IB => nx53675z365,
      SEL => rome2datao5_s_7_BXINV,
      O => rome2datao5_s_7_F5MUX
    );
  rome2datao5_s_7_BXINV_5016 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao5_s_7_BXINV
    );
  rome2datao5_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_7_F6MUX,
      O => rome2datao5_s(7)
    );
  rome2datao5_s_7_F6MUX_5017 : X_MUX2
    port map (
      IA => nx53675z360,
      IB => nx53675z363,
      SEL => rome2datao5_s_7_BYINV,
      O => rome2datao5_s_7_F6MUX
    );
  rome2datao5_s_7_BYINV_5018 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao5_s_7_BYINV
    );
  nx53675z360_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z360_F5MUX,
      O => nx53675z360
    );
  nx53675z360_F5MUX_5019 : X_MUX2
    port map (
      IA => nx53675z361,
      IB => nx53675z362,
      SEL => nx53675z360_BXINV,
      O => nx53675z360_F5MUX
    );
  nx53675z360_BXINV_5020 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z360_BXINV
    );
  rome2datao5_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_6_F5MUX,
      O => nx53675z369
    );
  rome2datao5_s_6_F5MUX_5021 : X_MUX2
    port map (
      IA => nx53675z370,
      IB => nx53675z371,
      SEL => rome2datao5_s_6_BXINV,
      O => rome2datao5_s_6_F5MUX
    );
  rome2datao5_s_6_BXINV_5022 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao5_s_6_BXINV
    );
  rome2datao5_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao5_s_6_F6MUX,
      O => rome2datao5_s(6)
    );
  rome2datao5_s_6_F6MUX_5023 : X_MUX2
    port map (
      IA => nx53675z366,
      IB => nx53675z369,
      SEL => rome2datao5_s_6_BYINV,
      O => rome2datao5_s_6_F6MUX
    );
  rome2datao5_s_6_BYINV_5024 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao5_s_6_BYINV
    );
  nx53675z366_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z366_F5MUX,
      O => nx53675z366
    );
  nx53675z366_F5MUX_5025 : X_MUX2
    port map (
      IA => nx53675z367,
      IB => nx53675z368,
      SEL => nx53675z366_BXINV,
      O => nx53675z366_F5MUX
    );
  nx53675z366_BXINV_5026 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z366_BXINV
    );
  rome2datao7_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_10_F5MUX,
      O => nx53675z475
    );
  rome2datao7_s_10_F5MUX_5027 : X_MUX2
    port map (
      IA => nx53675z476,
      IB => nx53675z477,
      SEL => rome2datao7_s_10_BXINV,
      O => rome2datao7_s_10_F5MUX
    );
  rome2datao7_s_10_BXINV_5028 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao7_s_10_BXINV
    );
  rome2datao7_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_10_F6MUX,
      O => rome2datao7_s(10)
    );
  rome2datao7_s_10_F6MUX_5029 : X_MUX2
    port map (
      IA => nx53675z472,
      IB => nx53675z475,
      SEL => rome2datao7_s_10_BYINV,
      O => rome2datao7_s_10_F6MUX
    );
  rome2datao7_s_10_BYINV_5030 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao7_s_10_BYINV
    );
  nx53675z472_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z472_F5MUX,
      O => nx53675z472
    );
  nx53675z472_F5MUX_5031 : X_MUX2
    port map (
      IA => nx53675z473,
      IB => nx53675z474,
      SEL => nx53675z472_BXINV,
      O => nx53675z472_F5MUX
    );
  nx53675z472_BXINV_5032 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z472_BXINV
    );
  rome2datao7_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_9_F5MUX,
      O => nx53675z481
    );
  rome2datao7_s_9_F5MUX_5033 : X_MUX2
    port map (
      IA => nx53675z482,
      IB => nx53675z483,
      SEL => rome2datao7_s_9_BXINV,
      O => rome2datao7_s_9_F5MUX
    );
  rome2datao7_s_9_BXINV_5034 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao7_s_9_BXINV
    );
  rome2datao7_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_9_F6MUX,
      O => rome2datao7_s(9)
    );
  rome2datao7_s_9_F6MUX_5035 : X_MUX2
    port map (
      IA => nx53675z478,
      IB => nx53675z481,
      SEL => rome2datao7_s_9_BYINV,
      O => rome2datao7_s_9_F6MUX
    );
  rome2datao7_s_9_BYINV_5036 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao7_s_9_BYINV
    );
  nx53675z478_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z478_F5MUX,
      O => nx53675z478
    );
  nx53675z478_F5MUX_5037 : X_MUX2
    port map (
      IA => nx53675z479,
      IB => nx53675z480,
      SEL => nx53675z478_BXINV,
      O => nx53675z478_F5MUX
    );
  nx53675z478_BXINV_5038 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z478_BXINV
    );
  rome2datao7_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_8_F5MUX,
      O => nx53675z487
    );
  rome2datao7_s_8_F5MUX_5039 : X_MUX2
    port map (
      IA => nx53675z488,
      IB => nx53675z489,
      SEL => rome2datao7_s_8_BXINV,
      O => rome2datao7_s_8_F5MUX
    );
  rome2datao7_s_8_BXINV_5040 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao7_s_8_BXINV
    );
  rome2datao7_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_8_F6MUX,
      O => rome2datao7_s(8)
    );
  rome2datao7_s_8_F6MUX_5041 : X_MUX2
    port map (
      IA => nx53675z484,
      IB => nx53675z487,
      SEL => rome2datao7_s_8_BYINV,
      O => rome2datao7_s_8_F6MUX
    );
  rome2datao7_s_8_BYINV_5042 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao7_s_8_BYINV
    );
  nx53675z484_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z484_F5MUX,
      O => nx53675z484
    );
  nx53675z484_F5MUX_5043 : X_MUX2
    port map (
      IA => nx53675z485,
      IB => nx53675z486,
      SEL => nx53675z484_BXINV,
      O => nx53675z484_F5MUX
    );
  nx53675z484_BXINV_5044 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z484_BXINV
    );
  rome2datao7_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_7_F5MUX,
      O => nx53675z493
    );
  rome2datao7_s_7_F5MUX_5045 : X_MUX2
    port map (
      IA => nx53675z494,
      IB => nx53675z495,
      SEL => rome2datao7_s_7_BXINV,
      O => rome2datao7_s_7_F5MUX
    );
  rome2datao7_s_7_BXINV_5046 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao7_s_7_BXINV
    );
  rome2datao7_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_7_F6MUX,
      O => rome2datao7_s(7)
    );
  rome2datao7_s_7_F6MUX_5047 : X_MUX2
    port map (
      IA => nx53675z490,
      IB => nx53675z493,
      SEL => rome2datao7_s_7_BYINV,
      O => rome2datao7_s_7_F6MUX
    );
  rome2datao7_s_7_BYINV_5048 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao7_s_7_BYINV
    );
  nx53675z490_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z490_F5MUX,
      O => nx53675z490
    );
  nx53675z490_F5MUX_5049 : X_MUX2
    port map (
      IA => nx53675z491,
      IB => nx53675z492,
      SEL => nx53675z490_BXINV,
      O => nx53675z490_F5MUX
    );
  nx53675z490_BXINV_5050 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z490_BXINV
    );
  rome2datao7_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_6_F5MUX,
      O => nx53675z499
    );
  rome2datao7_s_6_F5MUX_5051 : X_MUX2
    port map (
      IA => nx53675z500,
      IB => nx53675z501,
      SEL => rome2datao7_s_6_BXINV,
      O => rome2datao7_s_6_F5MUX
    );
  rome2datao7_s_6_BXINV_5052 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao7_s_6_BXINV
    );
  rome2datao7_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_6_F6MUX,
      O => rome2datao7_s(6)
    );
  rome2datao7_s_6_F6MUX_5053 : X_MUX2
    port map (
      IA => nx53675z496,
      IB => nx53675z499,
      SEL => rome2datao7_s_6_BYINV,
      O => rome2datao7_s_6_F6MUX
    );
  rome2datao7_s_6_BYINV_5054 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao7_s_6_BYINV
    );
  nx53675z496_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z496_F5MUX,
      O => nx53675z496
    );
  nx53675z496_F5MUX_5055 : X_MUX2
    port map (
      IA => nx53675z497,
      IB => nx53675z498,
      SEL => nx53675z496_BXINV,
      O => nx53675z496_F5MUX
    );
  nx53675z496_BXINV_5056 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z496_BXINV
    );
  romo2datao9_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_12_F5MUX,
      O => nx53675z1432
    );
  romo2datao9_s_12_F5MUX_5057 : X_MUX2
    port map (
      IA => nx53675z1433,
      IB => nx53675z1434,
      SEL => romo2datao9_s_12_BXINV,
      O => romo2datao9_s_12_F5MUX
    );
  romo2datao9_s_12_BXINV_5058 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_12_BXINV
    );
  romo2datao9_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_12_F6MUX,
      O => romo2datao9_s(12)
    );
  romo2datao9_s_12_F6MUX_5059 : X_MUX2
    port map (
      IA => nx53675z1429,
      IB => nx53675z1432,
      SEL => romo2datao9_s_12_BYINV,
      O => romo2datao9_s_12_F6MUX
    );
  romo2datao9_s_12_BYINV_5060 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_12_BYINV
    );
  nx53675z1429_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1429_F5MUX,
      O => nx53675z1429
    );
  nx53675z1429_F5MUX_5061 : X_MUX2
    port map (
      IA => nx53675z1430,
      IB => nx53675z1431,
      SEL => nx53675z1429_BXINV,
      O => nx53675z1429_F5MUX
    );
  nx53675z1429_BXINV_5062 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1429_BXINV
    );
  romo2datao5_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_12_F5MUX,
      O => nx53675z1116
    );
  romo2datao5_s_12_F5MUX_5063 : X_MUX2
    port map (
      IA => nx53675z1117,
      IB => nx53675z1118,
      SEL => romo2datao5_s_12_BXINV,
      O => romo2datao5_s_12_F5MUX
    );
  romo2datao5_s_12_BXINV_5064 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_12_BXINV
    );
  romo2datao5_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_12_F6MUX,
      O => romo2datao5_s(12)
    );
  romo2datao5_s_12_F6MUX_5065 : X_MUX2
    port map (
      IA => nx53675z1113,
      IB => nx53675z1116,
      SEL => romo2datao5_s_12_BYINV,
      O => romo2datao5_s_12_F6MUX
    );
  romo2datao5_s_12_BYINV_5066 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_12_BYINV
    );
  nx53675z1113_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1113_F5MUX,
      O => nx53675z1113
    );
  nx53675z1113_F5MUX_5067 : X_MUX2
    port map (
      IA => nx53675z1114,
      IB => nx53675z1115,
      SEL => nx53675z1113_BXINV,
      O => nx53675z1113_F5MUX
    );
  nx53675z1113_BXINV_5068 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1113_BXINV
    );
  U_DCT2D_reg_databuf_reg_4_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_4_2_DXMUX,
      CE => U_DCT2D_databuf_reg_4_2_CEINV,
      CLK => U_DCT2D_databuf_reg_4_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_4_2_FFX_RST,
      O => U_DCT2D_databuf_reg_4_Q(2)
    );
  U_DCT2D_databuf_reg_4_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_4_2_FFX_RST
    );
  romo2datao4_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_2_F5MUX,
      O => nx53675z1097
    );
  romo2datao4_s_2_F5MUX_5069 : X_MUX2
    port map (
      IA => nx53675z1098,
      IB => nx53675z1099,
      SEL => romo2datao4_s_2_BXINV,
      O => romo2datao4_s_2_F5MUX
    );
  romo2datao4_s_2_BXINV_5070 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_2_BXINV
    );
  romo2datao4_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_2_F6MUX,
      O => romo2datao4_s(2)
    );
  romo2datao4_s_2_F6MUX_5071 : X_MUX2
    port map (
      IA => nx53675z1094,
      IB => nx53675z1097,
      SEL => romo2datao4_s_2_BYINV,
      O => romo2datao4_s_2_F6MUX
    );
  romo2datao4_s_2_BYINV_5072 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_2_BYINV
    );
  nx53675z1094_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1094_F5MUX,
      O => nx53675z1094
    );
  nx53675z1094_F5MUX_5073 : X_MUX2
    port map (
      IA => nx53675z1095,
      IB => nx53675z1096,
      SEL => nx53675z1094_BXINV,
      O => nx53675z1094_F5MUX
    );
  nx53675z1094_BXINV_5074 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1094_BXINV
    );
  rome2datao3_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_9_F5MUX,
      O => nx53675z221
    );
  rome2datao3_s_9_F5MUX_5075 : X_MUX2
    port map (
      IA => nx53675z222,
      IB => nx53675z223,
      SEL => rome2datao3_s_9_BXINV,
      O => rome2datao3_s_9_F5MUX
    );
  rome2datao3_s_9_BXINV_5076 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao3_s_9_BXINV
    );
  rome2datao3_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_9_F6MUX,
      O => rome2datao3_s(9)
    );
  rome2datao3_s_9_F6MUX_5077 : X_MUX2
    port map (
      IA => nx53675z218,
      IB => nx53675z221,
      SEL => rome2datao3_s_9_BYINV,
      O => rome2datao3_s_9_F6MUX
    );
  rome2datao3_s_9_BYINV_5078 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao3_s_9_BYINV
    );
  U_DCT2D_ix54537z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_0_5_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_7_5_Q,
      O => U_DCT2D_nx54537z1
    );
  nx53675z218_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z218_F5MUX,
      O => nx53675z218
    );
  nx53675z218_F5MUX_5079 : X_MUX2
    port map (
      IA => nx53675z219,
      IB => nx53675z220,
      SEL => nx53675z218_BXINV,
      O => nx53675z218_F5MUX
    );
  nx53675z218_BXINV_5080 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z218_BXINV
    );
  rome2datao3_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_5_F5MUX,
      O => nx53675z245
    );
  rome2datao3_s_5_F5MUX_5081 : X_MUX2
    port map (
      IA => nx53675z246,
      IB => nx53675z247,
      SEL => rome2datao3_s_5_BXINV,
      O => rome2datao3_s_5_F5MUX
    );
  rome2datao3_s_5_BXINV_5082 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao3_s_5_BXINV
    );
  rome2datao3_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_5_F6MUX,
      O => rome2datao3_s(5)
    );
  rome2datao3_s_5_F6MUX_5083 : X_MUX2
    port map (
      IA => nx53675z242,
      IB => nx53675z245,
      SEL => rome2datao3_s_5_BYINV,
      O => rome2datao3_s_5_F6MUX
    );
  rome2datao3_s_5_BYINV_5084 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao3_s_5_BYINV
    );
  nx53675z242_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z242_F5MUX,
      O => nx53675z242
    );
  nx53675z242_F5MUX_5085 : X_MUX2
    port map (
      IA => nx53675z243,
      IB => nx53675z244,
      SEL => nx53675z242_BXINV,
      O => nx53675z242_F5MUX
    );
  nx53675z242_BXINV_5086 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z242_BXINV
    );
  rome2datao3_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_3_F5MUX,
      O => nx53675z256
    );
  rome2datao3_s_3_F5MUX_5087 : X_MUX2
    port map (
      IA => nx53675z257,
      IB => nx53675z258,
      SEL => rome2datao3_s_3_BXINV,
      O => rome2datao3_s_3_F5MUX
    );
  rome2datao3_s_3_BXINV_5088 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao3_s_3_BXINV
    );
  rome2datao3_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao3_s_3_F6MUX,
      O => rome2datao3_s(3)
    );
  rome2datao3_s_3_F6MUX_5089 : X_MUX2
    port map (
      IA => nx53675z254,
      IB => nx53675z256,
      SEL => rome2datao3_s_3_BYINV,
      O => rome2datao3_s_3_F6MUX
    );
  rome2datao3_s_3_BYINV_5090 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao3_s_3_BYINV
    );
  nx53675z254_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z254_F5MUX,
      O => nx53675z254
    );
  nx53675z254_F5MUX_5091 : X_MUX2
    port map (
      IA => U2_ROME3_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx53675z255,
      SEL => nx53675z254_BXINV,
      O => nx53675z254_F5MUX
    );
  nx53675z254_BXINV_5092 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z254_BXINV
    );
  romo2datao4_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_10_F5MUX,
      O => nx53675z1049
    );
  romo2datao4_s_10_F5MUX_5093 : X_MUX2
    port map (
      IA => nx53675z1050,
      IB => nx53675z1051,
      SEL => romo2datao4_s_10_BXINV,
      O => romo2datao4_s_10_F5MUX
    );
  romo2datao4_s_10_BXINV_5094 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_10_BXINV
    );
  romo2datao4_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_10_F6MUX,
      O => romo2datao4_s(10)
    );
  romo2datao4_s_10_F6MUX_5095 : X_MUX2
    port map (
      IA => nx53675z1046,
      IB => nx53675z1049,
      SEL => romo2datao4_s_10_BYINV,
      O => romo2datao4_s_10_F6MUX
    );
  romo2datao4_s_10_BYINV_5096 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_10_BYINV
    );
  nx53675z1046_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1046_F5MUX,
      O => nx53675z1046
    );
  nx53675z1046_F5MUX_5097 : X_MUX2
    port map (
      IA => nx53675z1047,
      IB => nx53675z1048,
      SEL => nx53675z1046_BXINV,
      O => nx53675z1046_F5MUX
    );
  nx53675z1046_BXINV_5098 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1046_BXINV
    );
  romo2datao3_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_6_F5MUX,
      O => nx53675z994
    );
  romo2datao3_s_6_F5MUX_5099 : X_MUX2
    port map (
      IA => nx53675z995,
      IB => nx53675z996,
      SEL => romo2datao3_s_6_BXINV,
      O => romo2datao3_s_6_F5MUX
    );
  romo2datao3_s_6_BXINV_5100 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_6_BXINV
    );
  romo2datao3_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_6_F6MUX,
      O => romo2datao3_s(6)
    );
  romo2datao3_s_6_F6MUX_5101 : X_MUX2
    port map (
      IA => nx53675z991,
      IB => nx53675z994,
      SEL => romo2datao3_s_6_BYINV,
      O => romo2datao3_s_6_F6MUX
    );
  romo2datao3_s_6_BYINV_5102 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_6_BYINV
    );
  nx53675z991_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z991_F5MUX,
      O => nx53675z991
    );
  nx53675z991_F5MUX_5103 : X_MUX2
    port map (
      IA => nx53675z992,
      IB => nx53675z993,
      SEL => nx53675z991_BXINV,
      O => nx53675z991_F5MUX
    );
  nx53675z991_BXINV_5104 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z991_BXINV
    );
  romo2datao3_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_4_F5MUX,
      O => nx53675z1006
    );
  romo2datao3_s_4_F5MUX_5105 : X_MUX2
    port map (
      IA => nx53675z1007,
      IB => nx53675z1008,
      SEL => romo2datao3_s_4_BXINV,
      O => romo2datao3_s_4_F5MUX
    );
  romo2datao3_s_4_BXINV_5106 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_4_BXINV
    );
  romo2datao3_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_4_F6MUX,
      O => romo2datao3_s(4)
    );
  romo2datao3_s_4_F6MUX_5107 : X_MUX2
    port map (
      IA => nx53675z1003,
      IB => nx53675z1006,
      SEL => romo2datao3_s_4_BYINV,
      O => romo2datao3_s_4_F6MUX
    );
  romo2datao3_s_4_BYINV_5108 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_4_BYINV
    );
  nx53675z1003_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1003_F5MUX,
      O => nx53675z1003
    );
  nx53675z1003_F5MUX_5109 : X_MUX2
    port map (
      IA => nx53675z1004,
      IB => nx53675z1005,
      SEL => nx53675z1003_BXINV,
      O => nx53675z1003_F5MUX
    );
  nx53675z1003_BXINV_5110 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1003_BXINV
    );
  romo2datao10_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_4_F5MUX,
      O => nx53675z1559
    );
  romo2datao10_s_4_F5MUX_5111 : X_MUX2
    port map (
      IA => nx53675z1560,
      IB => nx53675z1561,
      SEL => romo2datao10_s_4_BXINV,
      O => romo2datao10_s_4_F5MUX
    );
  romo2datao10_s_4_BXINV_5112 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_4_BXINV
    );
  romo2datao10_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_4_F6MUX,
      O => romo2datao10_s(4)
    );
  romo2datao10_s_4_F6MUX_5113 : X_MUX2
    port map (
      IA => nx53675z1556,
      IB => nx53675z1559,
      SEL => romo2datao10_s_4_BYINV,
      O => romo2datao10_s_4_F6MUX
    );
  romo2datao10_s_4_BYINV_5114 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_4_BYINV
    );
  nx53675z1556_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1556_F5MUX,
      O => nx53675z1556
    );
  nx53675z1556_F5MUX_5115 : X_MUX2
    port map (
      IA => nx53675z1557,
      IB => nx53675z1558,
      SEL => nx53675z1556_BXINV,
      O => nx53675z1556_F5MUX
    );
  nx53675z1556_BXINV_5116 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1556_BXINV
    );
  romo2datao10_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_3_F5MUX,
      O => nx53675z1565
    );
  romo2datao10_s_3_F5MUX_5117 : X_MUX2
    port map (
      IA => nx53675z1566,
      IB => nx53675z1567,
      SEL => romo2datao10_s_3_BXINV,
      O => romo2datao10_s_3_F5MUX
    );
  romo2datao10_s_3_BXINV_5118 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_3_BXINV
    );
  romo2datao10_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_3_F6MUX,
      O => romo2datao10_s(3)
    );
  romo2datao10_s_3_F6MUX_5119 : X_MUX2
    port map (
      IA => nx53675z1562,
      IB => nx53675z1565,
      SEL => romo2datao10_s_3_BYINV,
      O => romo2datao10_s_3_F6MUX
    );
  romo2datao10_s_3_BYINV_5120 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_3_BYINV
    );
  nx53675z1562_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1562_F5MUX,
      O => nx53675z1562
    );
  nx53675z1562_F5MUX_5121 : X_MUX2
    port map (
      IA => nx53675z1563,
      IB => nx53675z1564,
      SEL => nx53675z1562_BXINV,
      O => nx53675z1562_F5MUX
    );
  nx53675z1562_BXINV_5122 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1562_BXINV
    );
  romo2datao4_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_9_F5MUX,
      O => nx53675z1055
    );
  romo2datao4_s_9_F5MUX_5123 : X_MUX2
    port map (
      IA => nx53675z1056,
      IB => nx53675z1057,
      SEL => romo2datao4_s_9_BXINV,
      O => romo2datao4_s_9_F5MUX
    );
  romo2datao4_s_9_BXINV_5124 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_9_BXINV
    );
  romo2datao4_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_9_F6MUX,
      O => romo2datao4_s(9)
    );
  romo2datao4_s_9_F6MUX_5125 : X_MUX2
    port map (
      IA => nx53675z1052,
      IB => nx53675z1055,
      SEL => romo2datao4_s_9_BYINV,
      O => romo2datao4_s_9_F6MUX
    );
  romo2datao4_s_9_BYINV_5126 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_9_BYINV
    );
  nx53675z1052_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1052_F5MUX,
      O => nx53675z1052
    );
  nx53675z1052_F5MUX_5127 : X_MUX2
    port map (
      IA => nx53675z1053,
      IB => nx53675z1054,
      SEL => nx53675z1052_BXINV,
      O => nx53675z1052_F5MUX
    );
  nx53675z1052_BXINV_5128 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1052_BXINV
    );
  romo2datao4_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_8_F5MUX,
      O => nx53675z1061
    );
  romo2datao4_s_8_F5MUX_5129 : X_MUX2
    port map (
      IA => nx53675z1062,
      IB => nx53675z1063,
      SEL => romo2datao4_s_8_BXINV,
      O => romo2datao4_s_8_F5MUX
    );
  romo2datao4_s_8_BXINV_5130 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_8_BXINV
    );
  romo2datao4_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_8_F6MUX,
      O => romo2datao4_s(8)
    );
  romo2datao4_s_8_F6MUX_5131 : X_MUX2
    port map (
      IA => nx53675z1058,
      IB => nx53675z1061,
      SEL => romo2datao4_s_8_BYINV,
      O => romo2datao4_s_8_F6MUX
    );
  romo2datao4_s_8_BYINV_5132 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_8_BYINV
    );
  nx53675z1058_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1058_F5MUX,
      O => nx53675z1058
    );
  nx53675z1058_F5MUX_5133 : X_MUX2
    port map (
      IA => nx53675z1059,
      IB => nx53675z1060,
      SEL => nx53675z1058_BXINV,
      O => nx53675z1058_F5MUX
    );
  nx53675z1058_BXINV_5134 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1058_BXINV
    );
  romo2datao4_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_7_F5MUX,
      O => nx53675z1067
    );
  romo2datao4_s_7_F5MUX_5135 : X_MUX2
    port map (
      IA => nx53675z1068,
      IB => nx53675z1069,
      SEL => romo2datao4_s_7_BXINV,
      O => romo2datao4_s_7_F5MUX
    );
  romo2datao4_s_7_BXINV_5136 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_7_BXINV
    );
  romo2datao4_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_7_F6MUX,
      O => romo2datao4_s(7)
    );
  romo2datao4_s_7_F6MUX_5137 : X_MUX2
    port map (
      IA => nx53675z1064,
      IB => nx53675z1067,
      SEL => romo2datao4_s_7_BYINV,
      O => romo2datao4_s_7_F6MUX
    );
  romo2datao4_s_7_BYINV_5138 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_7_BYINV
    );
  nx53675z1064_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1064_F5MUX,
      O => nx53675z1064
    );
  nx53675z1064_F5MUX_5139 : X_MUX2
    port map (
      IA => nx53675z1065,
      IB => nx53675z1066,
      SEL => nx53675z1064_BXINV,
      O => nx53675z1064_F5MUX
    );
  nx53675z1064_BXINV_5140 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1064_BXINV
    );
  romo2datao4_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_6_F5MUX,
      O => nx53675z1073
    );
  romo2datao4_s_6_F5MUX_5141 : X_MUX2
    port map (
      IA => nx53675z1074,
      IB => nx53675z1075,
      SEL => romo2datao4_s_6_BXINV,
      O => romo2datao4_s_6_F5MUX
    );
  romo2datao4_s_6_BXINV_5142 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao4_s_6_BXINV
    );
  romo2datao4_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao4_s_6_F6MUX,
      O => romo2datao4_s(6)
    );
  romo2datao4_s_6_F6MUX_5143 : X_MUX2
    port map (
      IA => nx53675z1070,
      IB => nx53675z1073,
      SEL => romo2datao4_s_6_BYINV,
      O => romo2datao4_s_6_F6MUX
    );
  romo2datao4_s_6_BYINV_5144 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao4_s_6_BYINV
    );
  nx53675z1070_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1070_F5MUX,
      O => nx53675z1070
    );
  nx53675z1070_F5MUX_5145 : X_MUX2
    port map (
      IA => nx53675z1071,
      IB => nx53675z1072,
      SEL => nx53675z1070_BXINV,
      O => nx53675z1070_F5MUX
    );
  nx53675z1070_BXINV_5146 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1070_BXINV
    );
  rome2datao6_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_6_F5MUX,
      O => nx53675z434
    );
  rome2datao6_s_6_F5MUX_5147 : X_MUX2
    port map (
      IA => nx53675z435,
      IB => nx53675z436,
      SEL => rome2datao6_s_6_BXINV,
      O => rome2datao6_s_6_F5MUX
    );
  rome2datao6_s_6_BXINV_5148 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao6_s_6_BXINV
    );
  rome2datao6_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_6_F6MUX,
      O => rome2datao6_s(6)
    );
  rome2datao6_s_6_F6MUX_5149 : X_MUX2
    port map (
      IA => nx53675z431,
      IB => nx53675z434,
      SEL => rome2datao6_s_6_BYINV,
      O => rome2datao6_s_6_F6MUX
    );
  rome2datao6_s_6_BYINV_5150 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao6_s_6_BYINV
    );
  nx53675z431_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z431_F5MUX,
      O => nx53675z431
    );
  nx53675z431_F5MUX_5151 : X_MUX2
    port map (
      IA => nx53675z432,
      IB => nx53675z433,
      SEL => nx53675z431_BXINV,
      O => nx53675z431_F5MUX
    );
  nx53675z431_BXINV_5152 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z431_BXINV
    );
  rome2datao6_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_5_F5MUX,
      O => nx53675z440
    );
  rome2datao6_s_5_F5MUX_5153 : X_MUX2
    port map (
      IA => nx53675z441,
      IB => nx53675z442,
      SEL => rome2datao6_s_5_BXINV,
      O => rome2datao6_s_5_F5MUX
    );
  rome2datao6_s_5_BXINV_5154 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao6_s_5_BXINV
    );
  rome2datao6_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao6_s_5_F6MUX,
      O => rome2datao6_s(5)
    );
  rome2datao6_s_5_F6MUX_5155 : X_MUX2
    port map (
      IA => nx53675z437,
      IB => nx53675z440,
      SEL => rome2datao6_s_5_BYINV,
      O => rome2datao6_s_5_F6MUX
    );
  rome2datao6_s_5_BYINV_5156 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao6_s_5_BYINV
    );
  nx53675z437_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z437_F5MUX,
      O => nx53675z437
    );
  nx53675z437_F5MUX_5157 : X_MUX2
    port map (
      IA => nx53675z438,
      IB => nx53675z439,
      SEL => nx53675z437_BXINV,
      O => nx53675z437_F5MUX
    );
  nx53675z437_BXINV_5158 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z437_BXINV
    );
  romo2datao5_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_11_F5MUX,
      O => nx53675z1122
    );
  romo2datao5_s_11_F5MUX_5159 : X_MUX2
    port map (
      IA => nx53675z1123,
      IB => nx53675z1124,
      SEL => romo2datao5_s_11_BXINV,
      O => romo2datao5_s_11_F5MUX
    );
  romo2datao5_s_11_BXINV_5160 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_11_BXINV
    );
  romo2datao5_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_11_F6MUX,
      O => romo2datao5_s(11)
    );
  romo2datao5_s_11_F6MUX_5161 : X_MUX2
    port map (
      IA => nx53675z1119,
      IB => nx53675z1122,
      SEL => romo2datao5_s_11_BYINV,
      O => romo2datao5_s_11_F6MUX
    );
  romo2datao5_s_11_BYINV_5162 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_11_BYINV
    );
  nx53675z1119_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1119_F5MUX,
      O => nx53675z1119
    );
  nx53675z1119_F5MUX_5163 : X_MUX2
    port map (
      IA => nx53675z1120,
      IB => nx53675z1121,
      SEL => nx53675z1119_BXINV,
      O => nx53675z1119_F5MUX
    );
  nx53675z1119_BXINV_5164 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1119_BXINV
    );
  romo2datao9_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_1_F5MUX,
      O => nx53675z1498
    );
  romo2datao9_s_1_F5MUX_5165 : X_MUX2
    port map (
      IA => nx53675z1499,
      IB => nx53675z1500,
      SEL => romo2datao9_s_1_BXINV,
      O => romo2datao9_s_1_F5MUX
    );
  romo2datao9_s_1_BXINV_5166 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao9_s_1_BXINV
    );
  romo2datao9_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao9_s_1_F6MUX,
      O => romo2datao9_s(1)
    );
  romo2datao9_s_1_F6MUX_5167 : X_MUX2
    port map (
      IA => nx53675z1495,
      IB => nx53675z1498,
      SEL => romo2datao9_s_1_BYINV,
      O => romo2datao9_s_1_F6MUX
    );
  romo2datao9_s_1_BYINV_5168 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao9_s_1_BYINV
    );
  nx53675z1495_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1495_F5MUX,
      O => nx53675z1495
    );
  nx53675z1495_F5MUX_5169 : X_MUX2
    port map (
      IA => nx53675z1496,
      IB => nx53675z1497,
      SEL => nx53675z1495_BXINV,
      O => nx53675z1495_F5MUX
    );
  nx53675z1495_BXINV_5170 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1495_BXINV
    );
  romo2datao6_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_13_F5MUX,
      O => nx53675z1189
    );
  romo2datao6_s_13_F5MUX_5171 : X_MUX2
    port map (
      IA => nx53675z1190,
      IB => nx53675z1191,
      SEL => romo2datao6_s_13_BXINV,
      O => romo2datao6_s_13_F5MUX
    );
  romo2datao6_s_13_BXINV_5172 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_13_BXINV
    );
  romo2datao6_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_13_F6MUX,
      O => romo2datao6_s(13)
    );
  romo2datao6_s_13_F6MUX_5173 : X_MUX2
    port map (
      IA => nx53675z1187,
      IB => nx53675z1189,
      SEL => romo2datao6_s_13_BYINV,
      O => romo2datao6_s_13_F6MUX
    );
  romo2datao6_s_13_BYINV_5174 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_13_BYINV
    );
  U_DCT2D_ix4406z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_6_5_Q,
      ADR1 => U_DCT2D_latchbuf_reg_1_5_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx4406z1
    );
  U_DCT2D_reg_databuf_reg_1_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_1_4_DYMUX,
      CE => U_DCT2D_databuf_reg_1_4_CEINV,
      CLK => U_DCT2D_databuf_reg_1_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_1_4_FFY_RST,
      O => U_DCT2D_databuf_reg_1_Q(5)
    );
  U_DCT2D_databuf_reg_1_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_1_4_FFY_RST
    );
  U_DCT2D_ix3409z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_1_4_Q,
      ADR1 => U_DCT2D_latchbuf_reg_6_4_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx3409z1
    );
  U_DCT2D_reg_databuf_reg_1_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_1_4_DXMUX,
      CE => U_DCT2D_databuf_reg_1_4_CEINV,
      CLK => U_DCT2D_databuf_reg_1_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_1_4_FFX_RST,
      O => U_DCT2D_databuf_reg_1_Q(4)
    );
  U_DCT2D_databuf_reg_1_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_1_4_FFX_RST
    );
  U_DCT2D_ix6400z1321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_1_7_Q,
      ADR2 => U_DCT2D_latchbuf_reg_6_7_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx6400z1
    );
  nx53675z1187_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1187_F5MUX,
      O => nx53675z1187
    );
  nx53675z1187_F5MUX_5175 : X_MUX2
    port map (
      IA => nx53675z1187_G,
      IB => nx53675z1188,
      SEL => nx53675z1187_BXINV,
      O => nx53675z1187_F5MUX
    );
  nx53675z1187_BXINV_5176 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1187_BXINV
    );
  romo2datao6_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_6_F5MUX,
      O => nx53675z1231
    );
  romo2datao6_s_6_F5MUX_5177 : X_MUX2
    port map (
      IA => nx53675z1232,
      IB => nx53675z1233,
      SEL => romo2datao6_s_6_BXINV,
      O => romo2datao6_s_6_F5MUX
    );
  romo2datao6_s_6_BXINV_5178 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_6_BXINV
    );
  romo2datao6_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_6_F6MUX,
      O => romo2datao6_s(6)
    );
  romo2datao6_s_6_F6MUX_5179 : X_MUX2
    port map (
      IA => nx53675z1228,
      IB => nx53675z1231,
      SEL => romo2datao6_s_6_BYINV,
      O => romo2datao6_s_6_F6MUX
    );
  romo2datao6_s_6_BYINV_5180 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_6_BYINV
    );
  nx53675z1228_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1228_F5MUX,
      O => nx53675z1228
    );
  nx53675z1228_F5MUX_5181 : X_MUX2
    port map (
      IA => nx53675z1229,
      IB => nx53675z1230,
      SEL => nx53675z1228_BXINV,
      O => nx53675z1228_F5MUX
    );
  nx53675z1228_BXINV_5182 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1228_BXINV
    );
  U_DCT2D_reg_databuf_reg_4_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_4_4_DYMUX,
      CE => U_DCT2D_databuf_reg_4_4_CEINV,
      CLK => U_DCT2D_databuf_reg_4_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_4_4_FFY_RST,
      O => U_DCT2D_databuf_reg_4_Q(5)
    );
  U_DCT2D_databuf_reg_4_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_4_4_FFY_RST
    );
  romo2datao6_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_5_F5MUX,
      O => nx53675z1237
    );
  romo2datao6_s_5_F5MUX_5183 : X_MUX2
    port map (
      IA => nx53675z1238,
      IB => nx53675z1239,
      SEL => romo2datao6_s_5_BXINV,
      O => romo2datao6_s_5_F5MUX
    );
  romo2datao6_s_5_BXINV_5184 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_5_BXINV
    );
  romo2datao6_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_5_F6MUX,
      O => romo2datao6_s(5)
    );
  romo2datao6_s_5_F6MUX_5185 : X_MUX2
    port map (
      IA => nx53675z1234,
      IB => nx53675z1237,
      SEL => romo2datao6_s_5_BYINV,
      O => romo2datao6_s_5_F6MUX
    );
  romo2datao6_s_5_BYINV_5186 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_5_BYINV
    );
  nx53675z1234_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1234_F5MUX,
      O => nx53675z1234
    );
  nx53675z1234_F5MUX_5187 : X_MUX2
    port map (
      IA => nx53675z1235,
      IB => nx53675z1236,
      SEL => nx53675z1234_BXINV,
      O => nx53675z1234_F5MUX
    );
  nx53675z1234_BXINV_5188 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1234_BXINV
    );
  romo2datao6_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_4_F5MUX,
      O => nx53675z1243
    );
  romo2datao6_s_4_F5MUX_5189 : X_MUX2
    port map (
      IA => nx53675z1244,
      IB => nx53675z1245,
      SEL => romo2datao6_s_4_BXINV,
      O => romo2datao6_s_4_F5MUX
    );
  romo2datao6_s_4_BXINV_5190 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_4_BXINV
    );
  romo2datao6_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_4_F6MUX,
      O => romo2datao6_s(4)
    );
  romo2datao6_s_4_F6MUX_5191 : X_MUX2
    port map (
      IA => nx53675z1240,
      IB => nx53675z1243,
      SEL => romo2datao6_s_4_BYINV,
      O => romo2datao6_s_4_F6MUX
    );
  romo2datao6_s_4_BYINV_5192 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_4_BYINV
    );
  nx53675z1240_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1240_F5MUX,
      O => nx53675z1240
    );
  nx53675z1240_F5MUX_5193 : X_MUX2
    port map (
      IA => nx53675z1241,
      IB => nx53675z1242,
      SEL => nx53675z1240_BXINV,
      O => nx53675z1240_F5MUX
    );
  nx53675z1240_BXINV_5194 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1240_BXINV
    );
  romo2datao6_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_3_F5MUX,
      O => nx53675z1249
    );
  romo2datao6_s_3_F5MUX_5195 : X_MUX2
    port map (
      IA => nx53675z1250,
      IB => nx53675z1251,
      SEL => romo2datao6_s_3_BXINV,
      O => romo2datao6_s_3_F5MUX
    );
  romo2datao6_s_3_BXINV_5196 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_3_BXINV
    );
  romo2datao6_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_3_F6MUX,
      O => romo2datao6_s(3)
    );
  romo2datao6_s_3_F6MUX_5197 : X_MUX2
    port map (
      IA => nx53675z1246,
      IB => nx53675z1249,
      SEL => romo2datao6_s_3_BYINV,
      O => romo2datao6_s_3_F6MUX
    );
  romo2datao6_s_3_BYINV_5198 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_3_BYINV
    );
  nx53675z1246_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1246_F5MUX,
      O => nx53675z1246
    );
  nx53675z1246_F5MUX_5199 : X_MUX2
    port map (
      IA => nx53675z1247,
      IB => nx53675z1248,
      SEL => nx53675z1246_BXINV,
      O => nx53675z1246_F5MUX
    );
  nx53675z1246_BXINV_5200 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1246_BXINV
    );
  romo2datao6_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_2_F5MUX,
      O => nx53675z1255
    );
  romo2datao6_s_2_F5MUX_5201 : X_MUX2
    port map (
      IA => nx53675z1256,
      IB => nx53675z1257,
      SEL => romo2datao6_s_2_BXINV,
      O => romo2datao6_s_2_F5MUX
    );
  romo2datao6_s_2_BXINV_5202 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_2_BXINV
    );
  romo2datao6_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_2_F6MUX,
      O => romo2datao6_s(2)
    );
  romo2datao6_s_2_F6MUX_5203 : X_MUX2
    port map (
      IA => nx53675z1252,
      IB => nx53675z1255,
      SEL => romo2datao6_s_2_BYINV,
      O => romo2datao6_s_2_F6MUX
    );
  romo2datao6_s_2_BYINV_5204 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_2_BYINV
    );
  nx53675z1252_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1252_F5MUX,
      O => nx53675z1252
    );
  nx53675z1252_F5MUX_5205 : X_MUX2
    port map (
      IA => nx53675z1253,
      IB => nx53675z1254,
      SEL => nx53675z1252_BXINV,
      O => nx53675z1252_F5MUX
    );
  nx53675z1252_BXINV_5206 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1252_BXINV
    );
  romo2datao5_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_10_F5MUX,
      O => nx53675z1128
    );
  romo2datao5_s_10_F5MUX_5207 : X_MUX2
    port map (
      IA => nx53675z1129,
      IB => nx53675z1130,
      SEL => romo2datao5_s_10_BXINV,
      O => romo2datao5_s_10_F5MUX
    );
  romo2datao5_s_10_BXINV_5208 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_10_BXINV
    );
  romo2datao5_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_10_F6MUX,
      O => romo2datao5_s(10)
    );
  romo2datao5_s_10_F6MUX_5209 : X_MUX2
    port map (
      IA => nx53675z1125,
      IB => nx53675z1128,
      SEL => romo2datao5_s_10_BYINV,
      O => romo2datao5_s_10_F6MUX
    );
  romo2datao5_s_10_BYINV_5210 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_10_BYINV
    );
  nx53675z1125_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1125_F5MUX,
      O => nx53675z1125
    );
  nx53675z1125_F5MUX_5211 : X_MUX2
    port map (
      IA => nx53675z1126,
      IB => nx53675z1127,
      SEL => nx53675z1125_BXINV,
      O => nx53675z1125_F5MUX
    );
  nx53675z1125_BXINV_5212 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1125_BXINV
    );
  U_DCT2D_ix53540z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_0_4_Q,
      ADR1 => U_DCT2D_latchbuf_reg_7_4_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx53540z1
    );
  romo2datao5_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_9_F5MUX,
      O => nx53675z1134
    );
  romo2datao5_s_9_F5MUX_5213 : X_MUX2
    port map (
      IA => nx53675z1135,
      IB => nx53675z1136,
      SEL => romo2datao5_s_9_BXINV,
      O => romo2datao5_s_9_F5MUX
    );
  romo2datao5_s_9_BXINV_5214 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_9_BXINV
    );
  romo2datao5_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_9_F6MUX,
      O => romo2datao5_s(9)
    );
  romo2datao5_s_9_F6MUX_5215 : X_MUX2
    port map (
      IA => nx53675z1131,
      IB => nx53675z1134,
      SEL => romo2datao5_s_9_BYINV,
      O => romo2datao5_s_9_F6MUX
    );
  romo2datao5_s_9_BYINV_5216 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_9_BYINV
    );
  nx53675z1131_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1131_F5MUX,
      O => nx53675z1131
    );
  nx53675z1131_F5MUX_5217 : X_MUX2
    port map (
      IA => nx53675z1132,
      IB => nx53675z1133,
      SEL => nx53675z1131_BXINV,
      O => nx53675z1131_F5MUX
    );
  nx53675z1131_BXINV_5218 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1131_BXINV
    );
  romo2datao5_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_8_F5MUX,
      O => nx53675z1140
    );
  romo2datao5_s_8_F5MUX_5219 : X_MUX2
    port map (
      IA => nx53675z1141,
      IB => nx53675z1142,
      SEL => romo2datao5_s_8_BXINV,
      O => romo2datao5_s_8_F5MUX
    );
  romo2datao5_s_8_BXINV_5220 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_8_BXINV
    );
  romo2datao5_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_8_F6MUX,
      O => romo2datao5_s(8)
    );
  romo2datao5_s_8_F6MUX_5221 : X_MUX2
    port map (
      IA => nx53675z1137,
      IB => nx53675z1140,
      SEL => romo2datao5_s_8_BYINV,
      O => romo2datao5_s_8_F6MUX
    );
  romo2datao5_s_8_BYINV_5222 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_8_BYINV
    );
  nx53675z1137_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1137_F5MUX,
      O => nx53675z1137
    );
  nx53675z1137_F5MUX_5223 : X_MUX2
    port map (
      IA => nx53675z1138,
      IB => nx53675z1139,
      SEL => nx53675z1137_BXINV,
      O => nx53675z1137_F5MUX
    );
  nx53675z1137_BXINV_5224 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1137_BXINV
    );
  romo2datao5_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_2_F5MUX,
      O => nx53675z1176
    );
  romo2datao5_s_2_F5MUX_5225 : X_MUX2
    port map (
      IA => nx53675z1177,
      IB => nx53675z1178,
      SEL => romo2datao5_s_2_BXINV,
      O => romo2datao5_s_2_F5MUX
    );
  romo2datao5_s_2_BXINV_5226 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_2_BXINV
    );
  romo2datao5_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_2_F6MUX,
      O => romo2datao5_s(2)
    );
  romo2datao5_s_2_F6MUX_5227 : X_MUX2
    port map (
      IA => nx53675z1173,
      IB => nx53675z1176,
      SEL => romo2datao5_s_2_BYINV,
      O => romo2datao5_s_2_F6MUX
    );
  romo2datao5_s_2_BYINV_5228 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_2_BYINV
    );
  nx53675z1173_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1173_F5MUX,
      O => nx53675z1173
    );
  nx53675z1173_F5MUX_5229 : X_MUX2
    port map (
      IA => nx53675z1174,
      IB => nx53675z1175,
      SEL => nx53675z1173_BXINV,
      O => nx53675z1173_F5MUX
    );
  nx53675z1173_BXINV_5230 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1173_BXINV
    );
  romo2datao5_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_1_F5MUX,
      O => nx53675z1182
    );
  romo2datao5_s_1_F5MUX_5231 : X_MUX2
    port map (
      IA => nx53675z1183,
      IB => nx53675z1184,
      SEL => romo2datao5_s_1_BXINV,
      O => romo2datao5_s_1_F5MUX
    );
  romo2datao5_s_1_BXINV_5232 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_1_BXINV
    );
  romo2datao5_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_1_F6MUX,
      O => romo2datao5_s(1)
    );
  romo2datao5_s_1_F6MUX_5233 : X_MUX2
    port map (
      IA => nx53675z1179,
      IB => nx53675z1182,
      SEL => romo2datao5_s_1_BYINV,
      O => romo2datao5_s_1_F6MUX
    );
  romo2datao5_s_1_BYINV_5234 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_1_BYINV
    );
  nx53675z1179_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1179_F5MUX,
      O => nx53675z1179
    );
  nx53675z1179_F5MUX_5235 : X_MUX2
    port map (
      IA => nx53675z1180,
      IB => nx53675z1181,
      SEL => nx53675z1179_BXINV,
      O => nx53675z1179_F5MUX
    );
  nx53675z1179_BXINV_5236 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1179_BXINV
    );
  romo2datao5_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_0_F5MUX,
      O => U2_ROMO5_modgen_rom_ix0_nx_ro64_32_l
    );
  romo2datao5_s_0_F5MUX_5237 : X_MUX2
    port map (
      IA => nx53675z1185,
      IB => nx53675z1186,
      SEL => romo2datao5_s_0_BXINV,
      O => romo2datao5_s_0_F5MUX
    );
  romo2datao5_s_0_BXINV_5238 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_0_BXINV
    );
  romo2datao5_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_0_F6MUX,
      O => romo2datao5_s(0)
    );
  romo2datao5_s_0_F6MUX_5239 : X_MUX2
    port map (
      IA => U2_ROMO5_modgen_rom_ix0_nx_ro64_32_u,
      IB => U2_ROMO5_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romo2datao5_s_0_BYINV,
      O => romo2datao5_s_0_F6MUX
    );
  romo2datao5_s_0_BYINV_5240 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_0_BYINV
    );
  U2_ROMO5_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROMO5_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U2_ROMO5_modgen_rom_ix0_nx_ro64_32_u
    );
  U2_ROMO5_modgen_rom_ix0_nx_ro64_32_u_F5MUX_5241 : X_MUX2
    port map (
      IA => U2_ROMO5_modgen_rom_ix0_nx_rm64_16_u,
      IB => U2_ROMO5_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U2_ROMO5_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U2_ROMO5_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U2_ROMO5_modgen_rom_ix0_nx_ro64_32_u_BXINV_5242 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => U2_ROMO5_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romo2datao3_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_11_F5MUX,
      O => nx53675z964
    );
  romo2datao3_s_11_F5MUX_5243 : X_MUX2
    port map (
      IA => nx53675z965,
      IB => nx53675z966,
      SEL => romo2datao3_s_11_BXINV,
      O => romo2datao3_s_11_F5MUX
    );
  romo2datao3_s_11_BXINV_5244 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_11_BXINV
    );
  romo2datao3_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_11_F6MUX,
      O => romo2datao3_s(11)
    );
  romo2datao3_s_11_F6MUX_5245 : X_MUX2
    port map (
      IA => nx53675z961,
      IB => nx53675z964,
      SEL => romo2datao3_s_11_BYINV,
      O => romo2datao3_s_11_F6MUX
    );
  romo2datao3_s_11_BYINV_5246 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_11_BYINV
    );
  nx53675z961_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z961_F5MUX,
      O => nx53675z961
    );
  nx53675z961_F5MUX_5247 : X_MUX2
    port map (
      IA => nx53675z962,
      IB => nx53675z963,
      SEL => nx53675z961_BXINV,
      O => nx53675z961_F5MUX
    );
  nx53675z961_BXINV_5248 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z961_BXINV
    );
  romo2datao2_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_3_F5MUX,
      O => nx53675z933
    );
  romo2datao2_s_3_F5MUX_5249 : X_MUX2
    port map (
      IA => nx53675z934,
      IB => nx53675z935,
      SEL => romo2datao2_s_3_BXINV,
      O => romo2datao2_s_3_F5MUX
    );
  romo2datao2_s_3_BXINV_5250 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao2_s_3_BXINV
    );
  romo2datao2_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao2_s_3_F6MUX,
      O => romo2datao2_s(3)
    );
  romo2datao2_s_3_F6MUX_5251 : X_MUX2
    port map (
      IA => nx53675z930,
      IB => nx53675z933,
      SEL => romo2datao2_s_3_BYINV,
      O => romo2datao2_s_3_F6MUX
    );
  romo2datao2_s_3_BYINV_5252 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao2_s_3_BYINV
    );
  nx53675z930_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z930_F5MUX,
      O => nx53675z930
    );
  nx53675z930_F5MUX_5253 : X_MUX2
    port map (
      IA => nx53675z931,
      IB => nx53675z932,
      SEL => nx53675z930_BXINV,
      O => nx53675z930_F5MUX
    );
  nx53675z930_BXINV_5254 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z930_BXINV
    );
  rome2datao8_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_8_F5MUX,
      O => nx53675z552
    );
  rome2datao8_s_8_F5MUX_5255 : X_MUX2
    port map (
      IA => nx53675z553,
      IB => nx53675z554,
      SEL => rome2datao8_s_8_BXINV,
      O => rome2datao8_s_8_F5MUX
    );
  rome2datao8_s_8_BXINV_5256 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao8_s_8_BXINV
    );
  rome2datao8_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_8_F6MUX,
      O => rome2datao8_s(8)
    );
  rome2datao8_s_8_F6MUX_5257 : X_MUX2
    port map (
      IA => nx53675z549,
      IB => nx53675z552,
      SEL => rome2datao8_s_8_BYINV,
      O => rome2datao8_s_8_F6MUX
    );
  rome2datao8_s_8_BYINV_5258 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao8_s_8_BYINV
    );
  nx53675z549_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z549_F5MUX,
      O => nx53675z549
    );
  nx53675z549_F5MUX_5259 : X_MUX2
    port map (
      IA => nx53675z550,
      IB => nx53675z551,
      SEL => nx53675z549_BXINV,
      O => nx53675z549_F5MUX
    );
  nx53675z549_BXINV_5260 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z549_BXINV
    );
  rome2datao8_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_7_F5MUX,
      O => nx53675z558
    );
  rome2datao8_s_7_F5MUX_5261 : X_MUX2
    port map (
      IA => nx53675z559,
      IB => nx53675z560,
      SEL => rome2datao8_s_7_BXINV,
      O => rome2datao8_s_7_F5MUX
    );
  rome2datao8_s_7_BXINV_5262 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao8_s_7_BXINV
    );
  rome2datao8_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_7_F6MUX,
      O => rome2datao8_s(7)
    );
  rome2datao8_s_7_F6MUX_5263 : X_MUX2
    port map (
      IA => nx53675z555,
      IB => nx53675z558,
      SEL => rome2datao8_s_7_BYINV,
      O => rome2datao8_s_7_F6MUX
    );
  rome2datao8_s_7_BYINV_5264 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao8_s_7_BYINV
    );
  nx53675z555_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z555_F5MUX,
      O => nx53675z555
    );
  nx53675z555_F5MUX_5265 : X_MUX2
    port map (
      IA => nx53675z556,
      IB => nx53675z557,
      SEL => nx53675z555_BXINV,
      O => nx53675z555_F5MUX
    );
  nx53675z555_BXINV_5266 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z555_BXINV
    );
  rome2datao8_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_6_F5MUX,
      O => nx53675z564
    );
  rome2datao8_s_6_F5MUX_5267 : X_MUX2
    port map (
      IA => nx53675z565,
      IB => nx53675z566,
      SEL => rome2datao8_s_6_BXINV,
      O => rome2datao8_s_6_F5MUX
    );
  rome2datao8_s_6_BXINV_5268 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao8_s_6_BXINV
    );
  rome2datao8_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_6_F6MUX,
      O => rome2datao8_s(6)
    );
  rome2datao8_s_6_F6MUX_5269 : X_MUX2
    port map (
      IA => nx53675z561,
      IB => nx53675z564,
      SEL => rome2datao8_s_6_BYINV,
      O => rome2datao8_s_6_F6MUX
    );
  rome2datao8_s_6_BYINV_5270 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao8_s_6_BYINV
    );
  nx53675z561_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z561_F5MUX,
      O => nx53675z561
    );
  nx53675z561_F5MUX_5271 : X_MUX2
    port map (
      IA => nx53675z562,
      IB => nx53675z563,
      SEL => nx53675z561_BXINV,
      O => nx53675z561_F5MUX
    );
  nx53675z561_BXINV_5272 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z561_BXINV
    );
  U_DCT2D_reg_databuf_reg_4_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_4_4_DXMUX,
      CE => U_DCT2D_databuf_reg_4_4_CEINV,
      CLK => U_DCT2D_databuf_reg_4_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_4_4_FFX_RST,
      O => U_DCT2D_databuf_reg_4_Q(4)
    );
  U_DCT2D_databuf_reg_4_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_4_4_FFX_RST
    );
  rome2datao8_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_5_F5MUX,
      O => nx53675z570
    );
  rome2datao8_s_5_F5MUX_5273 : X_MUX2
    port map (
      IA => nx53675z571,
      IB => nx53675z572,
      SEL => rome2datao8_s_5_BXINV,
      O => rome2datao8_s_5_F5MUX
    );
  rome2datao8_s_5_BXINV_5274 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao8_s_5_BXINV
    );
  rome2datao8_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_5_F6MUX,
      O => rome2datao8_s(5)
    );
  rome2datao8_s_5_F6MUX_5275 : X_MUX2
    port map (
      IA => nx53675z567,
      IB => nx53675z570,
      SEL => rome2datao8_s_5_BYINV,
      O => rome2datao8_s_5_F6MUX
    );
  rome2datao8_s_5_BYINV_5276 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao8_s_5_BYINV
    );
  nx53675z567_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z567_F5MUX,
      O => nx53675z567
    );
  nx53675z567_F5MUX_5277 : X_MUX2
    port map (
      IA => nx53675z568,
      IB => nx53675z569,
      SEL => nx53675z567_BXINV,
      O => nx53675z567_F5MUX
    );
  nx53675z567_BXINV_5278 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z567_BXINV
    );
  rome2datao8_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_4_F5MUX,
      O => nx53675z576
    );
  rome2datao8_s_4_F5MUX_5279 : X_MUX2
    port map (
      IA => nx53675z577,
      IB => nx53675z578,
      SEL => rome2datao8_s_4_BXINV,
      O => rome2datao8_s_4_F5MUX
    );
  rome2datao8_s_4_BXINV_5280 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao8_s_4_BXINV
    );
  rome2datao8_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_4_F6MUX,
      O => rome2datao8_s(4)
    );
  rome2datao8_s_4_F6MUX_5281 : X_MUX2
    port map (
      IA => nx53675z573,
      IB => nx53675z576,
      SEL => rome2datao8_s_4_BYINV,
      O => rome2datao8_s_4_F6MUX
    );
  rome2datao8_s_4_BYINV_5282 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao8_s_4_BYINV
    );
  U_DCT2D_ix56531z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_0_7_Q,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_7_7_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx56531z1
    );
  nx53675z573_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z573_F5MUX,
      O => nx53675z573
    );
  nx53675z573_F5MUX_5283 : X_MUX2
    port map (
      IA => nx53675z574,
      IB => nx53675z575,
      SEL => nx53675z573_BXINV,
      O => nx53675z573_F5MUX
    );
  nx53675z573_BXINV_5284 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z573_BXINV
    );
  rome2datao7_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_5_F5MUX,
      O => nx53675z505
    );
  rome2datao7_s_5_F5MUX_5285 : X_MUX2
    port map (
      IA => nx53675z506,
      IB => nx53675z507,
      SEL => rome2datao7_s_5_BXINV,
      O => rome2datao7_s_5_F5MUX
    );
  rome2datao7_s_5_BXINV_5286 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao7_s_5_BXINV
    );
  rome2datao7_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_5_F6MUX,
      O => rome2datao7_s(5)
    );
  rome2datao7_s_5_F6MUX_5287 : X_MUX2
    port map (
      IA => nx53675z502,
      IB => nx53675z505,
      SEL => rome2datao7_s_5_BYINV,
      O => rome2datao7_s_5_F6MUX
    );
  rome2datao7_s_5_BYINV_5288 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao7_s_5_BYINV
    );
  nx53675z502_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z502_F5MUX,
      O => nx53675z502
    );
  nx53675z502_F5MUX_5289 : X_MUX2
    port map (
      IA => nx53675z503,
      IB => nx53675z504,
      SEL => nx53675z502_BXINV,
      O => nx53675z502_F5MUX
    );
  nx53675z502_BXINV_5290 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z502_BXINV
    );
  rome2datao7_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_4_F5MUX,
      O => nx53675z511
    );
  rome2datao7_s_4_F5MUX_5291 : X_MUX2
    port map (
      IA => nx53675z512,
      IB => nx53675z513,
      SEL => rome2datao7_s_4_BXINV,
      O => rome2datao7_s_4_F5MUX
    );
  rome2datao7_s_4_BXINV_5292 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao7_s_4_BXINV
    );
  rome2datao7_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao7_s_4_F6MUX,
      O => rome2datao7_s(4)
    );
  rome2datao7_s_4_F6MUX_5293 : X_MUX2
    port map (
      IA => nx53675z508,
      IB => nx53675z511,
      SEL => rome2datao7_s_4_BYINV,
      O => rome2datao7_s_4_F6MUX
    );
  rome2datao7_s_4_BYINV_5294 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao7_s_4_BYINV
    );
  nx53675z508_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z508_F5MUX,
      O => nx53675z508
    );
  nx53675z508_F5MUX_5295 : X_MUX2
    port map (
      IA => nx53675z509,
      IB => nx53675z510,
      SEL => nx53675z508_BXINV,
      O => nx53675z508_F5MUX
    );
  nx53675z508_BXINV_5296 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z508_BXINV
    );
  romo2datao6_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_12_F5MUX,
      O => nx53675z1195
    );
  romo2datao6_s_12_F5MUX_5297 : X_MUX2
    port map (
      IA => nx53675z1196,
      IB => nx53675z1197,
      SEL => romo2datao6_s_12_BXINV,
      O => romo2datao6_s_12_F5MUX
    );
  romo2datao6_s_12_BXINV_5298 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_12_BXINV
    );
  romo2datao6_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_12_F6MUX,
      O => romo2datao6_s(12)
    );
  romo2datao6_s_12_F6MUX_5299 : X_MUX2
    port map (
      IA => nx53675z1192,
      IB => nx53675z1195,
      SEL => romo2datao6_s_12_BYINV,
      O => romo2datao6_s_12_F6MUX
    );
  romo2datao6_s_12_BYINV_5300 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_12_BYINV
    );
  nx53675z1192_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1192_F5MUX,
      O => nx53675z1192
    );
  nx53675z1192_F5MUX_5301 : X_MUX2
    port map (
      IA => nx53675z1193,
      IB => nx53675z1194,
      SEL => nx53675z1192_BXINV,
      O => nx53675z1192_F5MUX
    );
  nx53675z1192_BXINV_5302 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1192_BXINV
    );
  romo2datao7_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_12_F5MUX,
      O => nx53675z1274
    );
  romo2datao7_s_12_F5MUX_5303 : X_MUX2
    port map (
      IA => nx53675z1275,
      IB => nx53675z1276,
      SEL => romo2datao7_s_12_BXINV,
      O => romo2datao7_s_12_F5MUX
    );
  romo2datao7_s_12_BXINV_5304 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_12_BXINV
    );
  romo2datao7_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_12_F6MUX,
      O => romo2datao7_s(12)
    );
  romo2datao7_s_12_F6MUX_5305 : X_MUX2
    port map (
      IA => nx53675z1271,
      IB => nx53675z1274,
      SEL => romo2datao7_s_12_BYINV,
      O => romo2datao7_s_12_F6MUX
    );
  romo2datao7_s_12_BYINV_5306 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_12_BYINV
    );
  nx53675z1271_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1271_F5MUX,
      O => nx53675z1271
    );
  nx53675z1271_F5MUX_5307 : X_MUX2
    port map (
      IA => nx53675z1272,
      IB => nx53675z1273,
      SEL => nx53675z1271_BXINV,
      O => nx53675z1271_F5MUX
    );
  nx53675z1271_BXINV_5308 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1271_BXINV
    );
  romo2datao7_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_11_F5MUX,
      O => nx53675z1280
    );
  romo2datao7_s_11_F5MUX_5309 : X_MUX2
    port map (
      IA => nx53675z1281,
      IB => nx53675z1282,
      SEL => romo2datao7_s_11_BXINV,
      O => romo2datao7_s_11_F5MUX
    );
  romo2datao7_s_11_BXINV_5310 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_11_BXINV
    );
  romo2datao7_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_11_F6MUX,
      O => romo2datao7_s(11)
    );
  romo2datao7_s_11_F6MUX_5311 : X_MUX2
    port map (
      IA => nx53675z1277,
      IB => nx53675z1280,
      SEL => romo2datao7_s_11_BYINV,
      O => romo2datao7_s_11_F6MUX
    );
  romo2datao7_s_11_BYINV_5312 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_11_BYINV
    );
  nx53675z1277_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1277_F5MUX,
      O => nx53675z1277
    );
  nx53675z1277_F5MUX_5313 : X_MUX2
    port map (
      IA => nx53675z1278,
      IB => nx53675z1279,
      SEL => nx53675z1277_BXINV,
      O => nx53675z1277_F5MUX
    );
  nx53675z1277_BXINV_5314 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1277_BXINV
    );
  romo2datao6_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_11_F5MUX,
      O => nx53675z1201
    );
  romo2datao6_s_11_F5MUX_5315 : X_MUX2
    port map (
      IA => nx53675z1202,
      IB => nx53675z1203,
      SEL => romo2datao6_s_11_BXINV,
      O => romo2datao6_s_11_F5MUX
    );
  romo2datao6_s_11_BXINV_5316 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_11_BXINV
    );
  romo2datao6_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_11_F6MUX,
      O => romo2datao6_s(11)
    );
  romo2datao6_s_11_F6MUX_5317 : X_MUX2
    port map (
      IA => nx53675z1198,
      IB => nx53675z1201,
      SEL => romo2datao6_s_11_BYINV,
      O => romo2datao6_s_11_F6MUX
    );
  romo2datao6_s_11_BYINV_5318 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_11_BYINV
    );
  nx53675z1198_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1198_F5MUX,
      O => nx53675z1198
    );
  nx53675z1198_F5MUX_5319 : X_MUX2
    port map (
      IA => nx53675z1199,
      IB => nx53675z1200,
      SEL => nx53675z1198_BXINV,
      O => nx53675z1198_F5MUX
    );
  nx53675z1198_BXINV_5320 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1198_BXINV
    );
  romo2datao6_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_10_F5MUX,
      O => nx53675z1207
    );
  romo2datao6_s_10_F5MUX_5321 : X_MUX2
    port map (
      IA => nx53675z1208,
      IB => nx53675z1209,
      SEL => romo2datao6_s_10_BXINV,
      O => romo2datao6_s_10_F5MUX
    );
  romo2datao6_s_10_BXINV_5322 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_10_BXINV
    );
  romo2datao6_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_10_F6MUX,
      O => romo2datao6_s(10)
    );
  romo2datao6_s_10_F6MUX_5323 : X_MUX2
    port map (
      IA => nx53675z1204,
      IB => nx53675z1207,
      SEL => romo2datao6_s_10_BYINV,
      O => romo2datao6_s_10_F6MUX
    );
  romo2datao6_s_10_BYINV_5324 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_10_BYINV
    );
  nx53675z1204_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1204_F5MUX,
      O => nx53675z1204
    );
  nx53675z1204_F5MUX_5325 : X_MUX2
    port map (
      IA => nx53675z1205,
      IB => nx53675z1206,
      SEL => nx53675z1204_BXINV,
      O => nx53675z1204_F5MUX
    );
  nx53675z1204_BXINV_5326 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1204_BXINV
    );
  romo2datao6_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_9_F5MUX,
      O => nx53675z1213
    );
  romo2datao6_s_9_F5MUX_5327 : X_MUX2
    port map (
      IA => nx53675z1214,
      IB => nx53675z1215,
      SEL => romo2datao6_s_9_BXINV,
      O => romo2datao6_s_9_F5MUX
    );
  romo2datao6_s_9_BXINV_5328 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_9_BXINV
    );
  romo2datao6_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_9_F6MUX,
      O => romo2datao6_s(9)
    );
  romo2datao6_s_9_F6MUX_5329 : X_MUX2
    port map (
      IA => nx53675z1210,
      IB => nx53675z1213,
      SEL => romo2datao6_s_9_BYINV,
      O => romo2datao6_s_9_F6MUX
    );
  romo2datao6_s_9_BYINV_5330 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_9_BYINV
    );
  nx53675z1210_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1210_F5MUX,
      O => nx53675z1210
    );
  nx53675z1210_F5MUX_5331 : X_MUX2
    port map (
      IA => nx53675z1211,
      IB => nx53675z1212,
      SEL => nx53675z1210_BXINV,
      O => nx53675z1210_F5MUX
    );
  nx53675z1210_BXINV_5332 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1210_BXINV
    );
  romo2datao6_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_1_F5MUX,
      O => nx53675z1261
    );
  romo2datao6_s_1_F5MUX_5333 : X_MUX2
    port map (
      IA => nx53675z1262,
      IB => nx53675z1263,
      SEL => romo2datao6_s_1_BXINV,
      O => romo2datao6_s_1_F5MUX
    );
  romo2datao6_s_1_BXINV_5334 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_1_BXINV
    );
  romo2datao6_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_1_F6MUX,
      O => romo2datao6_s(1)
    );
  romo2datao6_s_1_F6MUX_5335 : X_MUX2
    port map (
      IA => nx53675z1258,
      IB => nx53675z1261,
      SEL => romo2datao6_s_1_BYINV,
      O => romo2datao6_s_1_F6MUX
    );
  romo2datao6_s_1_BYINV_5336 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_1_BYINV
    );
  nx53675z1258_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1258_F5MUX,
      O => nx53675z1258
    );
  nx53675z1258_F5MUX_5337 : X_MUX2
    port map (
      IA => nx53675z1259,
      IB => nx53675z1260,
      SEL => nx53675z1258_BXINV,
      O => nx53675z1258_F5MUX
    );
  nx53675z1258_BXINV_5338 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1258_BXINV
    );
  romo2datao5_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_7_F5MUX,
      O => nx53675z1146
    );
  romo2datao5_s_7_F5MUX_5339 : X_MUX2
    port map (
      IA => nx53675z1147,
      IB => nx53675z1148,
      SEL => romo2datao5_s_7_BXINV,
      O => romo2datao5_s_7_F5MUX
    );
  romo2datao5_s_7_BXINV_5340 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao5_s_7_BXINV
    );
  romo2datao5_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao5_s_7_F6MUX,
      O => romo2datao5_s(7)
    );
  romo2datao5_s_7_F6MUX_5341 : X_MUX2
    port map (
      IA => nx53675z1143,
      IB => nx53675z1146,
      SEL => romo2datao5_s_7_BYINV,
      O => romo2datao5_s_7_F6MUX
    );
  romo2datao5_s_7_BYINV_5342 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao5_s_7_BYINV
    );
  nx53675z1143_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1143_F5MUX,
      O => nx53675z1143
    );
  nx53675z1143_F5MUX_5343 : X_MUX2
    port map (
      IA => nx53675z1144,
      IB => nx53675z1145,
      SEL => nx53675z1143_BXINV,
      O => nx53675z1143_F5MUX
    );
  nx53675z1143_BXINV_5344 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1143_BXINV
    );
  romo2datao3_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_9_F5MUX,
      O => nx53675z976
    );
  romo2datao3_s_9_F5MUX_5345 : X_MUX2
    port map (
      IA => nx53675z977,
      IB => nx53675z978,
      SEL => romo2datao3_s_9_BXINV,
      O => romo2datao3_s_9_F5MUX
    );
  romo2datao3_s_9_BXINV_5346 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_9_BXINV
    );
  romo2datao3_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_9_F6MUX,
      O => romo2datao3_s(9)
    );
  romo2datao3_s_9_F6MUX_5347 : X_MUX2
    port map (
      IA => nx53675z973,
      IB => nx53675z976,
      SEL => romo2datao3_s_9_BYINV,
      O => romo2datao3_s_9_F6MUX
    );
  romo2datao3_s_9_BYINV_5348 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_9_BYINV
    );
  nx53675z973_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z973_F5MUX,
      O => nx53675z973
    );
  nx53675z973_F5MUX_5349 : X_MUX2
    port map (
      IA => nx53675z974,
      IB => nx53675z975,
      SEL => nx53675z973_BXINV,
      O => nx53675z973_F5MUX
    );
  nx53675z973_BXINV_5350 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z973_BXINV
    );
  rome2datao8_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_3_F5MUX,
      O => nx53675z581
    );
  rome2datao8_s_3_F5MUX_5351 : X_MUX2
    port map (
      IA => nx53675z582,
      IB => nx53675z583,
      SEL => rome2datao8_s_3_BXINV,
      O => rome2datao8_s_3_F5MUX
    );
  rome2datao8_s_3_BXINV_5352 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => rome2datao8_s_3_BXINV
    );
  rome2datao8_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2datao8_s_3_F6MUX,
      O => rome2datao8_s(3)
    );
  rome2datao8_s_3_F6MUX_5353 : X_MUX2
    port map (
      IA => nx53675z579,
      IB => nx53675z581,
      SEL => rome2datao8_s_3_BYINV,
      O => rome2datao8_s_3_F6MUX
    );
  rome2datao8_s_3_BYINV_5354 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(5),
      O => rome2datao8_s_3_BYINV
    );
  nx53675z579_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z579_F5MUX,
      O => nx53675z579
    );
  nx53675z579_F5MUX_5355 : X_MUX2
    port map (
      IA => U2_ROME8_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx53675z580,
      SEL => nx53675z579_BXINV,
      O => nx53675z579_F5MUX
    );
  nx53675z579_BXINV_5356 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rome2addro0_s(4),
      O => nx53675z579_BXINV
    );
  romo2datao6_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_0_F5MUX,
      O => U2_ROMO6_modgen_rom_ix0_nx_ro64_32_l
    );
  romo2datao6_s_0_F5MUX_5357 : X_MUX2
    port map (
      IA => nx53675z1264,
      IB => nx53675z1265,
      SEL => romo2datao6_s_0_BXINV,
      O => romo2datao6_s_0_F5MUX
    );
  romo2datao6_s_0_BXINV_5358 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao6_s_0_BXINV
    );
  romo2datao6_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao6_s_0_F6MUX,
      O => romo2datao6_s(0)
    );
  romo2datao6_s_0_F6MUX_5359 : X_MUX2
    port map (
      IA => U2_ROMO6_modgen_rom_ix0_nx_ro64_32_u,
      IB => U2_ROMO6_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romo2datao6_s_0_BYINV,
      O => romo2datao6_s_0_F6MUX
    );
  romo2datao6_s_0_BYINV_5360 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao6_s_0_BYINV
    );
  U2_ROMO6_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U2_ROMO6_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U2_ROMO6_modgen_rom_ix0_nx_ro64_32_u
    );
  U2_ROMO6_modgen_rom_ix0_nx_ro64_32_u_F5MUX_5361 : X_MUX2
    port map (
      IA => U2_ROMO6_modgen_rom_ix0_nx_rm64_16_u,
      IB => U2_ROMO6_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U2_ROMO6_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U2_ROMO6_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U2_ROMO6_modgen_rom_ix0_nx_ro64_32_u_BXINV_5362 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => U2_ROMO6_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romo2datao10_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_11_F5MUX,
      O => nx53675z1517
    );
  romo2datao10_s_11_F5MUX_5363 : X_MUX2
    port map (
      IA => nx53675z1518,
      IB => nx53675z1519,
      SEL => romo2datao10_s_11_BXINV,
      O => romo2datao10_s_11_F5MUX
    );
  romo2datao10_s_11_BXINV_5364 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao10_s_11_BXINV
    );
  romo2datao10_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao10_s_11_F6MUX,
      O => romo2datao10_s(11)
    );
  romo2datao10_s_11_F6MUX_5365 : X_MUX2
    port map (
      IA => nx53675z1514,
      IB => nx53675z1517,
      SEL => romo2datao10_s_11_BYINV,
      O => romo2datao10_s_11_F6MUX
    );
  romo2datao10_s_11_BYINV_5366 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao10_s_11_BYINV
    );
  nx53675z1514_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1514_F5MUX,
      O => nx53675z1514
    );
  nx53675z1514_F5MUX_5367 : X_MUX2
    port map (
      IA => nx53675z1515,
      IB => nx53675z1516,
      SEL => nx53675z1514_BXINV,
      O => nx53675z1514_F5MUX
    );
  nx53675z1514_BXINV_5368 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1514_BXINV
    );
  romo2datao7_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_13_F5MUX,
      O => nx53675z1268
    );
  romo2datao7_s_13_F5MUX_5369 : X_MUX2
    port map (
      IA => nx53675z1269,
      IB => nx53675z1270,
      SEL => romo2datao7_s_13_BXINV,
      O => romo2datao7_s_13_F5MUX
    );
  romo2datao7_s_13_BXINV_5370 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_13_BXINV
    );
  romo2datao7_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_13_F6MUX,
      O => romo2datao7_s(13)
    );
  romo2datao7_s_13_F6MUX_5371 : X_MUX2
    port map (
      IA => nx53675z1266,
      IB => nx53675z1268,
      SEL => romo2datao7_s_13_BYINV,
      O => romo2datao7_s_13_F6MUX
    );
  romo2datao7_s_13_BYINV_5372 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_13_BYINV
    );
  nx53675z1266_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1266_F5MUX,
      O => nx53675z1266
    );
  nx53675z1266_F5MUX_5373 : X_MUX2
    port map (
      IA => nx53675z1266_G,
      IB => nx53675z1267,
      SEL => nx53675z1266_BXINV,
      O => nx53675z1266_F5MUX
    );
  nx53675z1266_BXINV_5374 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1266_BXINV
    );
  romo2datao7_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_10_F5MUX,
      O => nx53675z1286
    );
  romo2datao7_s_10_F5MUX_5375 : X_MUX2
    port map (
      IA => nx53675z1287,
      IB => nx53675z1288,
      SEL => romo2datao7_s_10_BXINV,
      O => romo2datao7_s_10_F5MUX
    );
  romo2datao7_s_10_BXINV_5376 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao7_s_10_BXINV
    );
  romo2datao7_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao7_s_10_F6MUX,
      O => romo2datao7_s(10)
    );
  romo2datao7_s_10_F6MUX_5377 : X_MUX2
    port map (
      IA => nx53675z1283,
      IB => nx53675z1286,
      SEL => romo2datao7_s_10_BYINV,
      O => romo2datao7_s_10_F6MUX
    );
  romo2datao7_s_10_BYINV_5378 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao7_s_10_BYINV
    );
  nx53675z1283_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z1283_F5MUX,
      O => nx53675z1283
    );
  nx53675z1283_F5MUX_5379 : X_MUX2
    port map (
      IA => nx53675z1284,
      IB => nx53675z1285,
      SEL => nx53675z1283_BXINV,
      O => nx53675z1283_F5MUX
    );
  nx53675z1283_BXINV_5380 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z1283_BXINV
    );
  romo2datao3_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_7_F5MUX,
      O => nx53675z988
    );
  romo2datao3_s_7_F5MUX_5381 : X_MUX2
    port map (
      IA => nx53675z989,
      IB => nx53675z990,
      SEL => romo2datao3_s_7_BXINV,
      O => romo2datao3_s_7_F5MUX
    );
  romo2datao3_s_7_BXINV_5382 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_7_BXINV
    );
  romo2datao3_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_7_F6MUX,
      O => romo2datao3_s(7)
    );
  romo2datao3_s_7_F6MUX_5383 : X_MUX2
    port map (
      IA => nx53675z985,
      IB => nx53675z988,
      SEL => romo2datao3_s_7_BYINV,
      O => romo2datao3_s_7_F6MUX
    );
  romo2datao3_s_7_BYINV_5384 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_7_BYINV
    );
  nx53675z985_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z985_F5MUX,
      O => nx53675z985
    );
  nx53675z985_F5MUX_5385 : X_MUX2
    port map (
      IA => nx53675z986,
      IB => nx53675z987,
      SEL => nx53675z985_BXINV,
      O => nx53675z985_F5MUX
    );
  nx53675z985_BXINV_5386 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z985_BXINV
    );
  U_DCT2D_reg_databuf_reg_4_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_4_6_DYMUX,
      CE => U_DCT2D_databuf_reg_4_6_CEINV,
      CLK => U_DCT2D_databuf_reg_4_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_4_6_FFY_RST,
      O => U_DCT2D_databuf_reg_4_Q(7)
    );
  U_DCT2D_databuf_reg_4_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_4_6_FFY_RST
    );
  romo2datao3_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_5_F5MUX,
      O => nx53675z1000
    );
  romo2datao3_s_5_F5MUX_5387 : X_MUX2
    port map (
      IA => nx53675z1001,
      IB => nx53675z1002,
      SEL => romo2datao3_s_5_BXINV,
      O => romo2datao3_s_5_F5MUX
    );
  romo2datao3_s_5_BXINV_5388 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => romo2datao3_s_5_BXINV
    );
  romo2datao3_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2datao3_s_5_F6MUX,
      O => romo2datao3_s(5)
    );
  romo2datao3_s_5_F6MUX_5389 : X_MUX2
    port map (
      IA => nx53675z997,
      IB => nx53675z1000,
      SEL => romo2datao3_s_5_BYINV,
      O => romo2datao3_s_5_F6MUX
    );
  romo2datao3_s_5_BYINV_5390 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(5),
      O => romo2datao3_s_5_BYINV
    );
  nx53675z997_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx53675z997_F5MUX,
      O => nx53675z997
    );
  nx53675z997_F5MUX_5391 : X_MUX2
    port map (
      IA => nx53675z998,
      IB => nx53675z999,
      SEL => nx53675z997_BXINV,
      O => nx53675z997_F5MUX
    );
  nx53675z997_BXINV_5392 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romo2addro0_s(4),
      O => nx53675z997_BXINV
    );
  romedatao0_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_10_F5MUX,
      O => nx54672z21
    );
  romedatao0_s_10_F5MUX_5393 : X_MUX2
    port map (
      IA => nx54672z22,
      IB => nx54672z23,
      SEL => romedatao0_s_10_BXINV,
      O => romedatao0_s_10_F5MUX
    );
  romedatao0_s_10_BXINV_5394 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao0_s_10_BXINV
    );
  romedatao0_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_10_F6MUX,
      O => romedatao0_s(10)
    );
  romedatao0_s_10_F6MUX_5395 : X_MUX2
    port map (
      IA => nx54672z18,
      IB => nx54672z21,
      SEL => romedatao0_s_10_BYINV,
      O => romedatao0_s_10_F6MUX
    );
  romedatao0_s_10_BYINV_5396 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao0_s_10_BYINV
    );
  ix54672z34386 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(0),
      ADR3 => romeaddro0_s(3),
      O => nx54672z19
    );
  nx54672z18_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z18_F5MUX,
      O => nx54672z18
    );
  nx54672z18_F5MUX_5397 : X_MUX2
    port map (
      IA => nx54672z19,
      IB => nx54672z20,
      SEL => nx54672z18_BXINV,
      O => nx54672z18_F5MUX
    );
  nx54672z18_BXINV_5398 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z18_BXINV
    );
  romedatao0_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_9_F5MUX,
      O => nx54672z27
    );
  romedatao0_s_9_F5MUX_5399 : X_MUX2
    port map (
      IA => nx54672z28,
      IB => nx54672z29,
      SEL => romedatao0_s_9_BXINV,
      O => romedatao0_s_9_F5MUX
    );
  romedatao0_s_9_BXINV_5400 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao0_s_9_BXINV
    );
  romedatao0_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_9_F6MUX,
      O => romedatao0_s(9)
    );
  romedatao0_s_9_F6MUX_5401 : X_MUX2
    port map (
      IA => nx54672z24,
      IB => nx54672z27,
      SEL => romedatao0_s_9_BYINV,
      O => romedatao0_s_9_F6MUX
    );
  romedatao0_s_9_BYINV_5402 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao0_s_9_BYINV
    );
  nx54672z24_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z24_F5MUX,
      O => nx54672z24
    );
  nx54672z24_F5MUX_5403 : X_MUX2
    port map (
      IA => nx54672z25,
      IB => nx54672z26,
      SEL => nx54672z24_BXINV,
      O => nx54672z24_F5MUX
    );
  nx54672z24_BXINV_5404 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z24_BXINV
    );
  romodatao0_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_13_F5MUX,
      O => nx54672z587
    );
  romodatao0_s_13_F5MUX_5405 : X_MUX2
    port map (
      IA => nx54672z588,
      IB => nx54672z589,
      SEL => romodatao0_s_13_BXINV,
      O => romodatao0_s_13_F5MUX
    );
  romodatao0_s_13_BXINV_5406 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_13_BXINV
    );
  romodatao0_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_13_F6MUX,
      O => romodatao0_s(13)
    );
  romodatao0_s_13_F6MUX_5407 : X_MUX2
    port map (
      IA => nx54672z585,
      IB => nx54672z587,
      SEL => romodatao0_s_13_BYINV,
      O => romodatao0_s_13_F6MUX
    );
  romodatao0_s_13_BYINV_5408 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_13_BYINV
    );
  nx54672z585_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z585_F5MUX,
      O => nx54672z585
    );
  nx54672z585_F5MUX_5409 : X_MUX2
    port map (
      IA => nx54672z585_G,
      IB => nx54672z586,
      SEL => nx54672z585_BXINV,
      O => nx54672z585_F5MUX
    );
  nx54672z585_BXINV_5410 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z585_BXINV
    );
  romedatao8_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_2_F5MUX,
      O => U1_ROME8_modgen_rom_ix2_nx_ro64_32_l
    );
  romedatao8_s_2_F5MUX_5411 : X_MUX2
    port map (
      IA => romedatao8_s_2_G,
      IB => nx54672z584,
      SEL => romedatao8_s_2_BXINV,
      O => romedatao8_s_2_F5MUX
    );
  romedatao8_s_2_BXINV_5412 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao8_s_2_BXINV
    );
  romedatao8_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_2_F6MUX,
      O => romedatao8_s(2)
    );
  romedatao8_s_2_F6MUX_5413 : X_MUX2
    port map (
      IA => U1_ROME8_modgen_rom_ix2_nx_ro64_32_u,
      IB => U1_ROME8_modgen_rom_ix2_nx_ro64_32_l,
      SEL => romedatao8_s_2_BYINV,
      O => romedatao8_s_2_F6MUX
    );
  romedatao8_s_2_BYINV_5414 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao8_s_2_BYINV
    );
  U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U1_ROME8_modgen_rom_ix2_nx_ro64_32_u
    );
  U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_F5MUX_5415 : X_MUX2
    port map (
      IA => U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U1_ROME8_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_BXINV_5416 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  U_DCT2D_ix55534z1324 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_0_6_Q,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_7_6_Q,
      O => U_DCT2D_nx55534z1
    );
  romedatao2_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_8_F5MUX,
      O => nx54672z162
    );
  romedatao2_s_8_F5MUX_5417 : X_MUX2
    port map (
      IA => nx54672z163,
      IB => nx54672z164,
      SEL => romedatao2_s_8_BXINV,
      O => romedatao2_s_8_F5MUX
    );
  romedatao2_s_8_BXINV_5418 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao2_s_8_BXINV
    );
  romedatao2_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_8_F6MUX,
      O => romedatao2_s(8)
    );
  romedatao2_s_8_F6MUX_5419 : X_MUX2
    port map (
      IA => nx54672z159,
      IB => nx54672z162,
      SEL => romedatao2_s_8_BYINV,
      O => romedatao2_s_8_F6MUX
    );
  romedatao2_s_8_BYINV_5420 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao2_s_8_BYINV
    );
  ix54672z7552 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(2),
      O => nx54672z160
    );
  nx54672z159_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z159_F5MUX,
      O => nx54672z159
    );
  nx54672z159_F5MUX_5421 : X_MUX2
    port map (
      IA => nx54672z160,
      IB => nx54672z161,
      SEL => nx54672z159_BXINV,
      O => nx54672z159_F5MUX
    );
  nx54672z159_BXINV_5422 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z159_BXINV
    );
  romodatao1_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_12_F5MUX,
      O => nx54672z670
    );
  romodatao1_s_12_F5MUX_5423 : X_MUX2
    port map (
      IA => nx54672z671,
      IB => nx54672z672,
      SEL => romodatao1_s_12_BXINV,
      O => romodatao1_s_12_F5MUX
    );
  romodatao1_s_12_BXINV_5424 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_12_BXINV
    );
  romodatao1_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_12_F6MUX,
      O => romodatao1_s(12)
    );
  romodatao1_s_12_F6MUX_5425 : X_MUX2
    port map (
      IA => nx54672z667,
      IB => nx54672z670,
      SEL => romodatao1_s_12_BYINV,
      O => romodatao1_s_12_F6MUX
    );
  romodatao1_s_12_BYINV_5426 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_12_BYINV
    );
  ix54672z59604 : X_LUT4
    generic map(
      INIT => X"8880"
    )
    port map (
      ADR0 => romoaddro1_s(2),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(1),
      O => nx54672z668
    );
  nx54672z667_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z667_F5MUX,
      O => nx54672z667
    );
  nx54672z667_F5MUX_5427 : X_MUX2
    port map (
      IA => nx54672z668,
      IB => nx54672z669,
      SEL => nx54672z667_BXINV,
      O => nx54672z667_F5MUX
    );
  nx54672z667_BXINV_5428 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z667_BXINV
    );
  romodatao1_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_11_F5MUX,
      O => nx54672z676
    );
  romodatao1_s_11_F5MUX_5429 : X_MUX2
    port map (
      IA => nx54672z677,
      IB => nx54672z678,
      SEL => romodatao1_s_11_BXINV,
      O => romodatao1_s_11_F5MUX
    );
  romodatao1_s_11_BXINV_5430 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_11_BXINV
    );
  romodatao1_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_11_F6MUX,
      O => romodatao1_s(11)
    );
  romodatao1_s_11_F6MUX_5431 : X_MUX2
    port map (
      IA => nx54672z673,
      IB => nx54672z676,
      SEL => romodatao1_s_11_BYINV,
      O => romodatao1_s_11_F6MUX
    );
  romodatao1_s_11_BYINV_5432 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_11_BYINV
    );
  nx54672z673_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z673_F5MUX,
      O => nx54672z673
    );
  nx54672z673_F5MUX_5433 : X_MUX2
    port map (
      IA => nx54672z674,
      IB => nx54672z675,
      SEL => nx54672z673_BXINV,
      O => nx54672z673_F5MUX
    );
  nx54672z673_BXINV_5434 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z673_BXINV
    );
  romodatao1_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_2_F5MUX,
      O => nx54672z730
    );
  romodatao1_s_2_F5MUX_5435 : X_MUX2
    port map (
      IA => nx54672z731,
      IB => nx54672z732,
      SEL => romodatao1_s_2_BXINV,
      O => romodatao1_s_2_F5MUX
    );
  romodatao1_s_2_BXINV_5436 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_2_BXINV
    );
  romodatao1_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_2_F6MUX,
      O => romodatao1_s(2)
    );
  romodatao1_s_2_F6MUX_5437 : X_MUX2
    port map (
      IA => nx54672z727,
      IB => nx54672z730,
      SEL => romodatao1_s_2_BYINV,
      O => romodatao1_s_2_F6MUX
    );
  romodatao1_s_2_BYINV_5438 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_2_BYINV
    );
  nx54672z727_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z727_F5MUX,
      O => nx54672z727
    );
  nx54672z727_F5MUX_5439 : X_MUX2
    port map (
      IA => nx54672z728,
      IB => nx54672z729,
      SEL => nx54672z727_BXINV,
      O => nx54672z727_F5MUX
    );
  nx54672z727_BXINV_5440 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z727_BXINV
    );
  romodatao1_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_1_F5MUX,
      O => nx54672z736
    );
  romodatao1_s_1_F5MUX_5441 : X_MUX2
    port map (
      IA => nx54672z737,
      IB => nx54672z738,
      SEL => romodatao1_s_1_BXINV,
      O => romodatao1_s_1_F5MUX
    );
  romodatao1_s_1_BXINV_5442 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_1_BXINV
    );
  romodatao1_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_1_F6MUX,
      O => romodatao1_s(1)
    );
  romodatao1_s_1_F6MUX_5443 : X_MUX2
    port map (
      IA => nx54672z733,
      IB => nx54672z736,
      SEL => romodatao1_s_1_BYINV,
      O => romodatao1_s_1_F6MUX
    );
  romodatao1_s_1_BYINV_5444 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_1_BYINV
    );
  nx54672z733_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z733_F5MUX,
      O => nx54672z733
    );
  nx54672z733_F5MUX_5445 : X_MUX2
    port map (
      IA => nx54672z734,
      IB => nx54672z735,
      SEL => nx54672z733_BXINV,
      O => nx54672z733_F5MUX
    );
  nx54672z733_BXINV_5446 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z733_BXINV
    );
  romedatao1_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_8_F5MUX,
      O => nx54672z97
    );
  romedatao1_s_8_F5MUX_5447 : X_MUX2
    port map (
      IA => nx54672z98,
      IB => nx54672z99,
      SEL => romedatao1_s_8_BXINV,
      O => romedatao1_s_8_F5MUX
    );
  romedatao1_s_8_BXINV_5448 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao1_s_8_BXINV
    );
  romedatao1_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_8_F6MUX,
      O => romedatao1_s(8)
    );
  romedatao1_s_8_F6MUX_5449 : X_MUX2
    port map (
      IA => nx54672z94,
      IB => nx54672z97,
      SEL => romedatao1_s_8_BYINV,
      O => romedatao1_s_8_F6MUX
    );
  romedatao1_s_8_BYINV_5450 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao1_s_8_BYINV
    );
  ix54672z7458 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z95
    );
  nx54672z94_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z94_F5MUX,
      O => nx54672z94
    );
  nx54672z94_F5MUX_5451 : X_MUX2
    port map (
      IA => nx54672z95,
      IB => nx54672z96,
      SEL => nx54672z94_BXINV,
      O => nx54672z94_F5MUX
    );
  nx54672z94_BXINV_5452 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z94_BXINV
    );
  romedatao1_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_7_F5MUX,
      O => nx54672z103
    );
  romedatao1_s_7_F5MUX_5453 : X_MUX2
    port map (
      IA => nx54672z104,
      IB => nx54672z105,
      SEL => romedatao1_s_7_BXINV,
      O => romedatao1_s_7_F5MUX
    );
  romedatao1_s_7_BXINV_5454 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao1_s_7_BXINV
    );
  romedatao1_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_7_F6MUX,
      O => romedatao1_s(7)
    );
  romedatao1_s_7_F6MUX_5455 : X_MUX2
    port map (
      IA => nx54672z100,
      IB => nx54672z103,
      SEL => romedatao1_s_7_BYINV,
      O => romedatao1_s_7_F6MUX
    );
  romedatao1_s_7_BYINV_5456 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao1_s_7_BYINV
    );
  nx54672z100_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z100_F5MUX,
      O => nx54672z100
    );
  nx54672z100_F5MUX_5457 : X_MUX2
    port map (
      IA => nx54672z101,
      IB => nx54672z102,
      SEL => nx54672z100_BXINV,
      O => nx54672z100_F5MUX
    );
  nx54672z100_BXINV_5458 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z100_BXINV
    );
  romedatao1_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_6_F5MUX,
      O => nx54672z109
    );
  romedatao1_s_6_F5MUX_5459 : X_MUX2
    port map (
      IA => nx54672z110,
      IB => nx54672z111,
      SEL => romedatao1_s_6_BXINV,
      O => romedatao1_s_6_F5MUX
    );
  romedatao1_s_6_BXINV_5460 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao1_s_6_BXINV
    );
  romedatao1_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_6_F6MUX,
      O => romedatao1_s(6)
    );
  romedatao1_s_6_F6MUX_5461 : X_MUX2
    port map (
      IA => nx54672z106,
      IB => nx54672z109,
      SEL => romedatao1_s_6_BYINV,
      O => romedatao1_s_6_F6MUX
    );
  romedatao1_s_6_BYINV_5462 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao1_s_6_BYINV
    );
  nx54672z106_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z106_F5MUX,
      O => nx54672z106
    );
  nx54672z106_F5MUX_5463 : X_MUX2
    port map (
      IA => nx54672z107,
      IB => nx54672z108,
      SEL => nx54672z106_BXINV,
      O => nx54672z106_F5MUX
    );
  nx54672z106_BXINV_5464 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z106_BXINV
    );
  romedatao1_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_5_F5MUX,
      O => nx54672z115
    );
  romedatao1_s_5_F5MUX_5465 : X_MUX2
    port map (
      IA => nx54672z116,
      IB => nx54672z117,
      SEL => romedatao1_s_5_BXINV,
      O => romedatao1_s_5_F5MUX
    );
  romedatao1_s_5_BXINV_5466 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao1_s_5_BXINV
    );
  romedatao1_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_5_F6MUX,
      O => romedatao1_s(5)
    );
  romedatao1_s_5_F6MUX_5467 : X_MUX2
    port map (
      IA => nx54672z112,
      IB => nx54672z115,
      SEL => romedatao1_s_5_BYINV,
      O => romedatao1_s_5_F6MUX
    );
  romedatao1_s_5_BYINV_5468 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao1_s_5_BYINV
    );
  nx54672z112_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z112_F5MUX,
      O => nx54672z112
    );
  nx54672z112_F5MUX_5469 : X_MUX2
    port map (
      IA => nx54672z113,
      IB => nx54672z114,
      SEL => nx54672z112_BXINV,
      O => nx54672z112_F5MUX
    );
  nx54672z112_BXINV_5470 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z112_BXINV
    );
  romedatao0_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_8_F5MUX,
      O => nx54672z33
    );
  romedatao0_s_8_F5MUX_5471 : X_MUX2
    port map (
      IA => nx54672z34,
      IB => nx54672z35,
      SEL => romedatao0_s_8_BXINV,
      O => romedatao0_s_8_F5MUX
    );
  romedatao0_s_8_BXINV_5472 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao0_s_8_BXINV
    );
  romedatao0_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_8_F6MUX,
      O => romedatao0_s(8)
    );
  romedatao0_s_8_F6MUX_5473 : X_MUX2
    port map (
      IA => nx54672z30,
      IB => nx54672z33,
      SEL => romedatao0_s_8_BYINV,
      O => romedatao0_s_8_F6MUX
    );
  romedatao0_s_8_BYINV_5474 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao0_s_8_BYINV
    );
  nx54672z30_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z30_F5MUX,
      O => nx54672z30
    );
  nx54672z30_F5MUX_5475 : X_MUX2
    port map (
      IA => nx54672z31,
      IB => nx54672z32,
      SEL => nx54672z30_BXINV,
      O => nx54672z30_F5MUX
    );
  nx54672z30_BXINV_5476 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z30_BXINV
    );
  U_DCT2D_reg_databuf_reg_4_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_4_6_DXMUX,
      CE => U_DCT2D_databuf_reg_4_6_CEINV,
      CLK => U_DCT2D_databuf_reg_4_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_4_6_FFX_RST,
      O => U_DCT2D_databuf_reg_4_Q(6)
    );
  U_DCT2D_databuf_reg_4_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_4_6_FFX_RST
    );
  romedatao0_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_7_F5MUX,
      O => nx54672z39
    );
  romedatao0_s_7_F5MUX_5477 : X_MUX2
    port map (
      IA => nx54672z40,
      IB => nx54672z41,
      SEL => romedatao0_s_7_BXINV,
      O => romedatao0_s_7_F5MUX
    );
  romedatao0_s_7_BXINV_5478 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao0_s_7_BXINV
    );
  romedatao0_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_7_F6MUX,
      O => romedatao0_s(7)
    );
  romedatao0_s_7_F6MUX_5479 : X_MUX2
    port map (
      IA => nx54672z36,
      IB => nx54672z39,
      SEL => romedatao0_s_7_BYINV,
      O => romedatao0_s_7_F6MUX
    );
  romedatao0_s_7_BYINV_5480 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao0_s_7_BYINV
    );
  nx54672z36_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z36_F5MUX,
      O => nx54672z36
    );
  nx54672z36_F5MUX_5481 : X_MUX2
    port map (
      IA => nx54672z37,
      IB => nx54672z38,
      SEL => nx54672z36_BXINV,
      O => nx54672z36_F5MUX
    );
  nx54672z36_BXINV_5482 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z36_BXINV
    );
  romedatao0_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_6_F5MUX,
      O => nx54672z45
    );
  romedatao0_s_6_F5MUX_5483 : X_MUX2
    port map (
      IA => nx54672z46,
      IB => nx54672z47,
      SEL => romedatao0_s_6_BXINV,
      O => romedatao0_s_6_F5MUX
    );
  romedatao0_s_6_BXINV_5484 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao0_s_6_BXINV
    );
  romedatao0_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_6_F6MUX,
      O => romedatao0_s(6)
    );
  romedatao0_s_6_F6MUX_5485 : X_MUX2
    port map (
      IA => nx54672z42,
      IB => nx54672z45,
      SEL => romedatao0_s_6_BYINV,
      O => romedatao0_s_6_F6MUX
    );
  romedatao0_s_6_BYINV_5486 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao0_s_6_BYINV
    );
  U_DCT2D_ix58525z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_0_10_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_7_10_Q,
      O => U_DCT2D_nx58525z1
    );
  nx54672z42_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z42_F5MUX,
      O => nx54672z42
    );
  nx54672z42_F5MUX_5487 : X_MUX2
    port map (
      IA => nx54672z43,
      IB => nx54672z44,
      SEL => nx54672z42_BXINV,
      O => nx54672z42_F5MUX
    );
  nx54672z42_BXINV_5488 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z42_BXINV
    );
  romedatao0_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_5_F5MUX,
      O => nx54672z51
    );
  romedatao0_s_5_F5MUX_5489 : X_MUX2
    port map (
      IA => nx54672z52,
      IB => nx54672z53,
      SEL => romedatao0_s_5_BXINV,
      O => romedatao0_s_5_F5MUX
    );
  romedatao0_s_5_BXINV_5490 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao0_s_5_BXINV
    );
  romedatao0_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_5_F6MUX,
      O => romedatao0_s(5)
    );
  romedatao0_s_5_F6MUX_5491 : X_MUX2
    port map (
      IA => nx54672z48,
      IB => nx54672z51,
      SEL => romedatao0_s_5_BYINV,
      O => romedatao0_s_5_F6MUX
    );
  romedatao0_s_5_BYINV_5492 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao0_s_5_BYINV
    );
  nx54672z48_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z48_F5MUX,
      O => nx54672z48
    );
  nx54672z48_F5MUX_5493 : X_MUX2
    port map (
      IA => nx54672z49,
      IB => nx54672z50,
      SEL => nx54672z48_BXINV,
      O => nx54672z48_F5MUX
    );
  nx54672z48_BXINV_5494 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z48_BXINV
    );
  romedatao0_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_4_F5MUX,
      O => nx54672z57
    );
  romedatao0_s_4_F5MUX_5495 : X_MUX2
    port map (
      IA => nx54672z58,
      IB => nx54672z59,
      SEL => romedatao0_s_4_BXINV,
      O => romedatao0_s_4_F5MUX
    );
  romedatao0_s_4_BXINV_5496 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao0_s_4_BXINV
    );
  romedatao0_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_4_F6MUX,
      O => romedatao0_s(4)
    );
  romedatao0_s_4_F6MUX_5497 : X_MUX2
    port map (
      IA => nx54672z54,
      IB => nx54672z57,
      SEL => romedatao0_s_4_BYINV,
      O => romedatao0_s_4_F6MUX
    );
  romedatao0_s_4_BYINV_5498 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao0_s_4_BYINV
    );
  nx54672z54_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z54_F5MUX,
      O => nx54672z54
    );
  nx54672z54_F5MUX_5499 : X_MUX2
    port map (
      IA => nx54672z55,
      IB => nx54672z56,
      SEL => nx54672z54_BXINV,
      O => nx54672z54_F5MUX
    );
  nx54672z54_BXINV_5500 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z54_BXINV
    );
  romodatao8_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_0_F5MUX,
      O => U1_ROMO8_modgen_rom_ix0_nx_ro64_32_l
    );
  romodatao8_s_0_F5MUX_5501 : X_MUX2
    port map (
      IA => nx54672z1292,
      IB => nx54672z1293,
      SEL => romodatao8_s_0_BXINV,
      O => romodatao8_s_0_F5MUX
    );
  romodatao8_s_0_BXINV_5502 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_0_BXINV
    );
  romodatao8_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_0_F6MUX,
      O => romodatao8_s(0)
    );
  romodatao8_s_0_F6MUX_5503 : X_MUX2
    port map (
      IA => U1_ROMO8_modgen_rom_ix0_nx_ro64_32_u,
      IB => U1_ROMO8_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romodatao8_s_0_BYINV,
      O => romodatao8_s_0_F6MUX
    );
  romodatao8_s_0_BYINV_5504 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_0_BYINV
    );
  ix54672z7221 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romoaddro8_s(2),
      O => U1_ROMO8_modgen_rom_ix0_nx_rm64_16_u
    );
  U1_ROMO8_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROMO8_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U1_ROMO8_modgen_rom_ix0_nx_ro64_32_u
    );
  U1_ROMO8_modgen_rom_ix0_nx_ro64_32_u_F5MUX_5505 : X_MUX2
    port map (
      IA => U1_ROMO8_modgen_rom_ix0_nx_rm64_16_u,
      IB => U1_ROMO8_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U1_ROMO8_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U1_ROMO8_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U1_ROMO8_modgen_rom_ix0_nx_ro64_32_u_BXINV_5506 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => U1_ROMO8_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romodatao1_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_13_F5MUX,
      O => nx54672z664
    );
  romodatao1_s_13_F5MUX_5507 : X_MUX2
    port map (
      IA => nx54672z665,
      IB => nx54672z666,
      SEL => romodatao1_s_13_BXINV,
      O => romodatao1_s_13_F5MUX
    );
  romodatao1_s_13_BXINV_5508 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_13_BXINV
    );
  romodatao1_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_13_F6MUX,
      O => romodatao1_s(13)
    );
  romodatao1_s_13_F6MUX_5509 : X_MUX2
    port map (
      IA => nx54672z662,
      IB => nx54672z664,
      SEL => romodatao1_s_13_BYINV,
      O => romodatao1_s_13_F6MUX
    );
  romodatao1_s_13_BYINV_5510 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_13_BYINV
    );
  nx54672z662_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z662_F5MUX,
      O => nx54672z662
    );
  nx54672z662_F5MUX_5511 : X_MUX2
    port map (
      IA => nx54672z662_G,
      IB => nx54672z663,
      SEL => nx54672z662_BXINV,
      O => nx54672z662_F5MUX
    );
  nx54672z662_BXINV_5512 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z662_BXINV
    );
  romodatao0_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_12_F5MUX,
      O => nx54672z593
    );
  romodatao0_s_12_F5MUX_5513 : X_MUX2
    port map (
      IA => nx54672z594,
      IB => nx54672z595,
      SEL => romodatao0_s_12_BXINV,
      O => romodatao0_s_12_F5MUX
    );
  romodatao0_s_12_BXINV_5514 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_12_BXINV
    );
  romodatao0_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_12_F6MUX,
      O => romodatao0_s(12)
    );
  romodatao0_s_12_F6MUX_5515 : X_MUX2
    port map (
      IA => nx54672z590,
      IB => nx54672z593,
      SEL => romodatao0_s_12_BYINV,
      O => romodatao0_s_12_F6MUX
    );
  romodatao0_s_12_BYINV_5516 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_12_BYINV
    );
  nx54672z590_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z590_F5MUX,
      O => nx54672z590
    );
  nx54672z590_F5MUX_5517 : X_MUX2
    port map (
      IA => nx54672z591,
      IB => nx54672z592,
      SEL => nx54672z590_BXINV,
      O => nx54672z590_F5MUX
    );
  nx54672z590_BXINV_5518 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z590_BXINV
    );
  romodatao0_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_11_F5MUX,
      O => nx54672z599
    );
  romodatao0_s_11_F5MUX_5519 : X_MUX2
    port map (
      IA => nx54672z600,
      IB => nx54672z601,
      SEL => romodatao0_s_11_BXINV,
      O => romodatao0_s_11_F5MUX
    );
  romodatao0_s_11_BXINV_5520 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_11_BXINV
    );
  romodatao0_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_11_F6MUX,
      O => romodatao0_s(11)
    );
  romodatao0_s_11_F6MUX_5521 : X_MUX2
    port map (
      IA => nx54672z596,
      IB => nx54672z599,
      SEL => romodatao0_s_11_BYINV,
      O => romodatao0_s_11_F6MUX
    );
  romodatao0_s_11_BYINV_5522 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_11_BYINV
    );
  nx54672z596_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z596_F5MUX,
      O => nx54672z596
    );
  nx54672z596_F5MUX_5523 : X_MUX2
    port map (
      IA => nx54672z597,
      IB => nx54672z598,
      SEL => nx54672z596_BXINV,
      O => nx54672z596_F5MUX
    );
  nx54672z596_BXINV_5524 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z596_BXINV
    );
  romodatao0_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_10_F5MUX,
      O => nx54672z605
    );
  romodatao0_s_10_F5MUX_5525 : X_MUX2
    port map (
      IA => nx54672z606,
      IB => nx54672z607,
      SEL => romodatao0_s_10_BXINV,
      O => romodatao0_s_10_F5MUX
    );
  romodatao0_s_10_BXINV_5526 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_10_BXINV
    );
  romodatao0_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_10_F6MUX,
      O => romodatao0_s(10)
    );
  romodatao0_s_10_F6MUX_5527 : X_MUX2
    port map (
      IA => nx54672z602,
      IB => nx54672z605,
      SEL => romodatao0_s_10_BYINV,
      O => romodatao0_s_10_F6MUX
    );
  romodatao0_s_10_BYINV_5528 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_10_BYINV
    );
  nx54672z602_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z602_F5MUX,
      O => nx54672z602
    );
  nx54672z602_F5MUX_5529 : X_MUX2
    port map (
      IA => nx54672z603,
      IB => nx54672z604,
      SEL => nx54672z602_BXINV,
      O => nx54672z602_F5MUX
    );
  nx54672z602_BXINV_5530 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z602_BXINV
    );
  romodatao0_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_9_F5MUX,
      O => nx54672z611
    );
  romodatao0_s_9_F5MUX_5531 : X_MUX2
    port map (
      IA => nx54672z612,
      IB => nx54672z613,
      SEL => romodatao0_s_9_BXINV,
      O => romodatao0_s_9_F5MUX
    );
  romodatao0_s_9_BXINV_5532 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_9_BXINV
    );
  romodatao0_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_9_F6MUX,
      O => romodatao0_s(9)
    );
  romodatao0_s_9_F6MUX_5533 : X_MUX2
    port map (
      IA => nx54672z608,
      IB => nx54672z611,
      SEL => romodatao0_s_9_BYINV,
      O => romodatao0_s_9_F6MUX
    );
  romodatao0_s_9_BYINV_5534 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_9_BYINV
    );
  nx54672z608_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z608_F5MUX,
      O => nx54672z608
    );
  nx54672z608_F5MUX_5535 : X_MUX2
    port map (
      IA => nx54672z609,
      IB => nx54672z610,
      SEL => nx54672z608_BXINV,
      O => nx54672z608_F5MUX
    );
  nx54672z608_BXINV_5536 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z608_BXINV
    );
  romodatao0_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_8_F5MUX,
      O => nx54672z617
    );
  romodatao0_s_8_F5MUX_5537 : X_MUX2
    port map (
      IA => nx54672z618,
      IB => nx54672z619,
      SEL => romodatao0_s_8_BXINV,
      O => romodatao0_s_8_F5MUX
    );
  romodatao0_s_8_BXINV_5538 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_8_BXINV
    );
  romodatao0_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_8_F6MUX,
      O => romodatao0_s(8)
    );
  romodatao0_s_8_F6MUX_5539 : X_MUX2
    port map (
      IA => nx54672z614,
      IB => nx54672z617,
      SEL => romodatao0_s_8_BYINV,
      O => romodatao0_s_8_F6MUX
    );
  romodatao0_s_8_BYINV_5540 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_8_BYINV
    );
  nx54672z614_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z614_F5MUX,
      O => nx54672z614
    );
  nx54672z614_F5MUX_5541 : X_MUX2
    port map (
      IA => nx54672z615,
      IB => nx54672z616,
      SEL => nx54672z614_BXINV,
      O => nx54672z614_F5MUX
    );
  nx54672z614_BXINV_5542 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z614_BXINV
    );
  romodatao0_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_1_F5MUX,
      O => nx54672z659
    );
  romodatao0_s_1_F5MUX_5543 : X_MUX2
    port map (
      IA => nx54672z660,
      IB => nx54672z661,
      SEL => romodatao0_s_1_BXINV,
      O => romodatao0_s_1_F5MUX
    );
  romodatao0_s_1_BXINV_5544 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_1_BXINV
    );
  romodatao0_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_1_F6MUX,
      O => romodatao0_s(1)
    );
  romodatao0_s_1_F6MUX_5545 : X_MUX2
    port map (
      IA => nx54672z656,
      IB => nx54672z659,
      SEL => romodatao0_s_1_BYINV,
      O => romodatao0_s_1_F6MUX
    );
  romodatao0_s_1_BYINV_5546 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_1_BYINV
    );
  nx54672z656_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z656_F5MUX,
      O => nx54672z656
    );
  nx54672z656_F5MUX_5547 : X_MUX2
    port map (
      IA => nx54672z657,
      IB => nx54672z658,
      SEL => nx54672z656_BXINV,
      O => nx54672z656_F5MUX
    );
  nx54672z656_BXINV_5548 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z656_BXINV
    );
  romedatao2_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_7_F5MUX,
      O => nx54672z168
    );
  romedatao2_s_7_F5MUX_5549 : X_MUX2
    port map (
      IA => nx54672z169,
      IB => nx54672z170,
      SEL => romedatao2_s_7_BXINV,
      O => romedatao2_s_7_F5MUX
    );
  romedatao2_s_7_BXINV_5550 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao2_s_7_BXINV
    );
  romedatao2_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_7_F6MUX,
      O => romedatao2_s(7)
    );
  romedatao2_s_7_F6MUX_5551 : X_MUX2
    port map (
      IA => nx54672z165,
      IB => nx54672z168,
      SEL => romedatao2_s_7_BYINV,
      O => romedatao2_s_7_F6MUX
    );
  romedatao2_s_7_BYINV_5552 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao2_s_7_BYINV
    );
  nx54672z165_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z165_F5MUX,
      O => nx54672z165
    );
  nx54672z165_F5MUX_5553 : X_MUX2
    port map (
      IA => nx54672z166,
      IB => nx54672z167,
      SEL => nx54672z165_BXINV,
      O => nx54672z165_F5MUX
    );
  nx54672z165_BXINV_5554 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z165_BXINV
    );
  romedatao2_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_6_F5MUX,
      O => nx54672z174
    );
  romedatao2_s_6_F5MUX_5555 : X_MUX2
    port map (
      IA => nx54672z175,
      IB => nx54672z176,
      SEL => romedatao2_s_6_BXINV,
      O => romedatao2_s_6_F5MUX
    );
  romedatao2_s_6_BXINV_5556 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao2_s_6_BXINV
    );
  romedatao2_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_6_F6MUX,
      O => romedatao2_s(6)
    );
  romedatao2_s_6_F6MUX_5557 : X_MUX2
    port map (
      IA => nx54672z171,
      IB => nx54672z174,
      SEL => romedatao2_s_6_BYINV,
      O => romedatao2_s_6_F6MUX
    );
  romedatao2_s_6_BYINV_5558 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao2_s_6_BYINV
    );
  nx54672z171_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z171_F5MUX,
      O => nx54672z171
    );
  nx54672z171_F5MUX_5559 : X_MUX2
    port map (
      IA => nx54672z172,
      IB => nx54672z173,
      SEL => nx54672z171_BXINV,
      O => nx54672z171_F5MUX
    );
  nx54672z171_BXINV_5560 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z171_BXINV
    );
  romedatao2_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_5_F5MUX,
      O => nx54672z180
    );
  romedatao2_s_5_F5MUX_5561 : X_MUX2
    port map (
      IA => nx54672z181,
      IB => nx54672z182,
      SEL => romedatao2_s_5_BXINV,
      O => romedatao2_s_5_F5MUX
    );
  romedatao2_s_5_BXINV_5562 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao2_s_5_BXINV
    );
  romedatao2_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_5_F6MUX,
      O => romedatao2_s(5)
    );
  romedatao2_s_5_F6MUX_5563 : X_MUX2
    port map (
      IA => nx54672z177,
      IB => nx54672z180,
      SEL => romedatao2_s_5_BYINV,
      O => romedatao2_s_5_F6MUX
    );
  romedatao2_s_5_BYINV_5564 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao2_s_5_BYINV
    );
  nx54672z177_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z177_F5MUX,
      O => nx54672z177
    );
  nx54672z177_F5MUX_5565 : X_MUX2
    port map (
      IA => nx54672z178,
      IB => nx54672z179,
      SEL => nx54672z177_BXINV,
      O => nx54672z177_F5MUX
    );
  nx54672z177_BXINV_5566 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z177_BXINV
    );
  romedatao2_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_4_F5MUX,
      O => nx54672z186
    );
  romedatao2_s_4_F5MUX_5567 : X_MUX2
    port map (
      IA => nx54672z187,
      IB => nx54672z188,
      SEL => romedatao2_s_4_BXINV,
      O => romedatao2_s_4_F5MUX
    );
  romedatao2_s_4_BXINV_5568 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao2_s_4_BXINV
    );
  romedatao2_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_4_F6MUX,
      O => romedatao2_s(4)
    );
  romedatao2_s_4_F6MUX_5569 : X_MUX2
    port map (
      IA => nx54672z183,
      IB => nx54672z186,
      SEL => romedatao2_s_4_BYINV,
      O => romedatao2_s_4_F6MUX
    );
  romedatao2_s_4_BYINV_5570 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao2_s_4_BYINV
    );
  nx54672z183_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z183_F5MUX,
      O => nx54672z183
    );
  nx54672z183_F5MUX_5571 : X_MUX2
    port map (
      IA => nx54672z184,
      IB => nx54672z185,
      SEL => nx54672z183_BXINV,
      O => nx54672z183_F5MUX
    );
  nx54672z183_BXINV_5572 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z183_BXINV
    );
  romedatao2_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_3_F5MUX,
      O => nx54672z191
    );
  romedatao2_s_3_F5MUX_5573 : X_MUX2
    port map (
      IA => nx54672z192,
      IB => nx54672z193,
      SEL => romedatao2_s_3_BXINV,
      O => romedatao2_s_3_F5MUX
    );
  romedatao2_s_3_BXINV_5574 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao2_s_3_BXINV
    );
  romedatao2_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_3_F6MUX,
      O => romedatao2_s(3)
    );
  romedatao2_s_3_F6MUX_5575 : X_MUX2
    port map (
      IA => nx54672z189,
      IB => nx54672z191,
      SEL => romedatao2_s_3_BYINV,
      O => romedatao2_s_3_F6MUX
    );
  romedatao2_s_3_BYINV_5576 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao2_s_3_BYINV
    );
  nx54672z189_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z189_F5MUX,
      O => nx54672z189
    );
  nx54672z189_F5MUX_5577 : X_MUX2
    port map (
      IA => U1_ROME2_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx54672z190,
      SEL => nx54672z189_BXINV,
      O => nx54672z189_F5MUX
    );
  nx54672z189_BXINV_5578 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z189_BXINV
    );
  romodatao2_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_12_F5MUX,
      O => nx54672z749
    );
  romodatao2_s_12_F5MUX_5579 : X_MUX2
    port map (
      IA => nx54672z750,
      IB => nx54672z751,
      SEL => romodatao2_s_12_BXINV,
      O => romodatao2_s_12_F5MUX
    );
  romodatao2_s_12_BXINV_5580 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_12_BXINV
    );
  romodatao2_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_12_F6MUX,
      O => romodatao2_s(12)
    );
  romodatao2_s_12_F6MUX_5581 : X_MUX2
    port map (
      IA => nx54672z746,
      IB => nx54672z749,
      SEL => romodatao2_s_12_BYINV,
      O => romodatao2_s_12_F6MUX
    );
  romodatao2_s_12_BYINV_5582 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_12_BYINV
    );
  ix54672z59715 : X_LUT4
    generic map(
      INIT => X"8880"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(1),
      ADR3 => romoaddro2_s(0),
      O => nx54672z747
    );
  nx54672z746_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z746_F5MUX,
      O => nx54672z746
    );
  nx54672z746_F5MUX_5583 : X_MUX2
    port map (
      IA => nx54672z747,
      IB => nx54672z748,
      SEL => nx54672z746_BXINV,
      O => nx54672z746_F5MUX
    );
  nx54672z746_BXINV_5584 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z746_BXINV
    );
  romodatao2_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_11_F5MUX,
      O => nx54672z755
    );
  romodatao2_s_11_F5MUX_5585 : X_MUX2
    port map (
      IA => nx54672z756,
      IB => nx54672z757,
      SEL => romodatao2_s_11_BXINV,
      O => romodatao2_s_11_F5MUX
    );
  romodatao2_s_11_BXINV_5586 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_11_BXINV
    );
  romodatao2_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_11_F6MUX,
      O => romodatao2_s(11)
    );
  romodatao2_s_11_F6MUX_5587 : X_MUX2
    port map (
      IA => nx54672z752,
      IB => nx54672z755,
      SEL => romodatao2_s_11_BYINV,
      O => romodatao2_s_11_F6MUX
    );
  romodatao2_s_11_BYINV_5588 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_11_BYINV
    );
  nx54672z752_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z752_F5MUX,
      O => nx54672z752
    );
  nx54672z752_F5MUX_5589 : X_MUX2
    port map (
      IA => nx54672z753,
      IB => nx54672z754,
      SEL => nx54672z752_BXINV,
      O => nx54672z752_F5MUX
    );
  nx54672z752_BXINV_5590 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z752_BXINV
    );
  U_DCT2D_reg_databuf_reg_4_9_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_4_8_DYMUX,
      CE => U_DCT2D_databuf_reg_4_8_CEINV,
      CLK => U_DCT2D_databuf_reg_4_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_4_8_FFY_RST,
      O => U_DCT2D_databuf_reg_4_Q(9)
    );
  U_DCT2D_databuf_reg_4_8_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_4_8_FFY_RST
    );
  romedatao2_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_13_F5MUX,
      O => nx54672z132
    );
  romedatao2_s_13_F5MUX_5591 : X_MUX2
    port map (
      IA => nx54672z133,
      IB => nx54672z134,
      SEL => romedatao2_s_13_BXINV,
      O => romedatao2_s_13_F5MUX
    );
  romedatao2_s_13_BXINV_5592 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao2_s_13_BXINV
    );
  romedatao2_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_13_F6MUX,
      O => romedatao2_s(13)
    );
  romedatao2_s_13_F6MUX_5593 : X_MUX2
    port map (
      IA => nx54672z130,
      IB => nx54672z132,
      SEL => romedatao2_s_13_BYINV,
      O => romedatao2_s_13_F6MUX
    );
  romedatao2_s_13_BYINV_5594 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao2_s_13_BYINV
    );
  nx54672z130_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z130_F5MUX,
      O => nx54672z130
    );
  nx54672z130_F5MUX_5595 : X_MUX2
    port map (
      IA => nx54672z130_G,
      IB => nx54672z131,
      SEL => nx54672z130_BXINV,
      O => nx54672z130_F5MUX
    );
  nx54672z130_BXINV_5596 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z130_BXINV
    );
  romedatao1_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_12_F5MUX,
      O => nx54672z73
    );
  romedatao1_s_12_F5MUX_5597 : X_MUX2
    port map (
      IA => nx54672z74,
      IB => nx54672z75,
      SEL => romedatao1_s_12_BXINV,
      O => romedatao1_s_12_F5MUX
    );
  romedatao1_s_12_BXINV_5598 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao1_s_12_BXINV
    );
  romedatao1_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_12_F6MUX,
      O => romedatao1_s(12)
    );
  romedatao1_s_12_F6MUX_5599 : X_MUX2
    port map (
      IA => nx54672z70,
      IB => nx54672z73,
      SEL => romedatao1_s_12_BYINV,
      O => romedatao1_s_12_F6MUX
    );
  romedatao1_s_12_BYINV_5600 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao1_s_12_BYINV
    );
  nx54672z70_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z70_F5MUX,
      O => nx54672z70
    );
  nx54672z70_F5MUX_5601 : X_MUX2
    port map (
      IA => nx54672z71,
      IB => nx54672z72,
      SEL => nx54672z70_BXINV,
      O => nx54672z70_F5MUX
    );
  nx54672z70_BXINV_5602 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z70_BXINV
    );
  romodatao2_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_13_F5MUX,
      O => nx54672z743
    );
  romodatao2_s_13_F5MUX_5603 : X_MUX2
    port map (
      IA => nx54672z744,
      IB => nx54672z745,
      SEL => romodatao2_s_13_BXINV,
      O => romodatao2_s_13_F5MUX
    );
  romodatao2_s_13_BXINV_5604 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_13_BXINV
    );
  romodatao2_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_13_F6MUX,
      O => romodatao2_s(13)
    );
  romodatao2_s_13_F6MUX_5605 : X_MUX2
    port map (
      IA => nx54672z741,
      IB => nx54672z743,
      SEL => romodatao2_s_13_BYINV,
      O => romodatao2_s_13_F6MUX
    );
  romodatao2_s_13_BYINV_5606 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_13_BYINV
    );
  nx54672z741_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z741_F5MUX,
      O => nx54672z741
    );
  nx54672z741_F5MUX_5607 : X_MUX2
    port map (
      IA => nx54672z741_G,
      IB => nx54672z742,
      SEL => nx54672z741_BXINV,
      O => nx54672z741_F5MUX
    );
  nx54672z741_BXINV_5608 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z741_BXINV
    );
  romodatao2_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_2_F5MUX,
      O => nx54672z809
    );
  romodatao2_s_2_F5MUX_5609 : X_MUX2
    port map (
      IA => nx54672z810,
      IB => nx54672z811,
      SEL => romodatao2_s_2_BXINV,
      O => romodatao2_s_2_F5MUX
    );
  romodatao2_s_2_BXINV_5610 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_2_BXINV
    );
  romodatao2_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_2_F6MUX,
      O => romodatao2_s(2)
    );
  romodatao2_s_2_F6MUX_5611 : X_MUX2
    port map (
      IA => nx54672z806,
      IB => nx54672z809,
      SEL => romodatao2_s_2_BYINV,
      O => romodatao2_s_2_F6MUX
    );
  romodatao2_s_2_BYINV_5612 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_2_BYINV
    );
  nx54672z806_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z806_F5MUX,
      O => nx54672z806
    );
  nx54672z806_F5MUX_5613 : X_MUX2
    port map (
      IA => nx54672z807,
      IB => nx54672z808,
      SEL => nx54672z806_BXINV,
      O => nx54672z806_F5MUX
    );
  nx54672z806_BXINV_5614 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z806_BXINV
    );
  romodatao2_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_1_F5MUX,
      O => nx54672z815
    );
  romodatao2_s_1_F5MUX_5615 : X_MUX2
    port map (
      IA => nx54672z816,
      IB => nx54672z817,
      SEL => romodatao2_s_1_BXINV,
      O => romodatao2_s_1_F5MUX
    );
  romodatao2_s_1_BXINV_5616 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_1_BXINV
    );
  romodatao2_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_1_F6MUX,
      O => romodatao2_s(1)
    );
  romodatao2_s_1_F6MUX_5617 : X_MUX2
    port map (
      IA => nx54672z812,
      IB => nx54672z815,
      SEL => romodatao2_s_1_BYINV,
      O => romodatao2_s_1_F6MUX
    );
  romodatao2_s_1_BYINV_5618 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_1_BYINV
    );
  nx54672z812_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z812_F5MUX,
      O => nx54672z812
    );
  nx54672z812_F5MUX_5619 : X_MUX2
    port map (
      IA => nx54672z813,
      IB => nx54672z814,
      SEL => nx54672z812_BXINV,
      O => nx54672z812_F5MUX
    );
  nx54672z812_BXINV_5620 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z812_BXINV
    );
  U_DCT2D_ix57528z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_0_8_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_7_8_Q,
      O => U_DCT2D_nx57528z1
    );
  romodatao2_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_0_F5MUX,
      O => U1_ROMO2_modgen_rom_ix0_nx_ro64_32_l
    );
  romodatao2_s_0_F5MUX_5621 : X_MUX2
    port map (
      IA => nx54672z818,
      IB => nx54672z819,
      SEL => romodatao2_s_0_BXINV,
      O => romodatao2_s_0_F5MUX
    );
  romodatao2_s_0_BXINV_5622 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_0_BXINV
    );
  romodatao2_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_0_F6MUX,
      O => romodatao2_s(0)
    );
  romodatao2_s_0_F6MUX_5623 : X_MUX2
    port map (
      IA => U1_ROMO2_modgen_rom_ix0_nx_ro64_32_u,
      IB => U1_ROMO2_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romodatao2_s_0_BYINV,
      O => romodatao2_s_0_F6MUX
    );
  romodatao2_s_0_BYINV_5624 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_0_BYINV
    );
  U1_ROMO2_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROMO2_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U1_ROMO2_modgen_rom_ix0_nx_ro64_32_u
    );
  U1_ROMO2_modgen_rom_ix0_nx_ro64_32_u_F5MUX_5625 : X_MUX2
    port map (
      IA => U1_ROMO2_modgen_rom_ix0_nx_rm64_16_u,
      IB => U1_ROMO2_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U1_ROMO2_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U1_ROMO2_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U1_ROMO2_modgen_rom_ix0_nx_ro64_32_u_BXINV_5626 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => U1_ROMO2_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romodatao1_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_10_F5MUX,
      O => nx54672z682
    );
  romodatao1_s_10_F5MUX_5627 : X_MUX2
    port map (
      IA => nx54672z683,
      IB => nx54672z684,
      SEL => romodatao1_s_10_BXINV,
      O => romodatao1_s_10_F5MUX
    );
  romodatao1_s_10_BXINV_5628 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_10_BXINV
    );
  romodatao1_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_10_F6MUX,
      O => romodatao1_s(10)
    );
  romodatao1_s_10_F6MUX_5629 : X_MUX2
    port map (
      IA => nx54672z679,
      IB => nx54672z682,
      SEL => romodatao1_s_10_BYINV,
      O => romodatao1_s_10_F6MUX
    );
  romodatao1_s_10_BYINV_5630 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_10_BYINV
    );
  nx54672z679_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z679_F5MUX,
      O => nx54672z679
    );
  nx54672z679_F5MUX_5631 : X_MUX2
    port map (
      IA => nx54672z680,
      IB => nx54672z681,
      SEL => nx54672z679_BXINV,
      O => nx54672z679_F5MUX
    );
  nx54672z679_BXINV_5632 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z679_BXINV
    );
  romodatao1_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_9_F5MUX,
      O => nx54672z688
    );
  romodatao1_s_9_F5MUX_5633 : X_MUX2
    port map (
      IA => nx54672z689,
      IB => nx54672z690,
      SEL => romodatao1_s_9_BXINV,
      O => romodatao1_s_9_F5MUX
    );
  romodatao1_s_9_BXINV_5634 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_9_BXINV
    );
  romodatao1_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_9_F6MUX,
      O => romodatao1_s(9)
    );
  romodatao1_s_9_F6MUX_5635 : X_MUX2
    port map (
      IA => nx54672z685,
      IB => nx54672z688,
      SEL => romodatao1_s_9_BYINV,
      O => romodatao1_s_9_F6MUX
    );
  romodatao1_s_9_BYINV_5636 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_9_BYINV
    );
  nx54672z685_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z685_F5MUX,
      O => nx54672z685
    );
  nx54672z685_F5MUX_5637 : X_MUX2
    port map (
      IA => nx54672z686,
      IB => nx54672z687,
      SEL => nx54672z685_BXINV,
      O => nx54672z685_F5MUX
    );
  nx54672z685_BXINV_5638 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z685_BXINV
    );
  romodatao1_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_8_F5MUX,
      O => nx54672z694
    );
  romodatao1_s_8_F5MUX_5639 : X_MUX2
    port map (
      IA => nx54672z695,
      IB => nx54672z696,
      SEL => romodatao1_s_8_BXINV,
      O => romodatao1_s_8_F5MUX
    );
  romodatao1_s_8_BXINV_5640 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_8_BXINV
    );
  romodatao1_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_8_F6MUX,
      O => romodatao1_s(8)
    );
  romodatao1_s_8_F6MUX_5641 : X_MUX2
    port map (
      IA => nx54672z691,
      IB => nx54672z694,
      SEL => romodatao1_s_8_BYINV,
      O => romodatao1_s_8_F6MUX
    );
  romodatao1_s_8_BYINV_5642 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_8_BYINV
    );
  nx54672z691_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z691_F5MUX,
      O => nx54672z691
    );
  nx54672z691_F5MUX_5643 : X_MUX2
    port map (
      IA => nx54672z692,
      IB => nx54672z693,
      SEL => nx54672z691_BXINV,
      O => nx54672z691_F5MUX
    );
  nx54672z691_BXINV_5644 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z691_BXINV
    );
  romodatao1_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_7_F5MUX,
      O => nx54672z700
    );
  romodatao1_s_7_F5MUX_5645 : X_MUX2
    port map (
      IA => nx54672z701,
      IB => nx54672z702,
      SEL => romodatao1_s_7_BXINV,
      O => romodatao1_s_7_F5MUX
    );
  romodatao1_s_7_BXINV_5646 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_7_BXINV
    );
  romodatao1_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_7_F6MUX,
      O => romodatao1_s(7)
    );
  romodatao1_s_7_F6MUX_5647 : X_MUX2
    port map (
      IA => nx54672z697,
      IB => nx54672z700,
      SEL => romodatao1_s_7_BYINV,
      O => romodatao1_s_7_F6MUX
    );
  romodatao1_s_7_BYINV_5648 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_7_BYINV
    );
  nx54672z697_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z697_F5MUX,
      O => nx54672z697
    );
  nx54672z697_F5MUX_5649 : X_MUX2
    port map (
      IA => nx54672z698,
      IB => nx54672z699,
      SEL => nx54672z697_BXINV,
      O => nx54672z697_F5MUX
    );
  nx54672z697_BXINV_5650 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z697_BXINV
    );
  romodatao1_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_6_F5MUX,
      O => nx54672z706
    );
  romodatao1_s_6_F5MUX_5651 : X_MUX2
    port map (
      IA => nx54672z707,
      IB => nx54672z708,
      SEL => romodatao1_s_6_BXINV,
      O => romodatao1_s_6_F5MUX
    );
  romodatao1_s_6_BXINV_5652 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_6_BXINV
    );
  romodatao1_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_6_F6MUX,
      O => romodatao1_s(6)
    );
  romodatao1_s_6_F6MUX_5653 : X_MUX2
    port map (
      IA => nx54672z703,
      IB => nx54672z706,
      SEL => romodatao1_s_6_BYINV,
      O => romodatao1_s_6_F6MUX
    );
  romodatao1_s_6_BYINV_5654 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_6_BYINV
    );
  nx54672z703_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z703_F5MUX,
      O => nx54672z703
    );
  nx54672z703_F5MUX_5655 : X_MUX2
    port map (
      IA => nx54672z704,
      IB => nx54672z705,
      SEL => nx54672z703_BXINV,
      O => nx54672z703_F5MUX
    );
  nx54672z703_BXINV_5656 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z703_BXINV
    );
  romodatao1_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_0_F5MUX,
      O => U1_ROMO1_modgen_rom_ix0_nx_ro64_32_l
    );
  romodatao1_s_0_F5MUX_5657 : X_MUX2
    port map (
      IA => nx54672z739,
      IB => nx54672z740,
      SEL => romodatao1_s_0_BXINV,
      O => romodatao1_s_0_F5MUX
    );
  romodatao1_s_0_BXINV_5658 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao1_s_0_BXINV
    );
  romodatao1_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao1_s_0_F6MUX,
      O => romodatao1_s(0)
    );
  romodatao1_s_0_F6MUX_5659 : X_MUX2
    port map (
      IA => U1_ROMO1_modgen_rom_ix0_nx_ro64_32_u,
      IB => U1_ROMO1_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romodatao1_s_0_BYINV,
      O => romodatao1_s_0_F6MUX
    );
  romodatao1_s_0_BYINV_5660 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao1_s_0_BYINV
    );
  U1_ROMO1_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROMO1_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U1_ROMO1_modgen_rom_ix0_nx_ro64_32_u
    );
  U1_ROMO1_modgen_rom_ix0_nx_ro64_32_u_F5MUX_5661 : X_MUX2
    port map (
      IA => U1_ROMO1_modgen_rom_ix0_nx_rm64_16_u,
      IB => U1_ROMO1_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U1_ROMO1_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U1_ROMO1_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U1_ROMO1_modgen_rom_ix0_nx_ro64_32_u_BXINV_5662 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => U1_ROMO1_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romedatao4_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_6_F5MUX,
      O => nx54672z304
    );
  romedatao4_s_6_F5MUX_5663 : X_MUX2
    port map (
      IA => nx54672z305,
      IB => nx54672z306,
      SEL => romedatao4_s_6_BXINV,
      O => romedatao4_s_6_F5MUX
    );
  romedatao4_s_6_BXINV_5664 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao4_s_6_BXINV
    );
  romedatao4_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_6_F6MUX,
      O => romedatao4_s(6)
    );
  romedatao4_s_6_F6MUX_5665 : X_MUX2
    port map (
      IA => nx54672z301,
      IB => nx54672z304,
      SEL => romedatao4_s_6_BYINV,
      O => romedatao4_s_6_F6MUX
    );
  romedatao4_s_6_BYINV_5666 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao4_s_6_BYINV
    );
  ix54672z34228 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(3),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(1),
      O => nx54672z302
    );
  nx54672z301_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z301_F5MUX,
      O => nx54672z301
    );
  nx54672z301_F5MUX_5667 : X_MUX2
    port map (
      IA => nx54672z302,
      IB => nx54672z303,
      SEL => nx54672z301_BXINV,
      O => nx54672z301_F5MUX
    );
  nx54672z301_BXINV_5668 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z301_BXINV
    );
  romedatao4_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_5_F5MUX,
      O => nx54672z310
    );
  romedatao4_s_5_F5MUX_5669 : X_MUX2
    port map (
      IA => nx54672z311,
      IB => nx54672z312,
      SEL => romedatao4_s_5_BXINV,
      O => romedatao4_s_5_F5MUX
    );
  romedatao4_s_5_BXINV_5670 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao4_s_5_BXINV
    );
  romedatao4_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_5_F6MUX,
      O => romedatao4_s(5)
    );
  romedatao4_s_5_F6MUX_5671 : X_MUX2
    port map (
      IA => nx54672z307,
      IB => nx54672z310,
      SEL => romedatao4_s_5_BYINV,
      O => romedatao4_s_5_F6MUX
    );
  romedatao4_s_5_BYINV_5672 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao4_s_5_BYINV
    );
  nx54672z307_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z307_F5MUX,
      O => nx54672z307
    );
  nx54672z307_F5MUX_5673 : X_MUX2
    port map (
      IA => nx54672z308,
      IB => nx54672z309,
      SEL => nx54672z307_BXINV,
      O => nx54672z307_F5MUX
    );
  nx54672z307_BXINV_5674 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z307_BXINV
    );
  romedatao1_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_13_F5MUX,
      O => nx54672z67
    );
  romedatao1_s_13_F5MUX_5675 : X_MUX2
    port map (
      IA => nx54672z68,
      IB => nx54672z69,
      SEL => romedatao1_s_13_BXINV,
      O => romedatao1_s_13_F5MUX
    );
  romedatao1_s_13_BXINV_5676 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao1_s_13_BXINV
    );
  romedatao1_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_13_F6MUX,
      O => romedatao1_s(13)
    );
  romedatao1_s_13_F6MUX_5677 : X_MUX2
    port map (
      IA => nx54672z65,
      IB => nx54672z67,
      SEL => romedatao1_s_13_BYINV,
      O => romedatao1_s_13_F6MUX
    );
  romedatao1_s_13_BYINV_5678 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao1_s_13_BYINV
    );
  nx54672z65_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z65_F5MUX,
      O => nx54672z65
    );
  nx54672z65_F5MUX_5679 : X_MUX2
    port map (
      IA => nx54672z65_G,
      IB => nx54672z66,
      SEL => nx54672z65_BXINV,
      O => nx54672z65_F5MUX
    );
  nx54672z65_BXINV_5680 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z65_BXINV
    );
  U_DCT2D_reg_databuf_reg_4_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_4_8_DXMUX,
      CE => U_DCT2D_databuf_reg_4_8_CEINV,
      CLK => U_DCT2D_databuf_reg_4_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_4_8_FFX_RST,
      O => U_DCT2D_databuf_reg_4_Q(8)
    );
  U_DCT2D_databuf_reg_4_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_4_8_FFX_RST
    );
  romedatao1_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_11_F5MUX,
      O => nx54672z79
    );
  romedatao1_s_11_F5MUX_5681 : X_MUX2
    port map (
      IA => nx54672z80,
      IB => nx54672z81,
      SEL => romedatao1_s_11_BXINV,
      O => romedatao1_s_11_F5MUX
    );
  romedatao1_s_11_BXINV_5682 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao1_s_11_BXINV
    );
  romedatao1_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_11_F6MUX,
      O => romedatao1_s(11)
    );
  romedatao1_s_11_F6MUX_5683 : X_MUX2
    port map (
      IA => nx54672z76,
      IB => nx54672z79,
      SEL => romedatao1_s_11_BYINV,
      O => romedatao1_s_11_F6MUX
    );
  romedatao1_s_11_BYINV_5684 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao1_s_11_BYINV
    );
  nx54672z76_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z76_F5MUX,
      O => nx54672z76
    );
  nx54672z76_F5MUX_5685 : X_MUX2
    port map (
      IA => nx54672z77,
      IB => nx54672z78,
      SEL => nx54672z76_BXINV,
      O => nx54672z76_F5MUX
    );
  nx54672z76_BXINV_5686 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z76_BXINV
    );
  romedatao1_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_10_F5MUX,
      O => nx54672z85
    );
  romedatao1_s_10_F5MUX_5687 : X_MUX2
    port map (
      IA => nx54672z86,
      IB => nx54672z87,
      SEL => romedatao1_s_10_BXINV,
      O => romedatao1_s_10_F5MUX
    );
  romedatao1_s_10_BXINV_5688 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao1_s_10_BXINV
    );
  romedatao1_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_10_F6MUX,
      O => romedatao1_s(10)
    );
  romedatao1_s_10_F6MUX_5689 : X_MUX2
    port map (
      IA => nx54672z82,
      IB => nx54672z85,
      SEL => romedatao1_s_10_BYINV,
      O => romedatao1_s_10_F6MUX
    );
  romedatao1_s_10_BYINV_5690 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao1_s_10_BYINV
    );
  nx54672z82_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z82_F5MUX,
      O => nx54672z82
    );
  nx54672z82_F5MUX_5691 : X_MUX2
    port map (
      IA => nx54672z83,
      IB => nx54672z84,
      SEL => nx54672z82_BXINV,
      O => nx54672z82_F5MUX
    );
  nx54672z82_BXINV_5692 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z82_BXINV
    );
  romedatao1_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_4_F5MUX,
      O => nx54672z121
    );
  romedatao1_s_4_F5MUX_5693 : X_MUX2
    port map (
      IA => nx54672z122,
      IB => nx54672z123,
      SEL => romedatao1_s_4_BXINV,
      O => romedatao1_s_4_F5MUX
    );
  romedatao1_s_4_BXINV_5694 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao1_s_4_BXINV
    );
  romedatao1_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_4_F6MUX,
      O => romedatao1_s(4)
    );
  romedatao1_s_4_F6MUX_5695 : X_MUX2
    port map (
      IA => nx54672z118,
      IB => nx54672z121,
      SEL => romedatao1_s_4_BYINV,
      O => romedatao1_s_4_F6MUX
    );
  romedatao1_s_4_BYINV_5696 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao1_s_4_BYINV
    );
  nx54672z118_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z118_F5MUX,
      O => nx54672z118
    );
  nx54672z118_F5MUX_5697 : X_MUX2
    port map (
      IA => nx54672z119,
      IB => nx54672z120,
      SEL => nx54672z118_BXINV,
      O => nx54672z118_F5MUX
    );
  nx54672z118_BXINV_5698 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z118_BXINV
    );
  romedatao1_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_3_F5MUX,
      O => nx54672z126
    );
  romedatao1_s_3_F5MUX_5699 : X_MUX2
    port map (
      IA => nx54672z127,
      IB => nx54672z128,
      SEL => romedatao1_s_3_BXINV,
      O => romedatao1_s_3_F5MUX
    );
  romedatao1_s_3_BXINV_5700 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao1_s_3_BXINV
    );
  romedatao1_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_3_F6MUX,
      O => romedatao1_s(3)
    );
  romedatao1_s_3_F6MUX_5701 : X_MUX2
    port map (
      IA => nx54672z124,
      IB => nx54672z126,
      SEL => romedatao1_s_3_BYINV,
      O => romedatao1_s_3_F6MUX
    );
  romedatao1_s_3_BYINV_5702 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao1_s_3_BYINV
    );
  nx54672z124_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z124_F5MUX,
      O => nx54672z124
    );
  nx54672z124_F5MUX_5703 : X_MUX2
    port map (
      IA => U1_ROME1_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx54672z125,
      SEL => nx54672z124_BXINV,
      O => nx54672z124_F5MUX
    );
  nx54672z124_BXINV_5704 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z124_BXINV
    );
  romedatao1_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_2_F5MUX,
      O => U1_ROME1_modgen_rom_ix2_nx_ro64_32_l
    );
  romedatao1_s_2_F5MUX_5705 : X_MUX2
    port map (
      IA => romedatao1_s_2_G,
      IB => nx54672z129,
      SEL => romedatao1_s_2_BXINV,
      O => romedatao1_s_2_F5MUX
    );
  romedatao1_s_2_BXINV_5706 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao1_s_2_BXINV
    );
  romedatao1_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_2_F6MUX,
      O => romedatao1_s(2)
    );
  romedatao1_s_2_F6MUX_5707 : X_MUX2
    port map (
      IA => U1_ROME1_modgen_rom_ix2_nx_ro64_32_u,
      IB => U1_ROME1_modgen_rom_ix2_nx_ro64_32_l,
      SEL => romedatao1_s_2_BYINV,
      O => romedatao1_s_2_F6MUX
    );
  romedatao1_s_2_BYINV_5708 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao1_s_2_BYINV
    );
  U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U1_ROME1_modgen_rom_ix2_nx_ro64_32_u
    );
  U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_F5MUX_5709 : X_MUX2
    port map (
      IA => U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U1_ROME1_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_BXINV_5710 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  romedatao0_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_12_F5MUX,
      O => nx54672z9
    );
  romedatao0_s_12_F5MUX_5711 : X_MUX2
    port map (
      IA => nx54672z10,
      IB => nx54672z11,
      SEL => romedatao0_s_12_BXINV,
      O => romedatao0_s_12_F5MUX
    );
  romedatao0_s_12_BXINV_5712 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao0_s_12_BXINV
    );
  romedatao0_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_12_F6MUX,
      O => romedatao0_s(12)
    );
  romedatao0_s_12_F6MUX_5713 : X_MUX2
    port map (
      IA => nx54672z6,
      IB => nx54672z9,
      SEL => romedatao0_s_12_BYINV,
      O => romedatao0_s_12_F6MUX
    );
  romedatao0_s_12_BYINV_5714 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao0_s_12_BYINV
    );
  nx54672z6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z6_F5MUX,
      O => nx54672z6
    );
  nx54672z6_F5MUX_5715 : X_MUX2
    port map (
      IA => nx54672z7,
      IB => nx54672z8,
      SEL => nx54672z6_BXINV,
      O => nx54672z6_F5MUX
    );
  nx54672z6_BXINV_5716 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z6_BXINV
    );
  romedatao0_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_11_F5MUX,
      O => nx54672z15
    );
  romedatao0_s_11_F5MUX_5717 : X_MUX2
    port map (
      IA => nx54672z16,
      IB => nx54672z17,
      SEL => romedatao0_s_11_BXINV,
      O => romedatao0_s_11_F5MUX
    );
  romedatao0_s_11_BXINV_5718 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao0_s_11_BXINV
    );
  romedatao0_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_11_F6MUX,
      O => romedatao0_s(11)
    );
  romedatao0_s_11_F6MUX_5719 : X_MUX2
    port map (
      IA => nx54672z12,
      IB => nx54672z15,
      SEL => romedatao0_s_11_BYINV,
      O => romedatao0_s_11_F6MUX
    );
  romedatao0_s_11_BYINV_5720 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao0_s_11_BYINV
    );
  nx54672z12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z12_F5MUX,
      O => nx54672z12
    );
  nx54672z12_F5MUX_5721 : X_MUX2
    port map (
      IA => nx54672z13,
      IB => nx54672z14,
      SEL => nx54672z12_BXINV,
      O => nx54672z12_F5MUX
    );
  nx54672z12_BXINV_5722 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z12_BXINV
    );
  romedatao0_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_3_F5MUX,
      O => nx54672z62
    );
  romedatao0_s_3_F5MUX_5723 : X_MUX2
    port map (
      IA => nx54672z63,
      IB => nx54672z64,
      SEL => romedatao0_s_3_BXINV,
      O => romedatao0_s_3_F5MUX
    );
  romedatao0_s_3_BXINV_5724 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao0_s_3_BXINV
    );
  romedatao0_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_3_F6MUX,
      O => romedatao0_s(3)
    );
  romedatao0_s_3_F6MUX_5725 : X_MUX2
    port map (
      IA => nx54672z60,
      IB => nx54672z62,
      SEL => romedatao0_s_3_BYINV,
      O => romedatao0_s_3_F6MUX
    );
  romedatao0_s_3_BYINV_5726 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao0_s_3_BYINV
    );
  nx54672z60_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z60_F5MUX,
      O => nx54672z60
    );
  nx54672z60_F5MUX_5727 : X_MUX2
    port map (
      IA => U1_ROME0_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx54672z61,
      SEL => nx54672z60_BXINV,
      O => nx54672z60_F5MUX
    );
  nx54672z60_BXINV_5728 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z60_BXINV
    );
  romodatao0_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_7_F5MUX,
      O => nx54672z623
    );
  romodatao0_s_7_F5MUX_5729 : X_MUX2
    port map (
      IA => nx54672z624,
      IB => nx54672z625,
      SEL => romodatao0_s_7_BXINV,
      O => romodatao0_s_7_F5MUX
    );
  romodatao0_s_7_BXINV_5730 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_7_BXINV
    );
  romodatao0_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_7_F6MUX,
      O => romodatao0_s(7)
    );
  romodatao0_s_7_F6MUX_5731 : X_MUX2
    port map (
      IA => nx54672z620,
      IB => nx54672z623,
      SEL => romodatao0_s_7_BYINV,
      O => romodatao0_s_7_F6MUX
    );
  romodatao0_s_7_BYINV_5732 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_7_BYINV
    );
  nx54672z620_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z620_F5MUX,
      O => nx54672z620
    );
  nx54672z620_F5MUX_5733 : X_MUX2
    port map (
      IA => nx54672z621,
      IB => nx54672z622,
      SEL => nx54672z620_BXINV,
      O => nx54672z620_F5MUX
    );
  nx54672z620_BXINV_5734 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z620_BXINV
    );
  romodatao0_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_6_F5MUX,
      O => nx54672z629
    );
  romodatao0_s_6_F5MUX_5735 : X_MUX2
    port map (
      IA => nx54672z630,
      IB => nx54672z631,
      SEL => romodatao0_s_6_BXINV,
      O => romodatao0_s_6_F5MUX
    );
  romodatao0_s_6_BXINV_5736 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_6_BXINV
    );
  romodatao0_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_6_F6MUX,
      O => romodatao0_s(6)
    );
  romodatao0_s_6_F6MUX_5737 : X_MUX2
    port map (
      IA => nx54672z626,
      IB => nx54672z629,
      SEL => romodatao0_s_6_BYINV,
      O => romodatao0_s_6_F6MUX
    );
  romodatao0_s_6_BYINV_5738 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_6_BYINV
    );
  nx54672z626_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z626_F5MUX,
      O => nx54672z626
    );
  nx54672z626_F5MUX_5739 : X_MUX2
    port map (
      IA => nx54672z627,
      IB => nx54672z628,
      SEL => nx54672z626_BXINV,
      O => nx54672z626_F5MUX
    );
  nx54672z626_BXINV_5740 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z626_BXINV
    );
  romodatao0_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_5_F5MUX,
      O => nx54672z635
    );
  romodatao0_s_5_F5MUX_5741 : X_MUX2
    port map (
      IA => nx54672z636,
      IB => nx54672z637,
      SEL => romodatao0_s_5_BXINV,
      O => romodatao0_s_5_F5MUX
    );
  romodatao0_s_5_BXINV_5742 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_5_BXINV
    );
  romodatao0_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_5_F6MUX,
      O => romodatao0_s(5)
    );
  romodatao0_s_5_F6MUX_5743 : X_MUX2
    port map (
      IA => nx54672z632,
      IB => nx54672z635,
      SEL => romodatao0_s_5_BYINV,
      O => romodatao0_s_5_F6MUX
    );
  romodatao0_s_5_BYINV_5744 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_5_BYINV
    );
  nx54672z632_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z632_F5MUX,
      O => nx54672z632
    );
  nx54672z632_F5MUX_5745 : X_MUX2
    port map (
      IA => nx54672z633,
      IB => nx54672z634,
      SEL => nx54672z632_BXINV,
      O => nx54672z632_F5MUX
    );
  nx54672z632_BXINV_5746 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z632_BXINV
    );
  romodatao0_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_4_F5MUX,
      O => nx54672z641
    );
  romodatao0_s_4_F5MUX_5747 : X_MUX2
    port map (
      IA => nx54672z642,
      IB => nx54672z643,
      SEL => romodatao0_s_4_BXINV,
      O => romodatao0_s_4_F5MUX
    );
  romodatao0_s_4_BXINV_5748 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_4_BXINV
    );
  romodatao0_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_4_F6MUX,
      O => romodatao0_s(4)
    );
  romodatao0_s_4_F6MUX_5749 : X_MUX2
    port map (
      IA => nx54672z638,
      IB => nx54672z641,
      SEL => romodatao0_s_4_BYINV,
      O => romodatao0_s_4_F6MUX
    );
  romodatao0_s_4_BYINV_5750 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_4_BYINV
    );
  U_DCT2D_reg_databuf_reg_4_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_4_10_DXMUX,
      CE => U_DCT2D_databuf_reg_4_10_CEINV,
      CLK => U_DCT2D_databuf_reg_4_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_4_10_FFX_RST,
      O => U_DCT2D_databuf_reg_4_Q(10)
    );
  U_DCT2D_databuf_reg_4_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_4_10_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_4_10_FFX_RST
    );
  U_DCT2D_databuf_reg_4_10_FFX_RSTAND_5751 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_4_10_FFX_RSTAND
    );
  nx54672z638_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z638_F5MUX,
      O => nx54672z638
    );
  nx54672z638_F5MUX_5752 : X_MUX2
    port map (
      IA => nx54672z639,
      IB => nx54672z640,
      SEL => nx54672z638_BXINV,
      O => nx54672z638_F5MUX
    );
  nx54672z638_BXINV_5753 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z638_BXINV
    );
  romodatao0_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_3_F5MUX,
      O => nx54672z647
    );
  romodatao0_s_3_F5MUX_5754 : X_MUX2
    port map (
      IA => nx54672z648,
      IB => nx54672z649,
      SEL => romodatao0_s_3_BXINV,
      O => romodatao0_s_3_F5MUX
    );
  romodatao0_s_3_BXINV_5755 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_3_BXINV
    );
  romodatao0_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_3_F6MUX,
      O => romodatao0_s(3)
    );
  romodatao0_s_3_F6MUX_5756 : X_MUX2
    port map (
      IA => nx54672z644,
      IB => nx54672z647,
      SEL => romodatao0_s_3_BYINV,
      O => romodatao0_s_3_F6MUX
    );
  romodatao0_s_3_BYINV_5757 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_3_BYINV
    );
  nx54672z644_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z644_F5MUX,
      O => nx54672z644
    );
  nx54672z644_F5MUX_5758 : X_MUX2
    port map (
      IA => nx54672z645,
      IB => nx54672z646,
      SEL => nx54672z644_BXINV,
      O => nx54672z644_F5MUX
    );
  nx54672z644_BXINV_5759 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z644_BXINV
    );
  romedatao0_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_13_F5MUX,
      O => nx54672z3
    );
  romedatao0_s_13_F5MUX_5760 : X_MUX2
    port map (
      IA => nx54672z4,
      IB => nx54672z5,
      SEL => romedatao0_s_13_BXINV,
      O => romedatao0_s_13_F5MUX
    );
  romedatao0_s_13_BXINV_5761 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao0_s_13_BXINV
    );
  romedatao0_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao0_s_13_F6MUX,
      O => romedatao0_s(13)
    );
  romedatao0_s_13_F6MUX_5762 : X_MUX2
    port map (
      IA => nx54672z1,
      IB => nx54672z3,
      SEL => romedatao0_s_13_BYINV,
      O => romedatao0_s_13_F6MUX
    );
  romedatao0_s_13_BYINV_5763 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao0_s_13_BYINV
    );
  nx54672z1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1_F5MUX,
      O => nx54672z1
    );
  nx54672z1_F5MUX_5764 : X_MUX2
    port map (
      IA => nx54672z1_G,
      IB => nx54672z2,
      SEL => nx54672z1_BXINV,
      O => nx54672z1_F5MUX
    );
  nx54672z1_BXINV_5765 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z1_BXINV
    );
  romedatao3_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_12_F5MUX,
      O => nx54672z203
    );
  romedatao3_s_12_F5MUX_5766 : X_MUX2
    port map (
      IA => nx54672z204,
      IB => nx54672z205,
      SEL => romedatao3_s_12_BXINV,
      O => romedatao3_s_12_F5MUX
    );
  romedatao3_s_12_BXINV_5767 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao3_s_12_BXINV
    );
  romedatao3_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_12_F6MUX,
      O => romedatao3_s(12)
    );
  romedatao3_s_12_F6MUX_5768 : X_MUX2
    port map (
      IA => nx54672z200,
      IB => nx54672z203,
      SEL => romedatao3_s_12_BYINV,
      O => romedatao3_s_12_F6MUX
    );
  romedatao3_s_12_BYINV_5769 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao3_s_12_BYINV
    );
  ix54672z61119 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z201
    );
  nx54672z200_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z200_F5MUX,
      O => nx54672z200
    );
  nx54672z200_F5MUX_5770 : X_MUX2
    port map (
      IA => nx54672z201,
      IB => nx54672z202,
      SEL => nx54672z200_BXINV,
      O => nx54672z200_F5MUX
    );
  nx54672z200_BXINV_5771 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z200_BXINV
    );
  romedatao3_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_6_F5MUX,
      O => nx54672z239
    );
  romedatao3_s_6_F5MUX_5772 : X_MUX2
    port map (
      IA => nx54672z240,
      IB => nx54672z241,
      SEL => romedatao3_s_6_BXINV,
      O => romedatao3_s_6_F5MUX
    );
  romedatao3_s_6_BXINV_5773 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao3_s_6_BXINV
    );
  romedatao3_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_6_F6MUX,
      O => romedatao3_s(6)
    );
  romedatao3_s_6_F6MUX_5774 : X_MUX2
    port map (
      IA => nx54672z236,
      IB => nx54672z239,
      SEL => romedatao3_s_6_BYINV,
      O => romedatao3_s_6_F6MUX
    );
  romedatao3_s_6_BYINV_5775 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao3_s_6_BYINV
    );
  nx54672z236_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z236_F5MUX,
      O => nx54672z236
    );
  nx54672z236_F5MUX_5776 : X_MUX2
    port map (
      IA => nx54672z237,
      IB => nx54672z238,
      SEL => nx54672z236_BXINV,
      O => nx54672z236_F5MUX
    );
  nx54672z236_BXINV_5777 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z236_BXINV
    );
  romedatao3_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_4_F5MUX,
      O => nx54672z251
    );
  romedatao3_s_4_F5MUX_5778 : X_MUX2
    port map (
      IA => nx54672z252,
      IB => nx54672z253,
      SEL => romedatao3_s_4_BXINV,
      O => romedatao3_s_4_F5MUX
    );
  romedatao3_s_4_BXINV_5779 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao3_s_4_BXINV
    );
  romedatao3_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_4_F6MUX,
      O => romedatao3_s(4)
    );
  romedatao3_s_4_F6MUX_5780 : X_MUX2
    port map (
      IA => nx54672z248,
      IB => nx54672z251,
      SEL => romedatao3_s_4_BYINV,
      O => romedatao3_s_4_F6MUX
    );
  romedatao3_s_4_BYINV_5781 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao3_s_4_BYINV
    );
  nx54672z248_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z248_F5MUX,
      O => nx54672z248
    );
  nx54672z248_F5MUX_5782 : X_MUX2
    port map (
      IA => nx54672z249,
      IB => nx54672z250,
      SEL => nx54672z248_BXINV,
      O => nx54672z248_F5MUX
    );
  nx54672z248_BXINV_5783 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z248_BXINV
    );
  romedatao3_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_2_F5MUX,
      O => U1_ROME3_modgen_rom_ix2_nx_ro64_32_l
    );
  romedatao3_s_2_F5MUX_5784 : X_MUX2
    port map (
      IA => romedatao3_s_2_G,
      IB => nx54672z259,
      SEL => romedatao3_s_2_BXINV,
      O => romedatao3_s_2_F5MUX
    );
  romedatao3_s_2_BXINV_5785 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao3_s_2_BXINV
    );
  romedatao3_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_2_F6MUX,
      O => romedatao3_s(2)
    );
  romedatao3_s_2_F6MUX_5786 : X_MUX2
    port map (
      IA => U1_ROME3_modgen_rom_ix2_nx_ro64_32_u,
      IB => U1_ROME3_modgen_rom_ix2_nx_ro64_32_l,
      SEL => romedatao3_s_2_BYINV,
      O => romedatao3_s_2_F6MUX
    );
  romedatao3_s_2_BYINV_5787 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao3_s_2_BYINV
    );
  U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U1_ROME3_modgen_rom_ix2_nx_ro64_32_u
    );
  U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_F5MUX_5788 : X_MUX2
    port map (
      IA => U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U1_ROME3_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_BXINV_5789 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  romedatao3_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_13_F5MUX,
      O => nx54672z197
    );
  romedatao3_s_13_F5MUX_5790 : X_MUX2
    port map (
      IA => nx54672z198,
      IB => nx54672z199,
      SEL => romedatao3_s_13_BXINV,
      O => romedatao3_s_13_F5MUX
    );
  romedatao3_s_13_BXINV_5791 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao3_s_13_BXINV
    );
  romedatao3_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_13_F6MUX,
      O => romedatao3_s(13)
    );
  romedatao3_s_13_F6MUX_5792 : X_MUX2
    port map (
      IA => nx54672z195,
      IB => nx54672z197,
      SEL => romedatao3_s_13_BYINV,
      O => romedatao3_s_13_F6MUX
    );
  romedatao3_s_13_BYINV_5793 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao3_s_13_BYINV
    );
  nx54672z195_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z195_F5MUX,
      O => nx54672z195
    );
  nx54672z195_F5MUX_5794 : X_MUX2
    port map (
      IA => nx54672z195_G,
      IB => nx54672z196,
      SEL => nx54672z195_BXINV,
      O => nx54672z195_F5MUX
    );
  nx54672z195_BXINV_5795 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z195_BXINV
    );
  U_DCT2D_ix35144z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_4_1_Q,
      ADR1 => U_DCT2D_latchbuf_reg_3_1_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx35144z1
    );
  romedatao5_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_5_F5MUX,
      O => nx54672z375
    );
  romedatao5_s_5_F5MUX_5796 : X_MUX2
    port map (
      IA => nx54672z376,
      IB => nx54672z377,
      SEL => romedatao5_s_5_BXINV,
      O => romedatao5_s_5_F5MUX
    );
  romedatao5_s_5_BXINV_5797 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao5_s_5_BXINV
    );
  romedatao5_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_5_F6MUX,
      O => romedatao5_s(5)
    );
  romedatao5_s_5_F6MUX_5798 : X_MUX2
    port map (
      IA => nx54672z372,
      IB => nx54672z375,
      SEL => romedatao5_s_5_BYINV,
      O => romedatao5_s_5_F6MUX
    );
  romedatao5_s_5_BYINV_5799 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao5_s_5_BYINV
    );
  ix54672z61639 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => romeaddro5_s(2),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(3),
      O => nx54672z373
    );
  nx54672z372_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z372_F5MUX,
      O => nx54672z372
    );
  nx54672z372_F5MUX_5800 : X_MUX2
    port map (
      IA => nx54672z373,
      IB => nx54672z374,
      SEL => nx54672z372_BXINV,
      O => nx54672z372_F5MUX
    );
  nx54672z372_BXINV_5801 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z372_BXINV
    );
  romedatao5_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_4_F5MUX,
      O => nx54672z381
    );
  romedatao5_s_4_F5MUX_5802 : X_MUX2
    port map (
      IA => nx54672z382,
      IB => nx54672z383,
      SEL => romedatao5_s_4_BXINV,
      O => romedatao5_s_4_F5MUX
    );
  romedatao5_s_4_BXINV_5803 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao5_s_4_BXINV
    );
  romedatao5_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_4_F6MUX,
      O => romedatao5_s(4)
    );
  romedatao5_s_4_F6MUX_5804 : X_MUX2
    port map (
      IA => nx54672z378,
      IB => nx54672z381,
      SEL => romedatao5_s_4_BYINV,
      O => romedatao5_s_4_F6MUX
    );
  romedatao5_s_4_BYINV_5805 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao5_s_4_BYINV
    );
  nx54672z378_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z378_F5MUX,
      O => nx54672z378
    );
  nx54672z378_F5MUX_5806 : X_MUX2
    port map (
      IA => nx54672z379,
      IB => nx54672z380,
      SEL => nx54672z378_BXINV,
      O => nx54672z378_F5MUX
    );
  nx54672z378_BXINV_5807 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z378_BXINV
    );
  romodatao5_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_8_F5MUX,
      O => nx54672z1010
    );
  romodatao5_s_8_F5MUX_5808 : X_MUX2
    port map (
      IA => nx54672z1011,
      IB => nx54672z1012,
      SEL => romodatao5_s_8_BXINV,
      O => romodatao5_s_8_F5MUX
    );
  romodatao5_s_8_BXINV_5809 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_8_BXINV
    );
  romodatao5_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_8_F6MUX,
      O => romodatao5_s(8)
    );
  romodatao5_s_8_F6MUX_5810 : X_MUX2
    port map (
      IA => nx54672z1007,
      IB => nx54672z1010,
      SEL => romodatao5_s_8_BYINV,
      O => romodatao5_s_8_F6MUX
    );
  romodatao5_s_8_BYINV_5811 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_8_BYINV
    );
  ix54672z5620 : X_LUT4
    generic map(
      INIT => X"2342"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(1),
      ADR3 => romoaddro5_s(0),
      O => nx54672z1008
    );
  nx54672z1007_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1007_F5MUX,
      O => nx54672z1007
    );
  nx54672z1007_F5MUX_5812 : X_MUX2
    port map (
      IA => nx54672z1008,
      IB => nx54672z1009,
      SEL => nx54672z1007_BXINV,
      O => nx54672z1007_F5MUX
    );
  nx54672z1007_BXINV_5813 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1007_BXINV
    );
  romedatao5_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_13_F5MUX,
      O => nx54672z327
    );
  romedatao5_s_13_F5MUX_5814 : X_MUX2
    port map (
      IA => nx54672z328,
      IB => nx54672z329,
      SEL => romedatao5_s_13_BXINV,
      O => romedatao5_s_13_F5MUX
    );
  romedatao5_s_13_BXINV_5815 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao5_s_13_BXINV
    );
  romedatao5_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_13_F6MUX,
      O => romedatao5_s(13)
    );
  romedatao5_s_13_F6MUX_5816 : X_MUX2
    port map (
      IA => nx54672z325,
      IB => nx54672z327,
      SEL => romedatao5_s_13_BYINV,
      O => romedatao5_s_13_F6MUX
    );
  romedatao5_s_13_BYINV_5817 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao5_s_13_BYINV
    );
  nx54672z325_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z325_F5MUX,
      O => nx54672z325
    );
  nx54672z325_F5MUX_5818 : X_MUX2
    port map (
      IA => nx54672z325_G,
      IB => nx54672z326,
      SEL => nx54672z325_BXINV,
      O => nx54672z325_F5MUX
    );
  nx54672z325_BXINV_5819 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z325_BXINV
    );
  romedatao2_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_12_F5MUX,
      O => nx54672z138
    );
  romedatao2_s_12_F5MUX_5820 : X_MUX2
    port map (
      IA => nx54672z139,
      IB => nx54672z140,
      SEL => romedatao2_s_12_BXINV,
      O => romedatao2_s_12_F5MUX
    );
  romedatao2_s_12_BXINV_5821 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao2_s_12_BXINV
    );
  romedatao2_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_12_F6MUX,
      O => romedatao2_s(12)
    );
  romedatao2_s_12_F6MUX_5822 : X_MUX2
    port map (
      IA => nx54672z135,
      IB => nx54672z138,
      SEL => romedatao2_s_12_BYINV,
      O => romedatao2_s_12_F6MUX
    );
  romedatao2_s_12_BYINV_5823 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao2_s_12_BYINV
    );
  nx54672z135_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z135_F5MUX,
      O => nx54672z135
    );
  nx54672z135_F5MUX_5824 : X_MUX2
    port map (
      IA => nx54672z136,
      IB => nx54672z137,
      SEL => nx54672z135_BXINV,
      O => nx54672z135_F5MUX
    );
  nx54672z135_BXINV_5825 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z135_BXINV
    );
  romedatao2_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_11_F5MUX,
      O => nx54672z144
    );
  romedatao2_s_11_F5MUX_5826 : X_MUX2
    port map (
      IA => nx54672z145,
      IB => nx54672z146,
      SEL => romedatao2_s_11_BXINV,
      O => romedatao2_s_11_F5MUX
    );
  romedatao2_s_11_BXINV_5827 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao2_s_11_BXINV
    );
  romedatao2_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_11_F6MUX,
      O => romedatao2_s(11)
    );
  romedatao2_s_11_F6MUX_5828 : X_MUX2
    port map (
      IA => nx54672z141,
      IB => nx54672z144,
      SEL => romedatao2_s_11_BYINV,
      O => romedatao2_s_11_F6MUX
    );
  romedatao2_s_11_BYINV_5829 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao2_s_11_BYINV
    );
  nx54672z141_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z141_F5MUX,
      O => nx54672z141
    );
  nx54672z141_F5MUX_5830 : X_MUX2
    port map (
      IA => nx54672z142,
      IB => nx54672z143,
      SEL => nx54672z141_BXINV,
      O => nx54672z141_F5MUX
    );
  nx54672z141_BXINV_5831 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z141_BXINV
    );
  romedatao2_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_10_F5MUX,
      O => nx54672z150
    );
  romedatao2_s_10_F5MUX_5832 : X_MUX2
    port map (
      IA => nx54672z151,
      IB => nx54672z152,
      SEL => romedatao2_s_10_BXINV,
      O => romedatao2_s_10_F5MUX
    );
  romedatao2_s_10_BXINV_5833 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao2_s_10_BXINV
    );
  romedatao2_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_10_F6MUX,
      O => romedatao2_s(10)
    );
  romedatao2_s_10_F6MUX_5834 : X_MUX2
    port map (
      IA => nx54672z147,
      IB => nx54672z150,
      SEL => romedatao2_s_10_BYINV,
      O => romedatao2_s_10_F6MUX
    );
  romedatao2_s_10_BYINV_5835 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao2_s_10_BYINV
    );
  nx54672z147_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z147_F5MUX,
      O => nx54672z147
    );
  nx54672z147_F5MUX_5836 : X_MUX2
    port map (
      IA => nx54672z148,
      IB => nx54672z149,
      SEL => nx54672z147_BXINV,
      O => nx54672z147_F5MUX
    );
  nx54672z147_BXINV_5837 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z147_BXINV
    );
  romedatao2_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_9_F5MUX,
      O => nx54672z156
    );
  romedatao2_s_9_F5MUX_5838 : X_MUX2
    port map (
      IA => nx54672z157,
      IB => nx54672z158,
      SEL => romedatao2_s_9_BXINV,
      O => romedatao2_s_9_F5MUX
    );
  romedatao2_s_9_BXINV_5839 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao2_s_9_BXINV
    );
  romedatao2_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_9_F6MUX,
      O => romedatao2_s(9)
    );
  romedatao2_s_9_F6MUX_5840 : X_MUX2
    port map (
      IA => nx54672z153,
      IB => nx54672z156,
      SEL => romedatao2_s_9_BYINV,
      O => romedatao2_s_9_F6MUX
    );
  romedatao2_s_9_BYINV_5841 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao2_s_9_BYINV
    );
  nx54672z153_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z153_F5MUX,
      O => nx54672z153
    );
  nx54672z153_F5MUX_5842 : X_MUX2
    port map (
      IA => nx54672z154,
      IB => nx54672z155,
      SEL => nx54672z153_BXINV,
      O => nx54672z153_F5MUX
    );
  nx54672z153_BXINV_5843 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z153_BXINV
    );
  romedatao2_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_2_F5MUX,
      O => U1_ROME2_modgen_rom_ix2_nx_ro64_32_l
    );
  romedatao2_s_2_F5MUX_5844 : X_MUX2
    port map (
      IA => romedatao2_s_2_G,
      IB => nx54672z194,
      SEL => romedatao2_s_2_BXINV,
      O => romedatao2_s_2_F5MUX
    );
  romedatao2_s_2_BXINV_5845 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao2_s_2_BXINV
    );
  romedatao2_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao2_s_2_F6MUX,
      O => romedatao2_s(2)
    );
  romedatao2_s_2_F6MUX_5846 : X_MUX2
    port map (
      IA => U1_ROME2_modgen_rom_ix2_nx_ro64_32_u,
      IB => U1_ROME2_modgen_rom_ix2_nx_ro64_32_l,
      SEL => romedatao2_s_2_BYINV,
      O => romedatao2_s_2_F6MUX
    );
  romedatao2_s_2_BYINV_5847 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao2_s_2_BYINV
    );
  U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U1_ROME2_modgen_rom_ix2_nx_ro64_32_u
    );
  U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_F5MUX_5848 : X_MUX2
    port map (
      IA => U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U1_ROME2_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_BXINV_5849 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  U_DCT2D_ix65206z24321 : X_LUT4
    generic map(
      INIT => X"3C66"
    )
    port map (
      ADR0 => rome2datao9_s(8),
      ADR1 => U_DCT2D_nx65206z589,
      ADR2 => romo2datao9_s(8),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z588
    );
  U_DCT2D_ix65206z24315 : X_LUT4
    generic map(
      INIT => X"56A6"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z583,
      ADR1 => rome2datao9_s(10),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao9_s(10),
      O => U_DCT2D_nx65206z582
    );
  U_DCT2D_nx65206z572_rt_5850 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_nx65206z572,
      O => U_DCT2D_nx65206z572_rt
    );
  nx54672z313_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z313_F5MUX,
      O => nx54672z313
    );
  nx54672z313_F5MUX_5851 : X_MUX2
    port map (
      IA => nx54672z314,
      IB => nx54672z315,
      SEL => nx54672z313_BXINV,
      O => nx54672z313_F5MUX
    );
  nx54672z313_BXINV_5852 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z313_BXINV
    );
  romedatao4_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_3_F5MUX,
      O => nx54672z321
    );
  romedatao4_s_3_F5MUX_5853 : X_MUX2
    port map (
      IA => nx54672z322,
      IB => nx54672z323,
      SEL => romedatao4_s_3_BXINV,
      O => romedatao4_s_3_F5MUX
    );
  romedatao4_s_3_BXINV_5854 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao4_s_3_BXINV
    );
  romedatao4_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_3_F6MUX,
      O => romedatao4_s(3)
    );
  romedatao4_s_3_F6MUX_5855 : X_MUX2
    port map (
      IA => nx54672z319,
      IB => nx54672z321,
      SEL => romedatao4_s_3_BYINV,
      O => romedatao4_s_3_F6MUX
    );
  romedatao4_s_3_BYINV_5856 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao4_s_3_BYINV
    );
  nx54672z319_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z319_F5MUX,
      O => nx54672z319
    );
  nx54672z319_F5MUX_5857 : X_MUX2
    port map (
      IA => U1_ROME4_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx54672z320,
      SEL => nx54672z319_BXINV,
      O => nx54672z319_F5MUX
    );
  nx54672z319_BXINV_5858 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z319_BXINV
    );
  romedatao4_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_2_F5MUX,
      O => U1_ROME4_modgen_rom_ix2_nx_ro64_32_l
    );
  romedatao4_s_2_F5MUX_5859 : X_MUX2
    port map (
      IA => romedatao4_s_2_G,
      IB => nx54672z324,
      SEL => romedatao4_s_2_BXINV,
      O => romedatao4_s_2_F5MUX
    );
  romedatao4_s_2_BXINV_5860 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao4_s_2_BXINV
    );
  romedatao4_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_2_F6MUX,
      O => romedatao4_s(2)
    );
  romedatao4_s_2_F6MUX_5861 : X_MUX2
    port map (
      IA => U1_ROME4_modgen_rom_ix2_nx_ro64_32_u,
      IB => U1_ROME4_modgen_rom_ix2_nx_ro64_32_l,
      SEL => romedatao4_s_2_BYINV,
      O => romedatao4_s_2_F6MUX
    );
  romedatao4_s_2_BYINV_5862 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao4_s_2_BYINV
    );
  U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U1_ROME4_modgen_rom_ix2_nx_ro64_32_u
    );
  U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_F5MUX_5863 : X_MUX2
    port map (
      IA => U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U1_ROME4_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_BXINV_5864 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  romedatao1_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_9_F5MUX,
      O => nx54672z91
    );
  romedatao1_s_9_F5MUX_5865 : X_MUX2
    port map (
      IA => nx54672z92,
      IB => nx54672z93,
      SEL => romedatao1_s_9_BXINV,
      O => romedatao1_s_9_F5MUX
    );
  romedatao1_s_9_BXINV_5866 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao1_s_9_BXINV
    );
  romedatao1_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao1_s_9_F6MUX,
      O => romedatao1_s(9)
    );
  romedatao1_s_9_F6MUX_5867 : X_MUX2
    port map (
      IA => nx54672z88,
      IB => nx54672z91,
      SEL => romedatao1_s_9_BYINV,
      O => romedatao1_s_9_F6MUX
    );
  romedatao1_s_9_BYINV_5868 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao1_s_9_BYINV
    );
  nx54672z88_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z88_F5MUX,
      O => nx54672z88
    );
  nx54672z88_F5MUX_5869 : X_MUX2
    port map (
      IA => nx54672z89,
      IB => nx54672z90,
      SEL => nx54672z88_BXINV,
      O => nx54672z88_F5MUX
    );
  nx54672z88_BXINV_5870 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z88_BXINV
    );
  romodatao0_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_2_F5MUX,
      O => nx54672z653
    );
  romodatao0_s_2_F5MUX_5871 : X_MUX2
    port map (
      IA => nx54672z654,
      IB => nx54672z655,
      SEL => romodatao0_s_2_BXINV,
      O => romodatao0_s_2_F5MUX
    );
  romodatao0_s_2_BXINV_5872 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao0_s_2_BXINV
    );
  romodatao0_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao0_s_2_F6MUX,
      O => romodatao0_s(2)
    );
  romodatao0_s_2_F6MUX_5873 : X_MUX2
    port map (
      IA => nx54672z650,
      IB => nx54672z653,
      SEL => romodatao0_s_2_BYINV,
      O => romodatao0_s_2_F6MUX
    );
  romodatao0_s_2_BYINV_5874 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao0_s_2_BYINV
    );
  nx54672z650_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z650_F5MUX,
      O => nx54672z650
    );
  nx54672z650_F5MUX_5875 : X_MUX2
    port map (
      IA => nx54672z651,
      IB => nx54672z652,
      SEL => nx54672z650_BXINV,
      O => nx54672z650_F5MUX
    );
  nx54672z650_BXINV_5876 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z650_BXINV
    );
  romedatao6_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_12_F5MUX,
      O => nx54672z398
    );
  romedatao6_s_12_F5MUX_5877 : X_MUX2
    port map (
      IA => nx54672z399,
      IB => nx54672z400,
      SEL => romedatao6_s_12_BXINV,
      O => romedatao6_s_12_F5MUX
    );
  romedatao6_s_12_BXINV_5878 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao6_s_12_BXINV
    );
  romedatao6_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_12_F6MUX,
      O => romedatao6_s(12)
    );
  romedatao6_s_12_F6MUX_5879 : X_MUX2
    port map (
      IA => nx54672z395,
      IB => nx54672z398,
      SEL => romedatao6_s_12_BYINV,
      O => romedatao6_s_12_F6MUX
    );
  romedatao6_s_12_BYINV_5880 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao6_s_12_BYINV
    );
  nx54672z395_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z395_F5MUX,
      O => nx54672z395
    );
  nx54672z395_F5MUX_5881 : X_MUX2
    port map (
      IA => nx54672z396,
      IB => nx54672z397,
      SEL => nx54672z395_BXINV,
      O => nx54672z395_F5MUX
    );
  nx54672z395_BXINV_5882 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z395_BXINV
    );
  romedatao6_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_4_F5MUX,
      O => nx54672z446
    );
  romedatao6_s_4_F5MUX_5883 : X_MUX2
    port map (
      IA => nx54672z447,
      IB => nx54672z448,
      SEL => romedatao6_s_4_BXINV,
      O => romedatao6_s_4_F5MUX
    );
  romedatao6_s_4_BXINV_5884 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao6_s_4_BXINV
    );
  romedatao6_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_4_F6MUX,
      O => romedatao6_s(4)
    );
  romedatao6_s_4_F6MUX_5885 : X_MUX2
    port map (
      IA => nx54672z443,
      IB => nx54672z446,
      SEL => romedatao6_s_4_BYINV,
      O => romedatao6_s_4_F6MUX
    );
  romedatao6_s_4_BYINV_5886 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao6_s_4_BYINV
    );
  nx54672z443_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z443_F5MUX,
      O => nx54672z443
    );
  nx54672z443_F5MUX_5887 : X_MUX2
    port map (
      IA => nx54672z444,
      IB => nx54672z445,
      SEL => nx54672z443_BXINV,
      O => nx54672z443_F5MUX
    );
  nx54672z443_BXINV_5888 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z443_BXINV
    );
  romedatao6_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_3_F5MUX,
      O => nx54672z451
    );
  romedatao6_s_3_F5MUX_5889 : X_MUX2
    port map (
      IA => nx54672z452,
      IB => nx54672z453,
      SEL => romedatao6_s_3_BXINV,
      O => romedatao6_s_3_F5MUX
    );
  romedatao6_s_3_BXINV_5890 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao6_s_3_BXINV
    );
  romedatao6_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_3_F6MUX,
      O => romedatao6_s(3)
    );
  romedatao6_s_3_F6MUX_5891 : X_MUX2
    port map (
      IA => nx54672z449,
      IB => nx54672z451,
      SEL => romedatao6_s_3_BYINV,
      O => romedatao6_s_3_F6MUX
    );
  romedatao6_s_3_BYINV_5892 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao6_s_3_BYINV
    );
  nx54672z449_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z449_F5MUX,
      O => nx54672z449
    );
  nx54672z449_F5MUX_5893 : X_MUX2
    port map (
      IA => U1_ROME6_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx54672z450,
      SEL => nx54672z449_BXINV,
      O => nx54672z449_F5MUX
    );
  nx54672z449_BXINV_5894 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z449_BXINV
    );
  romedatao6_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_2_F5MUX,
      O => U1_ROME6_modgen_rom_ix2_nx_ro64_32_l
    );
  romedatao6_s_2_F5MUX_5895 : X_MUX2
    port map (
      IA => romedatao6_s_2_G,
      IB => nx54672z454,
      SEL => romedatao6_s_2_BXINV,
      O => romedatao6_s_2_F5MUX
    );
  romedatao6_s_2_BXINV_5896 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao6_s_2_BXINV
    );
  romedatao6_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_2_F6MUX,
      O => romedatao6_s(2)
    );
  romedatao6_s_2_F6MUX_5897 : X_MUX2
    port map (
      IA => U1_ROME6_modgen_rom_ix2_nx_ro64_32_u,
      IB => U1_ROME6_modgen_rom_ix2_nx_ro64_32_l,
      SEL => romedatao6_s_2_BYINV,
      O => romedatao6_s_2_F6MUX
    );
  romedatao6_s_2_BYINV_5898 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao6_s_2_BYINV
    );
  U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U1_ROME6_modgen_rom_ix2_nx_ro64_32_u
    );
  U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_F5MUX_5899 : X_MUX2
    port map (
      IA => U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U1_ROME6_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_BXINV_5900 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  romedatao3_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_10_F5MUX,
      O => nx54672z215
    );
  romedatao3_s_10_F5MUX_5901 : X_MUX2
    port map (
      IA => nx54672z216,
      IB => nx54672z217,
      SEL => romedatao3_s_10_BXINV,
      O => romedatao3_s_10_F5MUX
    );
  romedatao3_s_10_BXINV_5902 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao3_s_10_BXINV
    );
  romedatao3_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_10_F6MUX,
      O => romedatao3_s(10)
    );
  romedatao3_s_10_F6MUX_5903 : X_MUX2
    port map (
      IA => nx54672z212,
      IB => nx54672z215,
      SEL => romedatao3_s_10_BYINV,
      O => romedatao3_s_10_F6MUX
    );
  romedatao3_s_10_BYINV_5904 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao3_s_10_BYINV
    );
  nx54672z212_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z212_F5MUX,
      O => nx54672z212
    );
  nx54672z212_F5MUX_5905 : X_MUX2
    port map (
      IA => nx54672z213,
      IB => nx54672z214,
      SEL => nx54672z212_BXINV,
      O => nx54672z212_F5MUX
    );
  nx54672z212_BXINV_5906 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z212_BXINV
    );
  romedatao3_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_8_F5MUX,
      O => nx54672z227
    );
  romedatao3_s_8_F5MUX_5907 : X_MUX2
    port map (
      IA => nx54672z228,
      IB => nx54672z229,
      SEL => romedatao3_s_8_BXINV,
      O => romedatao3_s_8_F5MUX
    );
  romedatao3_s_8_BXINV_5908 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao3_s_8_BXINV
    );
  romedatao3_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_8_F6MUX,
      O => romedatao3_s(8)
    );
  romedatao3_s_8_F6MUX_5909 : X_MUX2
    port map (
      IA => nx54672z224,
      IB => nx54672z227,
      SEL => romedatao3_s_8_BYINV,
      O => romedatao3_s_8_F6MUX
    );
  romedatao3_s_8_BYINV_5910 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao3_s_8_BYINV
    );
  nx54672z224_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z224_F5MUX,
      O => nx54672z224
    );
  nx54672z224_F5MUX_5911 : X_MUX2
    port map (
      IA => nx54672z225,
      IB => nx54672z226,
      SEL => nx54672z224_BXINV,
      O => nx54672z224_F5MUX
    );
  nx54672z224_BXINV_5912 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z224_BXINV
    );
  romedatao5_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_12_F5MUX,
      O => nx54672z333
    );
  romedatao5_s_12_F5MUX_5913 : X_MUX2
    port map (
      IA => nx54672z334,
      IB => nx54672z335,
      SEL => romedatao5_s_12_BXINV,
      O => romedatao5_s_12_F5MUX
    );
  romedatao5_s_12_BXINV_5914 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao5_s_12_BXINV
    );
  romedatao5_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_12_F6MUX,
      O => romedatao5_s(12)
    );
  romedatao5_s_12_F6MUX_5915 : X_MUX2
    port map (
      IA => nx54672z330,
      IB => nx54672z333,
      SEL => romedatao5_s_12_BYINV,
      O => romedatao5_s_12_F6MUX
    );
  romedatao5_s_12_BYINV_5916 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao5_s_12_BYINV
    );
  nx54672z330_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z330_F5MUX,
      O => nx54672z330
    );
  nx54672z330_F5MUX_5917 : X_MUX2
    port map (
      IA => nx54672z331,
      IB => nx54672z332,
      SEL => nx54672z330_BXINV,
      O => nx54672z330_F5MUX
    );
  nx54672z330_BXINV_5918 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z330_BXINV
    );
  romedatao5_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_11_F5MUX,
      O => nx54672z339
    );
  romedatao5_s_11_F5MUX_5919 : X_MUX2
    port map (
      IA => nx54672z340,
      IB => nx54672z341,
      SEL => romedatao5_s_11_BXINV,
      O => romedatao5_s_11_F5MUX
    );
  romedatao5_s_11_BXINV_5920 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao5_s_11_BXINV
    );
  romedatao5_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_11_F6MUX,
      O => romedatao5_s(11)
    );
  romedatao5_s_11_F6MUX_5921 : X_MUX2
    port map (
      IA => nx54672z336,
      IB => nx54672z339,
      SEL => romedatao5_s_11_BYINV,
      O => romedatao5_s_11_F6MUX
    );
  romedatao5_s_11_BYINV_5922 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao5_s_11_BYINV
    );
  nx54672z336_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z336_F5MUX,
      O => nx54672z336
    );
  nx54672z336_F5MUX_5923 : X_MUX2
    port map (
      IA => nx54672z337,
      IB => nx54672z338,
      SEL => nx54672z336_BXINV,
      O => nx54672z336_F5MUX
    );
  nx54672z336_BXINV_5924 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z336_BXINV
    );
  romedatao5_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_10_F5MUX,
      O => nx54672z345
    );
  romedatao5_s_10_F5MUX_5925 : X_MUX2
    port map (
      IA => nx54672z346,
      IB => nx54672z347,
      SEL => romedatao5_s_10_BXINV,
      O => romedatao5_s_10_F5MUX
    );
  romedatao5_s_10_BXINV_5926 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao5_s_10_BXINV
    );
  romedatao5_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_10_F6MUX,
      O => romedatao5_s(10)
    );
  romedatao5_s_10_F6MUX_5927 : X_MUX2
    port map (
      IA => nx54672z342,
      IB => nx54672z345,
      SEL => romedatao5_s_10_BYINV,
      O => romedatao5_s_10_F6MUX
    );
  romedatao5_s_10_BYINV_5928 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao5_s_10_BYINV
    );
  nx54672z342_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z342_F5MUX,
      O => nx54672z342
    );
  nx54672z342_F5MUX_5929 : X_MUX2
    port map (
      IA => nx54672z343,
      IB => nx54672z344,
      SEL => nx54672z342_BXINV,
      O => nx54672z342_F5MUX
    );
  nx54672z342_BXINV_5930 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z342_BXINV
    );
  romedatao5_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_9_F5MUX,
      O => nx54672z351
    );
  romedatao5_s_9_F5MUX_5931 : X_MUX2
    port map (
      IA => nx54672z352,
      IB => nx54672z353,
      SEL => romedatao5_s_9_BXINV,
      O => romedatao5_s_9_F5MUX
    );
  romedatao5_s_9_BXINV_5932 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao5_s_9_BXINV
    );
  romedatao5_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_9_F6MUX,
      O => romedatao5_s(9)
    );
  romedatao5_s_9_F6MUX_5933 : X_MUX2
    port map (
      IA => nx54672z348,
      IB => nx54672z351,
      SEL => romedatao5_s_9_BYINV,
      O => romedatao5_s_9_F6MUX
    );
  romedatao5_s_9_BYINV_5934 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao5_s_9_BYINV
    );
  U_DCT2D_reg_databuf_reg_7_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_7_2_DYMUX,
      CE => U_DCT2D_databuf_reg_7_2_CEINV,
      CLK => U_DCT2D_databuf_reg_7_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_7_2_FFY_RST,
      O => U_DCT2D_databuf_reg_7_Q(3)
    );
  U_DCT2D_databuf_reg_7_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_7_2_FFY_RST
    );
  nx54672z348_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z348_F5MUX,
      O => nx54672z348
    );
  nx54672z348_F5MUX_5935 : X_MUX2
    port map (
      IA => nx54672z349,
      IB => nx54672z350,
      SEL => nx54672z348_BXINV,
      O => nx54672z348_F5MUX
    );
  nx54672z348_BXINV_5936 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z348_BXINV
    );
  romedatao5_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_3_F5MUX,
      O => nx54672z386
    );
  romedatao5_s_3_F5MUX_5937 : X_MUX2
    port map (
      IA => nx54672z387,
      IB => nx54672z388,
      SEL => romedatao5_s_3_BXINV,
      O => romedatao5_s_3_F5MUX
    );
  romedatao5_s_3_BXINV_5938 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao5_s_3_BXINV
    );
  romedatao5_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_3_F6MUX,
      O => romedatao5_s(3)
    );
  romedatao5_s_3_F6MUX_5939 : X_MUX2
    port map (
      IA => nx54672z384,
      IB => nx54672z386,
      SEL => romedatao5_s_3_BYINV,
      O => romedatao5_s_3_F6MUX
    );
  romedatao5_s_3_BYINV_5940 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao5_s_3_BYINV
    );
  nx54672z384_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z384_F5MUX,
      O => nx54672z384
    );
  nx54672z384_F5MUX_5941 : X_MUX2
    port map (
      IA => U1_ROME5_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx54672z385,
      SEL => nx54672z384_BXINV,
      O => nx54672z384_F5MUX
    );
  nx54672z384_BXINV_5942 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z384_BXINV
    );
  romedatao5_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_2_F5MUX,
      O => U1_ROME5_modgen_rom_ix2_nx_ro64_32_l
    );
  romedatao5_s_2_F5MUX_5943 : X_MUX2
    port map (
      IA => romedatao5_s_2_G,
      IB => nx54672z389,
      SEL => romedatao5_s_2_BXINV,
      O => romedatao5_s_2_F5MUX
    );
  romedatao5_s_2_BXINV_5944 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao5_s_2_BXINV
    );
  romedatao5_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_2_F6MUX,
      O => romedatao5_s(2)
    );
  romedatao5_s_2_F6MUX_5945 : X_MUX2
    port map (
      IA => U1_ROME5_modgen_rom_ix2_nx_ro64_32_u,
      IB => U1_ROME5_modgen_rom_ix2_nx_ro64_32_l,
      SEL => romedatao5_s_2_BYINV,
      O => romedatao5_s_2_F6MUX
    );
  romedatao5_s_2_BYINV_5946 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao5_s_2_BYINV
    );
  U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U1_ROME5_modgen_rom_ix2_nx_ro64_32_u
    );
  U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_F5MUX_5947 : X_MUX2
    port map (
      IA => U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U1_ROME5_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_BXINV_5948 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  romodatao6_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_9_F5MUX,
      O => nx54672z1083
    );
  romodatao6_s_9_F5MUX_5949 : X_MUX2
    port map (
      IA => nx54672z1084,
      IB => nx54672z1085,
      SEL => romodatao6_s_9_BXINV,
      O => romodatao6_s_9_F5MUX
    );
  romodatao6_s_9_BXINV_5950 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_9_BXINV
    );
  romodatao6_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_9_F6MUX,
      O => romodatao6_s(9)
    );
  romodatao6_s_9_F6MUX_5951 : X_MUX2
    port map (
      IA => nx54672z1080,
      IB => nx54672z1083,
      SEL => romodatao6_s_9_BYINV,
      O => romodatao6_s_9_F6MUX
    );
  romodatao6_s_9_BYINV_5952 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_9_BYINV
    );
  ix54672z23666 : X_LUT4
    generic map(
      INIT => X"4564"
    )
    port map (
      ADR0 => romoaddro6_s(0),
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1081
    );
  nx54672z1080_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1080_F5MUX,
      O => nx54672z1080
    );
  nx54672z1080_F5MUX_5953 : X_MUX2
    port map (
      IA => nx54672z1081,
      IB => nx54672z1082,
      SEL => nx54672z1080_BXINV,
      O => nx54672z1080_F5MUX
    );
  nx54672z1080_BXINV_5954 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1080_BXINV
    );
  romodatao6_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_8_F5MUX,
      O => nx54672z1089
    );
  romodatao6_s_8_F5MUX_5955 : X_MUX2
    port map (
      IA => nx54672z1090,
      IB => nx54672z1091,
      SEL => romodatao6_s_8_BXINV,
      O => romodatao6_s_8_F5MUX
    );
  romodatao6_s_8_BXINV_5956 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_8_BXINV
    );
  romodatao6_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_8_F6MUX,
      O => romodatao6_s(8)
    );
  romodatao6_s_8_F6MUX_5957 : X_MUX2
    port map (
      IA => nx54672z1086,
      IB => nx54672z1089,
      SEL => romodatao6_s_8_BYINV,
      O => romodatao6_s_8_F6MUX
    );
  romodatao6_s_8_BYINV_5958 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_8_BYINV
    );
  nx54672z1086_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1086_F5MUX,
      O => nx54672z1086
    );
  nx54672z1086_F5MUX_5959 : X_MUX2
    port map (
      IA => nx54672z1087,
      IB => nx54672z1088,
      SEL => nx54672z1086_BXINV,
      O => nx54672z1086_F5MUX
    );
  nx54672z1086_BXINV_5960 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1086_BXINV
    );
  romodatao6_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_7_F5MUX,
      O => nx54672z1095
    );
  romodatao6_s_7_F5MUX_5961 : X_MUX2
    port map (
      IA => nx54672z1096,
      IB => nx54672z1097,
      SEL => romodatao6_s_7_BXINV,
      O => romodatao6_s_7_F5MUX
    );
  romodatao6_s_7_BXINV_5962 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_7_BXINV
    );
  romodatao6_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_7_F6MUX,
      O => romodatao6_s(7)
    );
  romodatao6_s_7_F6MUX_5963 : X_MUX2
    port map (
      IA => nx54672z1092,
      IB => nx54672z1095,
      SEL => romodatao6_s_7_BYINV,
      O => romodatao6_s_7_F6MUX
    );
  romodatao6_s_7_BYINV_5964 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_7_BYINV
    );
  U_DCT2D_ix36141z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_3_2_Q,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_4_2_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx36141z1
    );
  nx54672z1092_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1092_F5MUX,
      O => nx54672z1092
    );
  nx54672z1092_F5MUX_5965 : X_MUX2
    port map (
      IA => nx54672z1093,
      IB => nx54672z1094,
      SEL => nx54672z1092_BXINV,
      O => nx54672z1092_F5MUX
    );
  nx54672z1092_BXINV_5966 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1092_BXINV
    );
  romodatao5_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_7_F5MUX,
      O => nx54672z1016
    );
  romodatao5_s_7_F5MUX_5967 : X_MUX2
    port map (
      IA => nx54672z1017,
      IB => nx54672z1018,
      SEL => romodatao5_s_7_BXINV,
      O => romodatao5_s_7_F5MUX
    );
  romodatao5_s_7_BXINV_5968 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_7_BXINV
    );
  romodatao5_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_7_F6MUX,
      O => romodatao5_s(7)
    );
  romodatao5_s_7_F6MUX_5969 : X_MUX2
    port map (
      IA => nx54672z1013,
      IB => nx54672z1016,
      SEL => romodatao5_s_7_BYINV,
      O => romodatao5_s_7_F6MUX
    );
  romodatao5_s_7_BYINV_5970 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_7_BYINV
    );
  nx54672z1013_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1013_F5MUX,
      O => nx54672z1013
    );
  nx54672z1013_F5MUX_5971 : X_MUX2
    port map (
      IA => nx54672z1014,
      IB => nx54672z1015,
      SEL => nx54672z1013_BXINV,
      O => nx54672z1013_F5MUX
    );
  nx54672z1013_BXINV_5972 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1013_BXINV
    );
  romodatao5_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_6_F5MUX,
      O => nx54672z1022
    );
  romodatao5_s_6_F5MUX_5973 : X_MUX2
    port map (
      IA => nx54672z1023,
      IB => nx54672z1024,
      SEL => romodatao5_s_6_BXINV,
      O => romodatao5_s_6_F5MUX
    );
  romodatao5_s_6_BXINV_5974 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_6_BXINV
    );
  romodatao5_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_6_F6MUX,
      O => romodatao5_s(6)
    );
  romodatao5_s_6_F6MUX_5975 : X_MUX2
    port map (
      IA => nx54672z1019,
      IB => nx54672z1022,
      SEL => romodatao5_s_6_BYINV,
      O => romodatao5_s_6_F6MUX
    );
  romodatao5_s_6_BYINV_5976 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_6_BYINV
    );
  nx54672z1019_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1019_F5MUX,
      O => nx54672z1019
    );
  nx54672z1019_F5MUX_5977 : X_MUX2
    port map (
      IA => nx54672z1020,
      IB => nx54672z1021,
      SEL => nx54672z1019_BXINV,
      O => nx54672z1019_F5MUX
    );
  nx54672z1019_BXINV_5978 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1019_BXINV
    );
  romodatao5_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_5_F5MUX,
      O => nx54672z1028
    );
  romodatao5_s_5_F5MUX_5979 : X_MUX2
    port map (
      IA => nx54672z1029,
      IB => nx54672z1030,
      SEL => romodatao5_s_5_BXINV,
      O => romodatao5_s_5_F5MUX
    );
  romodatao5_s_5_BXINV_5980 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_5_BXINV
    );
  romodatao5_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_5_F6MUX,
      O => romodatao5_s(5)
    );
  romodatao5_s_5_F6MUX_5981 : X_MUX2
    port map (
      IA => nx54672z1025,
      IB => nx54672z1028,
      SEL => romodatao5_s_5_BYINV,
      O => romodatao5_s_5_F6MUX
    );
  romodatao5_s_5_BYINV_5982 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_5_BYINV
    );
  nx54672z1025_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1025_F5MUX,
      O => nx54672z1025
    );
  nx54672z1025_F5MUX_5983 : X_MUX2
    port map (
      IA => nx54672z1026,
      IB => nx54672z1027,
      SEL => nx54672z1025_BXINV,
      O => nx54672z1025_F5MUX
    );
  nx54672z1025_BXINV_5984 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1025_BXINV
    );
  romodatao5_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_4_F5MUX,
      O => nx54672z1034
    );
  romodatao5_s_4_F5MUX_5985 : X_MUX2
    port map (
      IA => nx54672z1035,
      IB => nx54672z1036,
      SEL => romodatao5_s_4_BXINV,
      O => romodatao5_s_4_F5MUX
    );
  romodatao5_s_4_BXINV_5986 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_4_BXINV
    );
  romodatao5_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_4_F6MUX,
      O => romodatao5_s(4)
    );
  romodatao5_s_4_F6MUX_5987 : X_MUX2
    port map (
      IA => nx54672z1031,
      IB => nx54672z1034,
      SEL => romodatao5_s_4_BYINV,
      O => romodatao5_s_4_F6MUX
    );
  romodatao5_s_4_BYINV_5988 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_4_BYINV
    );
  nx54672z1031_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1031_F5MUX,
      O => nx54672z1031
    );
  nx54672z1031_F5MUX_5989 : X_MUX2
    port map (
      IA => nx54672z1032,
      IB => nx54672z1033,
      SEL => nx54672z1031_BXINV,
      O => nx54672z1031_F5MUX
    );
  nx54672z1031_BXINV_5990 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1031_BXINV
    );
  romodatao5_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_3_F5MUX,
      O => nx54672z1040
    );
  romodatao5_s_3_F5MUX_5991 : X_MUX2
    port map (
      IA => nx54672z1041,
      IB => nx54672z1042,
      SEL => romodatao5_s_3_BXINV,
      O => romodatao5_s_3_F5MUX
    );
  romodatao5_s_3_BXINV_5992 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_3_BXINV
    );
  romodatao5_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_3_F6MUX,
      O => romodatao5_s(3)
    );
  romodatao5_s_3_F6MUX_5993 : X_MUX2
    port map (
      IA => nx54672z1037,
      IB => nx54672z1040,
      SEL => romodatao5_s_3_BYINV,
      O => romodatao5_s_3_F6MUX
    );
  romodatao5_s_3_BYINV_5994 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_3_BYINV
    );
  nx54672z1037_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1037_F5MUX,
      O => nx54672z1037
    );
  nx54672z1037_F5MUX_5995 : X_MUX2
    port map (
      IA => nx54672z1038,
      IB => nx54672z1039,
      SEL => nx54672z1037_BXINV,
      O => nx54672z1037_F5MUX
    );
  nx54672z1037_BXINV_5996 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1037_BXINV
    );
  romodatao5_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_13_F5MUX,
      O => nx54672z980
    );
  romodatao5_s_13_F5MUX_5997 : X_MUX2
    port map (
      IA => nx54672z981,
      IB => nx54672z982,
      SEL => romodatao5_s_13_BXINV,
      O => romodatao5_s_13_F5MUX
    );
  romodatao5_s_13_BXINV_5998 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_13_BXINV
    );
  romodatao5_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_13_F6MUX,
      O => romodatao5_s(13)
    );
  romodatao5_s_13_F6MUX_5999 : X_MUX2
    port map (
      IA => nx54672z978,
      IB => nx54672z980,
      SEL => romodatao5_s_13_BYINV,
      O => romodatao5_s_13_F6MUX
    );
  romodatao5_s_13_BYINV_6000 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_13_BYINV
    );
  nx54672z978_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z978_F5MUX,
      O => nx54672z978
    );
  nx54672z978_F5MUX_6001 : X_MUX2
    port map (
      IA => nx54672z978_G,
      IB => nx54672z979,
      SEL => nx54672z978_BXINV,
      O => nx54672z978_F5MUX
    );
  nx54672z978_BXINV_6002 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z978_BXINV
    );
  romodatao4_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_12_F5MUX,
      O => nx54672z907
    );
  romodatao4_s_12_F5MUX_6003 : X_MUX2
    port map (
      IA => nx54672z908,
      IB => nx54672z909,
      SEL => romodatao4_s_12_BXINV,
      O => romodatao4_s_12_F5MUX
    );
  romodatao4_s_12_BXINV_6004 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_12_BXINV
    );
  romodatao4_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_12_F6MUX,
      O => romodatao4_s(12)
    );
  romodatao4_s_12_F6MUX_6005 : X_MUX2
    port map (
      IA => nx54672z904,
      IB => nx54672z907,
      SEL => romodatao4_s_12_BYINV,
      O => romodatao4_s_12_F6MUX
    );
  romodatao4_s_12_BYINV_6006 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_12_BYINV
    );
  nx54672z904_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z904_F5MUX,
      O => nx54672z904
    );
  nx54672z904_F5MUX_6007 : X_MUX2
    port map (
      IA => nx54672z905,
      IB => nx54672z906,
      SEL => nx54672z904_BXINV,
      O => nx54672z904_F5MUX
    );
  nx54672z904_BXINV_6008 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z904_BXINV
    );
  romodatao4_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_10_F5MUX,
      O => nx54672z919
    );
  romodatao4_s_10_F5MUX_6009 : X_MUX2
    port map (
      IA => nx54672z920,
      IB => nx54672z921,
      SEL => romodatao4_s_10_BXINV,
      O => romodatao4_s_10_F5MUX
    );
  romodatao4_s_10_BXINV_6010 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_10_BXINV
    );
  romodatao4_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_10_F6MUX,
      O => romodatao4_s(10)
    );
  romodatao4_s_10_F6MUX_6011 : X_MUX2
    port map (
      IA => nx54672z916,
      IB => nx54672z919,
      SEL => romodatao4_s_10_BYINV,
      O => romodatao4_s_10_F6MUX
    );
  romodatao4_s_10_BYINV_6012 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_10_BYINV
    );
  nx54672z916_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z916_F5MUX,
      O => nx54672z916
    );
  nx54672z916_F5MUX_6013 : X_MUX2
    port map (
      IA => nx54672z917,
      IB => nx54672z918,
      SEL => nx54672z916_BXINV,
      O => nx54672z916_F5MUX
    );
  nx54672z916_BXINV_6014 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z916_BXINV
    );
  romodatao4_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_9_F5MUX,
      O => nx54672z925
    );
  romodatao4_s_9_F5MUX_6015 : X_MUX2
    port map (
      IA => nx54672z926,
      IB => nx54672z927,
      SEL => romodatao4_s_9_BXINV,
      O => romodatao4_s_9_F5MUX
    );
  romodatao4_s_9_BXINV_6016 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_9_BXINV
    );
  romodatao4_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_9_F6MUX,
      O => romodatao4_s(9)
    );
  romodatao4_s_9_F6MUX_6017 : X_MUX2
    port map (
      IA => nx54672z922,
      IB => nx54672z925,
      SEL => romodatao4_s_9_BYINV,
      O => romodatao4_s_9_F6MUX
    );
  romodatao4_s_9_BYINV_6018 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_9_BYINV
    );
  nx54672z922_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z922_F5MUX,
      O => nx54672z922
    );
  nx54672z922_F5MUX_6019 : X_MUX2
    port map (
      IA => nx54672z923,
      IB => nx54672z924,
      SEL => nx54672z922_BXINV,
      O => nx54672z922_F5MUX
    );
  nx54672z922_BXINV_6020 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z922_BXINV
    );
  romodatao4_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_3_F5MUX,
      O => nx54672z961
    );
  romodatao4_s_3_F5MUX_6021 : X_MUX2
    port map (
      IA => nx54672z962,
      IB => nx54672z963,
      SEL => romodatao4_s_3_BXINV,
      O => romodatao4_s_3_F5MUX
    );
  romodatao4_s_3_BXINV_6022 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_3_BXINV
    );
  romodatao4_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_3_F6MUX,
      O => romodatao4_s(3)
    );
  romodatao4_s_3_F6MUX_6023 : X_MUX2
    port map (
      IA => nx54672z958,
      IB => nx54672z961,
      SEL => romodatao4_s_3_BYINV,
      O => romodatao4_s_3_F6MUX
    );
  romodatao4_s_3_BYINV_6024 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_3_BYINV
    );
  U_DCT2D_reg_databuf_reg_7_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_7_2_DXMUX,
      CE => U_DCT2D_databuf_reg_7_2_CEINV,
      CLK => U_DCT2D_databuf_reg_7_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_7_2_FFX_RST,
      O => U_DCT2D_databuf_reg_7_Q(2)
    );
  U_DCT2D_databuf_reg_7_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_7_2_FFX_RST
    );
  nx54672z958_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z958_F5MUX,
      O => nx54672z958
    );
  nx54672z958_F5MUX_6025 : X_MUX2
    port map (
      IA => nx54672z959,
      IB => nx54672z960,
      SEL => nx54672z958_BXINV,
      O => nx54672z958_F5MUX
    );
  nx54672z958_BXINV_6026 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z958_BXINV
    );
  romodatao4_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_2_F5MUX,
      O => nx54672z967
    );
  romodatao4_s_2_F5MUX_6027 : X_MUX2
    port map (
      IA => nx54672z968,
      IB => nx54672z969,
      SEL => romodatao4_s_2_BXINV,
      O => romodatao4_s_2_F5MUX
    );
  romodatao4_s_2_BXINV_6028 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_2_BXINV
    );
  romodatao4_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_2_F6MUX,
      O => romodatao4_s(2)
    );
  romodatao4_s_2_F6MUX_6029 : X_MUX2
    port map (
      IA => nx54672z964,
      IB => nx54672z967,
      SEL => romodatao4_s_2_BYINV,
      O => romodatao4_s_2_F6MUX
    );
  romodatao4_s_2_BYINV_6030 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_2_BYINV
    );
  nx54672z964_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z964_F5MUX,
      O => nx54672z964
    );
  nx54672z964_F5MUX_6031 : X_MUX2
    port map (
      IA => nx54672z965,
      IB => nx54672z966,
      SEL => nx54672z964_BXINV,
      O => nx54672z964_F5MUX
    );
  nx54672z964_BXINV_6032 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z964_BXINV
    );
  U_DCT2D_ix39132z1324 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_3_5_Q,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_4_5_Q,
      O => U_DCT2D_nx39132z1
    );
  romodatao4_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_1_F5MUX,
      O => nx54672z973
    );
  romodatao4_s_1_F5MUX_6033 : X_MUX2
    port map (
      IA => nx54672z974,
      IB => nx54672z975,
      SEL => romodatao4_s_1_BXINV,
      O => romodatao4_s_1_F5MUX
    );
  romodatao4_s_1_BXINV_6034 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_1_BXINV
    );
  romodatao4_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_1_F6MUX,
      O => romodatao4_s(1)
    );
  romodatao4_s_1_F6MUX_6035 : X_MUX2
    port map (
      IA => nx54672z970,
      IB => nx54672z973,
      SEL => romodatao4_s_1_BYINV,
      O => romodatao4_s_1_F6MUX
    );
  romodatao4_s_1_BYINV_6036 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_1_BYINV
    );
  nx54672z970_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z970_F5MUX,
      O => nx54672z970
    );
  nx54672z970_F5MUX_6037 : X_MUX2
    port map (
      IA => nx54672z971,
      IB => nx54672z972,
      SEL => nx54672z970_BXINV,
      O => nx54672z970_F5MUX
    );
  nx54672z970_BXINV_6038 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z970_BXINV
    );
  romodatao4_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_0_F5MUX,
      O => U1_ROMO4_modgen_rom_ix0_nx_ro64_32_l
    );
  romodatao4_s_0_F5MUX_6039 : X_MUX2
    port map (
      IA => nx54672z976,
      IB => nx54672z977,
      SEL => romodatao4_s_0_BXINV,
      O => romodatao4_s_0_F5MUX
    );
  romodatao4_s_0_BXINV_6040 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_0_BXINV
    );
  romodatao4_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_0_F6MUX,
      O => romodatao4_s(0)
    );
  romodatao4_s_0_F6MUX_6041 : X_MUX2
    port map (
      IA => U1_ROMO4_modgen_rom_ix0_nx_ro64_32_u,
      IB => U1_ROMO4_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romodatao4_s_0_BYINV,
      O => romodatao4_s_0_F6MUX
    );
  romodatao4_s_0_BYINV_6042 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_0_BYINV
    );
  U1_ROMO4_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROMO4_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U1_ROMO4_modgen_rom_ix0_nx_ro64_32_u
    );
  U1_ROMO4_modgen_rom_ix0_nx_ro64_32_u_F5MUX_6043 : X_MUX2
    port map (
      IA => U1_ROMO4_modgen_rom_ix0_nx_rm64_16_u,
      IB => U1_ROMO4_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U1_ROMO4_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U1_ROMO4_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U1_ROMO4_modgen_rom_ix0_nx_ro64_32_u_BXINV_6044 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => U1_ROMO4_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romodatao3_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_8_F5MUX,
      O => nx54672z852
    );
  romodatao3_s_8_F5MUX_6045 : X_MUX2
    port map (
      IA => nx54672z853,
      IB => nx54672z854,
      SEL => romodatao3_s_8_BXINV,
      O => romodatao3_s_8_F5MUX
    );
  romodatao3_s_8_BXINV_6046 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_8_BXINV
    );
  romodatao3_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_8_F6MUX,
      O => romodatao3_s(8)
    );
  romodatao3_s_8_F6MUX_6047 : X_MUX2
    port map (
      IA => nx54672z849,
      IB => nx54672z852,
      SEL => romodatao3_s_8_BYINV,
      O => romodatao3_s_8_F6MUX
    );
  romodatao3_s_8_BYINV_6048 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_8_BYINV
    );
  nx54672z849_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z849_F5MUX,
      O => nx54672z849
    );
  nx54672z849_F5MUX_6049 : X_MUX2
    port map (
      IA => nx54672z850,
      IB => nx54672z851,
      SEL => nx54672z849_BXINV,
      O => nx54672z849_F5MUX
    );
  nx54672z849_BXINV_6050 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z849_BXINV
    );
  romodatao3_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_6_F5MUX,
      O => nx54672z864
    );
  romodatao3_s_6_F5MUX_6051 : X_MUX2
    port map (
      IA => nx54672z865,
      IB => nx54672z866,
      SEL => romodatao3_s_6_BXINV,
      O => romodatao3_s_6_F5MUX
    );
  romodatao3_s_6_BXINV_6052 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_6_BXINV
    );
  romodatao3_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_6_F6MUX,
      O => romodatao3_s(6)
    );
  romodatao3_s_6_F6MUX_6053 : X_MUX2
    port map (
      IA => nx54672z861,
      IB => nx54672z864,
      SEL => romodatao3_s_6_BYINV,
      O => romodatao3_s_6_F6MUX
    );
  romodatao3_s_6_BYINV_6054 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_6_BYINV
    );
  nx54672z861_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z861_F5MUX,
      O => nx54672z861
    );
  nx54672z861_F5MUX_6055 : X_MUX2
    port map (
      IA => nx54672z862,
      IB => nx54672z863,
      SEL => nx54672z861_BXINV,
      O => nx54672z861_F5MUX
    );
  nx54672z861_BXINV_6056 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z861_BXINV
    );
  romodatao2_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_5_F5MUX,
      O => nx54672z791
    );
  romodatao2_s_5_F5MUX_6057 : X_MUX2
    port map (
      IA => nx54672z792,
      IB => nx54672z793,
      SEL => romodatao2_s_5_BXINV,
      O => romodatao2_s_5_F5MUX
    );
  romodatao2_s_5_BXINV_6058 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_5_BXINV
    );
  romodatao2_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_5_F6MUX,
      O => romodatao2_s(5)
    );
  romodatao2_s_5_F6MUX_6059 : X_MUX2
    port map (
      IA => nx54672z788,
      IB => nx54672z791,
      SEL => romodatao2_s_5_BYINV,
      O => romodatao2_s_5_F6MUX
    );
  romodatao2_s_5_BYINV_6060 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_5_BYINV
    );
  nx54672z788_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z788_F5MUX,
      O => nx54672z788
    );
  nx54672z788_F5MUX_6061 : X_MUX2
    port map (
      IA => nx54672z789,
      IB => nx54672z790,
      SEL => nx54672z788_BXINV,
      O => nx54672z788_F5MUX
    );
  nx54672z788_BXINV_6062 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z788_BXINV
    );
  romodatao2_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_4_F5MUX,
      O => nx54672z797
    );
  romodatao2_s_4_F5MUX_6063 : X_MUX2
    port map (
      IA => nx54672z798,
      IB => nx54672z799,
      SEL => romodatao2_s_4_BXINV,
      O => romodatao2_s_4_F5MUX
    );
  romodatao2_s_4_BXINV_6064 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_4_BXINV
    );
  romodatao2_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_4_F6MUX,
      O => romodatao2_s(4)
    );
  romodatao2_s_4_F6MUX_6065 : X_MUX2
    port map (
      IA => nx54672z794,
      IB => nx54672z797,
      SEL => romodatao2_s_4_BYINV,
      O => romodatao2_s_4_F6MUX
    );
  romodatao2_s_4_BYINV_6066 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_4_BYINV
    );
  nx54672z794_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z794_F5MUX,
      O => nx54672z794
    );
  nx54672z794_F5MUX_6067 : X_MUX2
    port map (
      IA => nx54672z795,
      IB => nx54672z796,
      SEL => nx54672z794_BXINV,
      O => nx54672z794_F5MUX
    );
  nx54672z794_BXINV_6068 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z794_BXINV
    );
  romedatao7_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_12_F5MUX,
      O => nx54672z463
    );
  romedatao7_s_12_F5MUX_6069 : X_MUX2
    port map (
      IA => nx54672z464,
      IB => nx54672z465,
      SEL => romedatao7_s_12_BXINV,
      O => romedatao7_s_12_F5MUX
    );
  romedatao7_s_12_BXINV_6070 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao7_s_12_BXINV
    );
  romedatao7_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_12_F6MUX,
      O => romedatao7_s(12)
    );
  romedatao7_s_12_F6MUX_6071 : X_MUX2
    port map (
      IA => nx54672z460,
      IB => nx54672z463,
      SEL => romedatao7_s_12_BYINV,
      O => romedatao7_s_12_F6MUX
    );
  romedatao7_s_12_BYINV_6072 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao7_s_12_BYINV
    );
  ix54672z61491 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => romeaddro7_s(0),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(2),
      ADR3 => romeaddro7_s(1),
      O => nx54672z461
    );
  nx54672z460_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z460_F5MUX,
      O => nx54672z460
    );
  nx54672z460_F5MUX_6073 : X_MUX2
    port map (
      IA => nx54672z461,
      IB => nx54672z462,
      SEL => nx54672z460_BXINV,
      O => nx54672z460_F5MUX
    );
  nx54672z460_BXINV_6074 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z460_BXINV
    );
  romedatao7_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_11_F5MUX,
      O => nx54672z469
    );
  romedatao7_s_11_F5MUX_6075 : X_MUX2
    port map (
      IA => nx54672z470,
      IB => nx54672z471,
      SEL => romedatao7_s_11_BXINV,
      O => romedatao7_s_11_F5MUX
    );
  romedatao7_s_11_BXINV_6076 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao7_s_11_BXINV
    );
  romedatao7_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_11_F6MUX,
      O => romedatao7_s(11)
    );
  romedatao7_s_11_F6MUX_6077 : X_MUX2
    port map (
      IA => nx54672z466,
      IB => nx54672z469,
      SEL => romedatao7_s_11_BYINV,
      O => romedatao7_s_11_F6MUX
    );
  romedatao7_s_11_BYINV_6078 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao7_s_11_BYINV
    );
  nx54672z466_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z466_F5MUX,
      O => nx54672z466
    );
  nx54672z466_F5MUX_6079 : X_MUX2
    port map (
      IA => nx54672z467,
      IB => nx54672z468,
      SEL => nx54672z466_BXINV,
      O => nx54672z466_F5MUX
    );
  nx54672z466_BXINV_6080 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z466_BXINV
    );
  romedatao7_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_3_F5MUX,
      O => nx54672z516
    );
  romedatao7_s_3_F5MUX_6081 : X_MUX2
    port map (
      IA => nx54672z517,
      IB => nx54672z518,
      SEL => romedatao7_s_3_BXINV,
      O => romedatao7_s_3_F5MUX
    );
  romedatao7_s_3_BXINV_6082 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao7_s_3_BXINV
    );
  romedatao7_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_3_F6MUX,
      O => romedatao7_s(3)
    );
  romedatao7_s_3_F6MUX_6083 : X_MUX2
    port map (
      IA => nx54672z514,
      IB => nx54672z516,
      SEL => romedatao7_s_3_BYINV,
      O => romedatao7_s_3_F6MUX
    );
  romedatao7_s_3_BYINV_6084 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao7_s_3_BYINV
    );
  nx54672z514_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z514_F5MUX,
      O => nx54672z514
    );
  nx54672z514_F5MUX_6085 : X_MUX2
    port map (
      IA => U1_ROME7_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx54672z515,
      SEL => nx54672z514_BXINV,
      O => nx54672z514_F5MUX
    );
  nx54672z514_BXINV_6086 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z514_BXINV
    );
  romedatao7_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_2_F5MUX,
      O => U1_ROME7_modgen_rom_ix2_nx_ro64_32_l
    );
  romedatao7_s_2_F5MUX_6087 : X_MUX2
    port map (
      IA => romedatao7_s_2_G,
      IB => nx54672z519,
      SEL => romedatao7_s_2_BXINV,
      O => romedatao7_s_2_F5MUX
    );
  romedatao7_s_2_BXINV_6088 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao7_s_2_BXINV
    );
  romedatao7_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_2_F6MUX,
      O => romedatao7_s(2)
    );
  romedatao7_s_2_F6MUX_6089 : X_MUX2
    port map (
      IA => U1_ROME7_modgen_rom_ix2_nx_ro64_32_u,
      IB => U1_ROME7_modgen_rom_ix2_nx_ro64_32_l,
      SEL => romedatao7_s_2_BYINV,
      O => romedatao7_s_2_F6MUX
    );
  romedatao7_s_2_BYINV_6090 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao7_s_2_BYINV
    );
  U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_F5MUX,
      O => U1_ROME7_modgen_rom_ix2_nx_ro64_32_u
    );
  U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_F5MUX_6091 : X_MUX2
    port map (
      IA => U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_G,
      IB => U1_ROME7_modgen_rom_ix2_nx_rm64_16_l,
      SEL => U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_BXINV,
      O => U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_F5MUX
    );
  U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_BXINV_6092 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_BXINV
    );
  romodatao7_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_11_F5MUX,
      O => nx54672z1150
    );
  romodatao7_s_11_F5MUX_6093 : X_MUX2
    port map (
      IA => nx54672z1151,
      IB => nx54672z1152,
      SEL => romodatao7_s_11_BXINV,
      O => romodatao7_s_11_F5MUX
    );
  romodatao7_s_11_BXINV_6094 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_11_BXINV
    );
  romodatao7_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_11_F6MUX,
      O => romodatao7_s(11)
    );
  romodatao7_s_11_F6MUX_6095 : X_MUX2
    port map (
      IA => nx54672z1147,
      IB => nx54672z1150,
      SEL => romodatao7_s_11_BYINV,
      O => romodatao7_s_11_F6MUX
    );
  romodatao7_s_11_BYINV_6096 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_11_BYINV
    );
  ix54672z10844 : X_LUT4
    generic map(
      INIT => X"56A8"
    )
    port map (
      ADR0 => romoaddro7_s(2),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1148
    );
  nx54672z1147_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1147_F5MUX,
      O => nx54672z1147
    );
  nx54672z1147_F5MUX_6097 : X_MUX2
    port map (
      IA => nx54672z1148,
      IB => nx54672z1149,
      SEL => nx54672z1147_BXINV,
      O => nx54672z1147_F5MUX
    );
  nx54672z1147_BXINV_6098 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1147_BXINV
    );
  romodatao7_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_10_F5MUX,
      O => nx54672z1156
    );
  romodatao7_s_10_F5MUX_6099 : X_MUX2
    port map (
      IA => nx54672z1157,
      IB => nx54672z1158,
      SEL => romodatao7_s_10_BXINV,
      O => romodatao7_s_10_F5MUX
    );
  romodatao7_s_10_BXINV_6100 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_10_BXINV
    );
  romodatao7_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_10_F6MUX,
      O => romodatao7_s(10)
    );
  romodatao7_s_10_F6MUX_6101 : X_MUX2
    port map (
      IA => nx54672z1153,
      IB => nx54672z1156,
      SEL => romodatao7_s_10_BYINV,
      O => romodatao7_s_10_F6MUX
    );
  romodatao7_s_10_BYINV_6102 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_10_BYINV
    );
  nx54672z1153_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1153_F5MUX,
      O => nx54672z1153
    );
  nx54672z1153_F5MUX_6103 : X_MUX2
    port map (
      IA => nx54672z1154,
      IB => nx54672z1155,
      SEL => nx54672z1153_BXINV,
      O => nx54672z1153_F5MUX
    );
  nx54672z1153_BXINV_6104 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1153_BXINV
    );
  romodatao3_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_11_F5MUX,
      O => nx54672z834
    );
  romodatao3_s_11_F5MUX_6105 : X_MUX2
    port map (
      IA => nx54672z835,
      IB => nx54672z836,
      SEL => romodatao3_s_11_BXINV,
      O => romodatao3_s_11_F5MUX
    );
  romodatao3_s_11_BXINV_6106 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_11_BXINV
    );
  romodatao3_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_11_F6MUX,
      O => romodatao3_s(11)
    );
  romodatao3_s_11_F6MUX_6107 : X_MUX2
    port map (
      IA => nx54672z831,
      IB => nx54672z834,
      SEL => romodatao3_s_11_BYINV,
      O => romodatao3_s_11_F6MUX
    );
  romodatao3_s_11_BYINV_6108 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_11_BYINV
    );
  nx54672z831_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z831_F5MUX,
      O => nx54672z831
    );
  nx54672z831_F5MUX_6109 : X_MUX2
    port map (
      IA => nx54672z832,
      IB => nx54672z833,
      SEL => nx54672z831_BXINV,
      O => nx54672z831_F5MUX
    );
  nx54672z831_BXINV_6110 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z831_BXINV
    );
  romodatao2_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_3_F5MUX,
      O => nx54672z803
    );
  romodatao2_s_3_F5MUX_6111 : X_MUX2
    port map (
      IA => nx54672z804,
      IB => nx54672z805,
      SEL => romodatao2_s_3_BXINV,
      O => romodatao2_s_3_F5MUX
    );
  romodatao2_s_3_BXINV_6112 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao2_s_3_BXINV
    );
  romodatao2_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao2_s_3_F6MUX,
      O => romodatao2_s(3)
    );
  romodatao2_s_3_F6MUX_6113 : X_MUX2
    port map (
      IA => nx54672z800,
      IB => nx54672z803,
      SEL => romodatao2_s_3_BYINV,
      O => romodatao2_s_3_F6MUX
    );
  romodatao2_s_3_BYINV_6114 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao2_s_3_BYINV
    );
  nx54672z800_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z800_F5MUX,
      O => nx54672z800
    );
  nx54672z800_F5MUX_6115 : X_MUX2
    port map (
      IA => nx54672z801,
      IB => nx54672z802,
      SEL => nx54672z800_BXINV,
      O => nx54672z800_F5MUX
    );
  nx54672z800_BXINV_6116 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z800_BXINV
    );
  romedatao4_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_9_F5MUX,
      O => nx54672z286
    );
  romedatao4_s_9_F5MUX_6117 : X_MUX2
    port map (
      IA => nx54672z287,
      IB => nx54672z288,
      SEL => romedatao4_s_9_BXINV,
      O => romedatao4_s_9_F5MUX
    );
  romedatao4_s_9_BXINV_6118 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao4_s_9_BXINV
    );
  romedatao4_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_9_F6MUX,
      O => romedatao4_s(9)
    );
  romedatao4_s_9_F6MUX_6119 : X_MUX2
    port map (
      IA => nx54672z283,
      IB => nx54672z286,
      SEL => romedatao4_s_9_BYINV,
      O => romedatao4_s_9_F6MUX
    );
  romedatao4_s_9_BYINV_6120 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao4_s_9_BYINV
    );
  nx54672z283_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z283_F5MUX,
      O => nx54672z283
    );
  nx54672z283_F5MUX_6121 : X_MUX2
    port map (
      IA => nx54672z284,
      IB => nx54672z285,
      SEL => nx54672z283_BXINV,
      O => nx54672z283_F5MUX
    );
  nx54672z283_BXINV_6122 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z283_BXINV
    );
  romedatao4_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_8_F5MUX,
      O => nx54672z292
    );
  romedatao4_s_8_F5MUX_6123 : X_MUX2
    port map (
      IA => nx54672z293,
      IB => nx54672z294,
      SEL => romedatao4_s_8_BXINV,
      O => romedatao4_s_8_F5MUX
    );
  romedatao4_s_8_BXINV_6124 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao4_s_8_BXINV
    );
  romedatao4_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_8_F6MUX,
      O => romedatao4_s(8)
    );
  romedatao4_s_8_F6MUX_6125 : X_MUX2
    port map (
      IA => nx54672z289,
      IB => nx54672z292,
      SEL => romedatao4_s_8_BYINV,
      O => romedatao4_s_8_F6MUX
    );
  romedatao4_s_8_BYINV_6126 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao4_s_8_BYINV
    );
  nx54672z289_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z289_F5MUX,
      O => nx54672z289
    );
  nx54672z289_F5MUX_6127 : X_MUX2
    port map (
      IA => nx54672z290,
      IB => nx54672z291,
      SEL => nx54672z289_BXINV,
      O => nx54672z289_F5MUX
    );
  nx54672z289_BXINV_6128 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z289_BXINV
    );
  romedatao4_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_7_F5MUX,
      O => nx54672z298
    );
  romedatao4_s_7_F5MUX_6129 : X_MUX2
    port map (
      IA => nx54672z299,
      IB => nx54672z300,
      SEL => romedatao4_s_7_BXINV,
      O => romedatao4_s_7_F5MUX
    );
  romedatao4_s_7_BXINV_6130 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao4_s_7_BXINV
    );
  romedatao4_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_7_F6MUX,
      O => romedatao4_s(7)
    );
  romedatao4_s_7_F6MUX_6131 : X_MUX2
    port map (
      IA => nx54672z295,
      IB => nx54672z298,
      SEL => romedatao4_s_7_BYINV,
      O => romedatao4_s_7_F6MUX
    );
  romedatao4_s_7_BYINV_6132 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao4_s_7_BYINV
    );
  nx54672z295_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z295_F5MUX,
      O => nx54672z295
    );
  nx54672z295_F5MUX_6133 : X_MUX2
    port map (
      IA => nx54672z296,
      IB => nx54672z297,
      SEL => nx54672z295_BXINV,
      O => nx54672z295_F5MUX
    );
  nx54672z295_BXINV_6134 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z295_BXINV
    );
  romedatao3_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_11_F5MUX,
      O => nx54672z209
    );
  romedatao3_s_11_F5MUX_6135 : X_MUX2
    port map (
      IA => nx54672z210,
      IB => nx54672z211,
      SEL => romedatao3_s_11_BXINV,
      O => romedatao3_s_11_F5MUX
    );
  romedatao3_s_11_BXINV_6136 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao3_s_11_BXINV
    );
  romedatao3_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_11_F6MUX,
      O => romedatao3_s(11)
    );
  romedatao3_s_11_F6MUX_6137 : X_MUX2
    port map (
      IA => nx54672z206,
      IB => nx54672z209,
      SEL => romedatao3_s_11_BYINV,
      O => romedatao3_s_11_F6MUX
    );
  romedatao3_s_11_BYINV_6138 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao3_s_11_BYINV
    );
  U_DCT2D_reg_databuf_reg_7_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_7_4_DYMUX,
      CE => U_DCT2D_databuf_reg_7_4_CEINV,
      CLK => U_DCT2D_databuf_reg_7_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_7_4_FFY_RST,
      O => U_DCT2D_databuf_reg_7_Q(5)
    );
  U_DCT2D_databuf_reg_7_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_7_4_FFY_RST
    );
  nx54672z206_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z206_F5MUX,
      O => nx54672z206
    );
  nx54672z206_F5MUX_6139 : X_MUX2
    port map (
      IA => nx54672z207,
      IB => nx54672z208,
      SEL => nx54672z206_BXINV,
      O => nx54672z206_F5MUX
    );
  nx54672z206_BXINV_6140 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z206_BXINV
    );
  romedatao3_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_7_F5MUX,
      O => nx54672z233
    );
  romedatao3_s_7_F5MUX_6141 : X_MUX2
    port map (
      IA => nx54672z234,
      IB => nx54672z235,
      SEL => romedatao3_s_7_BXINV,
      O => romedatao3_s_7_F5MUX
    );
  romedatao3_s_7_BXINV_6142 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao3_s_7_BXINV
    );
  romedatao3_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_7_F6MUX,
      O => romedatao3_s(7)
    );
  romedatao3_s_7_F6MUX_6143 : X_MUX2
    port map (
      IA => nx54672z230,
      IB => nx54672z233,
      SEL => romedatao3_s_7_BYINV,
      O => romedatao3_s_7_F6MUX
    );
  romedatao3_s_7_BYINV_6144 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao3_s_7_BYINV
    );
  nx54672z230_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z230_F5MUX,
      O => nx54672z230
    );
  nx54672z230_F5MUX_6145 : X_MUX2
    port map (
      IA => nx54672z231,
      IB => nx54672z232,
      SEL => nx54672z230_BXINV,
      O => nx54672z230_F5MUX
    );
  nx54672z230_BXINV_6146 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z230_BXINV
    );
  romedatao7_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_13_F5MUX,
      O => nx54672z457
    );
  romedatao7_s_13_F5MUX_6147 : X_MUX2
    port map (
      IA => nx54672z458,
      IB => nx54672z459,
      SEL => romedatao7_s_13_BXINV,
      O => romedatao7_s_13_F5MUX
    );
  romedatao7_s_13_BXINV_6148 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao7_s_13_BXINV
    );
  romedatao7_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_13_F6MUX,
      O => romedatao7_s(13)
    );
  romedatao7_s_13_F6MUX_6149 : X_MUX2
    port map (
      IA => nx54672z455,
      IB => nx54672z457,
      SEL => romedatao7_s_13_BYINV,
      O => romedatao7_s_13_F6MUX
    );
  romedatao7_s_13_BYINV_6150 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao7_s_13_BYINV
    );
  nx54672z455_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z455_F5MUX,
      O => nx54672z455
    );
  nx54672z455_F5MUX_6151 : X_MUX2
    port map (
      IA => nx54672z455_G,
      IB => nx54672z456,
      SEL => nx54672z455_BXINV,
      O => nx54672z455_F5MUX
    );
  nx54672z455_BXINV_6152 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z455_BXINV
    );
  romedatao6_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_11_F5MUX,
      O => nx54672z404
    );
  romedatao6_s_11_F5MUX_6153 : X_MUX2
    port map (
      IA => nx54672z405,
      IB => nx54672z406,
      SEL => romedatao6_s_11_BXINV,
      O => romedatao6_s_11_F5MUX
    );
  romedatao6_s_11_BXINV_6154 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao6_s_11_BXINV
    );
  romedatao6_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_11_F6MUX,
      O => romedatao6_s(11)
    );
  romedatao6_s_11_F6MUX_6155 : X_MUX2
    port map (
      IA => nx54672z401,
      IB => nx54672z404,
      SEL => romedatao6_s_11_BYINV,
      O => romedatao6_s_11_F6MUX
    );
  romedatao6_s_11_BYINV_6156 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao6_s_11_BYINV
    );
  nx54672z401_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z401_F5MUX,
      O => nx54672z401
    );
  nx54672z401_F5MUX_6157 : X_MUX2
    port map (
      IA => nx54672z402,
      IB => nx54672z403,
      SEL => nx54672z401_BXINV,
      O => nx54672z401_F5MUX
    );
  nx54672z401_BXINV_6158 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z401_BXINV
    );
  romedatao6_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_10_F5MUX,
      O => nx54672z410
    );
  romedatao6_s_10_F5MUX_6159 : X_MUX2
    port map (
      IA => nx54672z411,
      IB => nx54672z412,
      SEL => romedatao6_s_10_BXINV,
      O => romedatao6_s_10_F5MUX
    );
  romedatao6_s_10_BXINV_6160 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao6_s_10_BXINV
    );
  romedatao6_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_10_F6MUX,
      O => romedatao6_s(10)
    );
  romedatao6_s_10_F6MUX_6161 : X_MUX2
    port map (
      IA => nx54672z407,
      IB => nx54672z410,
      SEL => romedatao6_s_10_BYINV,
      O => romedatao6_s_10_F6MUX
    );
  romedatao6_s_10_BYINV_6162 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao6_s_10_BYINV
    );
  nx54672z407_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z407_F5MUX,
      O => nx54672z407
    );
  nx54672z407_F5MUX_6163 : X_MUX2
    port map (
      IA => nx54672z408,
      IB => nx54672z409,
      SEL => nx54672z407_BXINV,
      O => nx54672z407_F5MUX
    );
  nx54672z407_BXINV_6164 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z407_BXINV
    );
  romedatao6_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_9_F5MUX,
      O => nx54672z416
    );
  romedatao6_s_9_F5MUX_6165 : X_MUX2
    port map (
      IA => nx54672z417,
      IB => nx54672z418,
      SEL => romedatao6_s_9_BXINV,
      O => romedatao6_s_9_F5MUX
    );
  romedatao6_s_9_BXINV_6166 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao6_s_9_BXINV
    );
  romedatao6_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_9_F6MUX,
      O => romedatao6_s(9)
    );
  romedatao6_s_9_F6MUX_6167 : X_MUX2
    port map (
      IA => nx54672z413,
      IB => nx54672z416,
      SEL => romedatao6_s_9_BYINV,
      O => romedatao6_s_9_F6MUX
    );
  romedatao6_s_9_BYINV_6168 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao6_s_9_BYINV
    );
  U_DCT2D_ix38135z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_3_4_Q,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_4_4_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx38135z1
    );
  nx54672z413_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z413_F5MUX,
      O => nx54672z413
    );
  nx54672z413_F5MUX_6169 : X_MUX2
    port map (
      IA => nx54672z414,
      IB => nx54672z415,
      SEL => nx54672z413_BXINV,
      O => nx54672z413_F5MUX
    );
  nx54672z413_BXINV_6170 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z413_BXINV
    );
  romedatao6_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_8_F5MUX,
      O => nx54672z422
    );
  romedatao6_s_8_F5MUX_6171 : X_MUX2
    port map (
      IA => nx54672z423,
      IB => nx54672z424,
      SEL => romedatao6_s_8_BXINV,
      O => romedatao6_s_8_F5MUX
    );
  romedatao6_s_8_BXINV_6172 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao6_s_8_BXINV
    );
  romedatao6_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_8_F6MUX,
      O => romedatao6_s(8)
    );
  romedatao6_s_8_F6MUX_6173 : X_MUX2
    port map (
      IA => nx54672z419,
      IB => nx54672z422,
      SEL => romedatao6_s_8_BYINV,
      O => romedatao6_s_8_F6MUX
    );
  romedatao6_s_8_BYINV_6174 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao6_s_8_BYINV
    );
  nx54672z419_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z419_F5MUX,
      O => nx54672z419
    );
  nx54672z419_F5MUX_6175 : X_MUX2
    port map (
      IA => nx54672z420,
      IB => nx54672z421,
      SEL => nx54672z419_BXINV,
      O => nx54672z419_F5MUX
    );
  nx54672z419_BXINV_6176 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z419_BXINV
    );
  romedatao6_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_7_F5MUX,
      O => nx54672z428
    );
  romedatao6_s_7_F5MUX_6177 : X_MUX2
    port map (
      IA => nx54672z429,
      IB => nx54672z430,
      SEL => romedatao6_s_7_BXINV,
      O => romedatao6_s_7_F5MUX
    );
  romedatao6_s_7_BXINV_6178 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao6_s_7_BXINV
    );
  romedatao6_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_7_F6MUX,
      O => romedatao6_s(7)
    );
  romedatao6_s_7_F6MUX_6179 : X_MUX2
    port map (
      IA => nx54672z425,
      IB => nx54672z428,
      SEL => romedatao6_s_7_BYINV,
      O => romedatao6_s_7_F6MUX
    );
  romedatao6_s_7_BYINV_6180 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao6_s_7_BYINV
    );
  nx54672z425_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z425_F5MUX,
      O => nx54672z425
    );
  nx54672z425_F5MUX_6181 : X_MUX2
    port map (
      IA => nx54672z426,
      IB => nx54672z427,
      SEL => nx54672z425_BXINV,
      O => nx54672z425_F5MUX
    );
  nx54672z425_BXINV_6182 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z425_BXINV
    );
  romedatao8_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_12_F5MUX,
      O => nx54672z528
    );
  romedatao8_s_12_F5MUX_6183 : X_MUX2
    port map (
      IA => nx54672z529,
      IB => nx54672z530,
      SEL => romedatao8_s_12_BXINV,
      O => romedatao8_s_12_F5MUX
    );
  romedatao8_s_12_BXINV_6184 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao8_s_12_BXINV
    );
  romedatao8_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_12_F6MUX,
      O => romedatao8_s(12)
    );
  romedatao8_s_12_F6MUX_6185 : X_MUX2
    port map (
      IA => nx54672z525,
      IB => nx54672z528,
      SEL => romedatao8_s_12_BYINV,
      O => romedatao8_s_12_F6MUX
    );
  romedatao8_s_12_BYINV_6186 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao8_s_12_BYINV
    );
  nx54672z525_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z525_F5MUX,
      O => nx54672z525
    );
  nx54672z525_F5MUX_6187 : X_MUX2
    port map (
      IA => nx54672z526,
      IB => nx54672z527,
      SEL => nx54672z525_BXINV,
      O => nx54672z525_F5MUX
    );
  nx54672z525_BXINV_6188 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z525_BXINV
    );
  romedatao8_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_11_F5MUX,
      O => nx54672z534
    );
  romedatao8_s_11_F5MUX_6189 : X_MUX2
    port map (
      IA => nx54672z535,
      IB => nx54672z536,
      SEL => romedatao8_s_11_BXINV,
      O => romedatao8_s_11_F5MUX
    );
  romedatao8_s_11_BXINV_6190 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao8_s_11_BXINV
    );
  romedatao8_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_11_F6MUX,
      O => romedatao8_s(11)
    );
  romedatao8_s_11_F6MUX_6191 : X_MUX2
    port map (
      IA => nx54672z531,
      IB => nx54672z534,
      SEL => romedatao8_s_11_BYINV,
      O => romedatao8_s_11_F6MUX
    );
  romedatao8_s_11_BYINV_6192 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao8_s_11_BYINV
    );
  nx54672z531_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z531_F5MUX,
      O => nx54672z531
    );
  nx54672z531_F5MUX_6193 : X_MUX2
    port map (
      IA => nx54672z532,
      IB => nx54672z533,
      SEL => nx54672z531_BXINV,
      O => nx54672z531_F5MUX
    );
  nx54672z531_BXINV_6194 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z531_BXINV
    );
  romedatao8_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_10_F5MUX,
      O => nx54672z540
    );
  romedatao8_s_10_F5MUX_6195 : X_MUX2
    port map (
      IA => nx54672z541,
      IB => nx54672z542,
      SEL => romedatao8_s_10_BXINV,
      O => romedatao8_s_10_F5MUX
    );
  romedatao8_s_10_BXINV_6196 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao8_s_10_BXINV
    );
  romedatao8_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_10_F6MUX,
      O => romedatao8_s(10)
    );
  romedatao8_s_10_F6MUX_6197 : X_MUX2
    port map (
      IA => nx54672z537,
      IB => nx54672z540,
      SEL => romedatao8_s_10_BYINV,
      O => romedatao8_s_10_F6MUX
    );
  romedatao8_s_10_BYINV_6198 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao8_s_10_BYINV
    );
  nx54672z537_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z537_F5MUX,
      O => nx54672z537
    );
  nx54672z537_F5MUX_6199 : X_MUX2
    port map (
      IA => nx54672z538,
      IB => nx54672z539,
      SEL => nx54672z537_BXINV,
      O => nx54672z537_F5MUX
    );
  nx54672z537_BXINV_6200 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z537_BXINV
    );
  romedatao8_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_9_F5MUX,
      O => nx54672z546
    );
  romedatao8_s_9_F5MUX_6201 : X_MUX2
    port map (
      IA => nx54672z547,
      IB => nx54672z548,
      SEL => romedatao8_s_9_BXINV,
      O => romedatao8_s_9_F5MUX
    );
  romedatao8_s_9_BXINV_6202 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao8_s_9_BXINV
    );
  romedatao8_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_9_F6MUX,
      O => romedatao8_s(9)
    );
  romedatao8_s_9_F6MUX_6203 : X_MUX2
    port map (
      IA => nx54672z543,
      IB => nx54672z546,
      SEL => romedatao8_s_9_BYINV,
      O => romedatao8_s_9_F6MUX
    );
  romedatao8_s_9_BYINV_6204 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao8_s_9_BYINV
    );
  nx54672z543_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z543_F5MUX,
      O => nx54672z543
    );
  nx54672z543_F5MUX_6205 : X_MUX2
    port map (
      IA => nx54672z544,
      IB => nx54672z545,
      SEL => nx54672z543_BXINV,
      O => nx54672z543_F5MUX
    );
  nx54672z543_BXINV_6206 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z543_BXINV
    );
  romedatao4_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_13_F5MUX,
      O => nx54672z262
    );
  romedatao4_s_13_F5MUX_6207 : X_MUX2
    port map (
      IA => nx54672z263,
      IB => nx54672z264,
      SEL => romedatao4_s_13_BXINV,
      O => romedatao4_s_13_F5MUX
    );
  romedatao4_s_13_BXINV_6208 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao4_s_13_BXINV
    );
  romedatao4_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao4_s_13_F6MUX,
      O => romedatao4_s(13)
    );
  romedatao4_s_13_F6MUX_6209 : X_MUX2
    port map (
      IA => nx54672z260,
      IB => nx54672z262,
      SEL => romedatao4_s_13_BYINV,
      O => romedatao4_s_13_F6MUX
    );
  romedatao4_s_13_BYINV_6210 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao4_s_13_BYINV
    );
  nx54672z260_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z260_F5MUX,
      O => nx54672z260
    );
  nx54672z260_F5MUX_6211 : X_MUX2
    port map (
      IA => nx54672z260_G,
      IB => nx54672z261,
      SEL => nx54672z260_BXINV,
      O => nx54672z260_F5MUX
    );
  nx54672z260_BXINV_6212 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z260_BXINV
    );
  romedatao8_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_13_F5MUX,
      O => nx54672z522
    );
  romedatao8_s_13_F5MUX_6213 : X_MUX2
    port map (
      IA => nx54672z523,
      IB => nx54672z524,
      SEL => romedatao8_s_13_BXINV,
      O => romedatao8_s_13_F5MUX
    );
  romedatao8_s_13_BXINV_6214 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao8_s_13_BXINV
    );
  romedatao8_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_13_F6MUX,
      O => romedatao8_s(13)
    );
  romedatao8_s_13_F6MUX_6215 : X_MUX2
    port map (
      IA => nx54672z520,
      IB => nx54672z522,
      SEL => romedatao8_s_13_BYINV,
      O => romedatao8_s_13_F6MUX
    );
  romedatao8_s_13_BYINV_6216 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao8_s_13_BYINV
    );
  nx54672z520_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z520_F5MUX,
      O => nx54672z520
    );
  nx54672z520_F5MUX_6217 : X_MUX2
    port map (
      IA => nx54672z520_G,
      IB => nx54672z521,
      SEL => nx54672z520_BXINV,
      O => nx54672z520_F5MUX
    );
  nx54672z520_BXINV_6218 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z520_BXINV
    );
  romedatao5_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_8_F5MUX,
      O => nx54672z357
    );
  romedatao5_s_8_F5MUX_6219 : X_MUX2
    port map (
      IA => nx54672z358,
      IB => nx54672z359,
      SEL => romedatao5_s_8_BXINV,
      O => romedatao5_s_8_F5MUX
    );
  romedatao5_s_8_BXINV_6220 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao5_s_8_BXINV
    );
  romedatao5_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_8_F6MUX,
      O => romedatao5_s(8)
    );
  romedatao5_s_8_F6MUX_6221 : X_MUX2
    port map (
      IA => nx54672z354,
      IB => nx54672z357,
      SEL => romedatao5_s_8_BYINV,
      O => romedatao5_s_8_F6MUX
    );
  romedatao5_s_8_BYINV_6222 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao5_s_8_BYINV
    );
  nx54672z354_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z354_F5MUX,
      O => nx54672z354
    );
  nx54672z354_F5MUX_6223 : X_MUX2
    port map (
      IA => nx54672z355,
      IB => nx54672z356,
      SEL => nx54672z354_BXINV,
      O => nx54672z354_F5MUX
    );
  nx54672z354_BXINV_6224 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z354_BXINV
    );
  romedatao5_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_7_F5MUX,
      O => nx54672z363
    );
  romedatao5_s_7_F5MUX_6225 : X_MUX2
    port map (
      IA => nx54672z364,
      IB => nx54672z365,
      SEL => romedatao5_s_7_BXINV,
      O => romedatao5_s_7_F5MUX
    );
  romedatao5_s_7_BXINV_6226 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao5_s_7_BXINV
    );
  romedatao5_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_7_F6MUX,
      O => romedatao5_s(7)
    );
  romedatao5_s_7_F6MUX_6227 : X_MUX2
    port map (
      IA => nx54672z360,
      IB => nx54672z363,
      SEL => romedatao5_s_7_BYINV,
      O => romedatao5_s_7_F6MUX
    );
  romedatao5_s_7_BYINV_6228 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao5_s_7_BYINV
    );
  U_DCT2D_reg_databuf_reg_7_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_7_4_DXMUX,
      CE => U_DCT2D_databuf_reg_7_4_CEINV,
      CLK => U_DCT2D_databuf_reg_7_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_7_4_FFX_RST,
      O => U_DCT2D_databuf_reg_7_Q(4)
    );
  U_DCT2D_databuf_reg_7_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_7_4_FFX_RST
    );
  nx54672z360_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z360_F5MUX,
      O => nx54672z360
    );
  nx54672z360_F5MUX_6229 : X_MUX2
    port map (
      IA => nx54672z361,
      IB => nx54672z362,
      SEL => nx54672z360_BXINV,
      O => nx54672z360_F5MUX
    );
  nx54672z360_BXINV_6230 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z360_BXINV
    );
  romedatao5_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_6_F5MUX,
      O => nx54672z369
    );
  romedatao5_s_6_F5MUX_6231 : X_MUX2
    port map (
      IA => nx54672z370,
      IB => nx54672z371,
      SEL => romedatao5_s_6_BXINV,
      O => romedatao5_s_6_F5MUX
    );
  romedatao5_s_6_BXINV_6232 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao5_s_6_BXINV
    );
  romedatao5_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao5_s_6_F6MUX,
      O => romedatao5_s(6)
    );
  romedatao5_s_6_F6MUX_6233 : X_MUX2
    port map (
      IA => nx54672z366,
      IB => nx54672z369,
      SEL => romedatao5_s_6_BYINV,
      O => romedatao5_s_6_F6MUX
    );
  romedatao5_s_6_BYINV_6234 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao5_s_6_BYINV
    );
  nx54672z366_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z366_F5MUX,
      O => nx54672z366
    );
  nx54672z366_F5MUX_6235 : X_MUX2
    port map (
      IA => nx54672z367,
      IB => nx54672z368,
      SEL => nx54672z366_BXINV,
      O => nx54672z366_F5MUX
    );
  nx54672z366_BXINV_6236 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z366_BXINV
    );
  romodatao6_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_12_F5MUX,
      O => nx54672z1065
    );
  romodatao6_s_12_F5MUX_6237 : X_MUX2
    port map (
      IA => nx54672z1066,
      IB => nx54672z1067,
      SEL => romodatao6_s_12_BXINV,
      O => romodatao6_s_12_F5MUX
    );
  romodatao6_s_12_BXINV_6238 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_12_BXINV
    );
  romodatao6_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_12_F6MUX,
      O => romodatao6_s(12)
    );
  romodatao6_s_12_F6MUX_6239 : X_MUX2
    port map (
      IA => nx54672z1062,
      IB => nx54672z1065,
      SEL => romodatao6_s_12_BYINV,
      O => romodatao6_s_12_F6MUX
    );
  romodatao6_s_12_BYINV_6240 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_12_BYINV
    );
  nx54672z1062_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1062_F5MUX,
      O => nx54672z1062
    );
  nx54672z1062_F5MUX_6241 : X_MUX2
    port map (
      IA => nx54672z1063,
      IB => nx54672z1064,
      SEL => nx54672z1062_BXINV,
      O => nx54672z1062_F5MUX
    );
  nx54672z1062_BXINV_6242 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1062_BXINV
    );
  romodatao6_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_6_F5MUX,
      O => nx54672z1101
    );
  romodatao6_s_6_F5MUX_6243 : X_MUX2
    port map (
      IA => nx54672z1102,
      IB => nx54672z1103,
      SEL => romodatao6_s_6_BXINV,
      O => romodatao6_s_6_F5MUX
    );
  romodatao6_s_6_BXINV_6244 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_6_BXINV
    );
  romodatao6_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_6_F6MUX,
      O => romodatao6_s(6)
    );
  romodatao6_s_6_F6MUX_6245 : X_MUX2
    port map (
      IA => nx54672z1098,
      IB => nx54672z1101,
      SEL => romodatao6_s_6_BYINV,
      O => romodatao6_s_6_F6MUX
    );
  romodatao6_s_6_BYINV_6246 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_6_BYINV
    );
  nx54672z1098_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1098_F5MUX,
      O => nx54672z1098
    );
  nx54672z1098_F5MUX_6247 : X_MUX2
    port map (
      IA => nx54672z1099,
      IB => nx54672z1100,
      SEL => nx54672z1098_BXINV,
      O => nx54672z1098_F5MUX
    );
  nx54672z1098_BXINV_6248 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1098_BXINV
    );
  romodatao6_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_5_F5MUX,
      O => nx54672z1107
    );
  romodatao6_s_5_F5MUX_6249 : X_MUX2
    port map (
      IA => nx54672z1108,
      IB => nx54672z1109,
      SEL => romodatao6_s_5_BXINV,
      O => romodatao6_s_5_F5MUX
    );
  romodatao6_s_5_BXINV_6250 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_5_BXINV
    );
  romodatao6_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_5_F6MUX,
      O => romodatao6_s(5)
    );
  romodatao6_s_5_F6MUX_6251 : X_MUX2
    port map (
      IA => nx54672z1104,
      IB => nx54672z1107,
      SEL => romodatao6_s_5_BYINV,
      O => romodatao6_s_5_F6MUX
    );
  romodatao6_s_5_BYINV_6252 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_5_BYINV
    );
  nx54672z1104_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1104_F5MUX,
      O => nx54672z1104
    );
  nx54672z1104_F5MUX_6253 : X_MUX2
    port map (
      IA => nx54672z1105,
      IB => nx54672z1106,
      SEL => nx54672z1104_BXINV,
      O => nx54672z1104_F5MUX
    );
  nx54672z1104_BXINV_6254 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1104_BXINV
    );
  U_DCT2D_ix41126z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_3_7_Q,
      ADR1 => U_DCT2D_latchbuf_reg_4_7_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx41126z1
    );
  romodatao6_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_4_F5MUX,
      O => nx54672z1113
    );
  romodatao6_s_4_F5MUX_6255 : X_MUX2
    port map (
      IA => nx54672z1114,
      IB => nx54672z1115,
      SEL => romodatao6_s_4_BXINV,
      O => romodatao6_s_4_F5MUX
    );
  romodatao6_s_4_BXINV_6256 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_4_BXINV
    );
  romodatao6_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_4_F6MUX,
      O => romodatao6_s(4)
    );
  romodatao6_s_4_F6MUX_6257 : X_MUX2
    port map (
      IA => nx54672z1110,
      IB => nx54672z1113,
      SEL => romodatao6_s_4_BYINV,
      O => romodatao6_s_4_F6MUX
    );
  romodatao6_s_4_BYINV_6258 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_4_BYINV
    );
  nx54672z1110_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1110_F5MUX,
      O => nx54672z1110
    );
  nx54672z1110_F5MUX_6259 : X_MUX2
    port map (
      IA => nx54672z1111,
      IB => nx54672z1112,
      SEL => nx54672z1110_BXINV,
      O => nx54672z1110_F5MUX
    );
  nx54672z1110_BXINV_6260 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1110_BXINV
    );
  romodatao6_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_3_F5MUX,
      O => nx54672z1119
    );
  romodatao6_s_3_F5MUX_6261 : X_MUX2
    port map (
      IA => nx54672z1120,
      IB => nx54672z1121,
      SEL => romodatao6_s_3_BXINV,
      O => romodatao6_s_3_F5MUX
    );
  romodatao6_s_3_BXINV_6262 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_3_BXINV
    );
  romodatao6_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_3_F6MUX,
      O => romodatao6_s(3)
    );
  romodatao6_s_3_F6MUX_6263 : X_MUX2
    port map (
      IA => nx54672z1116,
      IB => nx54672z1119,
      SEL => romodatao6_s_3_BYINV,
      O => romodatao6_s_3_F6MUX
    );
  romodatao6_s_3_BYINV_6264 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_3_BYINV
    );
  nx54672z1116_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1116_F5MUX,
      O => nx54672z1116
    );
  nx54672z1116_F5MUX_6265 : X_MUX2
    port map (
      IA => nx54672z1117,
      IB => nx54672z1118,
      SEL => nx54672z1116_BXINV,
      O => nx54672z1116_F5MUX
    );
  nx54672z1116_BXINV_6266 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1116_BXINV
    );
  romodatao6_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_2_F5MUX,
      O => nx54672z1125
    );
  romodatao6_s_2_F5MUX_6267 : X_MUX2
    port map (
      IA => nx54672z1126,
      IB => nx54672z1127,
      SEL => romodatao6_s_2_BXINV,
      O => romodatao6_s_2_F5MUX
    );
  romodatao6_s_2_BXINV_6268 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_2_BXINV
    );
  romodatao6_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_2_F6MUX,
      O => romodatao6_s(2)
    );
  romodatao6_s_2_F6MUX_6269 : X_MUX2
    port map (
      IA => nx54672z1122,
      IB => nx54672z1125,
      SEL => romodatao6_s_2_BYINV,
      O => romodatao6_s_2_F6MUX
    );
  romodatao6_s_2_BYINV_6270 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_2_BYINV
    );
  nx54672z1122_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1122_F5MUX,
      O => nx54672z1122
    );
  nx54672z1122_F5MUX_6271 : X_MUX2
    port map (
      IA => nx54672z1123,
      IB => nx54672z1124,
      SEL => nx54672z1122_BXINV,
      O => nx54672z1122_F5MUX
    );
  nx54672z1122_BXINV_6272 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1122_BXINV
    );
  romodatao5_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_12_F5MUX,
      O => nx54672z986
    );
  romodatao5_s_12_F5MUX_6273 : X_MUX2
    port map (
      IA => nx54672z987,
      IB => nx54672z988,
      SEL => romodatao5_s_12_BXINV,
      O => romodatao5_s_12_F5MUX
    );
  romodatao5_s_12_BXINV_6274 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_12_BXINV
    );
  romodatao5_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_12_F6MUX,
      O => romodatao5_s(12)
    );
  romodatao5_s_12_F6MUX_6275 : X_MUX2
    port map (
      IA => nx54672z983,
      IB => nx54672z986,
      SEL => romodatao5_s_12_BYINV,
      O => romodatao5_s_12_F6MUX
    );
  romodatao5_s_12_BYINV_6276 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_12_BYINV
    );
  nx54672z983_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z983_F5MUX,
      O => nx54672z983
    );
  nx54672z983_F5MUX_6277 : X_MUX2
    port map (
      IA => nx54672z984,
      IB => nx54672z985,
      SEL => nx54672z983_BXINV,
      O => nx54672z983_F5MUX
    );
  nx54672z983_BXINV_6278 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z983_BXINV
    );
  romodatao5_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_11_F5MUX,
      O => nx54672z992
    );
  romodatao5_s_11_F5MUX_6279 : X_MUX2
    port map (
      IA => nx54672z993,
      IB => nx54672z994,
      SEL => romodatao5_s_11_BXINV,
      O => romodatao5_s_11_F5MUX
    );
  romodatao5_s_11_BXINV_6280 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_11_BXINV
    );
  romodatao5_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_11_F6MUX,
      O => romodatao5_s(11)
    );
  romodatao5_s_11_F6MUX_6281 : X_MUX2
    port map (
      IA => nx54672z989,
      IB => nx54672z992,
      SEL => romodatao5_s_11_BYINV,
      O => romodatao5_s_11_F6MUX
    );
  romodatao5_s_11_BYINV_6282 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_11_BYINV
    );
  nx54672z989_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z989_F5MUX,
      O => nx54672z989
    );
  nx54672z989_F5MUX_6283 : X_MUX2
    port map (
      IA => nx54672z990,
      IB => nx54672z991,
      SEL => nx54672z989_BXINV,
      O => nx54672z989_F5MUX
    );
  nx54672z989_BXINV_6284 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z989_BXINV
    );
  romodatao5_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_10_F5MUX,
      O => nx54672z998
    );
  romodatao5_s_10_F5MUX_6285 : X_MUX2
    port map (
      IA => nx54672z999,
      IB => nx54672z1000,
      SEL => romodatao5_s_10_BXINV,
      O => romodatao5_s_10_F5MUX
    );
  romodatao5_s_10_BXINV_6286 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_10_BXINV
    );
  romodatao5_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_10_F6MUX,
      O => romodatao5_s(10)
    );
  romodatao5_s_10_F6MUX_6287 : X_MUX2
    port map (
      IA => nx54672z995,
      IB => nx54672z998,
      SEL => romodatao5_s_10_BYINV,
      O => romodatao5_s_10_F6MUX
    );
  romodatao5_s_10_BYINV_6288 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_10_BYINV
    );
  nx54672z995_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z995_F5MUX,
      O => nx54672z995
    );
  nx54672z995_F5MUX_6289 : X_MUX2
    port map (
      IA => nx54672z996,
      IB => nx54672z997,
      SEL => nx54672z995_BXINV,
      O => nx54672z995_F5MUX
    );
  nx54672z995_BXINV_6290 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z995_BXINV
    );
  romodatao5_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_9_F5MUX,
      O => nx54672z1004
    );
  romodatao5_s_9_F5MUX_6291 : X_MUX2
    port map (
      IA => nx54672z1005,
      IB => nx54672z1006,
      SEL => romodatao5_s_9_BXINV,
      O => romodatao5_s_9_F5MUX
    );
  romodatao5_s_9_BXINV_6292 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_9_BXINV
    );
  romodatao5_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_9_F6MUX,
      O => romodatao5_s(9)
    );
  romodatao5_s_9_F6MUX_6293 : X_MUX2
    port map (
      IA => nx54672z1001,
      IB => nx54672z1004,
      SEL => romodatao5_s_9_BYINV,
      O => romodatao5_s_9_F6MUX
    );
  romodatao5_s_9_BYINV_6294 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_9_BYINV
    );
  nx54672z1001_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1001_F5MUX,
      O => nx54672z1001
    );
  nx54672z1001_F5MUX_6295 : X_MUX2
    port map (
      IA => nx54672z1002,
      IB => nx54672z1003,
      SEL => nx54672z1001_BXINV,
      O => nx54672z1001_F5MUX
    );
  nx54672z1001_BXINV_6296 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1001_BXINV
    );
  romodatao5_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_2_F5MUX,
      O => nx54672z1046
    );
  romodatao5_s_2_F5MUX_6297 : X_MUX2
    port map (
      IA => nx54672z1047,
      IB => nx54672z1048,
      SEL => romodatao5_s_2_BXINV,
      O => romodatao5_s_2_F5MUX
    );
  romodatao5_s_2_BXINV_6298 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_2_BXINV
    );
  romodatao5_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_2_F6MUX,
      O => romodatao5_s(2)
    );
  romodatao5_s_2_F6MUX_6299 : X_MUX2
    port map (
      IA => nx54672z1043,
      IB => nx54672z1046,
      SEL => romodatao5_s_2_BYINV,
      O => romodatao5_s_2_F6MUX
    );
  romodatao5_s_2_BYINV_6300 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_2_BYINV
    );
  nx54672z1043_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1043_F5MUX,
      O => nx54672z1043
    );
  nx54672z1043_F5MUX_6301 : X_MUX2
    port map (
      IA => nx54672z1044,
      IB => nx54672z1045,
      SEL => nx54672z1043_BXINV,
      O => nx54672z1043_F5MUX
    );
  nx54672z1043_BXINV_6302 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1043_BXINV
    );
  romodatao5_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_1_F5MUX,
      O => nx54672z1052
    );
  romodatao5_s_1_F5MUX_6303 : X_MUX2
    port map (
      IA => nx54672z1053,
      IB => nx54672z1054,
      SEL => romodatao5_s_1_BXINV,
      O => romodatao5_s_1_F5MUX
    );
  romodatao5_s_1_BXINV_6304 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_1_BXINV
    );
  romodatao5_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_1_F6MUX,
      O => romodatao5_s(1)
    );
  romodatao5_s_1_F6MUX_6305 : X_MUX2
    port map (
      IA => nx54672z1049,
      IB => nx54672z1052,
      SEL => romodatao5_s_1_BYINV,
      O => romodatao5_s_1_F6MUX
    );
  romodatao5_s_1_BYINV_6306 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_1_BYINV
    );
  nx54672z1049_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1049_F5MUX,
      O => nx54672z1049
    );
  nx54672z1049_F5MUX_6307 : X_MUX2
    port map (
      IA => nx54672z1050,
      IB => nx54672z1051,
      SEL => nx54672z1049_BXINV,
      O => nx54672z1049_F5MUX
    );
  nx54672z1049_BXINV_6308 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1049_BXINV
    );
  romodatao8_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_12_F5MUX,
      O => nx54672z1223
    );
  romodatao8_s_12_F5MUX_6309 : X_MUX2
    port map (
      IA => nx54672z1224,
      IB => nx54672z1225,
      SEL => romodatao8_s_12_BXINV,
      O => romodatao8_s_12_F5MUX
    );
  romodatao8_s_12_BXINV_6310 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_12_BXINV
    );
  romodatao8_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_12_F6MUX,
      O => romodatao8_s(12)
    );
  romodatao8_s_12_F6MUX_6311 : X_MUX2
    port map (
      IA => nx54672z1220,
      IB => nx54672z1223,
      SEL => romodatao8_s_12_BYINV,
      O => romodatao8_s_12_F6MUX
    );
  romodatao8_s_12_BYINV_6312 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_12_BYINV
    );
  nx54672z1220_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1220_F5MUX,
      O => nx54672z1220
    );
  nx54672z1220_F5MUX_6313 : X_MUX2
    port map (
      IA => nx54672z1221,
      IB => nx54672z1222,
      SEL => nx54672z1220_BXINV,
      O => nx54672z1220_F5MUX
    );
  nx54672z1220_BXINV_6314 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1220_BXINV
    );
  romodatao8_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_11_F5MUX,
      O => nx54672z1229
    );
  romodatao8_s_11_F5MUX_6315 : X_MUX2
    port map (
      IA => nx54672z1230,
      IB => nx54672z1231,
      SEL => romodatao8_s_11_BXINV,
      O => romodatao8_s_11_F5MUX
    );
  romodatao8_s_11_BXINV_6316 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_11_BXINV
    );
  romodatao8_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_11_F6MUX,
      O => romodatao8_s(11)
    );
  romodatao8_s_11_F6MUX_6317 : X_MUX2
    port map (
      IA => nx54672z1226,
      IB => nx54672z1229,
      SEL => romodatao8_s_11_BYINV,
      O => romodatao8_s_11_F6MUX
    );
  romodatao8_s_11_BYINV_6318 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_11_BYINV
    );
  nx54672z1226_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1226_F5MUX,
      O => nx54672z1226
    );
  nx54672z1226_F5MUX_6319 : X_MUX2
    port map (
      IA => nx54672z1227,
      IB => nx54672z1228,
      SEL => nx54672z1226_BXINV,
      O => nx54672z1226_F5MUX
    );
  nx54672z1226_BXINV_6320 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1226_BXINV
    );
  romodatao6_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_13_F5MUX,
      O => nx54672z1059
    );
  romodatao6_s_13_F5MUX_6321 : X_MUX2
    port map (
      IA => nx54672z1060,
      IB => nx54672z1061,
      SEL => romodatao6_s_13_BXINV,
      O => romodatao6_s_13_F5MUX
    );
  romodatao6_s_13_BXINV_6322 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_13_BXINV
    );
  romodatao6_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_13_F6MUX,
      O => romodatao6_s(13)
    );
  romodatao6_s_13_F6MUX_6323 : X_MUX2
    port map (
      IA => nx54672z1057,
      IB => nx54672z1059,
      SEL => romodatao6_s_13_BYINV,
      O => romodatao6_s_13_F6MUX
    );
  romodatao6_s_13_BYINV_6324 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_13_BYINV
    );
  nx54672z1057_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1057_F5MUX,
      O => nx54672z1057
    );
  nx54672z1057_F5MUX_6325 : X_MUX2
    port map (
      IA => nx54672z1057_G,
      IB => nx54672z1058,
      SEL => nx54672z1057_BXINV,
      O => nx54672z1057_F5MUX
    );
  nx54672z1057_BXINV_6326 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1057_BXINV
    );
  romodatao5_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_0_F5MUX,
      O => U1_ROMO5_modgen_rom_ix0_nx_ro64_32_l
    );
  romodatao5_s_0_F5MUX_6327 : X_MUX2
    port map (
      IA => nx54672z1055,
      IB => nx54672z1056,
      SEL => romodatao5_s_0_BXINV,
      O => romodatao5_s_0_F5MUX
    );
  romodatao5_s_0_BXINV_6328 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao5_s_0_BXINV
    );
  romodatao5_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao5_s_0_F6MUX,
      O => romodatao5_s(0)
    );
  romodatao5_s_0_F6MUX_6329 : X_MUX2
    port map (
      IA => U1_ROMO5_modgen_rom_ix0_nx_ro64_32_u,
      IB => U1_ROMO5_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romodatao5_s_0_BYINV,
      O => romodatao5_s_0_F6MUX
    );
  romodatao5_s_0_BYINV_6330 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao5_s_0_BYINV
    );
  U1_ROMO5_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROMO5_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U1_ROMO5_modgen_rom_ix0_nx_ro64_32_u
    );
  U1_ROMO5_modgen_rom_ix0_nx_ro64_32_u_F5MUX_6331 : X_MUX2
    port map (
      IA => U1_ROMO5_modgen_rom_ix0_nx_rm64_16_u,
      IB => U1_ROMO5_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U1_ROMO5_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U1_ROMO5_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U1_ROMO5_modgen_rom_ix0_nx_ro64_32_u_BXINV_6332 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => U1_ROMO5_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romodatao4_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_8_F5MUX,
      O => nx54672z931
    );
  romodatao4_s_8_F5MUX_6333 : X_MUX2
    port map (
      IA => nx54672z932,
      IB => nx54672z933,
      SEL => romodatao4_s_8_BXINV,
      O => romodatao4_s_8_F5MUX
    );
  romodatao4_s_8_BXINV_6334 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_8_BXINV
    );
  romodatao4_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_8_F6MUX,
      O => romodatao4_s(8)
    );
  romodatao4_s_8_F6MUX_6335 : X_MUX2
    port map (
      IA => nx54672z928,
      IB => nx54672z931,
      SEL => romodatao4_s_8_BYINV,
      O => romodatao4_s_8_F6MUX
    );
  romodatao4_s_8_BYINV_6336 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_8_BYINV
    );
  nx54672z928_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z928_F5MUX,
      O => nx54672z928
    );
  nx54672z928_F5MUX_6337 : X_MUX2
    port map (
      IA => nx54672z929,
      IB => nx54672z930,
      SEL => nx54672z928_BXINV,
      O => nx54672z928_F5MUX
    );
  nx54672z928_BXINV_6338 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z928_BXINV
    );
  romodatao4_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_7_F5MUX,
      O => nx54672z937
    );
  romodatao4_s_7_F5MUX_6339 : X_MUX2
    port map (
      IA => nx54672z938,
      IB => nx54672z939,
      SEL => romodatao4_s_7_BXINV,
      O => romodatao4_s_7_F5MUX
    );
  romodatao4_s_7_BXINV_6340 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_7_BXINV
    );
  romodatao4_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_7_F6MUX,
      O => romodatao4_s(7)
    );
  romodatao4_s_7_F6MUX_6341 : X_MUX2
    port map (
      IA => nx54672z934,
      IB => nx54672z937,
      SEL => romodatao4_s_7_BYINV,
      O => romodatao4_s_7_F6MUX
    );
  romodatao4_s_7_BYINV_6342 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_7_BYINV
    );
  U_DCT2D_reg_databuf_reg_7_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_7_6_DYMUX,
      CE => U_DCT2D_databuf_reg_7_6_CEINV,
      CLK => U_DCT2D_databuf_reg_7_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_7_6_FFY_RST,
      O => U_DCT2D_databuf_reg_7_Q(7)
    );
  U_DCT2D_databuf_reg_7_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_7_6_FFY_RST
    );
  nx54672z934_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z934_F5MUX,
      O => nx54672z934
    );
  nx54672z934_F5MUX_6343 : X_MUX2
    port map (
      IA => nx54672z935,
      IB => nx54672z936,
      SEL => nx54672z934_BXINV,
      O => nx54672z934_F5MUX
    );
  nx54672z934_BXINV_6344 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z934_BXINV
    );
  romedatao7_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_10_F5MUX,
      O => nx54672z475
    );
  romedatao7_s_10_F5MUX_6345 : X_MUX2
    port map (
      IA => nx54672z476,
      IB => nx54672z477,
      SEL => romedatao7_s_10_BXINV,
      O => romedatao7_s_10_F5MUX
    );
  romedatao7_s_10_BXINV_6346 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao7_s_10_BXINV
    );
  romedatao7_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_10_F6MUX,
      O => romedatao7_s(10)
    );
  romedatao7_s_10_F6MUX_6347 : X_MUX2
    port map (
      IA => nx54672z472,
      IB => nx54672z475,
      SEL => romedatao7_s_10_BYINV,
      O => romedatao7_s_10_F6MUX
    );
  romedatao7_s_10_BYINV_6348 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao7_s_10_BYINV
    );
  nx54672z472_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z472_F5MUX,
      O => nx54672z472
    );
  nx54672z472_F5MUX_6349 : X_MUX2
    port map (
      IA => nx54672z473,
      IB => nx54672z474,
      SEL => nx54672z472_BXINV,
      O => nx54672z472_F5MUX
    );
  nx54672z472_BXINV_6350 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z472_BXINV
    );
  romedatao7_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_9_F5MUX,
      O => nx54672z481
    );
  romedatao7_s_9_F5MUX_6351 : X_MUX2
    port map (
      IA => nx54672z482,
      IB => nx54672z483,
      SEL => romedatao7_s_9_BXINV,
      O => romedatao7_s_9_F5MUX
    );
  romedatao7_s_9_BXINV_6352 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao7_s_9_BXINV
    );
  romedatao7_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_9_F6MUX,
      O => romedatao7_s(9)
    );
  romedatao7_s_9_F6MUX_6353 : X_MUX2
    port map (
      IA => nx54672z478,
      IB => nx54672z481,
      SEL => romedatao7_s_9_BYINV,
      O => romedatao7_s_9_F6MUX
    );
  romedatao7_s_9_BYINV_6354 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao7_s_9_BYINV
    );
  nx54672z478_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z478_F5MUX,
      O => nx54672z478
    );
  nx54672z478_F5MUX_6355 : X_MUX2
    port map (
      IA => nx54672z479,
      IB => nx54672z480,
      SEL => nx54672z478_BXINV,
      O => nx54672z478_F5MUX
    );
  nx54672z478_BXINV_6356 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z478_BXINV
    );
  romedatao7_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_8_F5MUX,
      O => nx54672z487
    );
  romedatao7_s_8_F5MUX_6357 : X_MUX2
    port map (
      IA => nx54672z488,
      IB => nx54672z489,
      SEL => romedatao7_s_8_BXINV,
      O => romedatao7_s_8_F5MUX
    );
  romedatao7_s_8_BXINV_6358 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao7_s_8_BXINV
    );
  romedatao7_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_8_F6MUX,
      O => romedatao7_s(8)
    );
  romedatao7_s_8_F6MUX_6359 : X_MUX2
    port map (
      IA => nx54672z484,
      IB => nx54672z487,
      SEL => romedatao7_s_8_BYINV,
      O => romedatao7_s_8_F6MUX
    );
  romedatao7_s_8_BYINV_6360 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao7_s_8_BYINV
    );
  nx54672z484_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z484_F5MUX,
      O => nx54672z484
    );
  nx54672z484_F5MUX_6361 : X_MUX2
    port map (
      IA => nx54672z485,
      IB => nx54672z486,
      SEL => nx54672z484_BXINV,
      O => nx54672z484_F5MUX
    );
  nx54672z484_BXINV_6362 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z484_BXINV
    );
  romedatao7_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_7_F5MUX,
      O => nx54672z493
    );
  romedatao7_s_7_F5MUX_6363 : X_MUX2
    port map (
      IA => nx54672z494,
      IB => nx54672z495,
      SEL => romedatao7_s_7_BXINV,
      O => romedatao7_s_7_F5MUX
    );
  romedatao7_s_7_BXINV_6364 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao7_s_7_BXINV
    );
  romedatao7_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_7_F6MUX,
      O => romedatao7_s(7)
    );
  romedatao7_s_7_F6MUX_6365 : X_MUX2
    port map (
      IA => nx54672z490,
      IB => nx54672z493,
      SEL => romedatao7_s_7_BYINV,
      O => romedatao7_s_7_F6MUX
    );
  romedatao7_s_7_BYINV_6366 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao7_s_7_BYINV
    );
  nx54672z490_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z490_F5MUX,
      O => nx54672z490
    );
  nx54672z490_F5MUX_6367 : X_MUX2
    port map (
      IA => nx54672z491,
      IB => nx54672z492,
      SEL => nx54672z490_BXINV,
      O => nx54672z490_F5MUX
    );
  nx54672z490_BXINV_6368 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z490_BXINV
    );
  romedatao7_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_6_F5MUX,
      O => nx54672z499
    );
  romedatao7_s_6_F5MUX_6369 : X_MUX2
    port map (
      IA => nx54672z500,
      IB => nx54672z501,
      SEL => romedatao7_s_6_BXINV,
      O => romedatao7_s_6_F5MUX
    );
  romedatao7_s_6_BXINV_6370 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao7_s_6_BXINV
    );
  romedatao7_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_6_F6MUX,
      O => romedatao7_s(6)
    );
  romedatao7_s_6_F6MUX_6371 : X_MUX2
    port map (
      IA => nx54672z496,
      IB => nx54672z499,
      SEL => romedatao7_s_6_BYINV,
      O => romedatao7_s_6_F6MUX
    );
  romedatao7_s_6_BYINV_6372 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao7_s_6_BYINV
    );
  U_DCT2D_ix40129z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_4_6_Q,
      ADR1 => U_DCT2D_latchbuf_reg_3_6_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx40129z1
    );
  nx54672z496_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z496_F5MUX,
      O => nx54672z496
    );
  nx54672z496_F5MUX_6373 : X_MUX2
    port map (
      IA => nx54672z497,
      IB => nx54672z498,
      SEL => nx54672z496_BXINV,
      O => nx54672z496_F5MUX
    );
  nx54672z496_BXINV_6374 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z496_BXINV
    );
  romodatao8_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_10_F5MUX,
      O => nx54672z1235
    );
  romodatao8_s_10_F5MUX_6375 : X_MUX2
    port map (
      IA => nx54672z1236,
      IB => nx54672z1237,
      SEL => romodatao8_s_10_BXINV,
      O => romodatao8_s_10_F5MUX
    );
  romodatao8_s_10_BXINV_6376 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_10_BXINV
    );
  romodatao8_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_10_F6MUX,
      O => romodatao8_s(10)
    );
  romodatao8_s_10_F6MUX_6377 : X_MUX2
    port map (
      IA => nx54672z1232,
      IB => nx54672z1235,
      SEL => romodatao8_s_10_BYINV,
      O => romodatao8_s_10_F6MUX
    );
  romodatao8_s_10_BYINV_6378 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_10_BYINV
    );
  nx54672z1232_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1232_F5MUX,
      O => nx54672z1232
    );
  nx54672z1232_F5MUX_6379 : X_MUX2
    port map (
      IA => nx54672z1233,
      IB => nx54672z1234,
      SEL => nx54672z1232_BXINV,
      O => nx54672z1232_F5MUX
    );
  nx54672z1232_BXINV_6380 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1232_BXINV
    );
  romodatao8_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_9_F5MUX,
      O => nx54672z1241
    );
  romodatao8_s_9_F5MUX_6381 : X_MUX2
    port map (
      IA => nx54672z1242,
      IB => nx54672z1243,
      SEL => romodatao8_s_9_BXINV,
      O => romodatao8_s_9_F5MUX
    );
  romodatao8_s_9_BXINV_6382 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_9_BXINV
    );
  romodatao8_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_9_F6MUX,
      O => romodatao8_s(9)
    );
  romodatao8_s_9_F6MUX_6383 : X_MUX2
    port map (
      IA => nx54672z1238,
      IB => nx54672z1241,
      SEL => romodatao8_s_9_BYINV,
      O => romodatao8_s_9_F6MUX
    );
  romodatao8_s_9_BYINV_6384 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_9_BYINV
    );
  nx54672z1238_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1238_F5MUX,
      O => nx54672z1238
    );
  nx54672z1238_F5MUX_6385 : X_MUX2
    port map (
      IA => nx54672z1239,
      IB => nx54672z1240,
      SEL => nx54672z1238_BXINV,
      O => nx54672z1238_F5MUX
    );
  nx54672z1238_BXINV_6386 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1238_BXINV
    );
  romodatao7_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_9_F5MUX,
      O => nx54672z1162
    );
  romodatao7_s_9_F5MUX_6387 : X_MUX2
    port map (
      IA => nx54672z1163,
      IB => nx54672z1164,
      SEL => romodatao7_s_9_BXINV,
      O => romodatao7_s_9_F5MUX
    );
  romodatao7_s_9_BXINV_6388 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_9_BXINV
    );
  romodatao7_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_9_F6MUX,
      O => romodatao7_s(9)
    );
  romodatao7_s_9_F6MUX_6389 : X_MUX2
    port map (
      IA => nx54672z1159,
      IB => nx54672z1162,
      SEL => romodatao7_s_9_BYINV,
      O => romodatao7_s_9_F6MUX
    );
  romodatao7_s_9_BYINV_6390 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_9_BYINV
    );
  U_DCT1D_ix59700z50254 : X_LUT4
    generic map(
      INIT => X"A3AC"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1348(16),
      ADR1 => U_DCT1D_rtlc5n1355(16),
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_rtlc5n1354(15),
      O => U_DCT1D_nx59700z214
    );
  U_DCT1D_ix59700z2163 : X_LUT4
    generic map(
      INIT => X"9955"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1350(9),
      ADR1 => romodatao8_s(1),
      ADR2 => VCC,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z526
    );
  U_DCT1D_ix59700z45375 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => romedatao8_s(3),
      ADR1 => U_DCT1D_rtlc5n1350(11),
      ADR2 => romodatao8_s(3),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z522
    );
  U_DCT1D_ix59700z2166 : X_LUT4
    generic map(
      INIT => X"9933"
    )
    port map (
      ADR0 => romodatao8_s(0),
      ADR1 => U_DCT1D_rtlc5n1350(8),
      ADR2 => VCC,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z528
    );
  U_DCT1D_ix59700z1548 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1345(11),
      ADR1 => U_DCT1D_rtlc5n1344(11),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z183
    );
  U_DCT1D_ix59700z1563 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1344(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1345(8),
      O => U_DCT1D_nx59700z192
    );
  U_DCT1D_ix59700z1537 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_rtlc5n1344(13),
      ADR2 => U_DCT1D_rtlc5n1345(13),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z177
    );
  U_DCT1D_ix59700z1553 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1345(10),
      ADR1 => U_DCT1D_rtlc5n1344(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z186
    );
  U_DCT1D_ix59700z50300 : X_LUT4
    generic map(
      INIT => X"B1E4"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => U_DCT1D_rtlc5n1354(8),
      ADR2 => U_DCT1D_rtlc5n1348(8),
      ADR3 => U_DCT1D_rtlc5n1355(8),
      O => U_DCT1D_nx59700z238
    );
  U_DCT1D_ix59700z50270 : X_LUT4
    generic map(
      INIT => X"DE12"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1355(13),
      ADR1 => U_DCT1D_state_reg(0),
      ADR2 => U_DCT1D_rtlc5n1354(13),
      ADR3 => U_DCT1D_rtlc5n1348(13),
      O => U_DCT1D_nx59700z223
    );
  U_DCT1D_ix59700z50282 : X_LUT4
    generic map(
      INIT => X"A3AC"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1348(11),
      ADR1 => U_DCT1D_rtlc5n1355(11),
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_rtlc5n1354(11),
      O => U_DCT1D_nx59700z229
    );
  U_DCT1D_ix59700z50288 : X_LUT4
    generic map(
      INIT => X"8DD8"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => U_DCT1D_rtlc5n1348(10),
      ADR2 => U_DCT1D_rtlc5n1355(10),
      ADR3 => U_DCT1D_rtlc5n1354(10),
      O => U_DCT1D_nx59700z232
    );
  ix53675z45507 : X_LUT4
    generic map(
      INIT => X"96C6"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(2),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1303
    );
  ix53675z53144 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro7_s(1),
      O => nx53675z1306
    );
  ix53675z44548 : X_LUT4
    generic map(
      INIT => X"C0C2"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => romo2addro7_s(2),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1311
    );
  ix53675z39057 : X_LUT4
    generic map(
      INIT => X"A244"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => romo2addro7_s(2),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1309
    );
  ix53675z62701 : X_LUT4
    generic map(
      INIT => X"F880"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => romo2addro7_s(2),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1312
    );
  ix53675z26404 : X_LUT4
    generic map(
      INIT => X"666C"
    )
    port map (
      ADR0 => romo2addro8_s(0),
      ADR1 => romo2addro8_s(2),
      ADR2 => romo2addro8_s(3),
      ADR3 => romo2addro8_s(1),
      O => nx53675z1360
    );
  ix53675z23396 : X_LUT4
    generic map(
      INIT => X"2B22"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => romo2addro7_s(2),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1308
    );
  ix53675z59862 : X_LUT4
    generic map(
      INIT => X"9A9A"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(0),
      ADR3 => VCC,
      O => nx53675z1366
    );
  ix53675z55520 : X_LUT4
    generic map(
      INIT => X"F10E"
    )
    port map (
      ADR0 => romo2addro8_s(0),
      ADR1 => romo2addro8_s(2),
      ADR2 => romo2addro8_s(3),
      ADR3 => romo2addro8_s(1),
      O => nx53675z1358
    );
  ix53675z41799 : X_LUT4
    generic map(
      INIT => X"9A66"
    )
    port map (
      ADR0 => romo2addro8_s(0),
      ADR1 => romo2addro8_s(2),
      ADR2 => romo2addro8_s(3),
      ADR3 => romo2addro8_s(1),
      O => nx53675z1361
    );
  U_DCT1D_reg_ramdatai_s_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramdatai_s_0_DXMUX,
      CE => ramdatai_s_0_CEINV,
      CLK => ramdatai_s_0_CLKINV,
      SET => GND,
      RST => ramdatai_s_0_FFX_RST,
      O => ramdatai_s(0)
    );
  ramdatai_s_0_FFX_RSTOR : X_OR2
    port map (
      I0 => ramdatai_s_0_SRINV,
      I1 => GSR,
      O => ramdatai_s_0_FFX_RST
    );
  U_DCT1D_ix59700z45348 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => romedatao8_s(9),
      ADR1 => U_DCT1D_rtlc5n1350(17),
      ADR2 => romodatao8_s(9),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z504
    );
  U_DCT1D_reg_ramdatai_s_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramdatai_s_2_DYMUX,
      CE => ramdatai_s_2_CEINV,
      CLK => ramdatai_s_2_CLKINV,
      SET => GND,
      RST => ramdatai_s_2_FFY_RST,
      O => ramdatai_s(3)
    );
  ramdatai_s_2_FFY_RSTOR : X_OR2
    port map (
      I0 => ramdatai_s_2_SRINV,
      I1 => GSR,
      O => ramdatai_s_2_FFY_RST
    );
  U_DCT1D_ix59700z45361 : X_LUT4
    generic map(
      INIT => X"A599"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1350(14),
      ADR1 => romedatao8_s(6),
      ADR2 => romodatao8_s(6),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z513
    );
  U_DCT1D_reg_ramdatai_s_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramdatai_s_2_DXMUX,
      CE => ramdatai_s_2_CEINV,
      CLK => ramdatai_s_2_CLKINV,
      SET => GND,
      RST => ramdatai_s_2_FFX_RST,
      O => ramdatai_s(2)
    );
  ramdatai_s_2_FFX_RSTOR : X_OR2
    port map (
      I0 => ramdatai_s_2_SRINV,
      I1 => GSR,
      O => ramdatai_s_2_FFX_RST
    );
  U_DCT1D_ix59700z2385 : X_LUT4
    generic map(
      INIT => X"2288"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => romodatao6_s(1),
      ADR2 => VCC,
      ADR3 => romodatao7_s(0),
      O => U_DCT1D_nx59700z374
    );
  U_DCT1D_ix59700z23988 : X_LUT4
    generic map(
      INIT => X"56A6"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z369,
      ADR1 => romedatao7_s(2),
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => romodatao7_s(2),
      O => U_DCT1D_nx59700z368
    );
  U_DCT1D_ix59700z1584 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1344(4),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1345(4),
      O => U_DCT1D_nx59700z204
    );
  U_DCT1D_ix59700z1558 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_rtlc5n1344(9),
      ADR2 => U_DCT1D_rtlc5n1345(9),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z189
    );
  U_DCT1D_ix59700z1573 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1345(6),
      ADR1 => U_DCT1D_rtlc5n1344(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z198
    );
  ix54672z8290 : X_LUT4
    generic map(
      INIT => X"1C86"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(0),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(2),
      O => nx54672z468
    );
  ix54672z29076 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(2),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(0),
      O => nx54672z517
    );
  ix54672z29073 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(2),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(0),
      O => U1_ROME7_modgen_rom_ix2_nx_rm64_16_u
    );
  ix54672z14383 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => VCC,
      ADR2 => romeaddro7_s(2),
      ADR3 => VCC,
      O => nx54672z518
    );
  ix54672z2214 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(0),
      O => nx54672z515
    );
  ix54672z17473 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romeaddro7_s(2),
      O => nx54672z519
    );
  ix54672z23981 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(3),
      O => U1_ROME7_modgen_rom_ix2_nx_rm64_16_l
    );
  nx54672z1159_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1159_F5MUX,
      O => nx54672z1159
    );
  nx54672z1159_F5MUX_6391 : X_MUX2
    port map (
      IA => nx54672z1160,
      IB => nx54672z1161,
      SEL => nx54672z1159_BXINV,
      O => nx54672z1159_F5MUX
    );
  nx54672z1159_BXINV_6392 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1159_BXINV
    );
  romodatao7_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_8_F5MUX,
      O => nx54672z1168
    );
  romodatao7_s_8_F5MUX_6393 : X_MUX2
    port map (
      IA => nx54672z1169,
      IB => nx54672z1170,
      SEL => romodatao7_s_8_BXINV,
      O => romodatao7_s_8_F5MUX
    );
  romodatao7_s_8_BXINV_6394 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_8_BXINV
    );
  romodatao7_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_8_F6MUX,
      O => romodatao7_s(8)
    );
  romodatao7_s_8_F6MUX_6395 : X_MUX2
    port map (
      IA => nx54672z1165,
      IB => nx54672z1168,
      SEL => romodatao7_s_8_BYINV,
      O => romodatao7_s_8_F6MUX
    );
  romodatao7_s_8_BYINV_6396 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_8_BYINV
    );
  nx54672z1165_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1165_F5MUX,
      O => nx54672z1165
    );
  nx54672z1165_F5MUX_6397 : X_MUX2
    port map (
      IA => nx54672z1166,
      IB => nx54672z1167,
      SEL => nx54672z1165_BXINV,
      O => nx54672z1165_F5MUX
    );
  nx54672z1165_BXINV_6398 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1165_BXINV
    );
  romodatao7_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_7_F5MUX,
      O => nx54672z1174
    );
  romodatao7_s_7_F5MUX_6399 : X_MUX2
    port map (
      IA => nx54672z1175,
      IB => nx54672z1176,
      SEL => romodatao7_s_7_BXINV,
      O => romodatao7_s_7_F5MUX
    );
  romodatao7_s_7_BXINV_6400 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_7_BXINV
    );
  romodatao7_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_7_F6MUX,
      O => romodatao7_s(7)
    );
  romodatao7_s_7_F6MUX_6401 : X_MUX2
    port map (
      IA => nx54672z1171,
      IB => nx54672z1174,
      SEL => romodatao7_s_7_BYINV,
      O => romodatao7_s_7_F6MUX
    );
  romodatao7_s_7_BYINV_6402 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_7_BYINV
    );
  nx54672z1171_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1171_F5MUX,
      O => nx54672z1171
    );
  nx54672z1171_F5MUX_6403 : X_MUX2
    port map (
      IA => nx54672z1172,
      IB => nx54672z1173,
      SEL => nx54672z1171_BXINV,
      O => nx54672z1171_F5MUX
    );
  nx54672z1171_BXINV_6404 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1171_BXINV
    );
  romodatao7_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_6_F5MUX,
      O => nx54672z1180
    );
  romodatao7_s_6_F5MUX_6405 : X_MUX2
    port map (
      IA => nx54672z1181,
      IB => nx54672z1182,
      SEL => romodatao7_s_6_BXINV,
      O => romodatao7_s_6_F5MUX
    );
  romodatao7_s_6_BXINV_6406 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_6_BXINV
    );
  romodatao7_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_6_F6MUX,
      O => romodatao7_s(6)
    );
  romodatao7_s_6_F6MUX_6407 : X_MUX2
    port map (
      IA => nx54672z1177,
      IB => nx54672z1180,
      SEL => romodatao7_s_6_BYINV,
      O => romodatao7_s_6_F6MUX
    );
  romodatao7_s_6_BYINV_6408 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_6_BYINV
    );
  nx54672z1177_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1177_F5MUX,
      O => nx54672z1177
    );
  nx54672z1177_F5MUX_6409 : X_MUX2
    port map (
      IA => nx54672z1178,
      IB => nx54672z1179,
      SEL => nx54672z1177_BXINV,
      O => nx54672z1177_F5MUX
    );
  nx54672z1177_BXINV_6410 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1177_BXINV
    );
  romodatao7_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_5_F5MUX,
      O => nx54672z1186
    );
  romodatao7_s_5_F5MUX_6411 : X_MUX2
    port map (
      IA => nx54672z1187,
      IB => nx54672z1188,
      SEL => romodatao7_s_5_BXINV,
      O => romodatao7_s_5_F5MUX
    );
  romodatao7_s_5_BXINV_6412 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_5_BXINV
    );
  romodatao7_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_5_F6MUX,
      O => romodatao7_s(5)
    );
  romodatao7_s_5_F6MUX_6413 : X_MUX2
    port map (
      IA => nx54672z1183,
      IB => nx54672z1186,
      SEL => romodatao7_s_5_BYINV,
      O => romodatao7_s_5_F6MUX
    );
  romodatao7_s_5_BYINV_6414 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_5_BYINV
    );
  nx54672z1183_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1183_F5MUX,
      O => nx54672z1183
    );
  nx54672z1183_F5MUX_6415 : X_MUX2
    port map (
      IA => nx54672z1184,
      IB => nx54672z1185,
      SEL => nx54672z1183_BXINV,
      O => nx54672z1183_F5MUX
    );
  nx54672z1183_BXINV_6416 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1183_BXINV
    );
  romodatao3_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_9_F5MUX,
      O => nx54672z846
    );
  romodatao3_s_9_F5MUX_6417 : X_MUX2
    port map (
      IA => nx54672z847,
      IB => nx54672z848,
      SEL => romodatao3_s_9_BXINV,
      O => romodatao3_s_9_F5MUX
    );
  romodatao3_s_9_BXINV_6418 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_9_BXINV
    );
  romodatao3_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_9_F6MUX,
      O => romodatao3_s(9)
    );
  romodatao3_s_9_F6MUX_6419 : X_MUX2
    port map (
      IA => nx54672z843,
      IB => nx54672z846,
      SEL => romodatao3_s_9_BYINV,
      O => romodatao3_s_9_F6MUX
    );
  romodatao3_s_9_BYINV_6420 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_9_BYINV
    );
  nx54672z843_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z843_F5MUX,
      O => nx54672z843
    );
  nx54672z843_F5MUX_6421 : X_MUX2
    port map (
      IA => nx54672z844,
      IB => nx54672z845,
      SEL => nx54672z843_BXINV,
      O => nx54672z843_F5MUX
    );
  nx54672z843_BXINV_6422 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z843_BXINV
    );
  romodatao3_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_5_F5MUX,
      O => nx54672z870
    );
  romodatao3_s_5_F5MUX_6423 : X_MUX2
    port map (
      IA => nx54672z871,
      IB => nx54672z872,
      SEL => romodatao3_s_5_BXINV,
      O => romodatao3_s_5_F5MUX
    );
  romodatao3_s_5_BXINV_6424 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_5_BXINV
    );
  romodatao3_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_5_F6MUX,
      O => romodatao3_s(5)
    );
  romodatao3_s_5_F6MUX_6425 : X_MUX2
    port map (
      IA => nx54672z867,
      IB => nx54672z870,
      SEL => romodatao3_s_5_BYINV,
      O => romodatao3_s_5_F6MUX
    );
  romodatao3_s_5_BYINV_6426 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_5_BYINV
    );
  nx54672z867_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z867_F5MUX,
      O => nx54672z867
    );
  nx54672z867_F5MUX_6427 : X_MUX2
    port map (
      IA => nx54672z868,
      IB => nx54672z869,
      SEL => nx54672z867_BXINV,
      O => nx54672z867_F5MUX
    );
  nx54672z867_BXINV_6428 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z867_BXINV
    );
  romedatao3_s_9_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_9_F5MUX,
      O => nx54672z221
    );
  romedatao3_s_9_F5MUX_6429 : X_MUX2
    port map (
      IA => nx54672z222,
      IB => nx54672z223,
      SEL => romedatao3_s_9_BXINV,
      O => romedatao3_s_9_F5MUX
    );
  romedatao3_s_9_BXINV_6430 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao3_s_9_BXINV
    );
  romedatao3_s_9_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_9_F6MUX,
      O => romedatao3_s(9)
    );
  romedatao3_s_9_F6MUX_6431 : X_MUX2
    port map (
      IA => nx54672z218,
      IB => nx54672z221,
      SEL => romedatao3_s_9_BYINV,
      O => romedatao3_s_9_F6MUX
    );
  romedatao3_s_9_BYINV_6432 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao3_s_9_BYINV
    );
  U_DCT2D_reg_databuf_reg_7_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_7_6_DXMUX,
      CE => U_DCT2D_databuf_reg_7_6_CEINV,
      CLK => U_DCT2D_databuf_reg_7_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_7_6_FFX_RST,
      O => U_DCT2D_databuf_reg_7_Q(6)
    );
  U_DCT2D_databuf_reg_7_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_7_6_FFX_RST
    );
  nx54672z218_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z218_F5MUX,
      O => nx54672z218
    );
  nx54672z218_F5MUX_6433 : X_MUX2
    port map (
      IA => nx54672z219,
      IB => nx54672z220,
      SEL => nx54672z218_BXINV,
      O => nx54672z218_F5MUX
    );
  nx54672z218_BXINV_6434 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z218_BXINV
    );
  romedatao3_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_5_F5MUX,
      O => nx54672z245
    );
  romedatao3_s_5_F5MUX_6435 : X_MUX2
    port map (
      IA => nx54672z246,
      IB => nx54672z247,
      SEL => romedatao3_s_5_BXINV,
      O => romedatao3_s_5_F5MUX
    );
  romedatao3_s_5_BXINV_6436 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao3_s_5_BXINV
    );
  romedatao3_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_5_F6MUX,
      O => romedatao3_s(5)
    );
  romedatao3_s_5_F6MUX_6437 : X_MUX2
    port map (
      IA => nx54672z242,
      IB => nx54672z245,
      SEL => romedatao3_s_5_BYINV,
      O => romedatao3_s_5_F6MUX
    );
  romedatao3_s_5_BYINV_6438 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao3_s_5_BYINV
    );
  nx54672z242_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z242_F5MUX,
      O => nx54672z242
    );
  nx54672z242_F5MUX_6439 : X_MUX2
    port map (
      IA => nx54672z243,
      IB => nx54672z244,
      SEL => nx54672z242_BXINV,
      O => nx54672z242_F5MUX
    );
  nx54672z242_BXINV_6440 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z242_BXINV
    );
  U_DCT2D_ix43120z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_3_10_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_4_10_Q,
      O => U_DCT2D_nx43120z1
    );
  romedatao3_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_3_F5MUX,
      O => nx54672z256
    );
  romedatao3_s_3_F5MUX_6441 : X_MUX2
    port map (
      IA => nx54672z257,
      IB => nx54672z258,
      SEL => romedatao3_s_3_BXINV,
      O => romedatao3_s_3_F5MUX
    );
  romedatao3_s_3_BXINV_6442 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao3_s_3_BXINV
    );
  romedatao3_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao3_s_3_F6MUX,
      O => romedatao3_s(3)
    );
  romedatao3_s_3_F6MUX_6443 : X_MUX2
    port map (
      IA => nx54672z254,
      IB => nx54672z256,
      SEL => romedatao3_s_3_BYINV,
      O => romedatao3_s_3_F6MUX
    );
  romedatao3_s_3_BYINV_6444 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao3_s_3_BYINV
    );
  nx54672z254_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z254_F5MUX,
      O => nx54672z254
    );
  nx54672z254_F5MUX_6445 : X_MUX2
    port map (
      IA => U1_ROME3_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx54672z255,
      SEL => nx54672z254_BXINV,
      O => nx54672z254_F5MUX
    );
  nx54672z254_BXINV_6446 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z254_BXINV
    );
  romedatao6_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_6_F5MUX,
      O => nx54672z434
    );
  romedatao6_s_6_F5MUX_6447 : X_MUX2
    port map (
      IA => nx54672z435,
      IB => nx54672z436,
      SEL => romedatao6_s_6_BXINV,
      O => romedatao6_s_6_F5MUX
    );
  romedatao6_s_6_BXINV_6448 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao6_s_6_BXINV
    );
  romedatao6_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_6_F6MUX,
      O => romedatao6_s(6)
    );
  romedatao6_s_6_F6MUX_6449 : X_MUX2
    port map (
      IA => nx54672z431,
      IB => nx54672z434,
      SEL => romedatao6_s_6_BYINV,
      O => romedatao6_s_6_F6MUX
    );
  romedatao6_s_6_BYINV_6450 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao6_s_6_BYINV
    );
  nx54672z431_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z431_F5MUX,
      O => nx54672z431
    );
  nx54672z431_F5MUX_6451 : X_MUX2
    port map (
      IA => nx54672z432,
      IB => nx54672z433,
      SEL => nx54672z431_BXINV,
      O => nx54672z431_F5MUX
    );
  nx54672z431_BXINV_6452 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z431_BXINV
    );
  romedatao6_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_5_F5MUX,
      O => nx54672z440
    );
  romedatao6_s_5_F5MUX_6453 : X_MUX2
    port map (
      IA => nx54672z441,
      IB => nx54672z442,
      SEL => romedatao6_s_5_BXINV,
      O => romedatao6_s_5_F5MUX
    );
  romedatao6_s_5_BXINV_6454 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao6_s_5_BXINV
    );
  romedatao6_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao6_s_5_F6MUX,
      O => romedatao6_s(5)
    );
  romedatao6_s_5_F6MUX_6455 : X_MUX2
    port map (
      IA => nx54672z437,
      IB => nx54672z440,
      SEL => romedatao6_s_5_BYINV,
      O => romedatao6_s_5_F6MUX
    );
  romedatao6_s_5_BYINV_6456 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao6_s_5_BYINV
    );
  nx54672z437_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z437_F5MUX,
      O => nx54672z437
    );
  nx54672z437_F5MUX_6457 : X_MUX2
    port map (
      IA => nx54672z438,
      IB => nx54672z439,
      SEL => nx54672z437_BXINV,
      O => nx54672z437_F5MUX
    );
  nx54672z437_BXINV_6458 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z437_BXINV
    );
  romedatao8_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_8_F5MUX,
      O => nx54672z552
    );
  romedatao8_s_8_F5MUX_6459 : X_MUX2
    port map (
      IA => nx54672z553,
      IB => nx54672z554,
      SEL => romedatao8_s_8_BXINV,
      O => romedatao8_s_8_F5MUX
    );
  romedatao8_s_8_BXINV_6460 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao8_s_8_BXINV
    );
  romedatao8_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_8_F6MUX,
      O => romedatao8_s(8)
    );
  romedatao8_s_8_F6MUX_6461 : X_MUX2
    port map (
      IA => nx54672z549,
      IB => nx54672z552,
      SEL => romedatao8_s_8_BYINV,
      O => romedatao8_s_8_F6MUX
    );
  romedatao8_s_8_BYINV_6462 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao8_s_8_BYINV
    );
  nx54672z549_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z549_F5MUX,
      O => nx54672z549
    );
  nx54672z549_F5MUX_6463 : X_MUX2
    port map (
      IA => nx54672z550,
      IB => nx54672z551,
      SEL => nx54672z549_BXINV,
      O => nx54672z549_F5MUX
    );
  nx54672z549_BXINV_6464 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z549_BXINV
    );
  romedatao8_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_7_F5MUX,
      O => nx54672z558
    );
  romedatao8_s_7_F5MUX_6465 : X_MUX2
    port map (
      IA => nx54672z559,
      IB => nx54672z560,
      SEL => romedatao8_s_7_BXINV,
      O => romedatao8_s_7_F5MUX
    );
  romedatao8_s_7_BXINV_6466 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao8_s_7_BXINV
    );
  romedatao8_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_7_F6MUX,
      O => romedatao8_s(7)
    );
  romedatao8_s_7_F6MUX_6467 : X_MUX2
    port map (
      IA => nx54672z555,
      IB => nx54672z558,
      SEL => romedatao8_s_7_BYINV,
      O => romedatao8_s_7_F6MUX
    );
  romedatao8_s_7_BYINV_6468 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao8_s_7_BYINV
    );
  nx54672z555_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z555_F5MUX,
      O => nx54672z555
    );
  nx54672z555_F5MUX_6469 : X_MUX2
    port map (
      IA => nx54672z556,
      IB => nx54672z557,
      SEL => nx54672z555_BXINV,
      O => nx54672z555_F5MUX
    );
  nx54672z555_BXINV_6470 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z555_BXINV
    );
  romedatao8_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_6_F5MUX,
      O => nx54672z564
    );
  romedatao8_s_6_F5MUX_6471 : X_MUX2
    port map (
      IA => nx54672z565,
      IB => nx54672z566,
      SEL => romedatao8_s_6_BXINV,
      O => romedatao8_s_6_F5MUX
    );
  romedatao8_s_6_BXINV_6472 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao8_s_6_BXINV
    );
  romedatao8_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_6_F6MUX,
      O => romedatao8_s(6)
    );
  romedatao8_s_6_F6MUX_6473 : X_MUX2
    port map (
      IA => nx54672z561,
      IB => nx54672z564,
      SEL => romedatao8_s_6_BYINV,
      O => romedatao8_s_6_F6MUX
    );
  romedatao8_s_6_BYINV_6474 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao8_s_6_BYINV
    );
  nx54672z561_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z561_F5MUX,
      O => nx54672z561
    );
  nx54672z561_F5MUX_6475 : X_MUX2
    port map (
      IA => nx54672z562,
      IB => nx54672z563,
      SEL => nx54672z561_BXINV,
      O => nx54672z561_F5MUX
    );
  nx54672z561_BXINV_6476 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z561_BXINV
    );
  romedatao8_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_5_F5MUX,
      O => nx54672z570
    );
  romedatao8_s_5_F5MUX_6477 : X_MUX2
    port map (
      IA => nx54672z571,
      IB => nx54672z572,
      SEL => romedatao8_s_5_BXINV,
      O => romedatao8_s_5_F5MUX
    );
  romedatao8_s_5_BXINV_6478 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao8_s_5_BXINV
    );
  romedatao8_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_5_F6MUX,
      O => romedatao8_s(5)
    );
  romedatao8_s_5_F6MUX_6479 : X_MUX2
    port map (
      IA => nx54672z567,
      IB => nx54672z570,
      SEL => romedatao8_s_5_BYINV,
      O => romedatao8_s_5_F6MUX
    );
  romedatao8_s_5_BYINV_6480 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao8_s_5_BYINV
    );
  nx54672z567_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z567_F5MUX,
      O => nx54672z567
    );
  nx54672z567_F5MUX_6481 : X_MUX2
    port map (
      IA => nx54672z568,
      IB => nx54672z569,
      SEL => nx54672z567_BXINV,
      O => nx54672z567_F5MUX
    );
  nx54672z567_BXINV_6482 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z567_BXINV
    );
  romedatao8_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_4_F5MUX,
      O => nx54672z576
    );
  romedatao8_s_4_F5MUX_6483 : X_MUX2
    port map (
      IA => nx54672z577,
      IB => nx54672z578,
      SEL => romedatao8_s_4_BXINV,
      O => romedatao8_s_4_F5MUX
    );
  romedatao8_s_4_BXINV_6484 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao8_s_4_BXINV
    );
  romedatao8_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_4_F6MUX,
      O => romedatao8_s(4)
    );
  romedatao8_s_4_F6MUX_6485 : X_MUX2
    port map (
      IA => nx54672z573,
      IB => nx54672z576,
      SEL => romedatao8_s_4_BYINV,
      O => romedatao8_s_4_F6MUX
    );
  romedatao8_s_4_BYINV_6486 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao8_s_4_BYINV
    );
  nx54672z573_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z573_F5MUX,
      O => nx54672z573
    );
  nx54672z573_F5MUX_6487 : X_MUX2
    port map (
      IA => nx54672z574,
      IB => nx54672z575,
      SEL => nx54672z573_BXINV,
      O => nx54672z573_F5MUX
    );
  nx54672z573_BXINV_6488 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z573_BXINV
    );
  romodatao6_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_11_F5MUX,
      O => nx54672z1071
    );
  romodatao6_s_11_F5MUX_6489 : X_MUX2
    port map (
      IA => nx54672z1072,
      IB => nx54672z1073,
      SEL => romodatao6_s_11_BXINV,
      O => romodatao6_s_11_F5MUX
    );
  romodatao6_s_11_BXINV_6490 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_11_BXINV
    );
  romodatao6_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_11_F6MUX,
      O => romodatao6_s(11)
    );
  romodatao6_s_11_F6MUX_6491 : X_MUX2
    port map (
      IA => nx54672z1068,
      IB => nx54672z1071,
      SEL => romodatao6_s_11_BYINV,
      O => romodatao6_s_11_F6MUX
    );
  romodatao6_s_11_BYINV_6492 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_11_BYINV
    );
  nx54672z1068_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1068_F5MUX,
      O => nx54672z1068
    );
  nx54672z1068_F5MUX_6493 : X_MUX2
    port map (
      IA => nx54672z1069,
      IB => nx54672z1070,
      SEL => nx54672z1068_BXINV,
      O => nx54672z1068_F5MUX
    );
  nx54672z1068_BXINV_6494 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1068_BXINV
    );
  romodatao6_s_10_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_10_F5MUX,
      O => nx54672z1077
    );
  romodatao6_s_10_F5MUX_6495 : X_MUX2
    port map (
      IA => nx54672z1078,
      IB => nx54672z1079,
      SEL => romodatao6_s_10_BXINV,
      O => romodatao6_s_10_F5MUX
    );
  romodatao6_s_10_BXINV_6496 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_10_BXINV
    );
  romodatao6_s_10_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_10_F6MUX,
      O => romodatao6_s(10)
    );
  romodatao6_s_10_F6MUX_6497 : X_MUX2
    port map (
      IA => nx54672z1074,
      IB => nx54672z1077,
      SEL => romodatao6_s_10_BYINV,
      O => romodatao6_s_10_F6MUX
    );
  romodatao6_s_10_BYINV_6498 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_10_BYINV
    );
  nx54672z1074_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1074_F5MUX,
      O => nx54672z1074
    );
  nx54672z1074_F5MUX_6499 : X_MUX2
    port map (
      IA => nx54672z1075,
      IB => nx54672z1076,
      SEL => nx54672z1074_BXINV,
      O => nx54672z1074_F5MUX
    );
  nx54672z1074_BXINV_6500 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1074_BXINV
    );
  romodatao6_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_1_F5MUX,
      O => nx54672z1131
    );
  romodatao6_s_1_F5MUX_6501 : X_MUX2
    port map (
      IA => nx54672z1132,
      IB => nx54672z1133,
      SEL => romodatao6_s_1_BXINV,
      O => romodatao6_s_1_F5MUX
    );
  romodatao6_s_1_BXINV_6502 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_1_BXINV
    );
  romodatao6_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_1_F6MUX,
      O => romodatao6_s(1)
    );
  romodatao6_s_1_F6MUX_6503 : X_MUX2
    port map (
      IA => nx54672z1128,
      IB => nx54672z1131,
      SEL => romodatao6_s_1_BYINV,
      O => romodatao6_s_1_F6MUX
    );
  romodatao6_s_1_BYINV_6504 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_1_BYINV
    );
  nx54672z1128_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1128_F5MUX,
      O => nx54672z1128
    );
  nx54672z1128_F5MUX_6505 : X_MUX2
    port map (
      IA => nx54672z1129,
      IB => nx54672z1130,
      SEL => nx54672z1128_BXINV,
      O => nx54672z1128_F5MUX
    );
  nx54672z1128_BXINV_6506 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1128_BXINV
    );
  romedatao7_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_5_F5MUX,
      O => nx54672z505
    );
  romedatao7_s_5_F5MUX_6507 : X_MUX2
    port map (
      IA => nx54672z506,
      IB => nx54672z507,
      SEL => romedatao7_s_5_BXINV,
      O => romedatao7_s_5_F5MUX
    );
  romedatao7_s_5_BXINV_6508 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao7_s_5_BXINV
    );
  romedatao7_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_5_F6MUX,
      O => romedatao7_s(5)
    );
  romedatao7_s_5_F6MUX_6509 : X_MUX2
    port map (
      IA => nx54672z502,
      IB => nx54672z505,
      SEL => romedatao7_s_5_BYINV,
      O => romedatao7_s_5_F6MUX
    );
  romedatao7_s_5_BYINV_6510 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao7_s_5_BYINV
    );
  nx54672z502_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z502_F5MUX,
      O => nx54672z502
    );
  nx54672z502_F5MUX_6511 : X_MUX2
    port map (
      IA => nx54672z503,
      IB => nx54672z504,
      SEL => nx54672z502_BXINV,
      O => nx54672z502_F5MUX
    );
  nx54672z502_BXINV_6512 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z502_BXINV
    );
  romedatao7_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_4_F5MUX,
      O => nx54672z511
    );
  romedatao7_s_4_F5MUX_6513 : X_MUX2
    port map (
      IA => nx54672z512,
      IB => nx54672z513,
      SEL => romedatao7_s_4_BXINV,
      O => romedatao7_s_4_F5MUX
    );
  romedatao7_s_4_BXINV_6514 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao7_s_4_BXINV
    );
  romedatao7_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao7_s_4_F6MUX,
      O => romedatao7_s(4)
    );
  romedatao7_s_4_F6MUX_6515 : X_MUX2
    port map (
      IA => nx54672z508,
      IB => nx54672z511,
      SEL => romedatao7_s_4_BYINV,
      O => romedatao7_s_4_F6MUX
    );
  romedatao7_s_4_BYINV_6516 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao7_s_4_BYINV
    );
  nx54672z508_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z508_F5MUX,
      O => nx54672z508
    );
  nx54672z508_F5MUX_6517 : X_MUX2
    port map (
      IA => nx54672z509,
      IB => nx54672z510,
      SEL => nx54672z508_BXINV,
      O => nx54672z508_F5MUX
    );
  nx54672z508_BXINV_6518 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z508_BXINV
    );
  romodatao8_s_8_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_8_F5MUX,
      O => nx54672z1247
    );
  romodatao8_s_8_F5MUX_6519 : X_MUX2
    port map (
      IA => nx54672z1248,
      IB => nx54672z1249,
      SEL => romodatao8_s_8_BXINV,
      O => romodatao8_s_8_F5MUX
    );
  romodatao8_s_8_BXINV_6520 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_8_BXINV
    );
  romodatao8_s_8_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_8_F6MUX,
      O => romodatao8_s(8)
    );
  romodatao8_s_8_F6MUX_6521 : X_MUX2
    port map (
      IA => nx54672z1244,
      IB => nx54672z1247,
      SEL => romodatao8_s_8_BYINV,
      O => romodatao8_s_8_F6MUX
    );
  romodatao8_s_8_BYINV_6522 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_8_BYINV
    );
  nx54672z1244_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1244_F5MUX,
      O => nx54672z1244
    );
  nx54672z1244_F5MUX_6523 : X_MUX2
    port map (
      IA => nx54672z1245,
      IB => nx54672z1246,
      SEL => nx54672z1244_BXINV,
      O => nx54672z1244_F5MUX
    );
  nx54672z1244_BXINV_6524 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1244_BXINV
    );
  romodatao8_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_7_F5MUX,
      O => nx54672z1253
    );
  romodatao8_s_7_F5MUX_6525 : X_MUX2
    port map (
      IA => nx54672z1254,
      IB => nx54672z1255,
      SEL => romodatao8_s_7_BXINV,
      O => romodatao8_s_7_F5MUX
    );
  romodatao8_s_7_BXINV_6526 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_7_BXINV
    );
  romodatao8_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_7_F6MUX,
      O => romodatao8_s(7)
    );
  romodatao8_s_7_F6MUX_6527 : X_MUX2
    port map (
      IA => nx54672z1250,
      IB => nx54672z1253,
      SEL => romodatao8_s_7_BYINV,
      O => romodatao8_s_7_F6MUX
    );
  romodatao8_s_7_BYINV_6528 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_7_BYINV
    );
  nx54672z1250_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1250_F5MUX,
      O => nx54672z1250
    );
  nx54672z1250_F5MUX_6529 : X_MUX2
    port map (
      IA => nx54672z1251,
      IB => nx54672z1252,
      SEL => nx54672z1250_BXINV,
      O => nx54672z1250_F5MUX
    );
  nx54672z1250_BXINV_6530 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1250_BXINV
    );
  romodatao8_s_6_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_6_F5MUX,
      O => nx54672z1259
    );
  romodatao8_s_6_F5MUX_6531 : X_MUX2
    port map (
      IA => nx54672z1260,
      IB => nx54672z1261,
      SEL => romodatao8_s_6_BXINV,
      O => romodatao8_s_6_F5MUX
    );
  romodatao8_s_6_BXINV_6532 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_6_BXINV
    );
  romodatao8_s_6_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_6_F6MUX,
      O => romodatao8_s(6)
    );
  romodatao8_s_6_F6MUX_6533 : X_MUX2
    port map (
      IA => nx54672z1256,
      IB => nx54672z1259,
      SEL => romodatao8_s_6_BYINV,
      O => romodatao8_s_6_F6MUX
    );
  romodatao8_s_6_BYINV_6534 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_6_BYINV
    );
  nx54672z1256_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1256_F5MUX,
      O => nx54672z1256
    );
  nx54672z1256_F5MUX_6535 : X_MUX2
    port map (
      IA => nx54672z1257,
      IB => nx54672z1258,
      SEL => nx54672z1256_BXINV,
      O => nx54672z1256_F5MUX
    );
  nx54672z1256_BXINV_6536 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1256_BXINV
    );
  romodatao8_s_5_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_5_F5MUX,
      O => nx54672z1265
    );
  romodatao8_s_5_F5MUX_6537 : X_MUX2
    port map (
      IA => nx54672z1266,
      IB => nx54672z1267,
      SEL => romodatao8_s_5_BXINV,
      O => romodatao8_s_5_F5MUX
    );
  romodatao8_s_5_BXINV_6538 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_5_BXINV
    );
  romodatao8_s_5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_5_F6MUX,
      O => romodatao8_s(5)
    );
  romodatao8_s_5_F6MUX_6539 : X_MUX2
    port map (
      IA => nx54672z1262,
      IB => nx54672z1265,
      SEL => romodatao8_s_5_BYINV,
      O => romodatao8_s_5_F6MUX
    );
  romodatao8_s_5_BYINV_6540 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_5_BYINV
    );
  nx54672z1262_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1262_F5MUX,
      O => nx54672z1262
    );
  nx54672z1262_F5MUX_6541 : X_MUX2
    port map (
      IA => nx54672z1263,
      IB => nx54672z1264,
      SEL => nx54672z1262_BXINV,
      O => nx54672z1262_F5MUX
    );
  nx54672z1262_BXINV_6542 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1262_BXINV
    );
  U_DCT2D_reg_databuf_reg_7_9_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_7_8_DYMUX,
      CE => U_DCT2D_databuf_reg_7_8_CEINV,
      CLK => U_DCT2D_databuf_reg_7_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_7_8_FFY_RST,
      O => U_DCT2D_databuf_reg_7_Q(9)
    );
  U_DCT2D_databuf_reg_7_8_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_7_8_FFY_RST
    );
  romodatao8_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_4_F5MUX,
      O => nx54672z1271
    );
  romodatao8_s_4_F5MUX_6543 : X_MUX2
    port map (
      IA => nx54672z1272,
      IB => nx54672z1273,
      SEL => romodatao8_s_4_BXINV,
      O => romodatao8_s_4_F5MUX
    );
  romodatao8_s_4_BXINV_6544 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_4_BXINV
    );
  romodatao8_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_4_F6MUX,
      O => romodatao8_s(4)
    );
  romodatao8_s_4_F6MUX_6545 : X_MUX2
    port map (
      IA => nx54672z1268,
      IB => nx54672z1271,
      SEL => romodatao8_s_4_BYINV,
      O => romodatao8_s_4_F6MUX
    );
  romodatao8_s_4_BYINV_6546 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_4_BYINV
    );
  nx54672z1268_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1268_F5MUX,
      O => nx54672z1268
    );
  nx54672z1268_F5MUX_6547 : X_MUX2
    port map (
      IA => nx54672z1269,
      IB => nx54672z1270,
      SEL => nx54672z1268_BXINV,
      O => nx54672z1268_F5MUX
    );
  nx54672z1268_BXINV_6548 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1268_BXINV
    );
  romodatao7_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_13_F5MUX,
      O => nx54672z1138
    );
  romodatao7_s_13_F5MUX_6549 : X_MUX2
    port map (
      IA => nx54672z1139,
      IB => nx54672z1140,
      SEL => romodatao7_s_13_BXINV,
      O => romodatao7_s_13_F5MUX
    );
  romodatao7_s_13_BXINV_6550 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_13_BXINV
    );
  romodatao7_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_13_F6MUX,
      O => romodatao7_s(13)
    );
  romodatao7_s_13_F6MUX_6551 : X_MUX2
    port map (
      IA => nx54672z1136,
      IB => nx54672z1138,
      SEL => romodatao7_s_13_BYINV,
      O => romodatao7_s_13_F6MUX
    );
  romodatao7_s_13_BYINV_6552 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_13_BYINV
    );
  nx54672z1136_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1136_F5MUX,
      O => nx54672z1136
    );
  nx54672z1136_F5MUX_6553 : X_MUX2
    port map (
      IA => nx54672z1136_G,
      IB => nx54672z1137,
      SEL => nx54672z1136_BXINV,
      O => nx54672z1136_F5MUX
    );
  nx54672z1136_BXINV_6554 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1136_BXINV
    );
  romodatao7_s_12_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_12_F5MUX,
      O => nx54672z1144
    );
  romodatao7_s_12_F5MUX_6555 : X_MUX2
    port map (
      IA => nx54672z1145,
      IB => nx54672z1146,
      SEL => romodatao7_s_12_BXINV,
      O => romodatao7_s_12_F5MUX
    );
  romodatao7_s_12_BXINV_6556 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_12_BXINV
    );
  romodatao7_s_12_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_12_F6MUX,
      O => romodatao7_s(12)
    );
  romodatao7_s_12_F6MUX_6557 : X_MUX2
    port map (
      IA => nx54672z1141,
      IB => nx54672z1144,
      SEL => romodatao7_s_12_BYINV,
      O => romodatao7_s_12_F6MUX
    );
  romodatao7_s_12_BYINV_6558 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_12_BYINV
    );
  nx54672z1141_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1141_F5MUX,
      O => nx54672z1141
    );
  nx54672z1141_F5MUX_6559 : X_MUX2
    port map (
      IA => nx54672z1142,
      IB => nx54672z1143,
      SEL => nx54672z1141_BXINV,
      O => nx54672z1141_F5MUX
    );
  nx54672z1141_BXINV_6560 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1141_BXINV
    );
  romodatao7_s_4_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_4_F5MUX,
      O => nx54672z1192
    );
  romodatao7_s_4_F5MUX_6561 : X_MUX2
    port map (
      IA => nx54672z1193,
      IB => nx54672z1194,
      SEL => romodatao7_s_4_BXINV,
      O => romodatao7_s_4_F5MUX
    );
  romodatao7_s_4_BXINV_6562 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_4_BXINV
    );
  romodatao7_s_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_4_F6MUX,
      O => romodatao7_s(4)
    );
  romodatao7_s_4_F6MUX_6563 : X_MUX2
    port map (
      IA => nx54672z1189,
      IB => nx54672z1192,
      SEL => romodatao7_s_4_BYINV,
      O => romodatao7_s_4_F6MUX
    );
  romodatao7_s_4_BYINV_6564 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_4_BYINV
    );
  nx54672z1189_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1189_F5MUX,
      O => nx54672z1189
    );
  nx54672z1189_F5MUX_6565 : X_MUX2
    port map (
      IA => nx54672z1190,
      IB => nx54672z1191,
      SEL => nx54672z1189_BXINV,
      O => nx54672z1189_F5MUX
    );
  nx54672z1189_BXINV_6566 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1189_BXINV
    );
  romodatao7_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_3_F5MUX,
      O => nx54672z1198
    );
  romodatao7_s_3_F5MUX_6567 : X_MUX2
    port map (
      IA => nx54672z1199,
      IB => nx54672z1200,
      SEL => romodatao7_s_3_BXINV,
      O => romodatao7_s_3_F5MUX
    );
  romodatao7_s_3_BXINV_6568 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_3_BXINV
    );
  romodatao7_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_3_F6MUX,
      O => romodatao7_s(3)
    );
  romodatao7_s_3_F6MUX_6569 : X_MUX2
    port map (
      IA => nx54672z1195,
      IB => nx54672z1198,
      SEL => romodatao7_s_3_BYINV,
      O => romodatao7_s_3_F6MUX
    );
  romodatao7_s_3_BYINV_6570 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_3_BYINV
    );
  nx54672z1195_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1195_F5MUX,
      O => nx54672z1195
    );
  nx54672z1195_F5MUX_6571 : X_MUX2
    port map (
      IA => nx54672z1196,
      IB => nx54672z1197,
      SEL => nx54672z1195_BXINV,
      O => nx54672z1195_F5MUX
    );
  nx54672z1195_BXINV_6572 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1195_BXINV
    );
  U_DCT2D_ix42123z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_3_8_Q,
      ADR1 => U_DCT2D_latchbuf_reg_4_8_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx42123z1
    );
  romodatao7_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_2_F5MUX,
      O => nx54672z1204
    );
  romodatao7_s_2_F5MUX_6573 : X_MUX2
    port map (
      IA => nx54672z1205,
      IB => nx54672z1206,
      SEL => romodatao7_s_2_BXINV,
      O => romodatao7_s_2_F5MUX
    );
  romodatao7_s_2_BXINV_6574 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_2_BXINV
    );
  romodatao7_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_2_F6MUX,
      O => romodatao7_s(2)
    );
  romodatao7_s_2_F6MUX_6575 : X_MUX2
    port map (
      IA => nx54672z1201,
      IB => nx54672z1204,
      SEL => romodatao7_s_2_BYINV,
      O => romodatao7_s_2_F6MUX
    );
  romodatao7_s_2_BYINV_6576 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_2_BYINV
    );
  nx54672z1201_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1201_F5MUX,
      O => nx54672z1201
    );
  nx54672z1201_F5MUX_6577 : X_MUX2
    port map (
      IA => nx54672z1202,
      IB => nx54672z1203,
      SEL => nx54672z1201_BXINV,
      O => nx54672z1201_F5MUX
    );
  nx54672z1201_BXINV_6578 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1201_BXINV
    );
  romodatao7_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_1_F5MUX,
      O => nx54672z1210
    );
  romodatao7_s_1_F5MUX_6579 : X_MUX2
    port map (
      IA => nx54672z1211,
      IB => nx54672z1212,
      SEL => romodatao7_s_1_BXINV,
      O => romodatao7_s_1_F5MUX
    );
  romodatao7_s_1_BXINV_6580 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_1_BXINV
    );
  romodatao7_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_1_F6MUX,
      O => romodatao7_s(1)
    );
  romodatao7_s_1_F6MUX_6581 : X_MUX2
    port map (
      IA => nx54672z1207,
      IB => nx54672z1210,
      SEL => romodatao7_s_1_BYINV,
      O => romodatao7_s_1_F6MUX
    );
  romodatao7_s_1_BYINV_6582 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_1_BYINV
    );
  nx54672z1207_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1207_F5MUX,
      O => nx54672z1207
    );
  nx54672z1207_F5MUX_6583 : X_MUX2
    port map (
      IA => nx54672z1208,
      IB => nx54672z1209,
      SEL => nx54672z1207_BXINV,
      O => nx54672z1207_F5MUX
    );
  nx54672z1207_BXINV_6584 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1207_BXINV
    );
  romodatao7_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_0_F5MUX,
      O => U1_ROMO7_modgen_rom_ix0_nx_ro64_32_l
    );
  romodatao7_s_0_F5MUX_6585 : X_MUX2
    port map (
      IA => nx54672z1213,
      IB => nx54672z1214,
      SEL => romodatao7_s_0_BXINV,
      O => romodatao7_s_0_F5MUX
    );
  romodatao7_s_0_BXINV_6586 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao7_s_0_BXINV
    );
  romodatao7_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao7_s_0_F6MUX,
      O => romodatao7_s(0)
    );
  romodatao7_s_0_F6MUX_6587 : X_MUX2
    port map (
      IA => U1_ROMO7_modgen_rom_ix0_nx_ro64_32_u,
      IB => U1_ROMO7_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romodatao7_s_0_BYINV,
      O => romodatao7_s_0_F6MUX
    );
  romodatao7_s_0_BYINV_6588 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao7_s_0_BYINV
    );
  U1_ROMO7_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROMO7_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U1_ROMO7_modgen_rom_ix0_nx_ro64_32_u
    );
  U1_ROMO7_modgen_rom_ix0_nx_ro64_32_u_F5MUX_6589 : X_MUX2
    port map (
      IA => U1_ROMO7_modgen_rom_ix0_nx_rm64_16_u,
      IB => U1_ROMO7_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U1_ROMO7_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U1_ROMO7_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U1_ROMO7_modgen_rom_ix0_nx_ro64_32_u_BXINV_6590 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => U1_ROMO7_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romodatao6_s_0_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_0_F5MUX,
      O => U1_ROMO6_modgen_rom_ix0_nx_ro64_32_l
    );
  romodatao6_s_0_F5MUX_6591 : X_MUX2
    port map (
      IA => nx54672z1134,
      IB => nx54672z1135,
      SEL => romodatao6_s_0_BXINV,
      O => romodatao6_s_0_F5MUX
    );
  romodatao6_s_0_BXINV_6592 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao6_s_0_BXINV
    );
  romodatao6_s_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao6_s_0_F6MUX,
      O => romodatao6_s(0)
    );
  romodatao6_s_0_F6MUX_6593 : X_MUX2
    port map (
      IA => U1_ROMO6_modgen_rom_ix0_nx_ro64_32_u,
      IB => U1_ROMO6_modgen_rom_ix0_nx_ro64_32_l,
      SEL => romodatao6_s_0_BYINV,
      O => romodatao6_s_0_F6MUX
    );
  romodatao6_s_0_BYINV_6594 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao6_s_0_BYINV
    );
  U1_ROMO6_modgen_rom_ix0_nx_ro64_32_u_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U1_ROMO6_modgen_rom_ix0_nx_ro64_32_u_F5MUX,
      O => U1_ROMO6_modgen_rom_ix0_nx_ro64_32_u
    );
  U1_ROMO6_modgen_rom_ix0_nx_ro64_32_u_F5MUX_6595 : X_MUX2
    port map (
      IA => U1_ROMO6_modgen_rom_ix0_nx_rm64_16_u,
      IB => U1_ROMO6_modgen_rom_ix0_nx_rm64_16_l,
      SEL => U1_ROMO6_modgen_rom_ix0_nx_ro64_32_u_BXINV,
      O => U1_ROMO6_modgen_rom_ix0_nx_ro64_32_u_F5MUX
    );
  U1_ROMO6_modgen_rom_ix0_nx_ro64_32_u_BXINV_6596 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => U1_ROMO6_modgen_rom_ix0_nx_ro64_32_u_BXINV
    );
  romodatao4_s_11_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_11_F5MUX,
      O => nx54672z913
    );
  romodatao4_s_11_F5MUX_6597 : X_MUX2
    port map (
      IA => nx54672z914,
      IB => nx54672z915,
      SEL => romodatao4_s_11_BXINV,
      O => romodatao4_s_11_F5MUX
    );
  romodatao4_s_11_BXINV_6598 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao4_s_11_BXINV
    );
  romodatao4_s_11_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao4_s_11_F6MUX,
      O => romodatao4_s(11)
    );
  romodatao4_s_11_F6MUX_6599 : X_MUX2
    port map (
      IA => nx54672z910,
      IB => nx54672z913,
      SEL => romodatao4_s_11_BYINV,
      O => romodatao4_s_11_F6MUX
    );
  romodatao4_s_11_BYINV_6600 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao4_s_11_BYINV
    );
  nx54672z910_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z910_F5MUX,
      O => nx54672z910
    );
  nx54672z910_F5MUX_6601 : X_MUX2
    port map (
      IA => nx54672z911,
      IB => nx54672z912,
      SEL => nx54672z910_BXINV,
      O => nx54672z910_F5MUX
    );
  nx54672z910_BXINV_6602 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z910_BXINV
    );
  romodatao3_s_7_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_7_F5MUX,
      O => nx54672z858
    );
  romodatao3_s_7_F5MUX_6603 : X_MUX2
    port map (
      IA => nx54672z859,
      IB => nx54672z860,
      SEL => romodatao3_s_7_BXINV,
      O => romodatao3_s_7_F5MUX
    );
  romodatao3_s_7_BXINV_6604 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_7_BXINV
    );
  romodatao3_s_7_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_7_F6MUX,
      O => romodatao3_s(7)
    );
  romodatao3_s_7_F6MUX_6605 : X_MUX2
    port map (
      IA => nx54672z855,
      IB => nx54672z858,
      SEL => romodatao3_s_7_BYINV,
      O => romodatao3_s_7_F6MUX
    );
  romodatao3_s_7_BYINV_6606 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_7_BYINV
    );
  nx54672z855_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z855_F5MUX,
      O => nx54672z855
    );
  nx54672z855_F5MUX_6607 : X_MUX2
    port map (
      IA => nx54672z856,
      IB => nx54672z857,
      SEL => nx54672z855_BXINV,
      O => nx54672z855_F5MUX
    );
  nx54672z855_BXINV_6608 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z855_BXINV
    );
  romodatao3_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_3_F5MUX,
      O => nx54672z882
    );
  romodatao3_s_3_F5MUX_6609 : X_MUX2
    port map (
      IA => nx54672z883,
      IB => nx54672z884,
      SEL => romodatao3_s_3_BXINV,
      O => romodatao3_s_3_F5MUX
    );
  romodatao3_s_3_BXINV_6610 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_3_BXINV
    );
  romodatao3_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_3_F6MUX,
      O => romodatao3_s(3)
    );
  romodatao3_s_3_F6MUX_6611 : X_MUX2
    port map (
      IA => nx54672z879,
      IB => nx54672z882,
      SEL => romodatao3_s_3_BYINV,
      O => romodatao3_s_3_F6MUX
    );
  romodatao3_s_3_BYINV_6612 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_3_BYINV
    );
  nx54672z879_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z879_F5MUX,
      O => nx54672z879
    );
  nx54672z879_F5MUX_6613 : X_MUX2
    port map (
      IA => nx54672z880,
      IB => nx54672z881,
      SEL => nx54672z879_BXINV,
      O => nx54672z879_F5MUX
    );
  nx54672z879_BXINV_6614 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z879_BXINV
    );
  romodatao3_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_1_F5MUX,
      O => nx54672z894
    );
  romodatao3_s_1_F5MUX_6615 : X_MUX2
    port map (
      IA => nx54672z895,
      IB => nx54672z896,
      SEL => romodatao3_s_1_BXINV,
      O => romodatao3_s_1_F5MUX
    );
  romodatao3_s_1_BXINV_6616 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao3_s_1_BXINV
    );
  romodatao3_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao3_s_1_F6MUX,
      O => romodatao3_s(1)
    );
  romodatao3_s_1_F6MUX_6617 : X_MUX2
    port map (
      IA => nx54672z891,
      IB => nx54672z894,
      SEL => romodatao3_s_1_BYINV,
      O => romodatao3_s_1_F6MUX
    );
  romodatao3_s_1_BYINV_6618 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao3_s_1_BYINV
    );
  nx54672z891_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z891_F5MUX,
      O => nx54672z891
    );
  nx54672z891_F5MUX_6619 : X_MUX2
    port map (
      IA => nx54672z892,
      IB => nx54672z893,
      SEL => nx54672z891_BXINV,
      O => nx54672z891_F5MUX
    );
  nx54672z891_BXINV_6620 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z891_BXINV
    );
  romedatao8_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_3_F5MUX,
      O => nx54672z581
    );
  romedatao8_s_3_F5MUX_6621 : X_MUX2
    port map (
      IA => nx54672z582,
      IB => nx54672z583,
      SEL => romedatao8_s_3_BXINV,
      O => romedatao8_s_3_F5MUX
    );
  romedatao8_s_3_BXINV_6622 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => romedatao8_s_3_BXINV
    );
  romedatao8_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romedatao8_s_3_F6MUX,
      O => romedatao8_s(3)
    );
  romedatao8_s_3_F6MUX_6623 : X_MUX2
    port map (
      IA => nx54672z579,
      IB => nx54672z581,
      SEL => romedatao8_s_3_BYINV,
      O => romedatao8_s_3_F6MUX
    );
  romedatao8_s_3_BYINV_6624 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(5),
      O => romedatao8_s_3_BYINV
    );
  nx54672z579_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z579_F5MUX,
      O => nx54672z579
    );
  nx54672z579_F5MUX_6625 : X_MUX2
    port map (
      IA => U1_ROME8_modgen_rom_ix2_nx_rm64_16_u,
      IB => nx54672z580,
      SEL => nx54672z579_BXINV,
      O => nx54672z579_F5MUX
    );
  nx54672z579_BXINV_6626 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romeaddro0_s(4),
      O => nx54672z579_BXINV
    );
  romodatao8_s_13_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_13_F5MUX,
      O => nx54672z1217
    );
  romodatao8_s_13_F5MUX_6627 : X_MUX2
    port map (
      IA => nx54672z1218,
      IB => nx54672z1219,
      SEL => romodatao8_s_13_BXINV,
      O => romodatao8_s_13_F5MUX
    );
  romodatao8_s_13_BXINV_6628 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_13_BXINV
    );
  romodatao8_s_13_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_13_F6MUX,
      O => romodatao8_s(13)
    );
  romodatao8_s_13_F6MUX_6629 : X_MUX2
    port map (
      IA => nx54672z1215,
      IB => nx54672z1217,
      SEL => romodatao8_s_13_BYINV,
      O => romodatao8_s_13_F6MUX
    );
  romodatao8_s_13_BYINV_6630 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_13_BYINV
    );
  nx54672z1215_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1215_F5MUX,
      O => nx54672z1215
    );
  nx54672z1215_F5MUX_6631 : X_MUX2
    port map (
      IA => nx54672z1215_G,
      IB => nx54672z1216,
      SEL => nx54672z1215_BXINV,
      O => nx54672z1215_F5MUX
    );
  nx54672z1215_BXINV_6632 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1215_BXINV
    );
  U_DCT2D_reg_databuf_reg_7_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_7_8_DXMUX,
      CE => U_DCT2D_databuf_reg_7_8_CEINV,
      CLK => U_DCT2D_databuf_reg_7_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_7_8_FFX_RST,
      O => U_DCT2D_databuf_reg_7_Q(8)
    );
  U_DCT2D_databuf_reg_7_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_7_8_FFX_RST
    );
  romodatao8_s_3_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_3_F5MUX,
      O => nx54672z1277
    );
  romodatao8_s_3_F5MUX_6633 : X_MUX2
    port map (
      IA => nx54672z1278,
      IB => nx54672z1279,
      SEL => romodatao8_s_3_BXINV,
      O => romodatao8_s_3_F5MUX
    );
  romodatao8_s_3_BXINV_6634 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_3_BXINV
    );
  romodatao8_s_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_3_F6MUX,
      O => romodatao8_s(3)
    );
  romodatao8_s_3_F6MUX_6635 : X_MUX2
    port map (
      IA => nx54672z1274,
      IB => nx54672z1277,
      SEL => romodatao8_s_3_BYINV,
      O => romodatao8_s_3_F6MUX
    );
  romodatao8_s_3_BYINV_6636 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_3_BYINV
    );
  nx54672z1274_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1274_F5MUX,
      O => nx54672z1274
    );
  nx54672z1274_F5MUX_6637 : X_MUX2
    port map (
      IA => nx54672z1275,
      IB => nx54672z1276,
      SEL => nx54672z1274_BXINV,
      O => nx54672z1274_F5MUX
    );
  nx54672z1274_BXINV_6638 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1274_BXINV
    );
  romodatao8_s_2_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_2_F5MUX,
      O => nx54672z1283
    );
  romodatao8_s_2_F5MUX_6639 : X_MUX2
    port map (
      IA => nx54672z1284,
      IB => nx54672z1285,
      SEL => romodatao8_s_2_BXINV,
      O => romodatao8_s_2_F5MUX
    );
  romodatao8_s_2_BXINV_6640 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_2_BXINV
    );
  romodatao8_s_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_2_F6MUX,
      O => romodatao8_s(2)
    );
  romodatao8_s_2_F6MUX_6641 : X_MUX2
    port map (
      IA => nx54672z1280,
      IB => nx54672z1283,
      SEL => romodatao8_s_2_BYINV,
      O => romodatao8_s_2_F6MUX
    );
  romodatao8_s_2_BYINV_6642 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_2_BYINV
    );
  nx54672z1280_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1280_F5MUX,
      O => nx54672z1280
    );
  nx54672z1280_F5MUX_6643 : X_MUX2
    port map (
      IA => nx54672z1281,
      IB => nx54672z1282,
      SEL => nx54672z1280_BXINV,
      O => nx54672z1280_F5MUX
    );
  nx54672z1280_BXINV_6644 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1280_BXINV
    );
  romodatao8_s_1_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_1_F5MUX,
      O => nx54672z1289
    );
  romodatao8_s_1_F5MUX_6645 : X_MUX2
    port map (
      IA => nx54672z1290,
      IB => nx54672z1291,
      SEL => romodatao8_s_1_BXINV,
      O => romodatao8_s_1_F5MUX
    );
  romodatao8_s_1_BXINV_6646 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => romodatao8_s_1_BXINV
    );
  romodatao8_s_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romodatao8_s_1_F6MUX,
      O => romodatao8_s(1)
    );
  romodatao8_s_1_F6MUX_6647 : X_MUX2
    port map (
      IA => nx54672z1286,
      IB => nx54672z1289,
      SEL => romodatao8_s_1_BYINV,
      O => romodatao8_s_1_F6MUX
    );
  romodatao8_s_1_BYINV_6648 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(5),
      O => romodatao8_s_1_BYINV
    );
  nx54672z1286_F5USED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx54672z1286_F5MUX,
      O => nx54672z1286
    );
  nx54672z1286_F5MUX_6649 : X_MUX2
    port map (
      IA => nx54672z1287,
      IB => nx54672z1288,
      SEL => nx54672z1286_BXINV,
      O => nx54672z1286_F5MUX
    );
  nx54672z1286_BXINV_6650 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => romoaddro0_s(4),
      O => nx54672z1286_BXINV
    );
  dcto1_obuf_10_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto1_10_O,
      CTL => dcto1_10_ENABLE,
      O => dcto1(10)
    );
  dcto1_10_ENABLEINV : X_INV
    port map (
      I => dcto1_10_GTS_OR_T,
      O => dcto1_10_ENABLE
    );
  dcto1_10_GTS_OR_T_6651 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto1_10_GTS_OR_T
    );
  dcto1_obuf_11_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto1_11_O,
      CTL => dcto1_11_ENABLE,
      O => dcto1(11)
    );
  dcto1_11_ENABLEINV : X_INV
    port map (
      I => dcto1_11_GTS_OR_T,
      O => dcto1_11_ENABLE
    );
  dcto1_11_GTS_OR_T_6652 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto1_11_GTS_OR_T
    );
  clk_ibuf_IBUFG_6653 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk,
      O => clk_INBUF
    );
  idv_ibuf : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => idv,
      O => idv_INBUF
    );
  odv_obuf : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => odv_O,
      CTL => odv_ENABLE,
      O => odv
    );
  odv_ENABLEINV : X_INV
    port map (
      I => odv_GTS_OR_T,
      O => odv_ENABLE
    );
  odv_GTS_OR_T_6654 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => odv_GTS_OR_T
    );
  rst_ibuf : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst,
      O => rst_INBUF
    );
  odv1_obuf : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => odv1_O,
      CTL => odv1_ENABLE,
      O => odv1
    );
  odv1_ENABLEINV : X_INV
    port map (
      I => odv1_GTS_OR_T,
      O => odv1_ENABLE
    );
  odv1_GTS_OR_T_6655 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => odv1_GTS_OR_T
    );
  dcti_ibuf_0_Q : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti(0),
      O => dcti_0_INBUF
    );
  dcti_ibuf_1_Q : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti(1),
      O => dcti_1_INBUF
    );
  dcti_ibuf_2_Q : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti(2),
      O => dcti_2_INBUF
    );
  dcti_ibuf_3_Q : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti(3),
      O => dcti_3_INBUF
    );
  dcti_ibuf_4_Q : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti(4),
      O => dcti_4_INBUF
    );
  dcti_ibuf_5_Q : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti(5),
      O => dcti_5_INBUF
    );
  dcti_ibuf_6_Q : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti(6),
      O => dcti_6_INBUF
    );
  dcti_ibuf_7_Q : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti(7),
      O => dcti_7_INBUF
    );
  dcto_obuf_0_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_0_O,
      CTL => dcto_0_ENABLE,
      O => dcto(0)
    );
  dcto_0_ENABLEINV : X_INV
    port map (
      I => dcto_0_GTS_OR_T,
      O => dcto_0_ENABLE
    );
  dcto_0_GTS_OR_T_6656 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto_0_GTS_OR_T
    );
  dcto_obuf_1_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_1_O,
      CTL => dcto_1_ENABLE,
      O => dcto(1)
    );
  dcto_1_ENABLEINV : X_INV
    port map (
      I => dcto_1_GTS_OR_T,
      O => dcto_1_ENABLE
    );
  dcto_1_GTS_OR_T_6657 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto_1_GTS_OR_T
    );
  U_DCT2D_reg_databuf_reg_7_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_7_10_DXMUX,
      CE => U_DCT2D_databuf_reg_7_10_CEINV,
      CLK => U_DCT2D_databuf_reg_7_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_7_10_FFX_RST,
      O => U_DCT2D_databuf_reg_7_Q(10)
    );
  U_DCT2D_databuf_reg_7_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_7_10_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_7_10_FFX_RST
    );
  U_DCT2D_databuf_reg_7_10_FFX_RSTAND_6658 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_7_10_FFX_RSTAND
    );
  dcto_obuf_2_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_2_O,
      CTL => dcto_2_ENABLE,
      O => dcto(2)
    );
  dcto_2_ENABLEINV : X_INV
    port map (
      I => dcto_2_GTS_OR_T,
      O => dcto_2_ENABLE
    );
  dcto_2_GTS_OR_T_6659 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto_2_GTS_OR_T
    );
  dcto_obuf_3_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_3_O,
      CTL => dcto_3_ENABLE,
      O => dcto(3)
    );
  dcto_3_ENABLEINV : X_INV
    port map (
      I => dcto_3_GTS_OR_T,
      O => dcto_3_ENABLE
    );
  dcto_3_GTS_OR_T_6660 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto_3_GTS_OR_T
    );
  dcto_obuf_4_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_4_O,
      CTL => dcto_4_ENABLE,
      O => dcto(4)
    );
  dcto_4_ENABLEINV : X_INV
    port map (
      I => dcto_4_GTS_OR_T,
      O => dcto_4_ENABLE
    );
  dcto_4_GTS_OR_T_6661 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto_4_GTS_OR_T
    );
  dcto_obuf_5_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_5_O,
      CTL => dcto_5_ENABLE,
      O => dcto(5)
    );
  dcto_5_ENABLEINV : X_INV
    port map (
      I => dcto_5_GTS_OR_T,
      O => dcto_5_ENABLE
    );
  dcto_5_GTS_OR_T_6662 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto_5_GTS_OR_T
    );
  dcto_obuf_6_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_6_O,
      CTL => dcto_6_ENABLE,
      O => dcto(6)
    );
  dcto_6_ENABLEINV : X_INV
    port map (
      I => dcto_6_GTS_OR_T,
      O => dcto_6_ENABLE
    );
  dcto_6_GTS_OR_T_6663 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto_6_GTS_OR_T
    );
  dcto_obuf_7_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_7_O,
      CTL => dcto_7_ENABLE,
      O => dcto(7)
    );
  dcto_7_ENABLEINV : X_INV
    port map (
      I => dcto_7_GTS_OR_T,
      O => dcto_7_ENABLE
    );
  dcto_7_GTS_OR_T_6664 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto_7_GTS_OR_T
    );
  dcto_obuf_8_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_8_O,
      CTL => dcto_8_ENABLE,
      O => dcto(8)
    );
  dcto_8_ENABLEINV : X_INV
    port map (
      I => dcto_8_GTS_OR_T,
      O => dcto_8_ENABLE
    );
  dcto_8_GTS_OR_T_6665 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto_8_GTS_OR_T
    );
  dcto_obuf_9_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_9_O,
      CTL => dcto_9_ENABLE,
      O => dcto(9)
    );
  dcto_9_ENABLEINV : X_INV
    port map (
      I => dcto_9_GTS_OR_T,
      O => dcto_9_ENABLE
    );
  dcto_9_GTS_OR_T_6666 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto_9_GTS_OR_T
    );
  ready_obuf : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ready_O,
      CTL => ready_ENABLE,
      O => ready
    );
  ready_ENABLEINV : X_INV
    port map (
      I => ready_GTS_OR_T,
      O => ready_ENABLE
    );
  ready_GTS_OR_T_6667 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => ready_GTS_OR_T
    );
  dcto_obuf_10_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_10_O,
      CTL => dcto_10_ENABLE,
      O => dcto(10)
    );
  dcto_10_ENABLEINV : X_INV
    port map (
      I => dcto_10_GTS_OR_T,
      O => dcto_10_ENABLE
    );
  dcto_10_GTS_OR_T_6668 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto_10_GTS_OR_T
    );
  dcto_obuf_11_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_11_O,
      CTL => dcto_11_ENABLE,
      O => dcto(11)
    );
  dcto_11_ENABLEINV : X_INV
    port map (
      I => dcto_11_GTS_OR_T,
      O => dcto_11_ENABLE
    );
  dcto_11_GTS_OR_T_6669 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto_11_GTS_OR_T
    );
  dcto1_obuf_0_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto1_0_O,
      CTL => dcto1_0_ENABLE,
      O => dcto1(0)
    );
  dcto1_0_ENABLEINV : X_INV
    port map (
      I => dcto1_0_GTS_OR_T,
      O => dcto1_0_ENABLE
    );
  dcto1_0_GTS_OR_T_6670 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto1_0_GTS_OR_T
    );
  dcto1_obuf_1_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto1_1_O,
      CTL => dcto1_1_ENABLE,
      O => dcto1(1)
    );
  dcto1_1_ENABLEINV : X_INV
    port map (
      I => dcto1_1_GTS_OR_T,
      O => dcto1_1_ENABLE
    );
  dcto1_1_GTS_OR_T_6671 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto1_1_GTS_OR_T
    );
  dcto1_obuf_2_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto1_2_O,
      CTL => dcto1_2_ENABLE,
      O => dcto1(2)
    );
  dcto1_2_ENABLEINV : X_INV
    port map (
      I => dcto1_2_GTS_OR_T,
      O => dcto1_2_ENABLE
    );
  dcto1_2_GTS_OR_T_6672 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto1_2_GTS_OR_T
    );
  dcto1_obuf_3_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto1_3_O,
      CTL => dcto1_3_ENABLE,
      O => dcto1(3)
    );
  dcto1_3_ENABLEINV : X_INV
    port map (
      I => dcto1_3_GTS_OR_T,
      O => dcto1_3_ENABLE
    );
  dcto1_3_GTS_OR_T_6673 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto1_3_GTS_OR_T
    );
  U_DCT1D_ix418z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_1_Q(1),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_6_Q(1),
      O => U_DCT1D_nx418z1
    );
  dcto1_obuf_4_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto1_4_O,
      CTL => dcto1_4_ENABLE,
      O => dcto1(4)
    );
  dcto1_4_ENABLEINV : X_INV
    port map (
      I => dcto1_4_GTS_OR_T,
      O => dcto1_4_ENABLE
    );
  dcto1_4_GTS_OR_T_6674 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto1_4_GTS_OR_T
    );
  dcto1_obuf_5_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto1_5_O,
      CTL => dcto1_5_ENABLE,
      O => dcto1(5)
    );
  dcto1_5_ENABLEINV : X_INV
    port map (
      I => dcto1_5_GTS_OR_T,
      O => dcto1_5_ENABLE
    );
  dcto1_5_GTS_OR_T_6675 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto1_5_GTS_OR_T
    );
  dcto1_obuf_6_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto1_6_O,
      CTL => dcto1_6_ENABLE,
      O => dcto1(6)
    );
  dcto1_6_ENABLEINV : X_INV
    port map (
      I => dcto1_6_GTS_OR_T,
      O => dcto1_6_ENABLE
    );
  dcto1_6_GTS_OR_T_6676 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto1_6_GTS_OR_T
    );
  dcto1_obuf_7_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto1_7_O,
      CTL => dcto1_7_ENABLE,
      O => dcto1(7)
    );
  dcto1_7_ENABLEINV : X_INV
    port map (
      I => dcto1_7_GTS_OR_T,
      O => dcto1_7_ENABLE
    );
  dcto1_7_GTS_OR_T_6677 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto1_7_GTS_OR_T
    );
  dcto1_obuf_8_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto1_8_O,
      CTL => dcto1_8_ENABLE,
      O => dcto1(8)
    );
  dcto1_8_ENABLEINV : X_INV
    port map (
      I => dcto1_8_GTS_OR_T,
      O => dcto1_8_ENABLE
    );
  dcto1_8_GTS_OR_T_6678 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto1_8_GTS_OR_T
    );
  dcto1_obuf_9_Q : X_TRI_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto1_9_O,
      CTL => dcto1_9_ENABLE,
      O => dcto1(9)
    );
  dcto1_9_ENABLEINV : X_INV
    port map (
      I => dcto1_9_GTS_OR_T,
      O => dcto1_9_ENABLE
    );
  dcto1_9_GTS_OR_T_6679 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => GTS,
      O => dcto1_9_GTS_OR_T
    );
  clk_ibuf_BUFG : X_BUFGMUX
    port map (
      I0 => clk_ibuf_IBUFG,
      I1 => GND,
      S => clk_ibuf_BUFG_S_INVNOT,
      O => clk_int,
      GSR => GSR
    );
  clk_ibuf_BUFG_SINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_19,
      O => clk_ibuf_BUFG_S_INVNOT
    );
  U2_RAM_mem_ix3035z34088_SSRBINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_41,
      O => U2_RAM_mem_ix3035z34088_SSRB_INTNOT
    );
  U2_RAM_mem_ix3035z34088_SSRAINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_41,
      O => U2_RAM_mem_ix3035z34088_SSRA_INTNOT
    );
  U2_RAM_mem_ix3035z34088_WEBINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_40,
      O => U2_RAM_mem_ix3035z34088_WEB_INTNOT
    );
  U2_RAM_mem_ix3035z34088 : X_RAMB16_S18_S18
    generic map(
      INIT_A => X"00000",
      INIT_B => X"00000",
      SRVAL_A => X"00000",
      SRVAL_B => X"00000",
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      SETUP_ALL => 484 ps,
      SETUP_READ_FIRST => 484 ps
    )
    port map (
      CLKA => clk_int,
      CLKB => clk_int,
      ENA => GLOBAL_LOGIC1_40,
      ENB => GLOBAL_LOGIC1_40,
      SSRA => U2_RAM_mem_ix3035z34088_SSRA_INTNOT,
      SSRB => U2_RAM_mem_ix3035z34088_SSRB_INTNOT,
      WEA => nx1552z1,
      WEB => U2_RAM_mem_ix3035z34088_WEB_INTNOT,
      GSR => GSR,
      ADDRA(9) => GLOBAL_LOGIC0_1,
      ADDRA(8) => GLOBAL_LOGIC0_1,
      ADDRA(7) => GLOBAL_LOGIC0_1,
      ADDRA(6) => GLOBAL_LOGIC0_1,
      ADDRA(5) => ramwaddro_s(5),
      ADDRA(4) => ramwaddro_s(4),
      ADDRA(3) => ramwaddro_s(3),
      ADDRA(2) => ramwaddro_s(2),
      ADDRA(1) => ramwaddro_s(1),
      ADDRA(0) => ramwaddro_s(0),
      ADDRB(9) => GLOBAL_LOGIC0_1,
      ADDRB(8) => GLOBAL_LOGIC0_1,
      ADDRB(7) => GLOBAL_LOGIC0_1,
      ADDRB(6) => GLOBAL_LOGIC0_1,
      ADDRB(5) => ramraddro_s(5),
      ADDRB(4) => ramraddro_s(4),
      ADDRB(3) => ramraddro_s(3),
      ADDRB(2) => ramraddro_s(2),
      ADDRB(1) => ramraddro_s(1),
      ADDRB(0) => ramraddro_s(0),
      DIA(15) => GLOBAL_LOGIC0_1,
      DIA(14) => GLOBAL_LOGIC0_1,
      DIA(13) => GLOBAL_LOGIC0_1,
      DIA(12) => GLOBAL_LOGIC0_1,
      DIA(11) => GLOBAL_LOGIC0_1,
      DIA(10) => GLOBAL_LOGIC0_1,
      DIA(9) => ramdatai_s(9),
      DIA(8) => ramdatai_s(8),
      DIA(7) => ramdatai_s(7),
      DIA(6) => ramdatai_s(6),
      DIA(5) => ramdatai_s(5),
      DIA(4) => ramdatai_s(4),
      DIA(3) => ramdatai_s(3),
      DIA(2) => ramdatai_s(2),
      DIA(1) => ramdatai_s(1),
      DIA(0) => ramdatai_s(0),
      DIPA(1) => GLOBAL_LOGIC0_2,
      DIPA(0) => GLOBAL_LOGIC0_3,
      DIB(15) => U2_RAM_mem_ix3035z34088_DIB15,
      DIB(14) => U2_RAM_mem_ix3035z34088_DIB14,
      DIB(13) => U2_RAM_mem_ix3035z34088_DIB13,
      DIB(12) => U2_RAM_mem_ix3035z34088_DIB12,
      DIB(11) => U2_RAM_mem_ix3035z34088_DIB11,
      DIB(10) => U2_RAM_mem_ix3035z34088_DIB10,
      DIB(9) => U2_RAM_mem_ix3035z34088_DIB9,
      DIB(8) => U2_RAM_mem_ix3035z34088_DIB8,
      DIB(7) => U2_RAM_mem_ix3035z34088_DIB7,
      DIB(6) => U2_RAM_mem_ix3035z34088_DIB6,
      DIB(5) => U2_RAM_mem_ix3035z34088_DIB5,
      DIB(4) => U2_RAM_mem_ix3035z34088_DIB4,
      DIB(3) => U2_RAM_mem_ix3035z34088_DIB3,
      DIB(2) => U2_RAM_mem_ix3035z34088_DIB2,
      DIB(1) => U2_RAM_mem_ix3035z34088_DIB1,
      DIB(0) => U2_RAM_mem_ix3035z34088_DIB0,
      DIPB(1) => U2_RAM_mem_ix3035z34088_DIPB1,
      DIPB(0) => U2_RAM_mem_ix3035z34088_DIPB0,
      DOA(15) => U2_RAM_mem_ix3035z34088_DOA15,
      DOA(14) => U2_RAM_mem_ix3035z34088_DOA14,
      DOA(13) => U2_RAM_mem_ix3035z34088_DOA13,
      DOA(12) => U2_RAM_mem_ix3035z34088_DOA12,
      DOA(11) => U2_RAM_mem_ix3035z34088_DOA11,
      DOA(10) => U2_RAM_mem_ix3035z34088_DOA10,
      DOA(9) => U2_RAM_mem_ix3035z34088_DOA9,
      DOA(8) => U2_RAM_mem_ix3035z34088_DOA8,
      DOA(7) => U2_RAM_mem_ix3035z34088_DOA7,
      DOA(6) => U2_RAM_mem_ix3035z34088_DOA6,
      DOA(5) => U2_RAM_mem_ix3035z34088_DOA5,
      DOA(4) => U2_RAM_mem_ix3035z34088_DOA4,
      DOA(3) => U2_RAM_mem_ix3035z34088_DOA3,
      DOA(2) => U2_RAM_mem_ix3035z34088_DOA2,
      DOA(1) => U2_RAM_mem_ix3035z34088_DOA1,
      DOA(0) => U2_RAM_mem_ix3035z34088_DOA0,
      DOPA(1) => U2_RAM_mem_ix3035z34088_DOPA1,
      DOPA(0) => U2_RAM_mem_ix3035z34088_DOPA0,
      DOB(15) => U2_RAM_mem_ix3035z34088_DOB15,
      DOB(14) => U2_RAM_mem_ix3035z34088_DOB14,
      DOB(13) => U2_RAM_mem_ix3035z34088_DOB13,
      DOB(12) => U2_RAM_mem_ix3035z34088_DOB12,
      DOB(11) => U2_RAM_mem_ix3035z34088_DOB11,
      DOB(10) => U2_RAM_mem_ix3035z34088_DOB10,
      DOB(9) => ramdatao2_s(9),
      DOB(8) => ramdatao2_s(8),
      DOB(7) => ramdatao2_s(7),
      DOB(6) => ramdatao2_s(6),
      DOB(5) => ramdatao2_s(5),
      DOB(4) => ramdatao2_s(4),
      DOB(3) => ramdatao2_s(3),
      DOB(2) => ramdatao2_s(2),
      DOB(1) => ramdatao2_s(1),
      DOB(0) => ramdatao2_s(0),
      DOPB(1) => U2_RAM_mem_ix3035z34088_DOPB1,
      DOPB(0) => U2_RAM_mem_ix3035z34088_DOPB0
    );
  U1_RAM_mem_ix3035z34088_SSRBINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_43,
      O => U1_RAM_mem_ix3035z34088_SSRB_INTNOT
    );
  U1_RAM_mem_ix3035z34088_SSRAINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_43,
      O => U1_RAM_mem_ix3035z34088_SSRA_INTNOT
    );
  U1_RAM_mem_ix3035z34088_WEBINV : X_INV
    port map (
      I => GLOBAL_LOGIC1_42,
      O => U1_RAM_mem_ix3035z34088_WEB_INTNOT
    );
  U1_RAM_mem_ix3035z34088 : X_RAMB16_S18_S18
    generic map(
      INIT_A => X"00000",
      INIT_B => X"00000",
      SRVAL_A => X"00000",
      SRVAL_B => X"00000",
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      SETUP_ALL => 484 ps,
      SETUP_READ_FIRST => 484 ps
    )
    port map (
      CLKA => clk_int,
      CLKB => clk_int,
      ENA => GLOBAL_LOGIC1_42,
      ENB => GLOBAL_LOGIC1_42,
      SSRA => U1_RAM_mem_ix3035z34088_SSRA_INTNOT,
      SSRB => U1_RAM_mem_ix3035z34088_SSRB_INTNOT,
      WEA => nx21201z1,
      WEB => U1_RAM_mem_ix3035z34088_WEB_INTNOT,
      GSR => GSR,
      ADDRA(9) => GLOBAL_LOGIC0,
      ADDRA(8) => GLOBAL_LOGIC0,
      ADDRA(7) => GLOBAL_LOGIC0,
      ADDRA(6) => GLOBAL_LOGIC0,
      ADDRA(5) => ramwaddro_s(5),
      ADDRA(4) => ramwaddro_s(4),
      ADDRA(3) => ramwaddro_s(3),
      ADDRA(2) => ramwaddro_s(2),
      ADDRA(1) => ramwaddro_s(1),
      ADDRA(0) => ramwaddro_s(0),
      ADDRB(9) => GLOBAL_LOGIC0,
      ADDRB(8) => GLOBAL_LOGIC0,
      ADDRB(7) => GLOBAL_LOGIC0,
      ADDRB(6) => GLOBAL_LOGIC0,
      ADDRB(5) => ramraddro_s(5),
      ADDRB(4) => ramraddro_s(4),
      ADDRB(3) => ramraddro_s(3),
      ADDRB(2) => ramraddro_s(2),
      ADDRB(1) => ramraddro_s(1),
      ADDRB(0) => ramraddro_s(0),
      DIA(15) => GLOBAL_LOGIC0,
      DIA(14) => GLOBAL_LOGIC0,
      DIA(13) => GLOBAL_LOGIC0,
      DIA(12) => GLOBAL_LOGIC0,
      DIA(11) => GLOBAL_LOGIC0,
      DIA(10) => GLOBAL_LOGIC0,
      DIA(9) => ramdatai_s(9),
      DIA(8) => ramdatai_s(8),
      DIA(7) => ramdatai_s(7),
      DIA(6) => ramdatai_s(6),
      DIA(5) => ramdatai_s(5),
      DIA(4) => ramdatai_s(4),
      DIA(3) => ramdatai_s(3),
      DIA(2) => ramdatai_s(2),
      DIA(1) => ramdatai_s(1),
      DIA(0) => ramdatai_s(0),
      DIPA(1) => GLOBAL_LOGIC0_0,
      DIPA(0) => GLOBAL_LOGIC0_1,
      DIB(15) => U1_RAM_mem_ix3035z34088_DIB15,
      DIB(14) => U1_RAM_mem_ix3035z34088_DIB14,
      DIB(13) => U1_RAM_mem_ix3035z34088_DIB13,
      DIB(12) => U1_RAM_mem_ix3035z34088_DIB12,
      DIB(11) => U1_RAM_mem_ix3035z34088_DIB11,
      DIB(10) => U1_RAM_mem_ix3035z34088_DIB10,
      DIB(9) => U1_RAM_mem_ix3035z34088_DIB9,
      DIB(8) => U1_RAM_mem_ix3035z34088_DIB8,
      DIB(7) => U1_RAM_mem_ix3035z34088_DIB7,
      DIB(6) => U1_RAM_mem_ix3035z34088_DIB6,
      DIB(5) => U1_RAM_mem_ix3035z34088_DIB5,
      DIB(4) => U1_RAM_mem_ix3035z34088_DIB4,
      DIB(3) => U1_RAM_mem_ix3035z34088_DIB3,
      DIB(2) => U1_RAM_mem_ix3035z34088_DIB2,
      DIB(1) => U1_RAM_mem_ix3035z34088_DIB1,
      DIB(0) => U1_RAM_mem_ix3035z34088_DIB0,
      DIPB(1) => U1_RAM_mem_ix3035z34088_DIPB1,
      DIPB(0) => U1_RAM_mem_ix3035z34088_DIPB0,
      DOA(15) => U1_RAM_mem_ix3035z34088_DOA15,
      DOA(14) => U1_RAM_mem_ix3035z34088_DOA14,
      DOA(13) => U1_RAM_mem_ix3035z34088_DOA13,
      DOA(12) => U1_RAM_mem_ix3035z34088_DOA12,
      DOA(11) => U1_RAM_mem_ix3035z34088_DOA11,
      DOA(10) => U1_RAM_mem_ix3035z34088_DOA10,
      DOA(9) => U1_RAM_mem_ix3035z34088_DOA9,
      DOA(8) => U1_RAM_mem_ix3035z34088_DOA8,
      DOA(7) => U1_RAM_mem_ix3035z34088_DOA7,
      DOA(6) => U1_RAM_mem_ix3035z34088_DOA6,
      DOA(5) => U1_RAM_mem_ix3035z34088_DOA5,
      DOA(4) => U1_RAM_mem_ix3035z34088_DOA4,
      DOA(3) => U1_RAM_mem_ix3035z34088_DOA3,
      DOA(2) => U1_RAM_mem_ix3035z34088_DOA2,
      DOA(1) => U1_RAM_mem_ix3035z34088_DOA1,
      DOA(0) => U1_RAM_mem_ix3035z34088_DOA0,
      DOPA(1) => U1_RAM_mem_ix3035z34088_DOPA1,
      DOPA(0) => U1_RAM_mem_ix3035z34088_DOPA0,
      DOB(15) => U1_RAM_mem_ix3035z34088_DOB15,
      DOB(14) => U1_RAM_mem_ix3035z34088_DOB14,
      DOB(13) => U1_RAM_mem_ix3035z34088_DOB13,
      DOB(12) => U1_RAM_mem_ix3035z34088_DOB12,
      DOB(11) => U1_RAM_mem_ix3035z34088_DOB11,
      DOB(10) => U1_RAM_mem_ix3035z34088_DOB10,
      DOB(9) => ramdatao1_s(9),
      DOB(8) => ramdatao1_s(8),
      DOB(7) => ramdatao1_s(7),
      DOB(6) => ramdatao1_s(6),
      DOB(5) => ramdatao1_s(5),
      DOB(4) => ramdatao1_s(4),
      DOB(3) => ramdatao1_s(3),
      DOB(2) => ramdatao1_s(2),
      DOB(1) => ramdatao1_s(1),
      DOB(0) => ramdatao1_s(0),
      DOPB(1) => U1_RAM_mem_ix3035z34088_DOPB1,
      DOPB(0) => U1_RAM_mem_ix3035z34088_DOPB0
    );
  U_DBUFCTL_rtlc4n377_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_rtlc4n377_F5MUX,
      O => U_DBUFCTL_rtlc4n377
    );
  U_DBUFCTL_rtlc4n377_F5MUX_6680 : X_MUX2
    port map (
      IA => nx31259z1,
      IB => nx31259z2,
      SEL => U_DBUFCTL_rtlc4n377_BXINV,
      O => U_DBUFCTL_rtlc4n377_F5MUX
    );
  U_DBUFCTL_rtlc4n377_BXINV_6681 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_mem1_lock_reg,
      O => U_DBUFCTL_rtlc4n377_BXINV
    );
  U_DCT2D_ix1822z45600 : X_LUT4
    generic map(
      INIT => X"DDF0"
    )
    port map (
      ADR0 => U_DCT2D_NOT_rtlcs2,
      ADR1 => reqrdfail_s,
      ADR2 => requestrd_s,
      ADR3 => U_DCT2D_istate_reg(1),
      O => U_DCT2D_nx1822z1
    );
  U_DCT2D_rtlc2n584_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n584_F5MUX,
      O => U_DCT2D_rtlc2n584
    );
  U_DCT2D_rtlc2n584_F5MUX_6682 : X_MUX2
    port map (
      IA => U_DCT2D_nx1822z1,
      IB => U_DCT2D_nx1822z2,
      SEL => U_DCT2D_rtlc2n584_BXINV,
      O => U_DCT2D_rtlc2n584_F5MUX
    );
  U_DCT2D_rtlc2n584_BXINV_6683 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_istate_reg(0),
      O => U_DCT2D_rtlc2n584_BXINV
    );
  U_DCT2D_istate_reg_1_DXMUX_6684 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcn348,
      O => U_DCT2D_istate_reg_1_DXMUX
    );
  U_DCT2D_istate_reg_1_DYMUX_6685 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2_istate_reg_fsm_SS9_n171(0),
      O => U_DCT2D_istate_reg_1_DYMUX
    );
  U_DCT2D_istate_reg_1_SRINV_6686 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_istate_reg_1_SRINV
    );
  U_DCT2D_istate_reg_1_CLKINV_6687 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_istate_reg_1_CLKINV
    );
  U_DCT2D_istate_reg_1_CEINV_6688 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n584,
      O => U_DCT2D_istate_reg_1_CEINV
    );
  memswitchrd_s_DXMUX_6689 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => memswitchrd_s_FXMUX,
      O => memswitchrd_s_DXMUX
    );
  memswitchrd_s_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => memswitchrd_s_FXMUX,
      O => NOT_U_DBUFCTL_rtlc0n25
    );
  memswitchrd_s_FXMUX_6690 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => memswitchrd_s_F,
      O => memswitchrd_s_FXMUX
    );
  memswitchrd_s_CLKINV_6691 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => memswitchrd_s_CLKINV
    );
  memswitchrd_s_CEINV_6692 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_rtlc4n374,
      O => memswitchrd_s_CEINV
    );
  ramraddro_s_5_DXMUX_6693 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx51407z1,
      O => ramraddro_s_5_DXMUX
    );
  ramraddro_s_5_DYMUX_6694 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx50410z1,
      O => ramraddro_s_5_DYMUX
    );
  ramraddro_s_5_SRINV_6695 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramraddro_s_5_SRINV
    );
  ramraddro_s_5_CLKINV_6696 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramraddro_s_5_CLKINV
    );
  ramraddro_s_5_CEINV_6697 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n446,
      O => ramraddro_s_5_CEINV
    );
  memswitchwr_s_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => memswitchwr_s_F,
      O => U_DBUFCTL_rtlc4n202
    );
  memswitchwr_s_DYMUX_6698 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => memswitchwr_s_GYMUX,
      O => memswitchwr_s_DYMUX
    );
  memswitchwr_s_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => memswitchwr_s_GYMUX,
      O => U_DBUFCTL_rtlcn1
    );
  memswitchwr_s_GYMUX_6699 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => memswitchwr_s_G,
      O => memswitchwr_s_GYMUX
    );
  memswitchwr_s_CLKINV_6700 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => memswitchwr_s_CLKINV
    );
  memswitchwr_s_CEINV_6701 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_rtlc4n373,
      O => memswitchwr_s_CEINV
    );
  U_DBUFCTL_mem1_full_reg_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_mem1_full_reg_F,
      O => nx24581z1
    );
  U_DBUFCTL_mem1_full_reg_DYMUX_6702 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_mem1_full_reg_GYMUX,
      O => U_DBUFCTL_mem1_full_reg_DYMUX
    );
  U_DBUFCTL_mem1_full_reg_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_mem1_full_reg_GYMUX,
      O => U_DBUFCTL_rtlcn38
    );
  U_DBUFCTL_mem1_full_reg_GYMUX_6703 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_mem1_full_reg_G,
      O => U_DBUFCTL_mem1_full_reg_GYMUX
    );
  U_DBUFCTL_mem1_full_reg_CLKINV_6704 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DBUFCTL_mem1_full_reg_CLKINV
    );
  U_DBUFCTL_mem1_full_reg_CEINV_6705 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx24581z1,
      O => U_DBUFCTL_mem1_full_reg_CEINV
    );
  ix31259z50210 : X_LUT4
    generic map(
      INIT => X"F070"
    )
    port map (
      ADR0 => releasewr_s,
      ADR1 => U_DBUFCTL_mem1_lock_reg,
      ADR2 => U_DBUFCTL_rtlcn38,
      ADR3 => memswitchwr_s,
      O => U_DBUFCTL_rtlcn35
    );
  U_DBUFCTL_mem1_lock_reg_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_mem1_lock_reg_F,
      O => nx1552z1
    );
  U_DBUFCTL_mem1_lock_reg_DYMUX_6706 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_rtlcn35,
      O => U_DBUFCTL_mem1_lock_reg_DYMUX
    );
  U_DBUFCTL_mem1_lock_reg_CLKINV_6707 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DBUFCTL_mem1_lock_reg_CLKINV
    );
  U_DBUFCTL_mem1_lock_reg_CEINV_6708 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_rtlc4n377,
      O => U_DBUFCTL_mem1_lock_reg_CEINV
    );
  U_DBUFCTL_mem2_full_reg_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_mem2_full_reg_F,
      O => nx43562z1
    );
  U_DBUFCTL_mem2_full_reg_DYMUX_6709 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_mem2_full_reg_GYMUX,
      O => U_DBUFCTL_mem2_full_reg_DYMUX
    );
  U_DBUFCTL_mem2_full_reg_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_mem2_full_reg_GYMUX,
      O => U_DBUFCTL_rtlcn42
    );
  U_DBUFCTL_mem2_full_reg_GYMUX_6710 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_mem2_full_reg_G,
      O => U_DBUFCTL_mem2_full_reg_GYMUX
    );
  U_DBUFCTL_mem2_full_reg_CLKINV_6711 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DBUFCTL_mem2_full_reg_CLKINV
    );
  U_DBUFCTL_mem2_full_reg_CEINV_6712 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => nx43562z1,
      O => U_DBUFCTL_mem2_full_reg_CEINV
    );
  U_DBUFCTL_mem2_lock_reg_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_mem2_lock_reg_F,
      O => nx21201z1
    );
  U_DBUFCTL_mem2_lock_reg_DYMUX_6713 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_rtlcn76,
      O => U_DBUFCTL_mem2_lock_reg_DYMUX
    );
  U_DBUFCTL_mem2_lock_reg_CLKINV_6714 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DBUFCTL_mem2_lock_reg_CLKINV
    );
  U_DBUFCTL_mem2_lock_reg_CEINV_6715 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_rtlc4n378,
      O => U_DBUFCTL_mem2_lock_reg_CEINV
    );
  U_DCT2D_col_reg_2_DYMUX_6716 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx35453z1,
      O => U_DCT2D_col_reg_2_DYMUX
    );
  U_DCT2D_col_reg_2_CLKINV_6717 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_col_reg_2_CLKINV
    );
  U_DCT2D_col_reg_2_CEINV_6718 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => U_DCT2D_col_reg_2_CEINV
    );
  U_DCT1D_reg_databuf_reg_1_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_1_0_DYMUX,
      CE => U_DCT1D_databuf_reg_1_0_CEINV,
      CLK => U_DCT1D_databuf_reg_1_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_1_0_FFY_RST,
      O => U_DCT1D_databuf_reg_1_Q(1)
    );
  U_DCT1D_databuf_reg_1_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_1_0_FFY_RST
    );
  U_DCT1D_col_reg_2_DYMUX_6719 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx35453z1,
      O => U_DCT1D_col_reg_2_DYMUX
    );
  U_DCT1D_col_reg_2_CLKINV_6720 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_col_reg_2_CLKINV
    );
  U_DCT1D_col_reg_2_CEINV_6721 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => U_DCT1D_col_reg_2_CEINV
    );
  U_DCT1D_ready_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ready_F,
      O => U_DCT1D_rtlc2n465
    );
  U_DCT1D_ready_DYMUX_6722 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ready_GYMUX,
      O => U_DCT1D_ready_DYMUX
    );
  U_DCT1D_ready_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ready_GYMUX,
      O => U_DCT1D_rtlcn339
    );
  U_DCT1D_ready_GYMUX_6723 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_ready_G,
      O => U_DCT1D_ready_GYMUX
    );
  U_DCT1D_ready_CLKINV_6724 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_ready_CLKINV
    );
  U_DCT1D_ready_CEINV_6725 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_istate_reg(0),
      O => U_DCT1D_ready_CEINV
    );
  U_DCT1D_row_reg_2_DYMUX_6726 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx53037z1,
      O => U_DCT1D_row_reg_2_DYMUX
    );
  U_DCT1D_row_reg_2_CLKINV_6727 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_row_reg_2_CLKINV
    );
  U_DCT1D_row_reg_2_CEINV_6728 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcn1047,
      O => U_DCT1D_row_reg_2_CEINV
    );
  rome2addro0_s_5_DXMUX_6729 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_romeaddro0_SS3_n342(5),
      O => rome2addro0_s_5_DXMUX
    );
  rome2addro0_s_5_DYMUX_6730 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_romeaddro0_SS3_n342(4),
      O => rome2addro0_s_5_DYMUX
    );
  rome2addro0_s_5_SRINV_6731 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro0_s_5_SRINV
    );
  rome2addro0_s_5_CLKINV_6732 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro0_s_5_CLKINV
    );
  rome2addro0_s_5_CEINV_6733 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro0_s_5_CEINV
    );
  romeaddro0_s_5_DXMUX_6734 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_romeaddro0_SS4_n350(5),
      O => romeaddro0_s_5_DXMUX
    );
  romeaddro0_s_5_DYMUX_6735 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_romeaddro0_SS4_n350(4),
      O => romeaddro0_s_5_DYMUX
    );
  romeaddro0_s_5_SRINV_6736 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro0_s_5_SRINV
    );
  romeaddro0_s_5_CLKINV_6737 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro0_s_5_CLKINV
    );
  romeaddro0_s_5_CEINV_6738 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro0_s_5_CEINV
    );
  U_DCT2D_ix38901z4913 : X_LUT4
    generic map(
      INIT => X"5455"
    )
    port map (
      ADR0 => ramraddro_s(0),
      ADR1 => ramraddro_s(1),
      ADR2 => ramraddro_s(2),
      ADR3 => U_DCT2D_colram_reg(3),
      O => U_DCT2D_nx38901z1
    );
  ramraddro_s_0_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramraddro_s_0_F,
      O => U_DCT2D_rtlc2n576
    );
  ramraddro_s_0_DYMUX_6739 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx38901z1,
      O => ramraddro_s_0_DYMUX
    );
  ramraddro_s_0_CLKINV_6740 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramraddro_s_0_CLKINV
    );
  ramraddro_s_0_CEINV_6741 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_NOT_rtlc2n488,
      O => ramraddro_s_0_CEINV
    );
  ramraddro_s_1_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramraddro_s_1_F,
      O => U_DCT2D_nx39898z2
    );
  ramraddro_s_1_DYMUX_6742 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx39898z1,
      O => ramraddro_s_1_DYMUX
    );
  ramraddro_s_1_CLKINV_6743 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramraddro_s_1_CLKINV
    );
  ramraddro_s_1_CEINV_6744 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx39898z2,
      O => ramraddro_s_1_CEINV
    );
  ramraddro_s_2_DYMUX_6745 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx40895z1,
      O => ramraddro_s_2_DYMUX
    );
  ramraddro_s_2_CLKINV_6746 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramraddro_s_2_CLKINV
    );
  ramraddro_s_2_CEINV_6747 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx40895z2,
      O => ramraddro_s_2_CEINV
    );
  U_DCT1D_istate_reg_1_DXMUX_6748 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcn403,
      O => U_DCT1D_istate_reg_1_DXMUX
    );
  U_DCT1D_istate_reg_1_DYMUX_6749 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcn349,
      O => U_DCT1D_istate_reg_1_DYMUX
    );
  U_DCT1D_istate_reg_1_SRINV_6750 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_istate_reg_1_SRINV
    );
  U_DCT1D_istate_reg_1_CLKINV_6751 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_istate_reg_1_CLKINV
    );
  U_DCT1D_istate_reg_1_CEINV_6752 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n471,
      O => U_DCT1D_istate_reg_1_CEINV
    );
  U_DCT1D_inpcnt_reg_2_DYMUX_6753 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59993z1,
      O => U_DCT1D_inpcnt_reg_2_DYMUX
    );
  U_DCT1D_inpcnt_reg_2_CLKINV_6754 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_inpcnt_reg_2_CLKINV
    );
  U_DCT1D_inpcnt_reg_2_CEINV_6755 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n365,
      O => U_DCT1D_inpcnt_reg_2_CEINV
    );
  reqrdfail_s_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => reqrdfail_s_F,
      O => U_DBUFCTL_rtlc4n373
    );
  reqrdfail_s_DYMUX_6756 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_rtlcn7,
      O => reqrdfail_s_DYMUX
    );
  reqrdfail_s_CLKINV_6757 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => reqrdfail_s_CLKINV
    );
  reqrdfail_s_CEINV_6758 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => requestrd_s,
      O => reqrdfail_s_CEINV
    );
  reqwrfail_s_DYMUX_6759 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_rtlc4n197,
      O => reqwrfail_s_DYMUX
    );
  reqwrfail_s_CLKINV_6760 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => reqwrfail_s_CLKINV
    );
  reqwrfail_s_CEINV_6761 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => requestwr_s,
      O => reqwrfail_s_CEINV
    );
  U_DCT2D_latchbuf_reg_7_1_DXMUX_6762 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatao_s(1),
      O => U_DCT2D_latchbuf_reg_7_1_DXMUX
    );
  U_DCT2D_latchbuf_reg_7_1_DYMUX_6763 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatao_s(0),
      O => U_DCT2D_latchbuf_reg_7_1_DYMUX
    );
  U_DCT2D_latchbuf_reg_7_1_SRINV_6764 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_7_1_SRINV
    );
  U_DCT2D_latchbuf_reg_7_1_CLKINV_6765 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_7_1_CLKINV
    );
  U_DCT2D_latchbuf_reg_7_1_CEINV_6766 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_7_1_CEINV
    );
  U_DCT2D_latchbuf_reg_7_3_DXMUX_6767 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatao_s(3),
      O => U_DCT2D_latchbuf_reg_7_3_DXMUX
    );
  U_DCT2D_latchbuf_reg_7_3_DYMUX_6768 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatao_s(2),
      O => U_DCT2D_latchbuf_reg_7_3_DYMUX
    );
  U_DCT2D_latchbuf_reg_7_3_SRINV_6769 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_7_3_SRINV
    );
  U_DCT2D_latchbuf_reg_7_3_CLKINV_6770 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_7_3_CLKINV
    );
  U_DCT2D_latchbuf_reg_7_3_CEINV_6771 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_7_3_CEINV
    );
  U_DCT2D_latchbuf_reg_7_5_DXMUX_6772 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatao_s(5),
      O => U_DCT2D_latchbuf_reg_7_5_DXMUX
    );
  U_DCT2D_latchbuf_reg_7_5_DYMUX_6773 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatao_s(4),
      O => U_DCT2D_latchbuf_reg_7_5_DYMUX
    );
  U_DCT2D_latchbuf_reg_7_5_SRINV_6774 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_7_5_SRINV
    );
  U_DCT2D_latchbuf_reg_7_5_CLKINV_6775 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_7_5_CLKINV
    );
  U_DCT2D_latchbuf_reg_7_5_CEINV_6776 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_7_5_CEINV
    );
  U_DCT1D_ix64957z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_1_Q(0),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_6_Q(0),
      O => U_DCT1D_nx64957z1
    );
  U_DCT2D_latchbuf_reg_7_7_DXMUX_6777 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatao_s(7),
      O => U_DCT2D_latchbuf_reg_7_7_DXMUX
    );
  U_DCT2D_latchbuf_reg_7_7_DYMUX_6778 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatao_s(6),
      O => U_DCT2D_latchbuf_reg_7_7_DYMUX
    );
  U_DCT2D_latchbuf_reg_7_7_SRINV_6779 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_7_7_SRINV
    );
  U_DCT2D_latchbuf_reg_7_7_CLKINV_6780 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_7_7_CLKINV
    );
  U_DCT2D_latchbuf_reg_7_7_CEINV_6781 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_7_7_CEINV
    );
  U_DCT2D_latchbuf_reg_7_10_DXMUX_6782 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatao_s(9),
      O => U_DCT2D_latchbuf_reg_7_10_DXMUX
    );
  U_DCT2D_latchbuf_reg_7_10_DYMUX_6783 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatao_s(8),
      O => U_DCT2D_latchbuf_reg_7_10_DYMUX
    );
  U_DCT2D_latchbuf_reg_7_10_SRINV_6784 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_7_10_SRINV
    );
  U_DCT2D_latchbuf_reg_7_10_CLKINV_6785 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_7_10_CLKINV
    );
  U_DCT2D_latchbuf_reg_7_10_CEINV_6786 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_7_10_CEINV
    );
  U_DCT2D_nx65206z252_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z252_G,
      O => U_DCT2D_nx65206z252
    );
  U_DCT2D_nx65206z571_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z571_G,
      O => U_DCT2D_nx65206z571
    );
  U_DCT1D_rtlc2n469_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n469_F,
      O => U_DCT1D_rtlc2n469
    );
  U_DCT1D_rtlc2n469_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n469_G,
      O => U_DCT1D_rtlc2n365
    );
  U_DCT2D_nx65206z251_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z251_F,
      O => U_DCT2D_nx65206z251
    );
  U_DCT2D_nx65206z251_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z251_G,
      O => U_DCT2D_nx65206z250
    );
  U_DCT2D_nx65206z218_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z218_F,
      O => U_DCT2D_nx65206z218
    );
  U_DCT2D_nx65206z218_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z218_G,
      O => U_DCT2D_nx65206z4
    );
  ramraddro_s_3_DYMUX_6787 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramraddro_s_3_BYINVNOT,
      O => ramraddro_s_3_DYMUX
    );
  ramraddro_s_3_BYINV : X_INV
    port map (
      I => ramraddro_s(3),
      O => ramraddro_s_3_BYINVNOT
    );
  ramraddro_s_3_CLKINV_6788 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramraddro_s_3_CLKINV
    );
  ramraddro_s_3_CEINV_6789 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n446,
      O => ramraddro_s_3_CEINV
    );
  requestwr_s_DYMUX_6790 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => requestwr_s_BYINVNOT,
      O => requestwr_s_DYMUX
    );
  requestwr_s_BYINV : X_INV
    port map (
      I => requestwr_s,
      O => requestwr_s_BYINVNOT
    );
  requestwr_s_CLKINV_6791 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => requestwr_s_CLKINV
    );
  requestwr_s_CEINV_6792 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n469,
      O => requestwr_s_CEINV
    );
  U_DBUFCTL_rtlc4n378_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_rtlc4n378_F,
      O => U_DBUFCTL_rtlc4n378
    );
  U_DBUFCTL_rtlc4n378_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_rtlc4n378_G,
      O => nx43562z2
    );
  U_DBUFCTL_rtlc4n374_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DBUFCTL_rtlc4n374_G,
      O => U_DBUFCTL_rtlc4n374
    );
  U_DCT2D_rtlc5n1702_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702_F,
      O => U_DCT2D_rtlc5n1702
    );
  U_DCT2D_rtlc5n1702_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1702_G,
      O => U_DCT2D_rtlcn1678
    );
  U_DCT1D_state_reg_1_DXMUX_6793 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5_state_reg_fsm_SS4_n374(1),
      O => U_DCT1D_state_reg_1_DXMUX
    );
  U_DCT1D_state_reg_1_DYMUX_6794 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg_1_BYINVNOT,
      O => U_DCT1D_state_reg_1_DYMUX
    );
  U_DCT1D_state_reg_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg_1_G,
      O => U_DCT1D_NOT_rtlcs7
    );
  U_DCT1D_state_reg_1_BYINV : X_INV
    port map (
      I => U_DCT1D_state_reg(0),
      O => U_DCT1D_state_reg_1_BYINVNOT
    );
  U_DCT1D_state_reg_1_SRINV_6795 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_state_reg_1_SRINV
    );
  U_DCT1D_state_reg_1_CLKINV_6796 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_state_reg_1_CLKINV
    );
  U_DCT1D_state_reg_1_CEINV_6797 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1690,
      O => U_DCT1D_state_reg_1_CEINV
    );
  U_DCT2D_rtlc2n581_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n581_F,
      O => U_DCT2D_rtlc2n581
    );
  U_DCT2D_rtlc2n581_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n581_G,
      O => nx53675z1582
    );
  U_DCT2D_nx64938z1_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx64938z1_F,
      O => U_DCT2D_nx64938z1
    );
  U_DCT2D_nx64938z1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx64938z1_G,
      O => U_DCT2D_nx30550z1
    );
  U_DCT2D_rtlcs5_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5_F,
      O => U_DCT2D_rtlcs5
    );
  U_DCT2D_rtlcs5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5_G,
      O => U_DCT2D_rtlcn65
    );
  U_DCT2D_rtlc2n580_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n580_F,
      O => U_DCT2D_rtlc2n580
    );
  U_DCT2D_rtlc2n580_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n580_G,
      O => U_DCT2D_rtlc2n582
    );
  U_DCT2D_nx14976z1_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx14976z1_F,
      O => U_DCT2D_nx14976z1
    );
  U_DCT2D_nx14976z1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx14976z1_G,
      O => U_DCT2D_nx16172z1
    );
  U_DCT1D_reg_databuf_reg_1_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_1_0_DXMUX,
      CE => U_DCT1D_databuf_reg_1_0_CEINV,
      CLK => U_DCT1D_databuf_reg_1_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_1_0_FFX_RST,
      O => U_DCT1D_databuf_reg_1_Q(0)
    );
  U_DCT1D_databuf_reg_1_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_1_0_FFX_RST
    );
  U_DCT2D_col_reg_0_DXMUX_6798 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_col_reg_0_BXINVNOT,
      O => U_DCT2D_col_reg_0_DXMUX
    );
  U_DCT2D_col_reg_0_BXINV : X_INV
    port map (
      I => U_DCT2D_col_reg(0),
      O => U_DCT2D_col_reg_0_BXINVNOT
    );
  U_DCT2D_col_reg_0_DYMUX_6799 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx36450z1,
      O => U_DCT2D_col_reg_0_DYMUX
    );
  U_DCT2D_col_reg_0_SRINV_6800 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_col_reg_0_SRINV
    );
  U_DCT2D_col_reg_0_CLKINV_6801 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_col_reg_0_CLKINV
    );
  U_DCT2D_col_reg_0_CEINV_6802 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => U_DCT2D_col_reg_0_CEINV
    );
  U_DCT1D_col_reg_0_DXMUX_6803 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_col_reg_0_BXINVNOT,
      O => U_DCT1D_col_reg_0_DXMUX
    );
  U_DCT1D_col_reg_0_BXINV : X_INV
    port map (
      I => U_DCT1D_col_reg(0),
      O => U_DCT1D_col_reg_0_BXINVNOT
    );
  U_DCT1D_col_reg_0_DYMUX_6804 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx36450z1,
      O => U_DCT1D_col_reg_0_DYMUX
    );
  U_DCT1D_col_reg_0_SRINV_6805 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_col_reg_0_SRINV
    );
  U_DCT1D_col_reg_0_CLKINV_6806 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_col_reg_0_CLKINV
    );
  U_DCT1D_col_reg_0_CEINV_6807 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => U_DCT1D_col_reg_0_CEINV
    );
  U_DCT2D_nx8385z1_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx8385z1_F,
      O => U_DCT2D_nx8385z1
    );
  U_DCT2D_nx8385z1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx8385z1_G,
      O => U_DCT2D_nx22763z1
    );
  U_DCT1D_completed_reg_DYMUX_6808 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => U_DCT1D_completed_reg_DYMUX
    );
  U_DCT1D_completed_reg_CLKINV_6809 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_completed_reg_CLKINV
    );
  U_DCT1D_completed_reg_CEINV_6810 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1685,
      O => U_DCT1D_completed_reg_CEINV
    );
  U_DCT2D_nx38337z1_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx38337z1_F,
      O => U_DCT2D_nx38337z1
    );
  U_DCT2D_nx38337z1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx38337z1_G,
      O => U_DCT2D_nx7189z1
    );
  U_DCT1D_nx47258z1_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx47258z1_F,
      O => U_DCT1D_nx47258z1
    );
  U_DCT1D_nx47258z1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx47258z1_G,
      O => U_DCT1D_nx2262z1
    );
  U_DCT1D_ix2412z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_1_Q(3),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_6_Q(3),
      O => U_DCT1D_nx2412z1
    );
  U_DCT1D_latchbuf_reg_0_1_DXMUX_6811 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(1),
      O => U_DCT1D_latchbuf_reg_0_1_DXMUX
    );
  U_DCT1D_latchbuf_reg_0_1_DYMUX_6812 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(0),
      O => U_DCT1D_latchbuf_reg_0_1_DYMUX
    );
  U_DCT1D_latchbuf_reg_0_1_SRINV_6813 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_0_1_SRINV
    );
  U_DCT1D_latchbuf_reg_0_1_CLKINV_6814 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_0_1_CLKINV
    );
  U_DCT1D_latchbuf_reg_0_1_CEINV_6815 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_0_1_CEINV
    );
  U_DCT1D_latchbuf_reg_0_3_DXMUX_6816 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(3),
      O => U_DCT1D_latchbuf_reg_0_3_DXMUX
    );
  U_DCT1D_latchbuf_reg_0_3_DYMUX_6817 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(2),
      O => U_DCT1D_latchbuf_reg_0_3_DYMUX
    );
  U_DCT1D_latchbuf_reg_0_3_SRINV_6818 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_0_3_SRINV
    );
  U_DCT1D_latchbuf_reg_0_3_CLKINV_6819 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_0_3_CLKINV
    );
  U_DCT1D_latchbuf_reg_0_3_CEINV_6820 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_0_3_CEINV
    );
  U_DCT1D_latchbuf_reg_0_5_DXMUX_6821 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(5),
      O => U_DCT1D_latchbuf_reg_0_5_DXMUX
    );
  U_DCT1D_latchbuf_reg_0_5_DYMUX_6822 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(4),
      O => U_DCT1D_latchbuf_reg_0_5_DYMUX
    );
  U_DCT1D_latchbuf_reg_0_5_SRINV_6823 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_0_5_SRINV
    );
  U_DCT1D_latchbuf_reg_0_5_CLKINV_6824 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_0_5_CLKINV
    );
  U_DCT1D_latchbuf_reg_0_5_CEINV_6825 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_0_5_CEINV
    );
  U_DCT1D_latchbuf_reg_0_7_DXMUX_6826 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(7),
      O => U_DCT1D_latchbuf_reg_0_7_DXMUX
    );
  U_DCT1D_latchbuf_reg_0_7_DYMUX_6827 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_Q(6),
      O => U_DCT1D_latchbuf_reg_0_7_DYMUX
    );
  U_DCT1D_latchbuf_reg_0_7_SRINV_6828 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_0_7_SRINV
    );
  U_DCT1D_latchbuf_reg_0_7_CLKINV_6829 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_0_7_CLKINV
    );
  U_DCT1D_latchbuf_reg_0_7_CEINV_6830 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_0_7_CEINV
    );
  U_DCT1D_latchbuf_reg_1_1_DXMUX_6831 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(1),
      O => U_DCT1D_latchbuf_reg_1_1_DXMUX
    );
  U_DCT1D_latchbuf_reg_1_1_DYMUX_6832 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(0),
      O => U_DCT1D_latchbuf_reg_1_1_DYMUX
    );
  U_DCT1D_latchbuf_reg_1_1_SRINV_6833 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_1_1_SRINV
    );
  U_DCT1D_latchbuf_reg_1_1_CLKINV_6834 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_1_1_CLKINV
    );
  U_DCT1D_latchbuf_reg_1_1_CEINV_6835 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_1_1_CEINV
    );
  U_DCT1D_latchbuf_reg_1_3_DXMUX_6836 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(3),
      O => U_DCT1D_latchbuf_reg_1_3_DXMUX
    );
  U_DCT1D_latchbuf_reg_1_3_DYMUX_6837 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(2),
      O => U_DCT1D_latchbuf_reg_1_3_DYMUX
    );
  U_DCT1D_latchbuf_reg_1_3_SRINV_6838 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_1_3_SRINV
    );
  U_DCT1D_latchbuf_reg_1_3_CLKINV_6839 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_1_3_CLKINV
    );
  U_DCT1D_latchbuf_reg_1_3_CEINV_6840 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_1_3_CEINV
    );
  U_DCT1D_latchbuf_reg_1_5_DXMUX_6841 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(5),
      O => U_DCT1D_latchbuf_reg_1_5_DXMUX
    );
  U_DCT1D_latchbuf_reg_1_5_DYMUX_6842 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(4),
      O => U_DCT1D_latchbuf_reg_1_5_DYMUX
    );
  U_DCT1D_latchbuf_reg_1_5_SRINV_6843 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_1_5_SRINV
    );
  U_DCT1D_latchbuf_reg_1_5_CLKINV_6844 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_1_5_CLKINV
    );
  U_DCT1D_latchbuf_reg_1_5_CEINV_6845 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_1_5_CEINV
    );
  U_DCT1D_latchbuf_reg_1_7_DXMUX_6846 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(7),
      O => U_DCT1D_latchbuf_reg_1_7_DXMUX
    );
  U_DCT1D_latchbuf_reg_1_7_DYMUX_6847 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_Q(6),
      O => U_DCT1D_latchbuf_reg_1_7_DYMUX
    );
  U_DCT1D_latchbuf_reg_1_7_SRINV_6848 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_1_7_SRINV
    );
  U_DCT1D_latchbuf_reg_1_7_CLKINV_6849 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_1_7_CLKINV
    );
  U_DCT1D_latchbuf_reg_1_7_CEINV_6850 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_1_7_CEINV
    );
  U_DCT1D_latchbuf_reg_2_1_DXMUX_6851 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(1),
      O => U_DCT1D_latchbuf_reg_2_1_DXMUX
    );
  U_DCT1D_latchbuf_reg_2_1_DYMUX_6852 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(0),
      O => U_DCT1D_latchbuf_reg_2_1_DYMUX
    );
  U_DCT1D_latchbuf_reg_2_1_SRINV_6853 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_2_1_SRINV
    );
  U_DCT1D_latchbuf_reg_2_1_CLKINV_6854 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_2_1_CLKINV
    );
  U_DCT1D_latchbuf_reg_2_1_CEINV_6855 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_2_1_CEINV
    );
  U_DCT1D_latchbuf_reg_2_3_DXMUX_6856 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(3),
      O => U_DCT1D_latchbuf_reg_2_3_DXMUX
    );
  U_DCT1D_latchbuf_reg_2_3_DYMUX_6857 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(2),
      O => U_DCT1D_latchbuf_reg_2_3_DYMUX
    );
  U_DCT1D_latchbuf_reg_2_3_SRINV_6858 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_2_3_SRINV
    );
  U_DCT1D_latchbuf_reg_2_3_CLKINV_6859 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_2_3_CLKINV
    );
  U_DCT1D_latchbuf_reg_2_3_CEINV_6860 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_2_3_CEINV
    );
  U_DCT1D_latchbuf_reg_2_5_DXMUX_6861 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(5),
      O => U_DCT1D_latchbuf_reg_2_5_DXMUX
    );
  U_DCT1D_latchbuf_reg_2_5_DYMUX_6862 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(4),
      O => U_DCT1D_latchbuf_reg_2_5_DYMUX
    );
  U_DCT1D_latchbuf_reg_2_5_SRINV_6863 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_2_5_SRINV
    );
  U_DCT1D_latchbuf_reg_2_5_CLKINV_6864 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_2_5_CLKINV
    );
  U_DCT1D_latchbuf_reg_2_5_CEINV_6865 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_2_5_CEINV
    );
  romo2addro0_s_1_DXMUX_6866 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_Q(0),
      O => romo2addro0_s_1_DXMUX
    );
  romo2addro0_s_1_DYMUX_6867 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_Q(0),
      O => romo2addro0_s_1_DYMUX
    );
  romo2addro0_s_1_SRINV_6868 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro0_s_1_SRINV
    );
  romo2addro0_s_1_CLKINV_6869 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro0_s_1_CLKINV
    );
  romo2addro0_s_1_CEINV_6870 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro0_s_1_CEINV
    );
  U_DCT1D_latchbuf_reg_2_7_DXMUX_6871 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(7),
      O => U_DCT1D_latchbuf_reg_2_7_DXMUX
    );
  U_DCT1D_latchbuf_reg_2_7_DYMUX_6872 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_Q(6),
      O => U_DCT1D_latchbuf_reg_2_7_DYMUX
    );
  U_DCT1D_latchbuf_reg_2_7_SRINV_6873 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_2_7_SRINV
    );
  U_DCT1D_latchbuf_reg_2_7_CLKINV_6874 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_2_7_CLKINV
    );
  U_DCT1D_latchbuf_reg_2_7_CEINV_6875 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_2_7_CEINV
    );
  romo2addro0_s_3_DXMUX_6876 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_Q(0),
      O => romo2addro0_s_3_DXMUX
    );
  romo2addro0_s_3_DYMUX_6877 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_Q(0),
      O => romo2addro0_s_3_DYMUX
    );
  romo2addro0_s_3_SRINV_6878 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro0_s_3_SRINV
    );
  romo2addro0_s_3_CLKINV_6879 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro0_s_3_CLKINV
    );
  romo2addro0_s_3_CEINV_6880 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro0_s_3_CEINV
    );
  U_DCT1D_latchbuf_reg_3_1_DXMUX_6881 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_Q(1),
      O => U_DCT1D_latchbuf_reg_3_1_DXMUX
    );
  U_DCT1D_latchbuf_reg_3_1_DYMUX_6882 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_Q(0),
      O => U_DCT1D_latchbuf_reg_3_1_DYMUX
    );
  U_DCT1D_latchbuf_reg_3_1_SRINV_6883 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_3_1_SRINV
    );
  U_DCT1D_latchbuf_reg_3_1_CLKINV_6884 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_3_1_CLKINV
    );
  U_DCT1D_latchbuf_reg_3_1_CEINV_6885 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_3_1_CEINV
    );
  romo2addro1_s_1_DXMUX_6886 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_Q(1),
      O => romo2addro1_s_1_DXMUX
    );
  romo2addro1_s_1_DYMUX_6887 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_Q(1),
      O => romo2addro1_s_1_DYMUX
    );
  romo2addro1_s_1_SRINV_6888 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro1_s_1_SRINV
    );
  romo2addro1_s_1_CLKINV_6889 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro1_s_1_CLKINV
    );
  romo2addro1_s_1_CEINV_6890 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro1_s_1_CEINV
    );
  U_DCT1D_latchbuf_reg_3_3_DXMUX_6891 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_Q(3),
      O => U_DCT1D_latchbuf_reg_3_3_DXMUX
    );
  U_DCT1D_latchbuf_reg_3_3_DYMUX_6892 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_Q(2),
      O => U_DCT1D_latchbuf_reg_3_3_DYMUX
    );
  U_DCT1D_latchbuf_reg_3_3_SRINV_6893 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_3_3_SRINV
    );
  U_DCT1D_latchbuf_reg_3_3_CLKINV_6894 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_3_3_CLKINV
    );
  U_DCT1D_latchbuf_reg_3_3_CEINV_6895 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_3_3_CEINV
    );
  romo2addro1_s_3_DXMUX_6896 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_Q(1),
      O => romo2addro1_s_3_DXMUX
    );
  romo2addro1_s_3_DYMUX_6897 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_Q(1),
      O => romo2addro1_s_3_DYMUX
    );
  romo2addro1_s_3_SRINV_6898 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro1_s_3_SRINV
    );
  romo2addro1_s_3_CLKINV_6899 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro1_s_3_CLKINV
    );
  romo2addro1_s_3_CEINV_6900 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro1_s_3_CEINV
    );
  U_DCT1D_latchbuf_reg_3_5_DXMUX_6901 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_Q(5),
      O => U_DCT1D_latchbuf_reg_3_5_DXMUX
    );
  U_DCT1D_latchbuf_reg_3_5_DYMUX_6902 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_Q(4),
      O => U_DCT1D_latchbuf_reg_3_5_DYMUX
    );
  U_DCT1D_latchbuf_reg_3_5_SRINV_6903 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_3_5_SRINV
    );
  U_DCT1D_latchbuf_reg_3_5_CLKINV_6904 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_3_5_CLKINV
    );
  U_DCT1D_latchbuf_reg_3_5_CEINV_6905 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_3_5_CEINV
    );
  romo2addro2_s_1_DXMUX_6906 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_Q(2),
      O => romo2addro2_s_1_DXMUX
    );
  romo2addro2_s_1_DYMUX_6907 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_Q(2),
      O => romo2addro2_s_1_DYMUX
    );
  romo2addro2_s_1_SRINV_6908 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro2_s_1_SRINV
    );
  romo2addro2_s_1_CLKINV_6909 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro2_s_1_CLKINV
    );
  romo2addro2_s_1_CEINV_6910 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro2_s_1_CEINV
    );
  U_DCT1D_latchbuf_reg_3_7_DXMUX_6911 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_Q(7),
      O => U_DCT1D_latchbuf_reg_3_7_DXMUX
    );
  U_DCT1D_latchbuf_reg_3_7_DYMUX_6912 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_Q(6),
      O => U_DCT1D_latchbuf_reg_3_7_DYMUX
    );
  U_DCT1D_latchbuf_reg_3_7_SRINV_6913 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_3_7_SRINV
    );
  U_DCT1D_latchbuf_reg_3_7_CLKINV_6914 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_3_7_CLKINV
    );
  U_DCT1D_latchbuf_reg_3_7_CEINV_6915 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_3_7_CEINV
    );
  romo2addro2_s_3_DXMUX_6916 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_Q(2),
      O => romo2addro2_s_3_DXMUX
    );
  romo2addro2_s_3_DYMUX_6917 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_Q(2),
      O => romo2addro2_s_3_DYMUX
    );
  romo2addro2_s_3_SRINV_6918 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro2_s_3_SRINV
    );
  romo2addro2_s_3_CLKINV_6919 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro2_s_3_CLKINV
    );
  romo2addro2_s_3_CEINV_6920 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro2_s_3_CEINV
    );
  U_DCT1D_latchbuf_reg_4_1_DXMUX_6921 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_Q(1),
      O => U_DCT1D_latchbuf_reg_4_1_DXMUX
    );
  U_DCT1D_latchbuf_reg_4_1_DYMUX_6922 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_Q(0),
      O => U_DCT1D_latchbuf_reg_4_1_DYMUX
    );
  U_DCT1D_latchbuf_reg_4_1_SRINV_6923 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_4_1_SRINV
    );
  U_DCT1D_latchbuf_reg_4_1_CLKINV_6924 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_4_1_CLKINV
    );
  U_DCT1D_latchbuf_reg_4_1_CEINV_6925 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_4_1_CEINV
    );
  romo2addro3_s_1_DXMUX_6926 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_Q(3),
      O => romo2addro3_s_1_DXMUX
    );
  romo2addro3_s_1_DYMUX_6927 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_Q(3),
      O => romo2addro3_s_1_DYMUX
    );
  romo2addro3_s_1_SRINV_6928 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro3_s_1_SRINV
    );
  romo2addro3_s_1_CLKINV_6929 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro3_s_1_CLKINV
    );
  romo2addro3_s_1_CEINV_6930 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro3_s_1_CEINV
    );
  U_DCT1D_latchbuf_reg_4_3_DXMUX_6931 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_Q(3),
      O => U_DCT1D_latchbuf_reg_4_3_DXMUX
    );
  U_DCT1D_latchbuf_reg_4_3_DYMUX_6932 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_Q(2),
      O => U_DCT1D_latchbuf_reg_4_3_DYMUX
    );
  U_DCT1D_latchbuf_reg_4_3_SRINV_6933 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_4_3_SRINV
    );
  U_DCT1D_latchbuf_reg_4_3_CLKINV_6934 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_4_3_CLKINV
    );
  U_DCT1D_latchbuf_reg_4_3_CEINV_6935 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_4_3_CEINV
    );
  romo2addro3_s_3_DXMUX_6936 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_Q(3),
      O => romo2addro3_s_3_DXMUX
    );
  romo2addro3_s_3_DYMUX_6937 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_Q(3),
      O => romo2addro3_s_3_DYMUX
    );
  romo2addro3_s_3_SRINV_6938 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro3_s_3_SRINV
    );
  romo2addro3_s_3_CLKINV_6939 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro3_s_3_CLKINV
    );
  romo2addro3_s_3_CEINV_6940 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro3_s_3_CEINV
    );
  U_DCT1D_latchbuf_reg_4_5_DXMUX_6941 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_Q(5),
      O => U_DCT1D_latchbuf_reg_4_5_DXMUX
    );
  U_DCT1D_latchbuf_reg_4_5_DYMUX_6942 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_Q(4),
      O => U_DCT1D_latchbuf_reg_4_5_DYMUX
    );
  U_DCT1D_latchbuf_reg_4_5_SRINV_6943 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_4_5_SRINV
    );
  U_DCT1D_latchbuf_reg_4_5_CLKINV_6944 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_4_5_CLKINV
    );
  U_DCT1D_latchbuf_reg_4_5_CEINV_6945 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_4_5_CEINV
    );
  romo2addro4_s_1_DXMUX_6946 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_Q(4),
      O => romo2addro4_s_1_DXMUX
    );
  romo2addro4_s_1_DYMUX_6947 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_Q(4),
      O => romo2addro4_s_1_DYMUX
    );
  romo2addro4_s_1_SRINV_6948 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro4_s_1_SRINV
    );
  romo2addro4_s_1_CLKINV_6949 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro4_s_1_CLKINV
    );
  romo2addro4_s_1_CEINV_6950 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro4_s_1_CEINV
    );
  U_DCT1D_latchbuf_reg_4_7_DXMUX_6951 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_Q(7),
      O => U_DCT1D_latchbuf_reg_4_7_DXMUX
    );
  U_DCT1D_latchbuf_reg_4_7_DYMUX_6952 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_Q(6),
      O => U_DCT1D_latchbuf_reg_4_7_DYMUX
    );
  U_DCT1D_latchbuf_reg_4_7_SRINV_6953 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_4_7_SRINV
    );
  U_DCT1D_latchbuf_reg_4_7_CLKINV_6954 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_4_7_CLKINV
    );
  U_DCT1D_latchbuf_reg_4_7_CEINV_6955 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_4_7_CEINV
    );
  romo2addro4_s_3_DXMUX_6956 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_Q(4),
      O => romo2addro4_s_3_DXMUX
    );
  romo2addro4_s_3_DYMUX_6957 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_Q(4),
      O => romo2addro4_s_3_DYMUX
    );
  romo2addro4_s_3_SRINV_6958 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro4_s_3_SRINV
    );
  romo2addro4_s_3_CLKINV_6959 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro4_s_3_CLKINV
    );
  romo2addro4_s_3_CEINV_6960 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro4_s_3_CEINV
    );
  U_DCT1D_latchbuf_reg_5_1_DXMUX_6961 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_Q(1),
      O => U_DCT1D_latchbuf_reg_5_1_DXMUX
    );
  U_DCT1D_latchbuf_reg_5_1_DYMUX_6962 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_Q(0),
      O => U_DCT1D_latchbuf_reg_5_1_DYMUX
    );
  U_DCT1D_latchbuf_reg_5_1_SRINV_6963 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_5_1_SRINV
    );
  U_DCT1D_latchbuf_reg_5_1_CLKINV_6964 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_5_1_CLKINV
    );
  U_DCT1D_latchbuf_reg_5_1_CEINV_6965 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_5_1_CEINV
    );
  romo2addro5_s_1_DXMUX_6966 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_Q(5),
      O => romo2addro5_s_1_DXMUX
    );
  romo2addro5_s_1_DYMUX_6967 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_Q(5),
      O => romo2addro5_s_1_DYMUX
    );
  romo2addro5_s_1_SRINV_6968 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro5_s_1_SRINV
    );
  romo2addro5_s_1_CLKINV_6969 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro5_s_1_CLKINV
    );
  romo2addro5_s_1_CEINV_6970 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro5_s_1_CEINV
    );
  U_DCT1D_reg_databuf_reg_1_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_1_2_DYMUX,
      CE => U_DCT1D_databuf_reg_1_2_CEINV,
      CLK => U_DCT1D_databuf_reg_1_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_1_2_FFY_RST,
      O => U_DCT1D_databuf_reg_1_Q(3)
    );
  U_DCT1D_databuf_reg_1_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_1_2_FFY_RST
    );
  U_DCT1D_latchbuf_reg_5_3_DXMUX_6971 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_Q(3),
      O => U_DCT1D_latchbuf_reg_5_3_DXMUX
    );
  U_DCT1D_latchbuf_reg_5_3_DYMUX_6972 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_Q(2),
      O => U_DCT1D_latchbuf_reg_5_3_DYMUX
    );
  U_DCT1D_latchbuf_reg_5_3_SRINV_6973 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_5_3_SRINV
    );
  U_DCT1D_latchbuf_reg_5_3_CLKINV_6974 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_5_3_CLKINV
    );
  U_DCT1D_latchbuf_reg_5_3_CEINV_6975 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_5_3_CEINV
    );
  romo2addro5_s_3_DXMUX_6976 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_Q(5),
      O => romo2addro5_s_3_DXMUX
    );
  romo2addro5_s_3_DYMUX_6977 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_Q(5),
      O => romo2addro5_s_3_DYMUX
    );
  romo2addro5_s_3_SRINV_6978 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro5_s_3_SRINV
    );
  romo2addro5_s_3_CLKINV_6979 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro5_s_3_CLKINV
    );
  romo2addro5_s_3_CEINV_6980 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro5_s_3_CEINV
    );
  U_DCT1D_latchbuf_reg_5_5_DXMUX_6981 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_Q(5),
      O => U_DCT1D_latchbuf_reg_5_5_DXMUX
    );
  U_DCT1D_latchbuf_reg_5_5_DYMUX_6982 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_Q(4),
      O => U_DCT1D_latchbuf_reg_5_5_DYMUX
    );
  U_DCT1D_latchbuf_reg_5_5_SRINV_6983 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_5_5_SRINV
    );
  U_DCT1D_latchbuf_reg_5_5_CLKINV_6984 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_5_5_CLKINV
    );
  U_DCT1D_latchbuf_reg_5_5_CEINV_6985 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_5_5_CEINV
    );
  romo2addro6_s_1_DXMUX_6986 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_Q(6),
      O => romo2addro6_s_1_DXMUX
    );
  romo2addro6_s_1_DYMUX_6987 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_Q(6),
      O => romo2addro6_s_1_DYMUX
    );
  romo2addro6_s_1_SRINV_6988 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro6_s_1_SRINV
    );
  romo2addro6_s_1_CLKINV_6989 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro6_s_1_CLKINV
    );
  romo2addro6_s_1_CEINV_6990 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro6_s_1_CEINV
    );
  U_DCT1D_latchbuf_reg_5_7_DXMUX_6991 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_Q(7),
      O => U_DCT1D_latchbuf_reg_5_7_DXMUX
    );
  U_DCT1D_latchbuf_reg_5_7_DYMUX_6992 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_Q(6),
      O => U_DCT1D_latchbuf_reg_5_7_DYMUX
    );
  U_DCT1D_latchbuf_reg_5_7_SRINV_6993 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_5_7_SRINV
    );
  U_DCT1D_latchbuf_reg_5_7_CLKINV_6994 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_5_7_CLKINV
    );
  U_DCT1D_latchbuf_reg_5_7_CEINV_6995 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_5_7_CEINV
    );
  romo2addro6_s_3_DXMUX_6996 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_Q(6),
      O => romo2addro6_s_3_DXMUX
    );
  romo2addro6_s_3_DYMUX_6997 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_Q(6),
      O => romo2addro6_s_3_DYMUX
    );
  romo2addro6_s_3_SRINV_6998 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro6_s_3_SRINV
    );
  romo2addro6_s_3_CLKINV_6999 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro6_s_3_CLKINV
    );
  romo2addro6_s_3_CEINV_7000 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro6_s_3_CEINV
    );
  U_DCT1D_latchbuf_reg_6_1_DXMUX_7001 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_7_Q(1),
      O => U_DCT1D_latchbuf_reg_6_1_DXMUX
    );
  U_DCT1D_latchbuf_reg_6_1_DYMUX_7002 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_7_Q(0),
      O => U_DCT1D_latchbuf_reg_6_1_DYMUX
    );
  U_DCT1D_latchbuf_reg_6_1_SRINV_7003 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_6_1_SRINV
    );
  U_DCT1D_latchbuf_reg_6_1_CLKINV_7004 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_6_1_CLKINV
    );
  U_DCT1D_latchbuf_reg_6_1_CEINV_7005 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_6_1_CEINV
    );
  romo2addro7_s_1_DXMUX_7006 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_Q(7),
      O => romo2addro7_s_1_DXMUX
    );
  romo2addro7_s_1_DYMUX_7007 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_Q(7),
      O => romo2addro7_s_1_DYMUX
    );
  romo2addro7_s_1_SRINV_7008 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro7_s_1_SRINV
    );
  romo2addro7_s_1_CLKINV_7009 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro7_s_1_CLKINV
    );
  romo2addro7_s_1_CEINV_7010 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro7_s_1_CEINV
    );
  U_DCT1D_latchbuf_reg_6_3_DXMUX_7011 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_7_Q(3),
      O => U_DCT1D_latchbuf_reg_6_3_DXMUX
    );
  U_DCT1D_latchbuf_reg_6_3_DYMUX_7012 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_7_Q(2),
      O => U_DCT1D_latchbuf_reg_6_3_DYMUX
    );
  U_DCT1D_latchbuf_reg_6_3_SRINV_7013 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_6_3_SRINV
    );
  U_DCT1D_latchbuf_reg_6_3_CLKINV_7014 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_6_3_CLKINV
    );
  U_DCT1D_latchbuf_reg_6_3_CEINV_7015 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_6_3_CEINV
    );
  romo2addro7_s_3_DXMUX_7016 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_Q(7),
      O => romo2addro7_s_3_DXMUX
    );
  romo2addro7_s_3_DYMUX_7017 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_Q(7),
      O => romo2addro7_s_3_DYMUX
    );
  romo2addro7_s_3_SRINV_7018 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro7_s_3_SRINV
    );
  romo2addro7_s_3_CLKINV_7019 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro7_s_3_CLKINV
    );
  romo2addro7_s_3_CEINV_7020 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro7_s_3_CEINV
    );
  U_DCT1D_latchbuf_reg_6_5_DXMUX_7021 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_7_Q(5),
      O => U_DCT1D_latchbuf_reg_6_5_DXMUX
    );
  U_DCT1D_latchbuf_reg_6_5_DYMUX_7022 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_7_Q(4),
      O => U_DCT1D_latchbuf_reg_6_5_DYMUX
    );
  U_DCT1D_latchbuf_reg_6_5_SRINV_7023 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_6_5_SRINV
    );
  U_DCT1D_latchbuf_reg_6_5_CLKINV_7024 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_6_5_CLKINV
    );
  U_DCT1D_latchbuf_reg_6_5_CEINV_7025 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_6_5_CEINV
    );
  romo2addro8_s_1_DXMUX_7026 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_Q(8),
      O => romo2addro8_s_1_DXMUX
    );
  romo2addro8_s_1_DYMUX_7027 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_Q(8),
      O => romo2addro8_s_1_DYMUX
    );
  romo2addro8_s_1_SRINV_7028 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro8_s_1_SRINV
    );
  romo2addro8_s_1_CLKINV_7029 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro8_s_1_CLKINV
    );
  romo2addro8_s_1_CEINV_7030 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro8_s_1_CEINV
    );
  U_DCT1D_ix1415z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_1_Q(2),
      ADR1 => U_DCT1D_latchbuf_reg_6_Q(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx1415z1
    );
  U_DCT1D_latchbuf_reg_6_7_DXMUX_7031 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_7_Q(7),
      O => U_DCT1D_latchbuf_reg_6_7_DXMUX
    );
  U_DCT1D_latchbuf_reg_6_7_DYMUX_7032 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_7_Q(6),
      O => U_DCT1D_latchbuf_reg_6_7_DYMUX
    );
  U_DCT1D_latchbuf_reg_6_7_SRINV_7033 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_6_7_SRINV
    );
  U_DCT1D_latchbuf_reg_6_7_CLKINV_7034 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_6_7_CLKINV
    );
  U_DCT1D_latchbuf_reg_6_7_CEINV_7035 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_6_7_CEINV
    );
  romo2addro8_s_3_DXMUX_7036 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_Q(8),
      O => romo2addro8_s_3_DXMUX
    );
  romo2addro8_s_3_DYMUX_7037 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_Q(8),
      O => romo2addro8_s_3_DYMUX
    );
  romo2addro8_s_3_SRINV_7038 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro8_s_3_SRINV
    );
  romo2addro8_s_3_CLKINV_7039 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro8_s_3_CLKINV
    );
  romo2addro8_s_3_CEINV_7040 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro8_s_3_CEINV
    );
  romo2addro9_s_1_DXMUX_7041 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_Q(9),
      O => romo2addro9_s_1_DXMUX
    );
  romo2addro9_s_1_DYMUX_7042 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_Q(9),
      O => romo2addro9_s_1_DYMUX
    );
  romo2addro9_s_1_SRINV_7043 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro9_s_1_SRINV
    );
  romo2addro9_s_1_CLKINV_7044 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro9_s_1_CLKINV
    );
  romo2addro9_s_1_CEINV_7045 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro9_s_1_CEINV
    );
  romo2addro9_s_3_DXMUX_7046 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_Q(9),
      O => romo2addro9_s_3_DXMUX
    );
  romo2addro9_s_3_DYMUX_7047 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_Q(9),
      O => romo2addro9_s_3_DYMUX
    );
  romo2addro9_s_3_SRINV_7048 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro9_s_3_SRINV
    );
  romo2addro9_s_3_CLKINV_7049 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro9_s_3_CLKINV
    );
  romo2addro9_s_3_CEINV_7050 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro9_s_3_CEINV
    );
  U_DCT1D_latchbuf_reg_7_7_DYMUX_7051 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latchbuf_reg_7_7_BYINVNOT,
      O => U_DCT1D_latchbuf_reg_7_7_DYMUX
    );
  U_DCT1D_latchbuf_reg_7_7_BYINV : X_INV
    port map (
      I => dcti_int(7),
      O => U_DCT1D_latchbuf_reg_7_7_BYINVNOT
    );
  U_DCT1D_latchbuf_reg_7_7_CLKINV_7052 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latchbuf_reg_7_7_CLKINV
    );
  U_DCT1D_latchbuf_reg_7_7_CEINV_7053 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => U_DCT1D_latchbuf_reg_7_7_CEINV
    );
  U_DCT2D_rtlc2n579_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n579_G,
      O => U_DCT2D_rtlc2n579
    );
  U_DCT2D_latch_done_reg_DYMUX_7054 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latch_done_reg_BYINVNOT,
      O => U_DCT2D_latch_done_reg_DYMUX
    );
  U_DCT2D_latch_done_reg_BYINV : X_INV
    port map (
      I => U_DCT2D_istate_reg(0),
      O => U_DCT2D_latch_done_reg_BYINVNOT
    );
  U_DCT2D_latch_done_reg_CLKINV_7055 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latch_done_reg_CLKINV
    );
  U_DCT2D_latch_done_reg_CEINV_7056 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n579,
      O => U_DCT2D_latch_done_reg_CEINV
    );
  U_DCT2D_nx6411z1_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx6411z1_F,
      O => U_DCT2D_nx6411z1
    );
  U_DCT2D_nx6411z1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx6411z1_G,
      O => U_DCT2D_NOT_rtlcs2
    );
  U_DCT2D_nx41892z2_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx41892z2_F,
      O => U_DCT2D_nx41892z2
    );
  U_DCT2D_nx41892z2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx41892z2_G,
      O => U_DCT2D_nx41892z3
    );
  U_DCT1D_row_reg_0_DXMUX_7057 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_row_reg_0_BXINVNOT,
      O => U_DCT1D_row_reg_0_DXMUX
    );
  U_DCT1D_row_reg_0_BXINV : X_INV
    port map (
      I => U_DCT1D_row_reg(0),
      O => U_DCT1D_row_reg_0_BXINVNOT
    );
  U_DCT1D_row_reg_0_DYMUX_7058 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx52040z1,
      O => U_DCT1D_row_reg_0_DYMUX
    );
  U_DCT1D_row_reg_0_SRINV_7059 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_row_reg_0_SRINV
    );
  U_DCT1D_row_reg_0_CLKINV_7060 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_row_reg_0_CLKINV
    );
  U_DCT1D_row_reg_0_CEINV_7061 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcn1047,
      O => U_DCT1D_row_reg_0_CEINV
    );
  U_DCT2D_state_reg_1_DXMUX_7062 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5_state_reg_fsm_SS3_n367(1),
      O => U_DCT2D_state_reg_1_DXMUX
    );
  U_DCT2D_state_reg_1_DYMUX_7063 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg_1_BYINVNOT,
      O => U_DCT2D_state_reg_1_DYMUX
    );
  U_DCT2D_state_reg_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg_1_G,
      O => U_DCT2D_NOT_rtlcs7
    );
  U_DCT2D_state_reg_1_BYINV : X_INV
    port map (
      I => U_DCT2D_state_reg(0),
      O => U_DCT2D_state_reg_1_BYINVNOT
    );
  U_DCT2D_state_reg_1_SRINV_7064 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_state_reg_1_SRINV
    );
  U_DCT2D_state_reg_1_CLKINV_7065 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_state_reg_1_CLKINV
    );
  U_DCT2D_state_reg_1_CEINV_7066 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcn1678,
      O => U_DCT2D_state_reg_1_CEINV
    );
  rome2addro10_s_1_DXMUX_7067 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_Q(10),
      O => rome2addro10_s_1_DXMUX
    );
  rome2addro10_s_1_DYMUX_7068 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_Q(10),
      O => rome2addro10_s_1_DYMUX
    );
  rome2addro10_s_1_SRINV_7069 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro10_s_1_SRINV
    );
  rome2addro10_s_1_CLKINV_7070 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro10_s_1_CLKINV
    );
  rome2addro10_s_1_CEINV_7071 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro10_s_1_CEINV
    );
  rome2addro10_s_3_DXMUX_7072 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_Q(10),
      O => rome2addro10_s_3_DXMUX
    );
  rome2addro10_s_3_DYMUX_7073 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_Q(10),
      O => rome2addro10_s_3_DYMUX
    );
  rome2addro10_s_3_SRINV_7074 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro10_s_3_SRINV
    );
  rome2addro10_s_3_CLKINV_7075 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro10_s_3_CLKINV
    );
  rome2addro10_s_3_CEINV_7076 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro10_s_3_CEINV
    );
  U_DCT1D_rtlc5n1684_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1684_F,
      O => U_DCT1D_rtlc5n1684
    );
  U_DCT1D_rtlc5n1684_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1684_G,
      O => U_DCT1D_rtlc5n1311
    );
  romeaddro0_s_1_DXMUX_7077 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_Q(0),
      O => romeaddro0_s_1_DXMUX
    );
  romeaddro0_s_1_DYMUX_7078 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_Q(0),
      O => romeaddro0_s_1_DYMUX
    );
  romeaddro0_s_1_SRINV_7079 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro0_s_1_SRINV
    );
  romeaddro0_s_1_CLKINV_7080 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro0_s_1_CLKINV
    );
  romeaddro0_s_1_CEINV_7081 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro0_s_1_CEINV
    );
  romeaddro0_s_3_DXMUX_7082 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_Q(0),
      O => romeaddro0_s_3_DXMUX
    );
  romeaddro0_s_3_DYMUX_7083 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_Q(0),
      O => romeaddro0_s_3_DYMUX
    );
  romeaddro0_s_3_SRINV_7084 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro0_s_3_SRINV
    );
  romeaddro0_s_3_CLKINV_7085 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro0_s_3_CLKINV
    );
  romeaddro0_s_3_CEINV_7086 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro0_s_3_CEINV
    );
  romeaddro1_s_1_DXMUX_7087 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_Q(1),
      O => romeaddro1_s_1_DXMUX
    );
  romeaddro1_s_1_DYMUX_7088 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_Q(1),
      O => romeaddro1_s_1_DYMUX
    );
  romeaddro1_s_1_SRINV_7089 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro1_s_1_SRINV
    );
  romeaddro1_s_1_CLKINV_7090 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro1_s_1_CLKINV
    );
  romeaddro1_s_1_CEINV_7091 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro1_s_1_CEINV
    );
  romeaddro1_s_3_DXMUX_7092 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_Q(1),
      O => romeaddro1_s_3_DXMUX
    );
  romeaddro1_s_3_DYMUX_7093 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_Q(1),
      O => romeaddro1_s_3_DYMUX
    );
  romeaddro1_s_3_SRINV_7094 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro1_s_3_SRINV
    );
  romeaddro1_s_3_CLKINV_7095 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro1_s_3_CLKINV
    );
  romeaddro1_s_3_CEINV_7096 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro1_s_3_CEINV
    );
  U_DCT1D_reg_databuf_reg_1_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_1_2_DXMUX,
      CE => U_DCT1D_databuf_reg_1_2_CEINV,
      CLK => U_DCT1D_databuf_reg_1_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_1_2_FFX_RST,
      O => U_DCT1D_databuf_reg_1_Q(2)
    );
  U_DCT1D_databuf_reg_1_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_1_2_FFX_RST
    );
  romeaddro2_s_1_DXMUX_7097 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_Q(2),
      O => romeaddro2_s_1_DXMUX
    );
  romeaddro2_s_1_DYMUX_7098 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_Q(2),
      O => romeaddro2_s_1_DYMUX
    );
  romeaddro2_s_1_SRINV_7099 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro2_s_1_SRINV
    );
  romeaddro2_s_1_CLKINV_7100 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro2_s_1_CLKINV
    );
  romeaddro2_s_1_CEINV_7101 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro2_s_1_CEINV
    );
  romeaddro2_s_3_DXMUX_7102 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_Q(2),
      O => romeaddro2_s_3_DXMUX
    );
  romeaddro2_s_3_DYMUX_7103 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_Q(2),
      O => romeaddro2_s_3_DYMUX
    );
  romeaddro2_s_3_SRINV_7104 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro2_s_3_SRINV
    );
  romeaddro2_s_3_CLKINV_7105 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro2_s_3_CLKINV
    );
  romeaddro2_s_3_CEINV_7106 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro2_s_3_CEINV
    );
  romeaddro3_s_1_DXMUX_7107 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_Q(3),
      O => romeaddro3_s_1_DXMUX
    );
  romeaddro3_s_1_DYMUX_7108 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_Q(3),
      O => romeaddro3_s_1_DYMUX
    );
  romeaddro3_s_1_SRINV_7109 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro3_s_1_SRINV
    );
  romeaddro3_s_1_CLKINV_7110 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro3_s_1_CLKINV
    );
  romeaddro3_s_1_CEINV_7111 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro3_s_1_CEINV
    );
  U_DCT1D_ix4406z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_1_Q(5),
      ADR1 => U_DCT1D_latchbuf_reg_6_Q(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx4406z1
    );
  romeaddro3_s_3_DXMUX_7112 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_Q(3),
      O => romeaddro3_s_3_DXMUX
    );
  romeaddro3_s_3_DYMUX_7113 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_Q(3),
      O => romeaddro3_s_3_DYMUX
    );
  romeaddro3_s_3_SRINV_7114 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro3_s_3_SRINV
    );
  romeaddro3_s_3_CLKINV_7115 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro3_s_3_CLKINV
    );
  romeaddro3_s_3_CEINV_7116 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro3_s_3_CEINV
    );
  romeaddro4_s_1_DXMUX_7117 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_Q(4),
      O => romeaddro4_s_1_DXMUX
    );
  romeaddro4_s_1_DYMUX_7118 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_Q(4),
      O => romeaddro4_s_1_DYMUX
    );
  romeaddro4_s_1_SRINV_7119 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro4_s_1_SRINV
    );
  romeaddro4_s_1_CLKINV_7120 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro4_s_1_CLKINV
    );
  romeaddro4_s_1_CEINV_7121 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro4_s_1_CEINV
    );
  romeaddro4_s_3_DXMUX_7122 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_Q(4),
      O => romeaddro4_s_3_DXMUX
    );
  romeaddro4_s_3_DYMUX_7123 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_Q(4),
      O => romeaddro4_s_3_DYMUX
    );
  romeaddro4_s_3_SRINV_7124 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro4_s_3_SRINV
    );
  romeaddro4_s_3_CLKINV_7125 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro4_s_3_CLKINV
    );
  romeaddro4_s_3_CEINV_7126 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro4_s_3_CEINV
    );
  romeaddro5_s_1_DXMUX_7127 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_Q(5),
      O => romeaddro5_s_1_DXMUX
    );
  romeaddro5_s_1_DYMUX_7128 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_Q(5),
      O => romeaddro5_s_1_DYMUX
    );
  romeaddro5_s_1_SRINV_7129 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro5_s_1_SRINV
    );
  romeaddro5_s_1_CLKINV_7130 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro5_s_1_CLKINV
    );
  romeaddro5_s_1_CEINV_7131 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro5_s_1_CEINV
    );
  romeaddro5_s_3_DXMUX_7132 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_Q(5),
      O => romeaddro5_s_3_DXMUX
    );
  romeaddro5_s_3_DYMUX_7133 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_Q(5),
      O => romeaddro5_s_3_DYMUX
    );
  romeaddro5_s_3_SRINV_7134 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro5_s_3_SRINV
    );
  romeaddro5_s_3_CLKINV_7135 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro5_s_3_CLKINV
    );
  romeaddro5_s_3_CEINV_7136 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro5_s_3_CEINV
    );
  romo2addro10_s_1_DXMUX_7137 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_6_Q(10),
      O => romo2addro10_s_1_DXMUX
    );
  romo2addro10_s_1_DYMUX_7138 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_7_Q(10),
      O => romo2addro10_s_1_DYMUX
    );
  romo2addro10_s_1_SRINV_7139 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro10_s_1_SRINV
    );
  romo2addro10_s_1_CLKINV_7140 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro10_s_1_CLKINV
    );
  romo2addro10_s_1_CEINV_7141 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro10_s_1_CEINV
    );
  romeaddro6_s_1_DXMUX_7142 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_Q(6),
      O => romeaddro6_s_1_DXMUX
    );
  romeaddro6_s_1_DYMUX_7143 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_Q(6),
      O => romeaddro6_s_1_DYMUX
    );
  romeaddro6_s_1_SRINV_7144 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro6_s_1_SRINV
    );
  romeaddro6_s_1_CLKINV_7145 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro6_s_1_CLKINV
    );
  romeaddro6_s_1_CEINV_7146 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro6_s_1_CEINV
    );
  romo2addro10_s_3_DXMUX_7147 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_4_Q(10),
      O => romo2addro10_s_3_DXMUX
    );
  romo2addro10_s_3_DYMUX_7148 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_5_Q(10),
      O => romo2addro10_s_3_DYMUX
    );
  romo2addro10_s_3_SRINV_7149 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro10_s_3_SRINV
    );
  romo2addro10_s_3_CLKINV_7150 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro10_s_3_CLKINV
    );
  romo2addro10_s_3_CEINV_7151 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro10_s_3_CEINV
    );
  romeaddro6_s_3_DXMUX_7152 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_Q(6),
      O => romeaddro6_s_3_DXMUX
    );
  romeaddro6_s_3_DYMUX_7153 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_Q(6),
      O => romeaddro6_s_3_DYMUX
    );
  romeaddro6_s_3_SRINV_7154 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro6_s_3_SRINV
    );
  romeaddro6_s_3_CLKINV_7155 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro6_s_3_CLKINV
    );
  romeaddro6_s_3_CEINV_7156 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro6_s_3_CEINV
    );
  romo2addro0_s_5_DXMUX_7157 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_col_reg(2),
      O => romo2addro0_s_5_DXMUX
    );
  romo2addro0_s_5_DYMUX_7158 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_col_reg(1),
      O => romo2addro0_s_5_DYMUX
    );
  romo2addro0_s_5_SRINV_7159 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romo2addro0_s_5_SRINV
    );
  romo2addro0_s_5_CLKINV_7160 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romo2addro0_s_5_CLKINV
    );
  romo2addro0_s_5_CEINV_7161 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => romo2addro0_s_5_CEINV
    );
  romeaddro7_s_1_DXMUX_7162 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_Q(7),
      O => romeaddro7_s_1_DXMUX
    );
  romeaddro7_s_1_DYMUX_7163 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_Q(7),
      O => romeaddro7_s_1_DYMUX
    );
  romeaddro7_s_1_SRINV_7164 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro7_s_1_SRINV
    );
  romeaddro7_s_1_CLKINV_7165 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro7_s_1_CLKINV
    );
  romeaddro7_s_1_CEINV_7166 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro7_s_1_CEINV
    );
  romeaddro7_s_3_DXMUX_7167 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_Q(7),
      O => romeaddro7_s_3_DXMUX
    );
  romeaddro7_s_3_DYMUX_7168 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_Q(7),
      O => romeaddro7_s_3_DYMUX
    );
  romeaddro7_s_3_SRINV_7169 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro7_s_3_SRINV
    );
  romeaddro7_s_3_CLKINV_7170 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro7_s_3_CLKINV
    );
  romeaddro7_s_3_CEINV_7171 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro7_s_3_CEINV
    );
  romeaddro8_s_1_DXMUX_7172 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_2_Q(8),
      O => romeaddro8_s_1_DXMUX
    );
  romeaddro8_s_1_DYMUX_7173 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_3_Q(8),
      O => romeaddro8_s_1_DYMUX
    );
  romeaddro8_s_1_SRINV_7174 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro8_s_1_SRINV
    );
  romeaddro8_s_1_CLKINV_7175 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro8_s_1_CLKINV
    );
  romeaddro8_s_1_CEINV_7176 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro8_s_1_CEINV
    );
  romeaddro8_s_3_DXMUX_7177 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_0_Q(8),
      O => romeaddro8_s_3_DXMUX
    );
  romeaddro8_s_3_DYMUX_7178 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_1_Q(8),
      O => romeaddro8_s_3_DYMUX
    );
  romeaddro8_s_3_SRINV_7179 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romeaddro8_s_3_SRINV
    );
  romeaddro8_s_3_CLKINV_7180 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romeaddro8_s_3_CLKINV
    );
  romeaddro8_s_3_CEINV_7181 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612,
      O => romeaddro8_s_3_CEINV
    );
  U_DCT2D_rtlc5n1854_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1854_F,
      O => U_DCT2D_rtlc5n1854
    );
  U_DCT2D_rtlc5n1854_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1854_G,
      O => U_DCT2D_rtlc5n1768
    );
  U_DCT2D_nx65206z1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z1_G,
      O => U_DCT2D_nx65206z1
    );
  U_DCT2D_nx65206z253_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z253_G,
      O => U_DCT2D_nx65206z253
    );
  U_DCT2D_nx65206z5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z5_G,
      O => U_DCT2D_nx65206z5
    );
  U_DCT2D_nx65206z78_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z78_G,
      O => U_DCT2D_nx65206z78
    );
  U_DCT2D_nx65206z79_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z79_G,
      O => U_DCT2D_nx65206z79
    );
  U_DCT2D_nx65206z42_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z42_G,
      O => U_DCT2D_nx65206z42
    );
  U_DCT2D_nx65206z572_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z572_F,
      O => U_DCT2D_nx65206z572
    );
  U_DCT2D_nx65206z572_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z572_G,
      O => U_DCT2D_nx65206z573
    );
  U_DCT2D_nx65206z583_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z583_F,
      O => U_DCT2D_nx65206z583
    );
  U_DCT2D_nx65206z296_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z296_G,
      O => U_DCT2D_nx65206z296
    );
  U_DCT2D_nx65206z586_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z586_F,
      O => U_DCT2D_nx65206z586
    );
  U_DCT2D_nx65206z215_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z215_F,
      O => U_DCT2D_nx65206z215
    );
  U_DCT2D_nx65206z215_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z215_G,
      O => U_DCT2D_nx65206z212
    );
  U_DCT2D_nx65206z297_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z297_G,
      O => U_DCT2D_nx65206z297
    );
  U_DCT2D_nx65206z121_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z121_G,
      O => U_DCT2D_nx65206z121
    );
  U_DCT2D_nx65206z595_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z595_F,
      O => U_DCT2D_nx65206z595
    );
  U_DCT2D_nx65206z604_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z604_F,
      O => U_DCT2D_nx65206z604
    );
  U_DCT2D_nx65206z580_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z580_F,
      O => U_DCT2D_nx65206z580
    );
  U_DCT2D_nx65206z589_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z589_F,
      O => U_DCT2D_nx65206z589
    );
  U_DCT2D_nx65206z598_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z598_F,
      O => U_DCT2D_nx65206z598
    );
  U_DCT2D_nx65206z607_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z607_F,
      O => U_DCT2D_nx65206z607
    );
  U_DCT2D_nx65206z413_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z413_G,
      O => U_DCT2D_nx65206z413
    );
  U_DCT1D_reg_databuf_reg_1_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_1_4_DYMUX,
      CE => U_DCT1D_databuf_reg_1_4_CEINV,
      CLK => U_DCT1D_databuf_reg_1_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_1_4_FFY_RST,
      O => U_DCT1D_databuf_reg_1_Q(5)
    );
  U_DCT1D_databuf_reg_1_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_1_4_FFY_RST
    );
  U_DCT2D_nx65206z592_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z592_F,
      O => U_DCT2D_nx65206z592
    );
  U_DCT2D_nx65206z224_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z224_G,
      O => U_DCT2D_nx65206z224
    );
  U_DCT2D_nx65206z601_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z601_F,
      O => U_DCT2D_nx65206z601
    );
  U_DCT2D_nx65206z233_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z233_G,
      O => U_DCT2D_nx65206z233
    );
  U_DCT2D_nx65206z221_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z221_G,
      O => U_DCT2D_nx65206z221
    );
  U_DCT2D_nx65206z230_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z230_G,
      O => U_DCT2D_nx65206z230
    );
  U_DCT2D_nx65206z239_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z239_G,
      O => U_DCT2D_nx65206z239
    );
  U_DCT2D_nx65206z227_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z227_G,
      O => U_DCT2D_nx65206z227
    );
  U_DCT2D_nx65206z334_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z334_G,
      O => U_DCT2D_nx65206z334
    );
  U_DCT2D_nx65206z248_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z248_G,
      O => U_DCT2D_nx65206z248
    );
  U_DCT1D_ix3409z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_1_Q(4),
      ADR1 => U_DCT1D_latchbuf_reg_6_Q(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx3409z1
    );
  U_DCT2D_nx65206z236_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z236_G,
      O => U_DCT2D_nx65206z236
    );
  U_DCT2D_nx65206z245_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z245_G,
      O => U_DCT2D_nx65206z245
    );
  U_DCT2D_nx65206z242_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx65206z242_G,
      O => U_DCT2D_nx65206z242
    );
  requestrd_s_DYMUX_7182 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => requestrd_s_BYINVNOT,
      O => requestrd_s_DYMUX
    );
  requestrd_s_BYINV : X_INV
    port map (
      I => requestrd_s,
      O => requestrd_s_BYINVNOT
    );
  requestrd_s_CLKINV_7183 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => requestrd_s_CLKINV
    );
  requestrd_s_CEINV_7184 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n581,
      O => requestrd_s_CEINV
    );
  U_DCT2D_rtlc2n446_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n446_F,
      O => U_DCT2D_rtlc2n446
    );
  U_DCT2D_rtlc2n446_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n446_G,
      O => U_DCT2D_nx49413z1
    );
  U_DCT2D_nx40895z2_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx40895z2_F,
      O => U_DCT2D_nx40895z2
    );
  U_DCT2D_nx40895z2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx40895z2_G,
      O => U_DCT2D_NOT_rtlc2n488
    );
  U_DCT1D_nx52393z1_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx52393z1_F,
      O => U_DCT1D_nx52393z1
    );
  U_DCT1D_nx52393z1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx52393z1_G,
      O => U_DCT1D_nx7397z1
    );
  U_DCT1D_rtlc2n293_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n293_F,
      O => U_DCT1D_rtlc2n293
    );
  U_DCT1D_rtlc2n293_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n293_G,
      O => U_DCT1D_NOT_rtlcs1
    );
  U_DCT1D_rtlc2n468_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n468_F,
      O => U_DCT1D_rtlc2n468
    );
  U_DCT1D_rtlc2n468_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n468_G,
      O => U_DCT1D_nx7599z1
    );
  U_DCT2D_colram_reg_3_DYMUX_7185 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_colram_reg_3_BYINVNOT,
      O => U_DCT2D_colram_reg_3_DYMUX
    );
  U_DCT2D_colram_reg_3_BYINV : X_INV
    port map (
      I => U_DCT2D_colram_reg(3),
      O => U_DCT2D_colram_reg_3_BYINVNOT
    );
  U_DCT2D_colram_reg_3_CLKINV_7186 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_colram_reg_3_CLKINV
    );
  U_DCT2D_colram_reg_3_CEINV_7187 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_nx41892z2,
      O => U_DCT2D_colram_reg_3_CEINV
    );
  U_DCT1D_rtlc5n1558_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558_F,
      O => U_DCT1D_rtlc5n1558
    );
  U_DCT1D_rtlc5n1558_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1558_G,
      O => U_DCT1D_rtlc5n1690
    );
  releasewr_s_DYMUX_7188 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => releasewr_s_DYMUX
    );
  releasewr_s_CLKINV_7189 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => releasewr_s_CLKINV
    );
  releasewr_s_CEINV_7190 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1684,
      O => releasewr_s_CEINV
    );
  U_DCT1D_latch_done_reg_DYMUX_7191 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_latch_done_reg_BYINVNOT,
      O => U_DCT1D_latch_done_reg_DYMUX
    );
  U_DCT1D_latch_done_reg_BYINV : X_INV
    port map (
      I => U_DCT1D_istate_reg(1),
      O => U_DCT1D_latch_done_reg_BYINVNOT
    );
  U_DCT1D_latch_done_reg_CLKINV_7192 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_latch_done_reg_CLKINV
    );
  U_DCT1D_latch_done_reg_CEINV_7193 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n468,
      O => U_DCT1D_latch_done_reg_CEINV
    );
  U_DCT1D_NOT_rtlcs2_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_NOT_rtlcs2_F,
      O => U_DCT1D_NOT_rtlcs2
    );
  U_DCT1D_NOT_rtlcs2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_NOT_rtlcs2_G,
      O => U_DCT1D_rtlcs3
    );
  U_DCT1D_nx62663z1_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx62663z1_F,
      O => U_DCT1D_nx62663z1
    );
  U_DCT1D_nx62663z1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx62663z1_G,
      O => U_DCT1D_nx42123z1
    );
  U_DCT1D_rtlc5n1612_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612_F,
      O => U_DCT1D_rtlc5n1612
    );
  U_DCT1D_rtlc5n1612_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1612_G,
      O => U_DCT1D_rtlcn1047
    );
  U_DCT2D_completed_reg_DYMUX_7194 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_completed_reg_BYINVNOT,
      O => U_DCT2D_completed_reg_DYMUX
    );
  U_DCT2D_completed_reg_BYINV : X_INV
    port map (
      I => U_DCT2D_istate_reg(0),
      O => U_DCT2D_completed_reg_BYINVNOT
    );
  U_DCT2D_completed_reg_CLKINV_7195 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_completed_reg_CLKINV
    );
  U_DCT2D_completed_reg_CEINV_7196 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n580,
      O => U_DCT2D_completed_reg_CEINV
    );
  U_DCT2D_col_tmp_reg_1_DXMUX_7197 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_col_tmp_reg_1_BXINVNOT,
      O => U_DCT2D_col_tmp_reg_1_DXMUX
    );
  U_DCT2D_col_tmp_reg_1_BXINV : X_INV
    port map (
      I => U_DCT2D_col_reg(1),
      O => U_DCT2D_col_tmp_reg_1_BXINVNOT
    );
  U_DCT2D_col_tmp_reg_1_DYMUX_7198 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n942(2),
      O => U_DCT2D_col_tmp_reg_1_DYMUX
    );
  U_DCT2D_col_tmp_reg_1_SRINV_7199 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_col_tmp_reg_1_SRINV
    );
  U_DCT2D_col_tmp_reg_1_CLKINV_7200 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_col_tmp_reg_1_CLKINV
    );
  U_DCT2D_col_tmp_reg_1_CEINV_7201 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlcs5,
      O => U_DCT2D_col_tmp_reg_1_CEINV
    );
  U_DCT1D_nx57528z1_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx57528z1_F,
      O => U_DCT1D_nx57528z1
    );
  U_DCT1D_nx57528z1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx57528z1_G,
      O => U_DCT1D_nx53004z1
    );
  ramwaddro_s_1_DXMUX_7202 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_row_reg(1),
      O => ramwaddro_s_1_DXMUX
    );
  ramwaddro_s_1_DYMUX_7203 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_row_reg(0),
      O => ramwaddro_s_1_DYMUX
    );
  ramwaddro_s_1_SRINV_7204 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramwaddro_s_1_SRINV
    );
  ramwaddro_s_1_CLKINV_7205 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramwaddro_s_1_CLKINV
    );
  ramwaddro_s_1_CEINV_7206 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => ramwaddro_s_1_CEINV
    );
  U_DCT1D_reg_databuf_reg_1_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_1_4_DXMUX,
      CE => U_DCT1D_databuf_reg_1_4_CEINV,
      CLK => U_DCT1D_databuf_reg_1_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_1_4_FFX_RST,
      O => U_DCT1D_databuf_reg_1_Q(4)
    );
  U_DCT1D_databuf_reg_1_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_1_4_FFX_RST
    );
  ramwaddro_s_3_DXMUX_7207 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_col_reg(0),
      O => ramwaddro_s_3_DXMUX
    );
  ramwaddro_s_3_DYMUX_7208 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_row_reg(2),
      O => ramwaddro_s_3_DYMUX
    );
  ramwaddro_s_3_SRINV_7209 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramwaddro_s_3_SRINV
    );
  ramwaddro_s_3_CLKINV_7210 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramwaddro_s_3_CLKINV
    );
  ramwaddro_s_3_CEINV_7211 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => ramwaddro_s_3_CEINV
    );
  ramwaddro_s_5_DXMUX_7212 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_col_reg(2),
      O => ramwaddro_s_5_DXMUX
    );
  ramwaddro_s_5_DYMUX_7213 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_col_reg(1),
      O => ramwaddro_s_5_DYMUX
    );
  ramwaddro_s_5_SRINV_7214 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramwaddro_s_5_SRINV
    );
  ramwaddro_s_5_CLKINV_7215 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramwaddro_s_5_CLKINV
    );
  ramwaddro_s_5_CEINV_7216 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => ramwaddro_s_5_CEINV
    );
  U_DCT1D_inpcnt_reg_0_DXMUX_7217 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_inpcnt_reg_0_BXINVNOT,
      O => U_DCT1D_inpcnt_reg_0_DXMUX
    );
  U_DCT1D_inpcnt_reg_0_BXINV : X_INV
    port map (
      I => U_DCT1D_inpcnt_reg(0),
      O => U_DCT1D_inpcnt_reg_0_BXINVNOT
    );
  U_DCT1D_inpcnt_reg_0_DYMUX_7218 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx58996z1,
      O => U_DCT1D_inpcnt_reg_0_DYMUX
    );
  U_DCT1D_inpcnt_reg_0_SRINV_7219 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_inpcnt_reg_0_SRINV
    );
  U_DCT1D_inpcnt_reg_0_CLKINV_7220 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_inpcnt_reg_0_CLKINV
    );
  U_DCT1D_inpcnt_reg_0_CEINV_7221 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n365,
      O => U_DCT1D_inpcnt_reg_0_CEINV
    );
  U_DCT1D_ix6400z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_1_Q(7),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_6_Q(7),
      O => U_DCT1D_nx6400z1
    );
  ramwe_s_DYMUX_7222 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => ramwe_s_DYMUX
    );
  ramwe_s_CLKINV_7223 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ramwe_s_CLKINV
    );
  ramwe_s_CEINV_7224 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_NOT_rtlcs2,
      O => ramwe_s_CEINV
    );
  rome2addro0_s_1_DXMUX_7225 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_Q(0),
      O => rome2addro0_s_1_DXMUX
    );
  rome2addro0_s_1_DYMUX_7226 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_Q(0),
      O => rome2addro0_s_1_DYMUX
    );
  rome2addro0_s_1_SRINV_7227 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro0_s_1_SRINV
    );
  rome2addro0_s_1_CLKINV_7228 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro0_s_1_CLKINV
    );
  rome2addro0_s_1_CEINV_7229 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro0_s_1_CEINV
    );
  rome2addro0_s_3_DXMUX_7230 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_Q(0),
      O => rome2addro0_s_3_DXMUX
    );
  rome2addro0_s_3_DYMUX_7231 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_Q(0),
      O => rome2addro0_s_3_DYMUX
    );
  rome2addro0_s_3_SRINV_7232 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro0_s_3_SRINV
    );
  rome2addro0_s_3_CLKINV_7233 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro0_s_3_CLKINV
    );
  rome2addro0_s_3_CEINV_7234 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro0_s_3_CEINV
    );
  rome2addro1_s_1_DXMUX_7235 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_Q(1),
      O => rome2addro1_s_1_DXMUX
    );
  rome2addro1_s_1_DYMUX_7236 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_Q(1),
      O => rome2addro1_s_1_DYMUX
    );
  rome2addro1_s_1_SRINV_7237 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro1_s_1_SRINV
    );
  rome2addro1_s_1_CLKINV_7238 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro1_s_1_CLKINV
    );
  rome2addro1_s_1_CEINV_7239 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro1_s_1_CEINV
    );
  rome2addro1_s_3_DXMUX_7240 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_Q(1),
      O => rome2addro1_s_3_DXMUX
    );
  rome2addro1_s_3_DYMUX_7241 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_Q(1),
      O => rome2addro1_s_3_DYMUX
    );
  rome2addro1_s_3_SRINV_7242 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro1_s_3_SRINV
    );
  rome2addro1_s_3_CLKINV_7243 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro1_s_3_CLKINV
    );
  rome2addro1_s_3_CEINV_7244 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro1_s_3_CEINV
    );
  rome2addro2_s_1_DXMUX_7245 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_Q(2),
      O => rome2addro2_s_1_DXMUX
    );
  rome2addro2_s_1_DYMUX_7246 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_Q(2),
      O => rome2addro2_s_1_DYMUX
    );
  rome2addro2_s_1_SRINV_7247 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro2_s_1_SRINV
    );
  rome2addro2_s_1_CLKINV_7248 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro2_s_1_CLKINV
    );
  rome2addro2_s_1_CEINV_7249 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro2_s_1_CEINV
    );
  rome2addro2_s_3_DXMUX_7250 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_Q(2),
      O => rome2addro2_s_3_DXMUX
    );
  rome2addro2_s_3_DYMUX_7251 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_Q(2),
      O => rome2addro2_s_3_DYMUX
    );
  rome2addro2_s_3_SRINV_7252 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro2_s_3_SRINV
    );
  rome2addro2_s_3_CLKINV_7253 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro2_s_3_CLKINV
    );
  rome2addro2_s_3_CEINV_7254 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro2_s_3_CEINV
    );
  rome2addro3_s_1_DXMUX_7255 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_Q(3),
      O => rome2addro3_s_1_DXMUX
    );
  rome2addro3_s_1_DYMUX_7256 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_Q(3),
      O => rome2addro3_s_1_DYMUX
    );
  rome2addro3_s_1_SRINV_7257 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro3_s_1_SRINV
    );
  rome2addro3_s_1_CLKINV_7258 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro3_s_1_CLKINV
    );
  rome2addro3_s_1_CEINV_7259 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro3_s_1_CEINV
    );
  rome2addro3_s_3_DXMUX_7260 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_Q(3),
      O => rome2addro3_s_3_DXMUX
    );
  rome2addro3_s_3_DYMUX_7261 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_Q(3),
      O => rome2addro3_s_3_DYMUX
    );
  rome2addro3_s_3_SRINV_7262 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro3_s_3_SRINV
    );
  rome2addro3_s_3_CLKINV_7263 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro3_s_3_CLKINV
    );
  rome2addro3_s_3_CEINV_7264 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro3_s_3_CEINV
    );
  rome2addro4_s_1_DXMUX_7265 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_Q(4),
      O => rome2addro4_s_1_DXMUX
    );
  rome2addro4_s_1_DYMUX_7266 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_Q(4),
      O => rome2addro4_s_1_DYMUX
    );
  rome2addro4_s_1_SRINV_7267 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro4_s_1_SRINV
    );
  rome2addro4_s_1_CLKINV_7268 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro4_s_1_CLKINV
    );
  rome2addro4_s_1_CEINV_7269 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro4_s_1_CEINV
    );
  rome2addro4_s_3_DXMUX_7270 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_Q(4),
      O => rome2addro4_s_3_DXMUX
    );
  rome2addro4_s_3_DYMUX_7271 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_Q(4),
      O => rome2addro4_s_3_DYMUX
    );
  rome2addro4_s_3_SRINV_7272 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro4_s_3_SRINV
    );
  rome2addro4_s_3_CLKINV_7273 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro4_s_3_CLKINV
    );
  rome2addro4_s_3_CEINV_7274 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro4_s_3_CEINV
    );
  rome2addro5_s_1_DXMUX_7275 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_Q(5),
      O => rome2addro5_s_1_DXMUX
    );
  rome2addro5_s_1_DYMUX_7276 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_Q(5),
      O => rome2addro5_s_1_DYMUX
    );
  rome2addro5_s_1_SRINV_7277 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro5_s_1_SRINV
    );
  rome2addro5_s_1_CLKINV_7278 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro5_s_1_CLKINV
    );
  rome2addro5_s_1_CEINV_7279 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro5_s_1_CEINV
    );
  rome2addro5_s_3_DXMUX_7280 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_Q(5),
      O => rome2addro5_s_3_DXMUX
    );
  rome2addro5_s_3_DYMUX_7281 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_Q(5),
      O => rome2addro5_s_3_DYMUX
    );
  rome2addro5_s_3_SRINV_7282 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro5_s_3_SRINV
    );
  rome2addro5_s_3_CLKINV_7283 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro5_s_3_CLKINV
    );
  rome2addro5_s_3_CEINV_7284 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro5_s_3_CEINV
    );
  rome2addro6_s_1_DXMUX_7285 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_Q(6),
      O => rome2addro6_s_1_DXMUX
    );
  rome2addro6_s_1_DYMUX_7286 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_Q(6),
      O => rome2addro6_s_1_DYMUX
    );
  rome2addro6_s_1_SRINV_7287 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro6_s_1_SRINV
    );
  rome2addro6_s_1_CLKINV_7288 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro6_s_1_CLKINV
    );
  rome2addro6_s_1_CEINV_7289 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro6_s_1_CEINV
    );
  rome2addro6_s_3_DXMUX_7290 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_Q(6),
      O => rome2addro6_s_3_DXMUX
    );
  rome2addro6_s_3_DYMUX_7291 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_Q(6),
      O => rome2addro6_s_3_DYMUX
    );
  rome2addro6_s_3_SRINV_7292 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro6_s_3_SRINV
    );
  rome2addro6_s_3_CLKINV_7293 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro6_s_3_CLKINV
    );
  rome2addro6_s_3_CEINV_7294 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro6_s_3_CEINV
    );
  rome2addro7_s_1_DXMUX_7295 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_Q(7),
      O => rome2addro7_s_1_DXMUX
    );
  rome2addro7_s_1_DYMUX_7296 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_Q(7),
      O => rome2addro7_s_1_DYMUX
    );
  rome2addro7_s_1_SRINV_7297 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro7_s_1_SRINV
    );
  rome2addro7_s_1_CLKINV_7298 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro7_s_1_CLKINV
    );
  rome2addro7_s_1_CEINV_7299 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro7_s_1_CEINV
    );
  rome2addro7_s_3_DXMUX_7300 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_Q(7),
      O => rome2addro7_s_3_DXMUX
    );
  rome2addro7_s_3_DYMUX_7301 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_Q(7),
      O => rome2addro7_s_3_DYMUX
    );
  rome2addro7_s_3_SRINV_7302 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro7_s_3_SRINV
    );
  rome2addro7_s_3_CLKINV_7303 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro7_s_3_CLKINV
    );
  rome2addro7_s_3_CEINV_7304 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro7_s_3_CEINV
    );
  rome2addro8_s_1_DXMUX_7305 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_Q(8),
      O => rome2addro8_s_1_DXMUX
    );
  rome2addro8_s_1_DYMUX_7306 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_Q(8),
      O => rome2addro8_s_1_DYMUX
    );
  rome2addro8_s_1_SRINV_7307 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro8_s_1_SRINV
    );
  rome2addro8_s_1_CLKINV_7308 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro8_s_1_CLKINV
    );
  rome2addro8_s_1_CEINV_7309 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro8_s_1_CEINV
    );
  rome2addro8_s_3_DXMUX_7310 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_Q(8),
      O => rome2addro8_s_3_DXMUX
    );
  rome2addro8_s_3_DYMUX_7311 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_Q(8),
      O => rome2addro8_s_3_DYMUX
    );
  rome2addro8_s_3_SRINV_7312 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro8_s_3_SRINV
    );
  rome2addro8_s_3_CLKINV_7313 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro8_s_3_CLKINV
    );
  rome2addro8_s_3_CEINV_7314 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro8_s_3_CEINV
    );
  rome2addro9_s_1_DXMUX_7315 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_2_Q(9),
      O => rome2addro9_s_1_DXMUX
    );
  rome2addro9_s_1_DYMUX_7316 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_3_Q(9),
      O => rome2addro9_s_1_DYMUX
    );
  rome2addro9_s_1_SRINV_7317 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro9_s_1_SRINV
    );
  rome2addro9_s_1_CLKINV_7318 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro9_s_1_CLKINV
    );
  rome2addro9_s_1_CEINV_7319 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro9_s_1_CEINV
    );
  rome2addro9_s_3_DXMUX_7320 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_0_Q(9),
      O => rome2addro9_s_3_DXMUX
    );
  rome2addro9_s_3_DYMUX_7321 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_databuf_reg_1_Q(9),
      O => rome2addro9_s_3_DYMUX
    );
  rome2addro9_s_3_SRINV_7322 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => rome2addro9_s_3_SRINV
    );
  rome2addro9_s_3_CLKINV_7323 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => rome2addro9_s_3_CLKINV
    );
  rome2addro9_s_3_CEINV_7324 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1768,
      O => rome2addro9_s_3_CEINV
    );
  U_DCT1D_rtlc2n471_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n471_F,
      O => U_DCT1D_rtlc2n471
    );
  U_DCT1D_rtlc2n471_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n471_G,
      O => U_DCT1D_nx2819z1
    );
  U_DCT2D_latchbuf_reg_0_1_DXMUX_7325 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_1_Q,
      O => U_DCT2D_latchbuf_reg_0_1_DXMUX
    );
  U_DCT2D_latchbuf_reg_0_1_DYMUX_7326 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_0_Q,
      O => U_DCT2D_latchbuf_reg_0_1_DYMUX
    );
  U_DCT2D_latchbuf_reg_0_1_SRINV_7327 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_0_1_SRINV
    );
  U_DCT2D_latchbuf_reg_0_1_CLKINV_7328 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_0_1_CLKINV
    );
  U_DCT2D_latchbuf_reg_0_1_CEINV_7329 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_0_1_CEINV
    );
  U_DCT2D_latchbuf_reg_0_3_DXMUX_7330 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_3_Q,
      O => U_DCT2D_latchbuf_reg_0_3_DXMUX
    );
  U_DCT2D_latchbuf_reg_0_3_DYMUX_7331 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_2_Q,
      O => U_DCT2D_latchbuf_reg_0_3_DYMUX
    );
  U_DCT2D_latchbuf_reg_0_3_SRINV_7332 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_0_3_SRINV
    );
  U_DCT2D_latchbuf_reg_0_3_CLKINV_7333 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_0_3_CLKINV
    );
  U_DCT2D_latchbuf_reg_0_3_CEINV_7334 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_0_3_CEINV
    );
  U_DCT2D_latchbuf_reg_0_5_DXMUX_7335 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_5_Q,
      O => U_DCT2D_latchbuf_reg_0_5_DXMUX
    );
  U_DCT2D_latchbuf_reg_0_5_DYMUX_7336 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_4_Q,
      O => U_DCT2D_latchbuf_reg_0_5_DYMUX
    );
  U_DCT2D_latchbuf_reg_0_5_SRINV_7337 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_0_5_SRINV
    );
  U_DCT2D_latchbuf_reg_0_5_CLKINV_7338 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_0_5_CLKINV
    );
  U_DCT2D_latchbuf_reg_0_5_CEINV_7339 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_0_5_CEINV
    );
  U_DCT1D_nx7397z1_rt_7340 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx7397z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx7397z1_rt
    );
  U_DCT2D_latchbuf_reg_0_7_DXMUX_7341 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_7_Q,
      O => U_DCT2D_latchbuf_reg_0_7_DXMUX
    );
  U_DCT2D_latchbuf_reg_0_7_DYMUX_7342 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_6_Q,
      O => U_DCT2D_latchbuf_reg_0_7_DYMUX
    );
  U_DCT2D_latchbuf_reg_0_7_SRINV_7343 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_0_7_SRINV
    );
  U_DCT2D_latchbuf_reg_0_7_CLKINV_7344 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_0_7_CLKINV
    );
  U_DCT2D_latchbuf_reg_0_7_CEINV_7345 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_0_7_CEINV
    );
  U_DCT2D_latchbuf_reg_0_10_DXMUX_7346 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_10_Q,
      O => U_DCT2D_latchbuf_reg_0_10_DXMUX
    );
  U_DCT2D_latchbuf_reg_0_10_DYMUX_7347 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_8_Q,
      O => U_DCT2D_latchbuf_reg_0_10_DYMUX
    );
  U_DCT2D_latchbuf_reg_0_10_SRINV_7348 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_0_10_SRINV
    );
  U_DCT2D_latchbuf_reg_0_10_CLKINV_7349 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_0_10_CLKINV
    );
  U_DCT2D_latchbuf_reg_0_10_CEINV_7350 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_0_10_CEINV
    );
  U_DCT2D_latchbuf_reg_1_1_DXMUX_7351 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_1_Q,
      O => U_DCT2D_latchbuf_reg_1_1_DXMUX
    );
  U_DCT2D_latchbuf_reg_1_1_DYMUX_7352 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_0_Q,
      O => U_DCT2D_latchbuf_reg_1_1_DYMUX
    );
  U_DCT2D_latchbuf_reg_1_1_SRINV_7353 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_1_1_SRINV
    );
  U_DCT2D_latchbuf_reg_1_1_CLKINV_7354 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_1_1_CLKINV
    );
  U_DCT2D_latchbuf_reg_1_1_CEINV_7355 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_1_1_CEINV
    );
  U_DCT2D_latchbuf_reg_1_3_DXMUX_7356 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_3_Q,
      O => U_DCT2D_latchbuf_reg_1_3_DXMUX
    );
  U_DCT2D_latchbuf_reg_1_3_DYMUX_7357 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_2_Q,
      O => U_DCT2D_latchbuf_reg_1_3_DYMUX
    );
  U_DCT2D_latchbuf_reg_1_3_SRINV_7358 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_1_3_SRINV
    );
  U_DCT2D_latchbuf_reg_1_3_CLKINV_7359 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_1_3_CLKINV
    );
  U_DCT2D_latchbuf_reg_1_3_CEINV_7360 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_1_3_CEINV
    );
  U_DCT2D_latchbuf_reg_1_5_DXMUX_7361 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_5_Q,
      O => U_DCT2D_latchbuf_reg_1_5_DXMUX
    );
  U_DCT2D_latchbuf_reg_1_5_DYMUX_7362 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_4_Q,
      O => U_DCT2D_latchbuf_reg_1_5_DYMUX
    );
  U_DCT2D_latchbuf_reg_1_5_SRINV_7363 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_1_5_SRINV
    );
  U_DCT2D_latchbuf_reg_1_5_CLKINV_7364 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_1_5_CLKINV
    );
  U_DCT2D_latchbuf_reg_1_5_CEINV_7365 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_1_5_CEINV
    );
  U_DCT2D_latchbuf_reg_1_7_DXMUX_7366 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_7_Q,
      O => U_DCT2D_latchbuf_reg_1_7_DXMUX
    );
  U_DCT2D_latchbuf_reg_1_7_DYMUX_7367 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_6_Q,
      O => U_DCT2D_latchbuf_reg_1_7_DYMUX
    );
  U_DCT2D_latchbuf_reg_1_7_SRINV_7368 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_1_7_SRINV
    );
  U_DCT2D_latchbuf_reg_1_7_CLKINV_7369 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_1_7_CLKINV
    );
  U_DCT2D_latchbuf_reg_1_7_CEINV_7370 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_1_7_CEINV
    );
  U_DCT2D_latchbuf_reg_1_10_DXMUX_7371 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_10_Q,
      O => U_DCT2D_latchbuf_reg_1_10_DXMUX
    );
  U_DCT2D_latchbuf_reg_1_10_DYMUX_7372 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_8_Q,
      O => U_DCT2D_latchbuf_reg_1_10_DYMUX
    );
  U_DCT2D_latchbuf_reg_1_10_SRINV_7373 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_1_10_SRINV
    );
  U_DCT2D_latchbuf_reg_1_10_CLKINV_7374 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_1_10_CLKINV
    );
  U_DCT2D_latchbuf_reg_1_10_CEINV_7375 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_1_10_CEINV
    );
  U_DCT2D_latchbuf_reg_2_1_DXMUX_7376 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_1_Q,
      O => U_DCT2D_latchbuf_reg_2_1_DXMUX
    );
  U_DCT2D_latchbuf_reg_2_1_DYMUX_7377 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_0_Q,
      O => U_DCT2D_latchbuf_reg_2_1_DYMUX
    );
  U_DCT2D_latchbuf_reg_2_1_SRINV_7378 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_2_1_SRINV
    );
  U_DCT2D_latchbuf_reg_2_1_CLKINV_7379 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_2_1_CLKINV
    );
  U_DCT2D_latchbuf_reg_2_1_CEINV_7380 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_2_1_CEINV
    );
  U_DCT2D_latchbuf_reg_2_3_DXMUX_7381 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_3_Q,
      O => U_DCT2D_latchbuf_reg_2_3_DXMUX
    );
  U_DCT2D_latchbuf_reg_2_3_DYMUX_7382 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_2_Q,
      O => U_DCT2D_latchbuf_reg_2_3_DYMUX
    );
  U_DCT2D_latchbuf_reg_2_3_SRINV_7383 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_2_3_SRINV
    );
  U_DCT2D_latchbuf_reg_2_3_CLKINV_7384 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_2_3_CLKINV
    );
  U_DCT2D_latchbuf_reg_2_3_CEINV_7385 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_2_3_CEINV
    );
  U_DCT2D_latchbuf_reg_2_5_DXMUX_7386 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_5_Q,
      O => U_DCT2D_latchbuf_reg_2_5_DXMUX
    );
  U_DCT2D_latchbuf_reg_2_5_DYMUX_7387 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_4_Q,
      O => U_DCT2D_latchbuf_reg_2_5_DYMUX
    );
  U_DCT2D_latchbuf_reg_2_5_SRINV_7388 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_2_5_SRINV
    );
  U_DCT2D_latchbuf_reg_2_5_CLKINV_7389 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_2_5_CLKINV
    );
  U_DCT2D_latchbuf_reg_2_5_CEINV_7390 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_2_5_CEINV
    );
  U_DCT1D_reg_databuf_reg_1_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_1_6_DYMUX,
      CE => U_DCT1D_databuf_reg_1_6_CEINV,
      CLK => U_DCT1D_databuf_reg_1_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_1_6_FFY_RST,
      O => U_DCT1D_databuf_reg_1_Q(7)
    );
  U_DCT1D_databuf_reg_1_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_1_6_FFY_RST
    );
  U_DCT2D_latchbuf_reg_2_7_DXMUX_7391 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_7_Q,
      O => U_DCT2D_latchbuf_reg_2_7_DXMUX
    );
  U_DCT2D_latchbuf_reg_2_7_DYMUX_7392 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_6_Q,
      O => U_DCT2D_latchbuf_reg_2_7_DYMUX
    );
  U_DCT2D_latchbuf_reg_2_7_SRINV_7393 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_2_7_SRINV
    );
  U_DCT2D_latchbuf_reg_2_7_CLKINV_7394 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_2_7_CLKINV
    );
  U_DCT2D_latchbuf_reg_2_7_CEINV_7395 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_2_7_CEINV
    );
  U_DCT2D_latchbuf_reg_2_10_DXMUX_7396 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_10_Q,
      O => U_DCT2D_latchbuf_reg_2_10_DXMUX
    );
  U_DCT2D_latchbuf_reg_2_10_DYMUX_7397 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_8_Q,
      O => U_DCT2D_latchbuf_reg_2_10_DYMUX
    );
  U_DCT2D_latchbuf_reg_2_10_SRINV_7398 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_2_10_SRINV
    );
  U_DCT2D_latchbuf_reg_2_10_CLKINV_7399 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_2_10_CLKINV
    );
  U_DCT2D_latchbuf_reg_2_10_CEINV_7400 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_2_10_CEINV
    );
  U_DCT2D_latchbuf_reg_3_1_DXMUX_7401 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_1_Q,
      O => U_DCT2D_latchbuf_reg_3_1_DXMUX
    );
  U_DCT2D_latchbuf_reg_3_1_DYMUX_7402 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_0_Q,
      O => U_DCT2D_latchbuf_reg_3_1_DYMUX
    );
  U_DCT2D_latchbuf_reg_3_1_SRINV_7403 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_3_1_SRINV
    );
  U_DCT2D_latchbuf_reg_3_1_CLKINV_7404 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_3_1_CLKINV
    );
  U_DCT2D_latchbuf_reg_3_1_CEINV_7405 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_3_1_CEINV
    );
  U_DCT2D_latchbuf_reg_3_3_DXMUX_7406 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_3_Q,
      O => U_DCT2D_latchbuf_reg_3_3_DXMUX
    );
  U_DCT2D_latchbuf_reg_3_3_DYMUX_7407 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_2_Q,
      O => U_DCT2D_latchbuf_reg_3_3_DYMUX
    );
  U_DCT2D_latchbuf_reg_3_3_SRINV_7408 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_3_3_SRINV
    );
  U_DCT2D_latchbuf_reg_3_3_CLKINV_7409 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_3_3_CLKINV
    );
  U_DCT2D_latchbuf_reg_3_3_CEINV_7410 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_3_3_CEINV
    );
  U_DCT2D_latchbuf_reg_3_5_DXMUX_7411 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_5_Q,
      O => U_DCT2D_latchbuf_reg_3_5_DXMUX
    );
  U_DCT2D_latchbuf_reg_3_5_DYMUX_7412 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_4_Q,
      O => U_DCT2D_latchbuf_reg_3_5_DYMUX
    );
  U_DCT2D_latchbuf_reg_3_5_SRINV_7413 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_3_5_SRINV
    );
  U_DCT2D_latchbuf_reg_3_5_CLKINV_7414 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_3_5_CLKINV
    );
  U_DCT2D_latchbuf_reg_3_5_CEINV_7415 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_3_5_CEINV
    );
  U_DCT2D_latchbuf_reg_3_7_DXMUX_7416 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_7_Q,
      O => U_DCT2D_latchbuf_reg_3_7_DXMUX
    );
  U_DCT2D_latchbuf_reg_3_7_DYMUX_7417 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_6_Q,
      O => U_DCT2D_latchbuf_reg_3_7_DYMUX
    );
  U_DCT2D_latchbuf_reg_3_7_SRINV_7418 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_3_7_SRINV
    );
  U_DCT2D_latchbuf_reg_3_7_CLKINV_7419 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_3_7_CLKINV
    );
  U_DCT2D_latchbuf_reg_3_7_CEINV_7420 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_3_7_CEINV
    );
  U_DCT2D_latchbuf_reg_3_10_DXMUX_7421 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_10_Q,
      O => U_DCT2D_latchbuf_reg_3_10_DXMUX
    );
  U_DCT2D_latchbuf_reg_3_10_DYMUX_7422 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_8_Q,
      O => U_DCT2D_latchbuf_reg_3_10_DYMUX
    );
  U_DCT2D_latchbuf_reg_3_10_SRINV_7423 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_3_10_SRINV
    );
  U_DCT2D_latchbuf_reg_3_10_CLKINV_7424 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_3_10_CLKINV
    );
  U_DCT2D_latchbuf_reg_3_10_CEINV_7425 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_3_10_CEINV
    );
  U_DCT2D_latchbuf_reg_4_1_DXMUX_7426 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_1_Q,
      O => U_DCT2D_latchbuf_reg_4_1_DXMUX
    );
  U_DCT2D_latchbuf_reg_4_1_DYMUX_7427 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_0_Q,
      O => U_DCT2D_latchbuf_reg_4_1_DYMUX
    );
  U_DCT2D_latchbuf_reg_4_1_SRINV_7428 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_4_1_SRINV
    );
  U_DCT2D_latchbuf_reg_4_1_CLKINV_7429 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_4_1_CLKINV
    );
  U_DCT2D_latchbuf_reg_4_1_CEINV_7430 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_4_1_CEINV
    );
  U_DCT2D_latchbuf_reg_4_3_DXMUX_7431 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_3_Q,
      O => U_DCT2D_latchbuf_reg_4_3_DXMUX
    );
  U_DCT2D_latchbuf_reg_4_3_DYMUX_7432 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_2_Q,
      O => U_DCT2D_latchbuf_reg_4_3_DYMUX
    );
  U_DCT2D_latchbuf_reg_4_3_SRINV_7433 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_4_3_SRINV
    );
  U_DCT2D_latchbuf_reg_4_3_CLKINV_7434 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_4_3_CLKINV
    );
  U_DCT2D_latchbuf_reg_4_3_CEINV_7435 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_4_3_CEINV
    );
  U_DCT2D_latchbuf_reg_4_5_DXMUX_7436 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_5_Q,
      O => U_DCT2D_latchbuf_reg_4_5_DXMUX
    );
  U_DCT2D_latchbuf_reg_4_5_DYMUX_7437 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_4_Q,
      O => U_DCT2D_latchbuf_reg_4_5_DYMUX
    );
  U_DCT2D_latchbuf_reg_4_5_SRINV_7438 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_4_5_SRINV
    );
  U_DCT2D_latchbuf_reg_4_5_CLKINV_7439 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_4_5_CLKINV
    );
  U_DCT2D_latchbuf_reg_4_5_CEINV_7440 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_4_5_CEINV
    );
  U_DCT1D_ix5403z1321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_1_Q(6),
      ADR2 => U_DCT1D_latchbuf_reg_6_Q(6),
      ADR3 => VCC,
      O => U_DCT1D_nx5403z1
    );
  U_DCT2D_latchbuf_reg_4_7_DXMUX_7441 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_7_Q,
      O => U_DCT2D_latchbuf_reg_4_7_DXMUX
    );
  U_DCT2D_latchbuf_reg_4_7_DYMUX_7442 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_6_Q,
      O => U_DCT2D_latchbuf_reg_4_7_DYMUX
    );
  U_DCT2D_latchbuf_reg_4_7_SRINV_7443 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_4_7_SRINV
    );
  U_DCT2D_latchbuf_reg_4_7_CLKINV_7444 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_4_7_CLKINV
    );
  U_DCT2D_latchbuf_reg_4_7_CEINV_7445 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_4_7_CEINV
    );
  U_DCT2D_latchbuf_reg_4_10_DXMUX_7446 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_10_Q,
      O => U_DCT2D_latchbuf_reg_4_10_DXMUX
    );
  U_DCT2D_latchbuf_reg_4_10_DYMUX_7447 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_8_Q,
      O => U_DCT2D_latchbuf_reg_4_10_DYMUX
    );
  U_DCT2D_latchbuf_reg_4_10_SRINV_7448 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_4_10_SRINV
    );
  U_DCT2D_latchbuf_reg_4_10_CLKINV_7449 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_4_10_CLKINV
    );
  U_DCT2D_latchbuf_reg_4_10_CEINV_7450 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_4_10_CEINV
    );
  U_DCT2D_latchbuf_reg_5_1_DXMUX_7451 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_1_Q,
      O => U_DCT2D_latchbuf_reg_5_1_DXMUX
    );
  U_DCT2D_latchbuf_reg_5_1_DYMUX_7452 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_0_Q,
      O => U_DCT2D_latchbuf_reg_5_1_DYMUX
    );
  U_DCT2D_latchbuf_reg_5_1_SRINV_7453 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_5_1_SRINV
    );
  U_DCT2D_latchbuf_reg_5_1_CLKINV_7454 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_5_1_CLKINV
    );
  U_DCT2D_latchbuf_reg_5_1_CEINV_7455 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_5_1_CEINV
    );
  U_DCT2D_latchbuf_reg_5_3_DXMUX_7456 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_3_Q,
      O => U_DCT2D_latchbuf_reg_5_3_DXMUX
    );
  U_DCT2D_latchbuf_reg_5_3_DYMUX_7457 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_2_Q,
      O => U_DCT2D_latchbuf_reg_5_3_DYMUX
    );
  U_DCT2D_latchbuf_reg_5_3_SRINV_7458 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_5_3_SRINV
    );
  U_DCT2D_latchbuf_reg_5_3_CLKINV_7459 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_5_3_CLKINV
    );
  U_DCT2D_latchbuf_reg_5_3_CEINV_7460 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_5_3_CEINV
    );
  U_DCT2D_latchbuf_reg_5_5_DXMUX_7461 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_5_Q,
      O => U_DCT2D_latchbuf_reg_5_5_DXMUX
    );
  U_DCT2D_latchbuf_reg_5_5_DYMUX_7462 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_4_Q,
      O => U_DCT2D_latchbuf_reg_5_5_DYMUX
    );
  U_DCT2D_latchbuf_reg_5_5_SRINV_7463 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_5_5_SRINV
    );
  U_DCT2D_latchbuf_reg_5_5_CLKINV_7464 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_5_5_CLKINV
    );
  U_DCT2D_latchbuf_reg_5_5_CEINV_7465 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_5_5_CEINV
    );
  U_DCT2D_latchbuf_reg_5_7_DXMUX_7466 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_7_Q,
      O => U_DCT2D_latchbuf_reg_5_7_DXMUX
    );
  U_DCT2D_latchbuf_reg_5_7_DYMUX_7467 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_6_Q,
      O => U_DCT2D_latchbuf_reg_5_7_DYMUX
    );
  U_DCT2D_latchbuf_reg_5_7_SRINV_7468 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_5_7_SRINV
    );
  U_DCT2D_latchbuf_reg_5_7_CLKINV_7469 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_5_7_CLKINV
    );
  U_DCT2D_latchbuf_reg_5_7_CEINV_7470 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_5_7_CEINV
    );
  U_DCT2D_latchbuf_reg_5_10_DXMUX_7471 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_10_Q,
      O => U_DCT2D_latchbuf_reg_5_10_DXMUX
    );
  U_DCT2D_latchbuf_reg_5_10_DYMUX_7472 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_8_Q,
      O => U_DCT2D_latchbuf_reg_5_10_DYMUX
    );
  U_DCT2D_latchbuf_reg_5_10_SRINV_7473 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_5_10_SRINV
    );
  U_DCT2D_latchbuf_reg_5_10_CLKINV_7474 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_5_10_CLKINV
    );
  U_DCT2D_latchbuf_reg_5_10_CEINV_7475 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_5_10_CEINV
    );
  U_DCT2D_latchbuf_reg_6_1_DXMUX_7476 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_1_Q,
      O => U_DCT2D_latchbuf_reg_6_1_DXMUX
    );
  U_DCT2D_latchbuf_reg_6_1_DYMUX_7477 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_0_Q,
      O => U_DCT2D_latchbuf_reg_6_1_DYMUX
    );
  U_DCT2D_latchbuf_reg_6_1_SRINV_7478 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_6_1_SRINV
    );
  U_DCT2D_latchbuf_reg_6_1_CLKINV_7479 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_6_1_CLKINV
    );
  U_DCT2D_latchbuf_reg_6_1_CEINV_7480 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_6_1_CEINV
    );
  U_DCT2D_latchbuf_reg_6_3_DXMUX_7481 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_3_Q,
      O => U_DCT2D_latchbuf_reg_6_3_DXMUX
    );
  U_DCT2D_latchbuf_reg_6_3_DYMUX_7482 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_2_Q,
      O => U_DCT2D_latchbuf_reg_6_3_DYMUX
    );
  U_DCT2D_latchbuf_reg_6_3_SRINV_7483 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_6_3_SRINV
    );
  U_DCT2D_latchbuf_reg_6_3_CLKINV_7484 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_6_3_CLKINV
    );
  U_DCT2D_latchbuf_reg_6_3_CEINV_7485 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_6_3_CEINV
    );
  U_DCT2D_latchbuf_reg_6_5_DXMUX_7486 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_5_Q,
      O => U_DCT2D_latchbuf_reg_6_5_DXMUX
    );
  U_DCT2D_latchbuf_reg_6_5_DYMUX_7487 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_4_Q,
      O => U_DCT2D_latchbuf_reg_6_5_DYMUX
    );
  U_DCT2D_latchbuf_reg_6_5_SRINV_7488 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_6_5_SRINV
    );
  U_DCT2D_latchbuf_reg_6_5_CLKINV_7489 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_6_5_CLKINV
    );
  U_DCT2D_latchbuf_reg_6_5_CEINV_7490 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_6_5_CEINV
    );
  U_DCT2D_latchbuf_reg_6_7_DXMUX_7491 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_7_Q,
      O => U_DCT2D_latchbuf_reg_6_7_DXMUX
    );
  U_DCT2D_latchbuf_reg_6_7_DYMUX_7492 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_6_Q,
      O => U_DCT2D_latchbuf_reg_6_7_DYMUX
    );
  U_DCT2D_latchbuf_reg_6_7_SRINV_7493 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_6_7_SRINV
    );
  U_DCT2D_latchbuf_reg_6_7_CLKINV_7494 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_6_7_CLKINV
    );
  U_DCT2D_latchbuf_reg_6_7_CEINV_7495 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_6_7_CEINV
    );
  U_DCT2D_latchbuf_reg_6_10_DXMUX_7496 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_10_Q,
      O => U_DCT2D_latchbuf_reg_6_10_DXMUX
    );
  U_DCT2D_latchbuf_reg_6_10_DYMUX_7497 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_8_Q,
      O => U_DCT2D_latchbuf_reg_6_10_DYMUX
    );
  U_DCT2D_latchbuf_reg_6_10_SRINV_7498 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latchbuf_reg_6_10_SRINV
    );
  U_DCT2D_latchbuf_reg_6_10_CLKINV_7499 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT2D_latchbuf_reg_6_10_CLKINV
    );
  U_DCT2D_latchbuf_reg_6_10_CEINV_7500 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n576,
      O => U_DCT2D_latchbuf_reg_6_10_CEINV
    );
  U_DCT1D_rtlc5n1685_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n1685_G,
      O => U_DCT1D_rtlc5n1685
    );
  U_DCT1D_nx59700z303_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z303_F,
      O => U_DCT1D_nx59700z303
    );
  U_DCT1D_nx59700z303_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z303_G,
      O => U_DCT1D_nx59700z254
    );
  U_DCT1D_nx59700z1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z1_G,
      O => U_DCT1D_nx59700z1
    );
  U_DCT1D_col_tmp_reg_1_DXMUX_7501 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_col_tmp_reg_1_BXINVNOT,
      O => U_DCT1D_col_tmp_reg_1_DXMUX
    );
  U_DCT1D_col_tmp_reg_1_BXINV : X_INV
    port map (
      I => U_DCT1D_col_reg(1),
      O => U_DCT1D_col_tmp_reg_1_BXINVNOT
    );
  U_DCT1D_col_tmp_reg_1_DYMUX_7502 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n875(2),
      O => U_DCT1D_col_tmp_reg_1_DYMUX
    );
  U_DCT1D_col_tmp_reg_1_SRINV_7503 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_col_tmp_reg_1_SRINV
    );
  U_DCT1D_col_tmp_reg_1_CLKINV_7504 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => U_DCT1D_col_tmp_reg_1_CLKINV
    );
  U_DCT1D_col_tmp_reg_1_CEINV_7505 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => U_DCT1D_col_tmp_reg_1_CEINV
    );
  U_DCT1D_nx59700z333_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z333_F,
      O => U_DCT1D_nx59700z333
    );
  U_DCT1D_nx59700z333_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z333_G,
      O => U_DCT1D_nx59700z332
    );
  U_DCT1D_nx59700z251_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z251_F,
      O => U_DCT1D_nx59700z251
    );
  U_DCT1D_nx59700z251_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z251_G,
      O => U_DCT1D_nx59700z250
    );
  U_DCT1D_nx59700z218_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z218_F,
      O => U_DCT1D_nx59700z218
    );
  U_DCT1D_nx59700z218_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z218_G,
      O => U_DCT1D_nx59700z4
    );
  U_DCT1D_nx59700z348_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z348_F,
      O => U_DCT1D_nx59700z348
    );
  U_DCT1D_reg_databuf_reg_1_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_1_6_DXMUX,
      CE => U_DCT1D_databuf_reg_1_6_CEINV,
      CLK => U_DCT1D_databuf_reg_1_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_1_6_FFX_RST,
      O => U_DCT1D_databuf_reg_1_Q(6)
    );
  U_DCT1D_databuf_reg_1_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_1_6_FFX_RST
    );
  U_DCT1D_nx59700z357_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z357_F,
      O => U_DCT1D_nx59700z357
    );
  U_DCT1D_nx59700z366_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z366_F,
      O => U_DCT1D_nx59700z366
    );
  U_DCT1D_nx59700z342_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z342_F,
      O => U_DCT1D_nx59700z342
    );
  U_DCT1D_nx59700z351_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z351_F,
      O => U_DCT1D_nx59700z351
    );
  U_DCT1D_nx59700z360_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z360_F,
      O => U_DCT1D_nx59700z360
    );
  U_DCT1D_nx59700z369_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z369_F,
      O => U_DCT1D_nx59700z369
    );
  U_DCT1D_nx59700z345_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z345_F,
      O => U_DCT1D_nx59700z345
    );
  U_DCT1D_nx59700z354_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z354_F,
      O => U_DCT1D_nx59700z354
    );
  U_DCT1D_nx59700z363_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z363_F,
      O => U_DCT1D_nx59700z363
    );
  U_DCT1D_nx59700z5_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z5_G,
      O => U_DCT1D_nx59700z5
    );
  U_DCT1D_nx59700z78_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z78_G,
      O => U_DCT1D_nx59700z78
    );
  U_DCT1D_nx59700z79_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z79_G,
      O => U_DCT1D_nx59700z79
    );
  U_DCT1D_nx59700z42_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z42_G,
      O => U_DCT1D_nx59700z42
    );
  U_DCT1D_nx59700z215_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z215_F,
      O => U_DCT1D_nx59700z215
    );
  U_DCT1D_nx59700z215_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z215_G,
      O => U_DCT1D_nx59700z212
    );
  U_DCT1D_nx59700z121_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z121_G,
      O => U_DCT1D_nx59700z121
    );
  U_DCT1D_nx59700z224_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z224_G,
      O => U_DCT1D_nx59700z224
    );
  U_DCT1D_nx59700z233_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z233_G,
      O => U_DCT1D_nx59700z233
    );
  U_DCT1D_nx59700z221_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z221_G,
      O => U_DCT1D_nx59700z221
    );
  U_DCT1D_nx59700z230_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z230_G,
      O => U_DCT1D_nx59700z230
    );
  U_DCT1D_nx59700z306_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z306_G,
      O => U_DCT1D_nx59700z306
    );
  U_DCT1D_nx59700z300_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z300_G,
      O => U_DCT1D_nx59700z300
    );
  U_DCT1D_nx59700z255_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z255_G,
      O => U_DCT1D_nx59700z255
    );
  U_DCT1D_nx59700z239_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z239_G,
      O => U_DCT1D_nx59700z239
    );
  U_DCT1D_reg_databuf_reg_1_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_1_8_DXMUX,
      CE => U_DCT1D_databuf_reg_1_8_CEINV,
      CLK => U_DCT1D_databuf_reg_1_8_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_1_8_FFX_RST,
      O => U_DCT1D_databuf_reg_1_Q(8)
    );
  U_DCT1D_databuf_reg_1_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_1_8_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_1_8_FFX_RST
    );
  U_DCT1D_databuf_reg_1_8_FFX_RSTAND_7506 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_1_8_FFX_RSTAND
    );
  U_DCT1D_nx59700z227_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z227_G,
      O => U_DCT1D_nx59700z227
    );
  U_DCT1D_nx59700z248_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z248_G,
      O => U_DCT1D_nx59700z248
    );
  U_DCT1D_nx59700z236_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z236_G,
      O => U_DCT1D_nx59700z236
    );
  U_DCT1D_nx59700z321_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z321_G,
      O => U_DCT1D_nx59700z321
    );
  U_DCT1D_nx59700z315_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z315_G,
      O => U_DCT1D_nx59700z315
    );
  U_DCT1D_nx59700z309_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z309_G,
      O => U_DCT1D_nx59700z309
    );
  U_DCT1D_nx59700z245_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z245_G,
      O => U_DCT1D_nx59700z245
    );
  U_DCT1D_nx59700z242_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z242_G,
      O => U_DCT1D_nx59700z242
    );
  U_DCT1D_nx59700z330_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z330_G,
      O => U_DCT1D_nx59700z330
    );
  U_DCT1D_nx59700z324_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z324_G,
      O => U_DCT1D_nx59700z324
    );
  U_DCT1D_nx59700z318_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z318_G,
      O => U_DCT1D_nx59700z318
    );
  U_DCT1D_nx59700z312_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z312_G,
      O => U_DCT1D_nx59700z312
    );
  U_DCT1D_nx59700z327_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z327_G,
      O => U_DCT1D_nx59700z327
    );
  U_DCT1D_nx59700z334_XUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z334_F,
      O => U_DCT1D_nx59700z334
    );
  U_DCT1D_nx59700z334_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_nx59700z334_G,
      O => U_DCT1D_nx59700z335
    );
  releaserd_s_DYMUX_7507 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => releaserd_s_BYINVNOT,
      O => releaserd_s_DYMUX
    );
  releaserd_s_BYINV : X_INV
    port map (
      I => U_DCT2D_istate_reg(0),
      O => releaserd_s_BYINVNOT
    );
  releaserd_s_CLKINV_7508 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => releaserd_s_CLKINV
    );
  releaserd_s_CEINV_7509 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc2n582,
      O => releaserd_s_CEINV
    );
  romoaddro0_s_1_DXMUX_7510 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_Q(0),
      O => romoaddro0_s_1_DXMUX
    );
  romoaddro0_s_1_DYMUX_7511 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_Q(0),
      O => romoaddro0_s_1_DYMUX
    );
  romoaddro0_s_1_SRINV_7512 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro0_s_1_SRINV
    );
  romoaddro0_s_1_CLKINV_7513 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro0_s_1_CLKINV
    );
  romoaddro0_s_1_CEINV_7514 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro0_s_1_CEINV
    );
  romoaddro0_s_3_DXMUX_7515 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_Q(0),
      O => romoaddro0_s_3_DXMUX
    );
  romoaddro0_s_3_DYMUX_7516 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_Q(0),
      O => romoaddro0_s_3_DYMUX
    );
  romoaddro0_s_3_SRINV_7517 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro0_s_3_SRINV
    );
  romoaddro0_s_3_CLKINV_7518 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro0_s_3_CLKINV
    );
  romoaddro0_s_3_CEINV_7519 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro0_s_3_CEINV
    );
  romoaddro1_s_1_DXMUX_7520 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_Q(1),
      O => romoaddro1_s_1_DXMUX
    );
  romoaddro1_s_1_DYMUX_7521 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_Q(1),
      O => romoaddro1_s_1_DYMUX
    );
  romoaddro1_s_1_SRINV_7522 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro1_s_1_SRINV
    );
  romoaddro1_s_1_CLKINV_7523 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro1_s_1_CLKINV
    );
  romoaddro1_s_1_CEINV_7524 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro1_s_1_CEINV
    );
  romoaddro1_s_3_DXMUX_7525 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_Q(1),
      O => romoaddro1_s_3_DXMUX
    );
  romoaddro1_s_3_DYMUX_7526 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_Q(1),
      O => romoaddro1_s_3_DYMUX
    );
  romoaddro1_s_3_SRINV_7527 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro1_s_3_SRINV
    );
  romoaddro1_s_3_CLKINV_7528 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro1_s_3_CLKINV
    );
  romoaddro1_s_3_CEINV_7529 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro1_s_3_CEINV
    );
  romoaddro2_s_1_DXMUX_7530 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_Q(2),
      O => romoaddro2_s_1_DXMUX
    );
  romoaddro2_s_1_DYMUX_7531 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_Q(2),
      O => romoaddro2_s_1_DYMUX
    );
  romoaddro2_s_1_SRINV_7532 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro2_s_1_SRINV
    );
  romoaddro2_s_1_CLKINV_7533 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro2_s_1_CLKINV
    );
  romoaddro2_s_1_CEINV_7534 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro2_s_1_CEINV
    );
  romoaddro2_s_3_DXMUX_7535 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_Q(2),
      O => romoaddro2_s_3_DXMUX
    );
  romoaddro2_s_3_DYMUX_7536 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_Q(2),
      O => romoaddro2_s_3_DYMUX
    );
  romoaddro2_s_3_SRINV_7537 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro2_s_3_SRINV
    );
  romoaddro2_s_3_CLKINV_7538 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro2_s_3_CLKINV
    );
  romoaddro2_s_3_CEINV_7539 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro2_s_3_CEINV
    );
  romoaddro3_s_1_DXMUX_7540 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_Q(3),
      O => romoaddro3_s_1_DXMUX
    );
  romoaddro3_s_1_DYMUX_7541 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_Q(3),
      O => romoaddro3_s_1_DYMUX
    );
  romoaddro3_s_1_SRINV_7542 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro3_s_1_SRINV
    );
  romoaddro3_s_1_CLKINV_7543 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro3_s_1_CLKINV
    );
  romoaddro3_s_1_CEINV_7544 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro3_s_1_CEINV
    );
  romoaddro3_s_3_DXMUX_7545 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_Q(3),
      O => romoaddro3_s_3_DXMUX
    );
  romoaddro3_s_3_DYMUX_7546 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_Q(3),
      O => romoaddro3_s_3_DYMUX
    );
  romoaddro3_s_3_SRINV_7547 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro3_s_3_SRINV
    );
  romoaddro3_s_3_CLKINV_7548 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro3_s_3_CLKINV
    );
  romoaddro3_s_3_CEINV_7549 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro3_s_3_CEINV
    );
  romoaddro4_s_1_DXMUX_7550 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_Q(4),
      O => romoaddro4_s_1_DXMUX
    );
  romoaddro4_s_1_DYMUX_7551 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_Q(4),
      O => romoaddro4_s_1_DYMUX
    );
  romoaddro4_s_1_SRINV_7552 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro4_s_1_SRINV
    );
  romoaddro4_s_1_CLKINV_7553 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro4_s_1_CLKINV
    );
  romoaddro4_s_1_CEINV_7554 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro4_s_1_CEINV
    );
  romoaddro4_s_3_DXMUX_7555 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_Q(4),
      O => romoaddro4_s_3_DXMUX
    );
  romoaddro4_s_3_DYMUX_7556 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_Q(4),
      O => romoaddro4_s_3_DYMUX
    );
  romoaddro4_s_3_SRINV_7557 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro4_s_3_SRINV
    );
  romoaddro4_s_3_CLKINV_7558 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro4_s_3_CLKINV
    );
  romoaddro4_s_3_CEINV_7559 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro4_s_3_CEINV
    );
  romoaddro5_s_1_DXMUX_7560 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_Q(5),
      O => romoaddro5_s_1_DXMUX
    );
  romoaddro5_s_1_DYMUX_7561 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_Q(5),
      O => romoaddro5_s_1_DYMUX
    );
  romoaddro5_s_1_SRINV_7562 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro5_s_1_SRINV
    );
  romoaddro5_s_1_CLKINV_7563 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro5_s_1_CLKINV
    );
  romoaddro5_s_1_CEINV_7564 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro5_s_1_CEINV
    );
  romoaddro5_s_3_DXMUX_7565 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_Q(5),
      O => romoaddro5_s_3_DXMUX
    );
  romoaddro5_s_3_DYMUX_7566 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_Q(5),
      O => romoaddro5_s_3_DYMUX
    );
  romoaddro5_s_3_SRINV_7567 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro5_s_3_SRINV
    );
  romoaddro5_s_3_CLKINV_7568 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro5_s_3_CLKINV
    );
  romoaddro5_s_3_CEINV_7569 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro5_s_3_CEINV
    );
  romoaddro6_s_1_DXMUX_7570 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_Q(6),
      O => romoaddro6_s_1_DXMUX
    );
  romoaddro6_s_1_DYMUX_7571 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_Q(6),
      O => romoaddro6_s_1_DYMUX
    );
  romoaddro6_s_1_SRINV_7572 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro6_s_1_SRINV
    );
  romoaddro6_s_1_CLKINV_7573 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro6_s_1_CLKINV
    );
  romoaddro6_s_1_CEINV_7574 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro6_s_1_CEINV
    );
  romoaddro6_s_3_DXMUX_7575 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_Q(6),
      O => romoaddro6_s_3_DXMUX
    );
  romoaddro6_s_3_DYMUX_7576 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_Q(6),
      O => romoaddro6_s_3_DYMUX
    );
  romoaddro6_s_3_SRINV_7577 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro6_s_3_SRINV
    );
  romoaddro6_s_3_CLKINV_7578 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro6_s_3_CLKINV
    );
  romoaddro6_s_3_CEINV_7579 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro6_s_3_CEINV
    );
  romoaddro7_s_1_DXMUX_7580 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_Q(7),
      O => romoaddro7_s_1_DXMUX
    );
  romoaddro7_s_1_DYMUX_7581 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_Q(7),
      O => romoaddro7_s_1_DYMUX
    );
  romoaddro7_s_1_SRINV_7582 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro7_s_1_SRINV
    );
  romoaddro7_s_1_CLKINV_7583 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro7_s_1_CLKINV
    );
  romoaddro7_s_1_CEINV_7584 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro7_s_1_CEINV
    );
  romoaddro7_s_3_DXMUX_7585 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_Q(7),
      O => romoaddro7_s_3_DXMUX
    );
  romoaddro7_s_3_DYMUX_7586 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_Q(7),
      O => romoaddro7_s_3_DYMUX
    );
  romoaddro7_s_3_SRINV_7587 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro7_s_3_SRINV
    );
  romoaddro7_s_3_CLKINV_7588 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro7_s_3_CLKINV
    );
  romoaddro7_s_3_CEINV_7589 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro7_s_3_CEINV
    );
  romoaddro8_s_1_DXMUX_7590 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_6_Q(8),
      O => romoaddro8_s_1_DXMUX
    );
  romoaddro8_s_1_DYMUX_7591 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_7_Q(8),
      O => romoaddro8_s_1_DYMUX
    );
  romoaddro8_s_1_SRINV_7592 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro8_s_1_SRINV
    );
  romoaddro8_s_1_CLKINV_7593 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro8_s_1_CLKINV
    );
  romoaddro8_s_1_CEINV_7594 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro8_s_1_CEINV
    );
  U_DCT2D_ix65206z2349 : X_LUT4
    generic map(
      INIT => X"9393"
    )
    port map (
      ADR0 => romo2datao10_s(0),
      ADR1 => U_DCT2D_rtlc5n1484(10),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z651
    );
  romoaddro8_s_3_DXMUX_7595 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_4_Q(8),
      O => romoaddro8_s_3_DXMUX
    );
  romoaddro8_s_3_DYMUX_7596 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_databuf_reg_5_Q(8),
      O => romoaddro8_s_3_DYMUX
    );
  romoaddro8_s_3_SRINV_7597 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro8_s_3_SRINV
    );
  romoaddro8_s_3_CLKINV_7598 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro8_s_3_CLKINV
    );
  romoaddro8_s_3_CEINV_7599 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro8_s_3_CEINV
    );
  romoaddro0_s_5_DXMUX_7600 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_col_reg(2),
      O => romoaddro0_s_5_DXMUX
    );
  romoaddro0_s_5_DYMUX_7601 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_col_reg(1),
      O => romoaddro0_s_5_DYMUX
    );
  romoaddro0_s_5_SRINV_7602 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => romoaddro0_s_5_SRINV
    );
  romoaddro0_s_5_CLKINV_7603 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => romoaddro0_s_5_CLKINV
    );
  romoaddro0_s_5_CEINV_7604 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcs3,
      O => romoaddro0_s_5_CEINV
    );
  U_DCT2D_ix65206z45559 : X_LUT4
    generic map(
      INIT => X"C939"
    )
    port map (
      ADR0 => rome2datao10_s(2),
      ADR1 => U_DCT2D_rtlc5n1484(12),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao10_s(2),
      O => U_DCT2D_nx65206z645
    );
  U_DCT2D_ix7397z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_6_8_Q,
      ADR1 => U_DCT2D_latchbuf_reg_1_8_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx7397z1
    );
  U_DCT2D_reg_databuf_reg_1_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_1_8_DXMUX,
      CE => U_DCT2D_databuf_reg_1_8_CEINV,
      CLK => U_DCT2D_databuf_reg_1_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_1_8_FFX_RST,
      O => U_DCT2D_databuf_reg_1_Q(8)
    );
  U_DCT2D_databuf_reg_1_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_1_8_FFX_RST
    );
  U_DCT2D_reg_databuf_reg_1_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_1_10_DXMUX,
      CE => U_DCT2D_databuf_reg_1_10_CEINV,
      CLK => U_DCT2D_databuf_reg_1_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_1_10_FFX_RST,
      O => U_DCT2D_databuf_reg_1_Q(10)
    );
  U_DCT2D_databuf_reg_1_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_10_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_1_10_FFX_RST
    );
  U_DCT2D_databuf_reg_1_10_FFX_RSTAND_7605 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_1_10_FFX_RSTAND
    );
  U_DCT1D_ix50549z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_0_Q(1),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_7_Q(1),
      O => U_DCT1D_nx50549z1
    );
  U_DCT1D_reg_databuf_reg_4_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_4_0_DYMUX,
      CE => U_DCT1D_databuf_reg_4_0_CEINV,
      CLK => U_DCT1D_databuf_reg_4_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_4_0_FFY_RST,
      O => U_DCT1D_databuf_reg_4_Q(1)
    );
  U_DCT1D_databuf_reg_4_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_4_0_FFY_RST
    );
  U_DCT1D_reg_databuf_reg_7_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_7_4_DYMUX,
      CE => U_DCT1D_databuf_reg_7_4_CEINV,
      CLK => U_DCT1D_databuf_reg_7_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_7_4_FFY_RST,
      O => U_DCT1D_databuf_reg_7_Q(5)
    );
  U_DCT1D_databuf_reg_7_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_7_4_FFY_RST
    );
  U_DCT1D_ix38135z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_3_Q(4),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_4_Q(4),
      ADR3 => VCC,
      O => U_DCT1D_nx38135z1
    );
  U_DCT1D_reg_databuf_reg_7_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_7_4_DXMUX,
      CE => U_DCT1D_databuf_reg_7_4_CEINV,
      CLK => U_DCT1D_databuf_reg_7_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_7_4_FFX_RST,
      O => U_DCT1D_databuf_reg_7_Q(4)
    );
  U_DCT1D_databuf_reg_7_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_7_4_FFX_RST
    );
  U_DCT1D_ix41126z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_4_Q(7),
      ADR1 => U_DCT1D_latchbuf_reg_3_Q(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx41126z1
    );
  U_DCT2D_reg_databuf_reg_0_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_0_2_DXMUX,
      CE => U_DCT2D_databuf_reg_0_2_CEINV,
      CLK => U_DCT2D_databuf_reg_0_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_0_2_FFX_RST,
      O => U_DCT2D_databuf_reg_0_Q(2)
    );
  U_DCT2D_databuf_reg_0_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_0_2_FFX_RST
    );
  U_DCT2D_ix55995z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_0_5_Q,
      ADR1 => U_DCT2D_latchbuf_reg_7_5_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx55995z1
    );
  U_DCT2D_reg_databuf_reg_0_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_0_4_DYMUX,
      CE => U_DCT2D_databuf_reg_0_4_CEINV,
      CLK => U_DCT2D_databuf_reg_0_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_0_4_FFY_RST,
      O => U_DCT2D_databuf_reg_0_Q(5)
    );
  U_DCT2D_databuf_reg_0_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_0_4_FFY_RST
    );
  U_DCT2D_ix56992z1321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_0_4_Q,
      ADR2 => U_DCT2D_latchbuf_reg_7_4_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx56992z1
    );
  U_DCT2D_reg_databuf_reg_0_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_0_4_DXMUX,
      CE => U_DCT2D_databuf_reg_0_4_CEINV,
      CLK => U_DCT2D_databuf_reg_0_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_0_4_FFX_RST,
      O => U_DCT2D_databuf_reg_0_Q(4)
    );
  U_DCT2D_databuf_reg_0_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_0_4_FFX_RST
    );
  U_DCT2D_ix65206z24310 : X_LUT4
    generic map(
      INIT => X"5A66"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z573,
      ADR1 => rome2datao9_s(12),
      ADR2 => romo2datao9_s(12),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z577
    );
  U_DCT2D_ix418z1321 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_1_1_Q,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_6_1_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx418z1
    );
  U_DCT2D_reg_databuf_reg_1_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_1_0_DYMUX,
      CE => U_DCT2D_databuf_reg_1_0_CEINV,
      CLK => U_DCT2D_databuf_reg_1_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_1_0_FFY_RST,
      O => U_DCT2D_databuf_reg_1_Q(1)
    );
  U_DCT2D_databuf_reg_1_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_1_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_1_0_FFY_RST
    );
  U_DCT2D_ix64957z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_1_0_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_6_0_Q,
      O => U_DCT2D_nx64957z1
    );
  U_DCT2D_ix65206z45535 : X_LUT4
    generic map(
      INIT => X"A599"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1484(18),
      ADR1 => rome2datao10_s(8),
      ADR2 => romo2datao10_s(8),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z627
    );
  U_DCT2D_ix65206z45527 : X_LUT4
    generic map(
      INIT => X"A959"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1484(20),
      ADR1 => rome2datao10_s(10),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao10_s(10),
      O => U_DCT2D_nx65206z621
    );
  U_DCT2D_ix65206z45519 : X_LUT4
    generic map(
      INIT => X"C939"
    )
    port map (
      ADR0 => rome2datao10_s(12),
      ADR1 => U_DCT2D_rtlc5n1484(22),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao10_s(12),
      O => U_DCT2D_nx65206z615
    );
  U_DCT2D_ix65206z1726 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2datao6_s(1),
      ADR1 => VCC,
      ADR2 => romo2datao7_s(0),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z294
    );
  U_DCT2D_ix65206z1709 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao6_s(6),
      ADR2 => romo2datao7_s(5),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z279
    );
  U_DCT2D_ix65206z2121 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2datao6_s(3),
      ADR1 => VCC,
      ADR2 => romo2datao7_s(2),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z288
    );
  U_DCT2D_ix65206z1702 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao6_s(8),
      ADR2 => romo2datao7_s(7),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z273
    );
  U_DCT2D_reg_databuf_reg_0_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_0_0_DYMUX,
      CE => U_DCT2D_databuf_reg_0_0_CEINV,
      CLK => U_DCT2D_databuf_reg_0_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_0_0_FFY_RST,
      O => U_DCT2D_databuf_reg_0_Q(1)
    );
  U_DCT2D_databuf_reg_0_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_0_0_FFY_RST
    );
  U_DCT2D_ix60980z1321 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_0_0_Q,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_7_0_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx60980z1
    );
  U_DCT2D_reg_databuf_reg_0_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_0_0_DXMUX,
      CE => U_DCT2D_databuf_reg_0_0_CEINV,
      CLK => U_DCT2D_databuf_reg_0_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_0_0_FFX_RST,
      O => U_DCT2D_databuf_reg_0_Q(0)
    );
  U_DCT2D_databuf_reg_0_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_0_0_FFX_RST
    );
  U_DCT2D_ix57989z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_0_3_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_7_3_Q,
      O => U_DCT2D_nx57989z1
    );
  U_DCT2D_reg_databuf_reg_0_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_0_2_DYMUX,
      CE => U_DCT2D_databuf_reg_0_2_CEINV,
      CLK => U_DCT2D_databuf_reg_0_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_0_2_FFY_RST,
      O => U_DCT2D_databuf_reg_0_Q(3)
    );
  U_DCT2D_databuf_reg_0_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_0_2_FFY_RST
    );
  U_DCT2D_ix58986z1321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_0_2_Q,
      ADR2 => U_DCT2D_latchbuf_reg_7_2_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx58986z1
    );
  U_DCT2D_ix65206z1423 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao0_s(13),
      ADR1 => romo2datao1_s(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z84
    );
  U_DCT1D_ix35144z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_3_Q(1),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_4_Q(1),
      ADR3 => VCC,
      O => U_DCT1D_nx35144z1
    );
  U_DCT1D_reg_databuf_reg_7_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_7_0_DYMUX,
      CE => U_DCT1D_databuf_reg_7_0_CEINV,
      CLK => U_DCT1D_databuf_reg_7_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_7_0_FFY_RST,
      O => U_DCT1D_databuf_reg_7_Q(1)
    );
  U_DCT1D_databuf_reg_7_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_7_0_FFY_RST
    );
  U_DCT1D_ix34147z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_4_Q(0),
      ADR1 => U_DCT1D_latchbuf_reg_3_Q(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx34147z1
    );
  U_DCT1D_ix54537z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_7_Q(5),
      ADR1 => U_DCT1D_latchbuf_reg_0_Q(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx54537z1
    );
  U_DCT1D_reg_databuf_reg_4_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_4_4_DYMUX,
      CE => U_DCT1D_databuf_reg_4_4_CEINV,
      CLK => U_DCT1D_databuf_reg_4_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_4_4_FFY_RST,
      O => U_DCT1D_databuf_reg_4_Q(5)
    );
  U_DCT1D_databuf_reg_4_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_4_4_FFY_RST
    );
  U_DCT1D_ix53540z1324 : X_LUT4
    generic map(
      INIT => X"C3C3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_0_Q(4),
      ADR2 => U_DCT1D_latchbuf_reg_7_Q(4),
      ADR3 => VCC,
      O => U_DCT1D_nx53540z1
    );
  U_DCT1D_reg_databuf_reg_4_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_4_4_DXMUX,
      CE => U_DCT1D_databuf_reg_4_4_CEINV,
      CLK => U_DCT1D_databuf_reg_4_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_4_4_FFX_RST,
      O => U_DCT1D_databuf_reg_4_Q(4)
    );
  U_DCT1D_databuf_reg_4_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_4_4_FFX_RST
    );
  U_DCT1D_ix56531z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_0_Q(7),
      ADR1 => U_DCT1D_latchbuf_reg_7_Q(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx56531z1
    );
  U_DCT1D_nx57528z1_rt_7606 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx57528z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx57528z1_rt
    );
  U_DCT1D_reg_databuf_reg_4_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_4_6_DYMUX,
      CE => U_DCT1D_databuf_reg_4_6_CEINV,
      CLK => U_DCT1D_databuf_reg_4_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_4_6_FFY_RST,
      O => U_DCT1D_databuf_reg_4_Q(7)
    );
  U_DCT1D_databuf_reg_4_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_4_6_FFY_RST
    );
  U_DCT1D_ix55534z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_7_Q(6),
      ADR1 => U_DCT1D_latchbuf_reg_0_Q(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx55534z1
    );
  U_DCT1D_reg_databuf_reg_4_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_4_6_DXMUX,
      CE => U_DCT1D_databuf_reg_4_6_CEINV,
      CLK => U_DCT1D_databuf_reg_4_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_4_6_FFX_RST,
      O => U_DCT1D_databuf_reg_4_Q(6)
    );
  U_DCT1D_databuf_reg_4_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_4_6_FFX_RST
    );
  U_DCT1D_reg_databuf_reg_4_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_4_8_DXMUX,
      CE => U_DCT1D_databuf_reg_4_8_CEINV,
      CLK => U_DCT1D_databuf_reg_4_8_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_4_8_FFX_RST,
      O => U_DCT1D_databuf_reg_4_Q(8)
    );
  U_DCT1D_databuf_reg_4_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_8_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_4_8_FFX_RST
    );
  U_DCT1D_databuf_reg_4_8_FFX_RSTAND_7607 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_4_8_FFX_RSTAND
    );
  U_DCT2D_ix65206z1687 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao6_s(12),
      ADR1 => romo2datao7_s(11),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z261
    );
  U_DCT2D_ix65206z1698 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao6_s(9),
      ADR2 => VCC,
      ADR3 => romo2datao7_s(8),
      O => U_DCT2D_nx65206z270
    );
  U_DCT2D_ix65206z1680 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romo2datao6_s(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romo2datao7_s(13),
      O => U_DCT2D_nx65206z255
    );
  U_DCT2D_ix65206z2065 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao6_s(11),
      ADR2 => VCC,
      ADR3 => romo2datao7_s(10),
      O => U_DCT2D_nx65206z264
    );
  U_DCT2D_reg_databuf_reg_0_9_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_0_8_DYMUX,
      CE => U_DCT2D_databuf_reg_0_8_CEINV,
      CLK => U_DCT2D_databuf_reg_0_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_0_8_FFY_RST,
      O => U_DCT2D_databuf_reg_0_Q(9)
    );
  U_DCT2D_databuf_reg_0_8_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_0_8_FFY_RST
    );
  U_DCT2D_ix53004z1321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_0_8_Q,
      ADR2 => U_DCT2D_latchbuf_reg_7_8_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx53004z1
    );
  U_DCT2D_nx38337z1_rt_7608 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_nx38337z1,
      O => U_DCT2D_nx38337z1_rt
    );
  U_DCT2D_reg_databuf_reg_0_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_0_8_DXMUX,
      CE => U_DCT2D_databuf_reg_0_8_CEINV,
      CLK => U_DCT2D_databuf_reg_0_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_0_8_FFX_RST,
      O => U_DCT2D_databuf_reg_0_Q(8)
    );
  U_DCT2D_databuf_reg_0_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_0_8_FFX_RST
    );
  U_DCT2D_reg_databuf_reg_0_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_0_10_DXMUX,
      CE => U_DCT2D_databuf_reg_0_10_CEINV,
      CLK => U_DCT2D_databuf_reg_0_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_0_10_FFX_RST,
      O => U_DCT2D_databuf_reg_0_Q(10)
    );
  U_DCT2D_databuf_reg_0_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_10_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_0_10_FFX_RST
    );
  U_DCT2D_databuf_reg_0_10_FFX_RSTAND_7609 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_0_10_FFX_RSTAND
    );
  U_DCT2D_ix65206z1589 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1480(3),
      ADR2 => VCC,
      ADR3 => U_DCT2D_rtlc5n1481(3),
      O => U_DCT2D_nx65206z207
    );
  U_DCT2D_ix65206z1578 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1480(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_rtlc5n1481(5),
      O => U_DCT2D_nx65206z201
    );
  U_DCT2D_ix65206z1593 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1480(2),
      ADR2 => romo2datao2_s(0),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z209
    );
  U_DCT2D_ix65206z45551 : X_LUT4
    generic map(
      INIT => X"C939"
    )
    port map (
      ADR0 => rome2datao10_s(4),
      ADR1 => U_DCT2D_rtlc5n1484(14),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao10_s(4),
      O => U_DCT2D_nx65206z639
    );
  U_DCT2D_ix65206z45543 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => rome2datao10_s(6),
      ADR1 => U_DCT2D_rtlc5n1484(16),
      ADR2 => romo2datao10_s(6),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z633
    );
  U_DCT2D_ix65206z1558 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1480(9),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_rtlc5n1481(9),
      O => U_DCT2D_nx65206z189
    );
  U_DCT2D_ix65206z1584 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1480(4),
      ADR1 => VCC,
      ADR2 => U_DCT2D_rtlc5n1481(4),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z204
    );
  U_DCT2D_ix65206z1568 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1480(7),
      ADR2 => VCC,
      ADR3 => U_DCT2D_rtlc5n1481(7),
      O => U_DCT2D_nx65206z195
    );
  U_DCT2D_ix65206z1573 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1480(6),
      ADR2 => U_DCT2D_rtlc5n1481(6),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z198
    );
  U_DCT1D_reg_databuf_reg_3_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_3_6_DXMUX,
      CE => U_DCT1D_databuf_reg_3_6_CEINV,
      CLK => U_DCT1D_databuf_reg_3_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_3_6_FFX_RST,
      O => U_DCT1D_databuf_reg_3_Q(6)
    );
  U_DCT1D_databuf_reg_3_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_3_6_FFX_RST
    );
  U_DCT1D_reg_databuf_reg_3_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_3_8_DXMUX,
      CE => U_DCT1D_databuf_reg_3_8_CEINV,
      CLK => U_DCT1D_databuf_reg_3_8_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_3_8_FFX_RST,
      O => U_DCT1D_databuf_reg_3_Q(8)
    );
  U_DCT1D_databuf_reg_3_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_8_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_3_8_FFX_RST
    );
  U_DCT1D_databuf_reg_3_8_FFX_RSTAND_7610 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_3_8_FFX_RSTAND
    );
  U_DCT2D_ix65206z1403 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao1_s(5),
      ADR1 => rome2datao0_s(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z68
    );
  U_DCT2D_ix65206z1414 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao0_s(3),
      ADR1 => rome2datao1_s(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z77
    );
  U_DCT2D_ix65206z24333 : X_LUT4
    generic map(
      INIT => X"5A66"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z601,
      ADR1 => rome2datao9_s(4),
      ADR2 => romo2datao9_s(4),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z600
    );
  U_DCT2D_ix65206z24327 : X_LUT4
    generic map(
      INIT => X"3C66"
    )
    port map (
      ADR0 => rome2datao9_s(6),
      ADR1 => U_DCT2D_nx65206z595,
      ADR2 => romo2datao9_s(6),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z594
    );
  U_DCT2D_reg_databuf_reg_3_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_3_0_DXMUX,
      CE => U_DCT2D_databuf_reg_3_0_CEINV,
      CLK => U_DCT2D_databuf_reg_3_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_3_0_FFX_RST,
      O => U_DCT2D_databuf_reg_3_Q(0)
    );
  U_DCT2D_databuf_reg_3_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_3_0_FFX_RST
    );
  U_DCT2D_ix57678z1321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_3_3_Q,
      ADR2 => U_DCT2D_latchbuf_reg_4_3_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx57678z1
    );
  U_DCT2D_reg_databuf_reg_3_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_3_2_DYMUX,
      CE => U_DCT2D_databuf_reg_3_2_CEINV,
      CLK => U_DCT2D_databuf_reg_3_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_3_2_FFY_RST,
      O => U_DCT2D_databuf_reg_3_Q(3)
    );
  U_DCT2D_databuf_reg_3_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_3_2_FFY_RST
    );
  U_DCT2D_ix56681z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_4_2_Q,
      ADR1 => U_DCT2D_latchbuf_reg_3_2_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx56681z1
    );
  U_DCT2D_reg_databuf_reg_3_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_3_2_DXMUX,
      CE => U_DCT2D_databuf_reg_3_2_CEINV,
      CLK => U_DCT2D_databuf_reg_3_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_3_2_FFX_RST,
      O => U_DCT2D_databuf_reg_3_Q(2)
    );
  U_DCT2D_databuf_reg_3_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_3_2_FFX_RST
    );
  U_DCT2D_ix65206z2100 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_nx115_bus(5),
      ADR1 => U_DCT2D_nx65206z553,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z552
    );
  U_DCT2D_ix65206z2116 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z564,
      ADR1 => U_DCT2D_nx115_bus(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z563
    );
  U_DCT2D_ix65206z2089 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z545,
      ADR1 => VCC,
      ADR2 => U_DCT2D_nx115_bus(7),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z544
    );
  U_DCT2D_ix65206z2893 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z557,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_nx115_bus(4),
      O => U_DCT2D_nx65206z556
    );
  U_DCT2D_ix65206z1542 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1480(12),
      ADR1 => VCC,
      ADR2 => U_DCT2D_rtlc5n1481(12),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z180
    );
  U_DCT2D_ix65206z1737 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1480(15),
      ADR1 => U_DCT2D_rtlc5n1481(15),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z171
    );
  U_DCT2D_ix65206z1519 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1480(15),
      ADR1 => U_DCT2D_rtlc5n1481(17),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z165
    );
  U_DCT2D_ix65206z1532 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1480(14),
      ADR2 => U_DCT2D_rtlc5n1481(14),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z174
    );
  U_DCT2D_ix65206z2078 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_nx115_bus(9),
      ADR1 => U_DCT2D_nx65206z537,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z536
    );
  U_DCT2D_ix65206z2094 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z549,
      ADR1 => U_DCT2D_nx115_bus(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z548
    );
  U_DCT2D_ix65206z2068 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z529,
      ADR1 => VCC,
      ADR2 => U_DCT2D_nx115_bus(11),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z528
    );
  U_DCT2D_ix65206z2084 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z541,
      ADR1 => U_DCT2D_nx115_bus(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z540
    );
  U_DCT2D_ix65206z1437 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao0_s(9),
      ADR2 => romo2datao1_s(8),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z96
    );
  U_DCT2D_ix65206z1420 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao0_s(13),
      ADR2 => romo2datao1_s(13),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z81
    );
  U_DCT2D_ix65206z1430 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2datao0_s(11),
      ADR1 => VCC,
      ADR2 => romo2datao1_s(10),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z90
    );
  U_DCT1D_ix49552z1324 : X_LUT4
    generic map(
      INIT => X"C3C3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_0_Q(0),
      ADR2 => U_DCT1D_latchbuf_reg_7_Q(0),
      ADR3 => VCC,
      O => U_DCT1D_nx49552z1
    );
  U_DCT1D_reg_databuf_reg_4_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_4_0_DXMUX,
      CE => U_DCT1D_databuf_reg_4_0_CEINV,
      CLK => U_DCT1D_databuf_reg_4_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_4_0_FFX_RST,
      O => U_DCT1D_databuf_reg_4_Q(0)
    );
  U_DCT1D_databuf_reg_4_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_4_0_FFX_RST
    );
  U_DCT1D_ix52543z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_0_Q(3),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_7_Q(3),
      O => U_DCT1D_nx52543z1
    );
  U_DCT1D_reg_databuf_reg_4_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_4_2_DYMUX,
      CE => U_DCT1D_databuf_reg_4_2_CEINV,
      CLK => U_DCT1D_databuf_reg_4_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_4_2_FFY_RST,
      O => U_DCT1D_databuf_reg_4_Q(3)
    );
  U_DCT1D_databuf_reg_4_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_4_2_FFY_RST
    );
  U_DCT1D_ix51546z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_0_Q(2),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_7_Q(2),
      ADR3 => VCC,
      O => U_DCT1D_nx51546z1
    );
  U_DCT1D_reg_databuf_reg_4_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_4_2_DXMUX,
      CE => U_DCT1D_databuf_reg_4_2_CEINV,
      CLK => U_DCT1D_databuf_reg_4_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_4_2_FFX_RST,
      O => U_DCT1D_databuf_reg_4_Q(2)
    );
  U_DCT1D_databuf_reg_4_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_4_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_4_2_FFX_RST
    );
  U_DCT2D_ix65206z1537 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1480(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_rtlc5n1481(13),
      O => U_DCT2D_nx65206z177
    );
  U_DCT2D_ix65206z1563 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1480(8),
      ADR1 => VCC,
      ADR2 => U_DCT2D_rtlc5n1481(8),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z192
    );
  U_DCT2D_ix65206z1548 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1481(11),
      ADR1 => U_DCT2D_rtlc5n1480(11),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z183
    );
  U_DCT2D_ix65206z1553 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1480(10),
      ADR2 => U_DCT2D_rtlc5n1481(10),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z186
    );
  U_DCT2D_reg_databuf_reg_6_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_6_6_DYMUX,
      CE => U_DCT2D_databuf_reg_6_6_CEINV,
      CLK => U_DCT2D_databuf_reg_6_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_6_6_FFY_RST,
      O => U_DCT2D_databuf_reg_6_Q(7)
    );
  U_DCT2D_databuf_reg_6_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_6_6_FFY_RST
    );
  U_DCT2D_ix45264z1324 : X_LUT4
    generic map(
      INIT => X"C3C3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_2_6_Q,
      ADR2 => U_DCT2D_latchbuf_reg_5_6_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx45264z1
    );
  U_DCT2D_reg_databuf_reg_6_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_6_6_DXMUX,
      CE => U_DCT2D_databuf_reg_6_6_CEINV,
      CLK => U_DCT2D_databuf_reg_6_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_6_6_FFX_RST,
      O => U_DCT2D_databuf_reg_6_Q(6)
    );
  U_DCT2D_databuf_reg_6_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_6_6_FFX_RST
    );
  U_DCT2D_ix48255z1324 : X_LUT4
    generic map(
      INIT => X"C3C3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_2_10_Q,
      ADR2 => U_DCT2D_latchbuf_reg_5_10_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx48255z1
    );
  U_DCT2D_reg_databuf_reg_6_9_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_6_8_DYMUX,
      CE => U_DCT2D_databuf_reg_6_8_CEINV,
      CLK => U_DCT2D_databuf_reg_6_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_6_8_FFY_RST,
      O => U_DCT2D_databuf_reg_6_Q(9)
    );
  U_DCT2D_databuf_reg_6_8_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_6_8_FFY_RST
    );
  U_DCT2D_ix39282z1324 : X_LUT4
    generic map(
      INIT => X"C3C3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_2_0_Q,
      ADR2 => U_DCT2D_latchbuf_reg_5_0_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx39282z1
    );
  U_DCT2D_reg_databuf_reg_6_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_6_0_DXMUX,
      CE => U_DCT2D_databuf_reg_6_0_CEINV,
      CLK => U_DCT2D_databuf_reg_6_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_6_0_FFX_RST,
      O => U_DCT2D_databuf_reg_6_Q(0)
    );
  U_DCT2D_databuf_reg_6_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_6_0_FFX_RST
    );
  U_DCT2D_ix42273z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_2_3_Q,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_5_3_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx42273z1
    );
  U_DCT2D_reg_databuf_reg_6_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_6_2_DYMUX,
      CE => U_DCT2D_databuf_reg_6_2_CEINV,
      CLK => U_DCT2D_databuf_reg_6_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_6_2_FFY_RST,
      O => U_DCT2D_databuf_reg_6_Q(3)
    );
  U_DCT2D_databuf_reg_6_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_6_2_FFY_RST
    );
  U_DCT2D_ix41276z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_2_2_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_5_2_Q,
      O => U_DCT2D_nx41276z1
    );
  U_DCT2D_ix65206z1523 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1480(15),
      ADR2 => U_DCT2D_rtlc5n1481(16),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z168
    );
  U_DCT2D_ix65206z1723 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao6_s(2),
      ADR2 => VCC,
      ADR3 => romo2datao7_s(1),
      O => U_DCT2D_nx65206z291
    );
  U_DCT1D_ix59700z1873 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z412,
      ADR1 => U_DCT1D_rtlc5n1347(11),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z411
    );
  U_DCT1D_ix59700z1891 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z424,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1347(8),
      O => U_DCT1D_nx59700z423
    );
  U_DCT1D_ix59700z1861 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z404,
      ADR1 => U_DCT1D_rtlc5n1347(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z403
    );
  U_DCT1D_reg_databuf_reg_7_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_7_0_DXMUX,
      CE => U_DCT1D_databuf_reg_7_0_CEINV,
      CLK => U_DCT1D_databuf_reg_7_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_7_0_FFX_RST,
      O => U_DCT1D_databuf_reg_7_Q(0)
    );
  U_DCT1D_databuf_reg_7_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_7_0_FFX_RST
    );
  U_DCT1D_ix37138z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_3_Q(3),
      ADR1 => U_DCT1D_latchbuf_reg_4_Q(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx37138z1
    );
  U_DCT1D_reg_databuf_reg_7_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_7_2_DYMUX,
      CE => U_DCT1D_databuf_reg_7_2_CEINV,
      CLK => U_DCT1D_databuf_reg_7_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_7_2_FFY_RST,
      O => U_DCT1D_databuf_reg_7_Q(3)
    );
  U_DCT1D_databuf_reg_7_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_7_2_FFY_RST
    );
  U_DCT1D_ix36141z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_3_Q(2),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_4_Q(2),
      O => U_DCT1D_nx36141z1
    );
  U_DCT1D_reg_databuf_reg_7_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_7_2_DXMUX,
      CE => U_DCT1D_databuf_reg_7_2_CEINV,
      CLK => U_DCT1D_databuf_reg_7_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_7_2_FFX_RST,
      O => U_DCT1D_databuf_reg_7_Q(2)
    );
  U_DCT1D_databuf_reg_7_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_7_2_FFX_RST
    );
  U_DCT1D_ix39132z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_3_Q(5),
      ADR1 => U_DCT1D_latchbuf_reg_4_Q(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx39132z1
    );
  U_DCT2D_ix54001z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_0_7_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_7_7_Q,
      O => U_DCT2D_nx54001z1
    );
  U_DCT2D_reg_databuf_reg_0_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_0_6_DYMUX,
      CE => U_DCT2D_databuf_reg_0_6_CEINV,
      CLK => U_DCT2D_databuf_reg_0_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_0_6_FFY_RST,
      O => U_DCT2D_databuf_reg_0_Q(7)
    );
  U_DCT2D_databuf_reg_0_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_0_6_FFY_RST
    );
  U_DCT2D_ix54998z1321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_0_6_Q,
      ADR2 => U_DCT2D_latchbuf_reg_7_6_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx54998z1
    );
  U_DCT2D_reg_databuf_reg_0_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_0_6_DXMUX,
      CE => U_DCT2D_databuf_reg_0_6_CEINV,
      CLK => U_DCT2D_databuf_reg_0_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_0_6_FFX_RST,
      O => U_DCT2D_databuf_reg_0_Q(6)
    );
  U_DCT2D_databuf_reg_0_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_0_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_0_6_FFX_RST
    );
  U_DCT2D_ix52007z1321 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_0_10_Q,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_7_10_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx52007z1
    );
  U_DCT1D_reg_databuf_reg_7_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_7_6_DYMUX,
      CE => U_DCT1D_databuf_reg_7_6_CEINV,
      CLK => U_DCT1D_databuf_reg_7_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_7_6_FFY_RST,
      O => U_DCT1D_databuf_reg_7_Q(7)
    );
  U_DCT1D_databuf_reg_7_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_7_6_FFY_RST
    );
  U_DCT1D_ix40129z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_3_Q(6),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_4_Q(6),
      ADR3 => VCC,
      O => U_DCT1D_nx40129z1
    );
  U_DCT1D_reg_databuf_reg_7_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_7_6_DXMUX,
      CE => U_DCT1D_databuf_reg_7_6_CEINV,
      CLK => U_DCT1D_databuf_reg_7_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_7_6_FFX_RST,
      O => U_DCT1D_databuf_reg_7_Q(6)
    );
  U_DCT1D_databuf_reg_7_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_7_6_FFX_RST
    );
  U_DCT1D_reg_databuf_reg_7_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_7_8_DXMUX,
      CE => U_DCT1D_databuf_reg_7_8_CEINV,
      CLK => U_DCT1D_databuf_reg_7_8_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_7_8_FFX_RST,
      O => U_DCT1D_databuf_reg_7_Q(8)
    );
  U_DCT1D_databuf_reg_7_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_7_8_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_7_8_FFX_RST
    );
  U_DCT1D_databuf_reg_7_8_FFX_RSTAND_7611 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_7_8_FFX_RSTAND
    );
  U_DCT2D_ix59983z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_0_1_Q,
      ADR1 => U_DCT2D_latchbuf_reg_7_1_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx59983z1
    );
  U_DCT2D_ix65206z1332 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao2_s(13),
      ADR2 => VCC,
      ADR3 => rome2datao3_s(12),
      O => U_DCT2D_nx65206z10
    );
  U_DCT1D_ix59700z1897 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z428,
      ADR1 => U_DCT1D_rtlc5n1347(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z427
    );
  U_DCT1D_ix59700z33456 : X_LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => romodatao6_s(0),
      ADR2 => U_DCT1D_rtlc5n1346(6),
      ADR3 => romedatao4_s(2),
      O => U_DCT1D_nx59700z431
    );
  U_DCT1D_ix59700z1323 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_rtlc5n1359(21),
      ADR2 => VCC,
      ADR3 => U_DCT1D_nx59700z3,
      O => U_DCT1D_nx59700z2
    );
  U_DCT1D_ix59700z1914 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z3,
      ADR2 => U_DCT1D_rtlc5n1359(18),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z440
    );
  U_DCT1D_ix59700z1906 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z3,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1359(20),
      O => U_DCT1D_nx59700z434
    );
  U_DCT1D_ix59700z1364 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao2_s(4),
      ADR2 => VCC,
      ADR3 => romedatao3_s(3),
      O => U_DCT1D_nx59700z37
    );
  U_DCT2D_ix65206z1350 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2datao2_s(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2datao3_s(7),
      O => U_DCT2D_nx65206z25
    );
  U_DCT2D_ix65206z1360 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao2_s(5),
      ADR2 => rome2datao3_s(4),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z34
    );
  U_DCT2D_ix65206z1343 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao2_s(10),
      ADR2 => rome2datao3_s(9),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z19
    );
  U_DCT2D_ix65206z1353 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao3_s(6),
      ADR1 => rome2datao2_s(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z28
    );
  U_DCT2D_ix65206z1684 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao6_s(13),
      ADR1 => romo2datao7_s(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z258
    );
  U_DCT2D_ix55684z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_3_1_Q,
      ADR1 => U_DCT2D_latchbuf_reg_4_1_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx55684z1
    );
  U_DCT2D_reg_databuf_reg_3_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_3_0_DYMUX,
      CE => U_DCT2D_databuf_reg_3_0_CEINV,
      CLK => U_DCT2D_databuf_reg_3_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_3_0_FFY_RST,
      O => U_DCT2D_databuf_reg_3_Q(1)
    );
  U_DCT2D_databuf_reg_3_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_3_0_FFY_RST
    );
  U_DCT2D_ix54687z1321 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_3_0_Q,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_4_0_Q,
      O => U_DCT2D_nx54687z1
    );
  U_DCT1D_reg_databuf_reg_0_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_0_2_DXMUX,
      CE => U_DCT1D_databuf_reg_0_2_CEINV,
      CLK => U_DCT1D_databuf_reg_0_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_0_2_FFX_RST,
      O => U_DCT1D_databuf_reg_0_Q(2)
    );
  U_DCT1D_databuf_reg_0_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_0_2_FFX_RST
    );
  U_DCT1D_ix55995z1321 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_0_Q(5),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_7_Q(5),
      O => U_DCT1D_nx55995z1
    );
  U_DCT1D_reg_databuf_reg_0_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_0_4_DYMUX,
      CE => U_DCT1D_databuf_reg_0_4_CEINV,
      CLK => U_DCT1D_databuf_reg_0_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_0_4_FFY_RST,
      O => U_DCT1D_databuf_reg_0_Q(5)
    );
  U_DCT1D_databuf_reg_0_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_0_4_FFY_RST
    );
  U_DCT1D_ix56992z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_0_Q(4),
      ADR1 => U_DCT1D_latchbuf_reg_7_Q(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx56992z1
    );
  U_DCT1D_reg_databuf_reg_0_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_0_4_DXMUX,
      CE => U_DCT1D_databuf_reg_0_4_CEINV,
      CLK => U_DCT1D_databuf_reg_0_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_0_4_FFX_RST,
      O => U_DCT1D_databuf_reg_0_Q(4)
    );
  U_DCT1D_databuf_reg_0_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_0_4_FFX_RST
    );
  U_DCT1D_ix54001z1321 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_0_Q(7),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_7_Q(7),
      ADR3 => VCC,
      O => U_DCT1D_nx54001z1
    );
  U_DCT2D_reg_databuf_reg_5_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_5_6_DXMUX,
      CE => U_DCT2D_databuf_reg_5_6_CEINV,
      CLK => U_DCT2D_databuf_reg_5_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_5_6_FFX_RST,
      O => U_DCT2D_databuf_reg_5_Q(6)
    );
  U_DCT2D_databuf_reg_5_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_5_6_FFX_RST
    );
  U_DCT2D_ix53390z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_6_10_Q,
      ADR1 => U_DCT2D_latchbuf_reg_1_10_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx53390z1
    );
  U_DCT2D_reg_databuf_reg_5_9_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_5_8_DYMUX,
      CE => U_DCT2D_databuf_reg_5_8_CEINV,
      CLK => U_DCT2D_databuf_reg_5_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_5_8_FFY_RST,
      O => U_DCT2D_databuf_reg_5_Q(9)
    );
  U_DCT2D_databuf_reg_5_8_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_5_8_FFY_RST
    );
  U_DCT2D_ix52393z1324 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_1_8_Q,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_6_8_Q,
      O => U_DCT2D_nx52393z1
    );
  U_DCT2D_nx64938z1_rt_7612 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_nx64938z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx64938z1_rt
    );
  U_DCT2D_reg_databuf_reg_5_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_5_8_DXMUX,
      CE => U_DCT2D_databuf_reg_5_8_CEINV,
      CLK => U_DCT2D_databuf_reg_5_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_5_8_FFX_RST,
      O => U_DCT2D_databuf_reg_5_Q(8)
    );
  U_DCT2D_databuf_reg_5_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_5_8_FFX_RST
    );
  U_DCT1D_reg_databuf_reg_5_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_5_8_DXMUX,
      CE => U_DCT1D_databuf_reg_5_8_CEINV,
      CLK => U_DCT1D_databuf_reg_5_8_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_5_8_FFX_RST,
      O => U_DCT1D_databuf_reg_5_Q(8)
    );
  U_DCT1D_databuf_reg_5_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_8_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_5_8_FFX_RST
    );
  U_DCT1D_databuf_reg_5_8_FFX_RSTAND_7613 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_5_8_FFX_RSTAND
    );
  U_DCT2D_ix45414z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_6_1_Q,
      ADR1 => U_DCT2D_latchbuf_reg_1_1_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx45414z1
    );
  U_DCT2D_reg_databuf_reg_5_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_5_0_DYMUX,
      CE => U_DCT2D_databuf_reg_5_0_CEINV,
      CLK => U_DCT2D_databuf_reg_5_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_5_0_FFY_RST,
      O => U_DCT2D_databuf_reg_5_Q(1)
    );
  U_DCT2D_databuf_reg_5_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_5_0_FFY_RST
    );
  U_DCT2D_ix44417z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_1_0_Q,
      ADR1 => U_DCT2D_latchbuf_reg_6_0_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx44417z1
    );
  U_DCT2D_reg_databuf_reg_5_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_5_0_DXMUX,
      CE => U_DCT2D_databuf_reg_5_0_CEINV,
      CLK => U_DCT2D_databuf_reg_5_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_5_0_FFX_RST,
      O => U_DCT2D_databuf_reg_5_Q(0)
    );
  U_DCT2D_databuf_reg_5_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_5_0_FFX_RST
    );
  U_DCT2D_ix47408z1324 : X_LUT4
    generic map(
      INIT => X"C3C3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_1_3_Q,
      ADR2 => U_DCT2D_latchbuf_reg_6_3_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx47408z1
    );
  U_DCT1D_ix59700z1879 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1347(10),
      ADR1 => U_DCT1D_nx59700z416,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z415
    );
  U_DCT1D_ix59700z1849 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z396,
      ADR1 => U_DCT1D_rtlc5n1347(15),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z395
    );
  U_DCT1D_ix59700z1867 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z408,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1347(12),
      O => U_DCT1D_nx59700z407
    );
  U_DCT1D_ix59700z1837 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z388,
      ADR1 => U_DCT1D_rtlc5n1347(17),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z387
    );
  U_DCT1D_reg_databuf_reg_0_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_0_6_DYMUX,
      CE => U_DCT1D_databuf_reg_0_6_CEINV,
      CLK => U_DCT1D_databuf_reg_0_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_0_6_FFY_RST,
      O => U_DCT1D_databuf_reg_0_Q(7)
    );
  U_DCT1D_databuf_reg_0_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_0_6_FFY_RST
    );
  U_DCT1D_ix54998z1321 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_0_Q(6),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_7_Q(6),
      O => U_DCT1D_nx54998z1
    );
  U_DCT1D_nx53004z1_rt_7614 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx53004z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx53004z1_rt
    );
  U_DCT1D_reg_databuf_reg_0_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_0_6_DXMUX,
      CE => U_DCT1D_databuf_reg_0_6_CEINV,
      CLK => U_DCT1D_databuf_reg_0_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_0_6_FFX_RST,
      O => U_DCT1D_databuf_reg_0_Q(6)
    );
  U_DCT1D_databuf_reg_0_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_0_6_FFX_RST
    );
  U_DCT1D_reg_databuf_reg_0_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_0_8_DXMUX,
      CE => U_DCT1D_databuf_reg_0_8_CEINV,
      CLK => U_DCT1D_databuf_reg_0_8_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_0_8_FFX_RST,
      O => U_DCT1D_databuf_reg_0_Q(8)
    );
  U_DCT1D_databuf_reg_0_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_8_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_0_8_FFX_RST
    );
  U_DCT1D_databuf_reg_0_8_FFX_RSTAND_7615 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_0_8_FFX_RSTAND
    );
  U_DCT1D_ix45414z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_1_Q(1),
      ADR1 => U_DCT1D_latchbuf_reg_6_Q(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx45414z1
    );
  U_DCT2D_ix65206z1712 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao6_s(5),
      ADR2 => VCC,
      ADR3 => romo2datao7_s(4),
      O => U_DCT2D_nx65206z282
    );
  U_DCT2D_ix65206z1695 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao6_s(10),
      ADR2 => VCC,
      ADR3 => romo2datao7_s(9),
      O => U_DCT2D_nx65206z267
    );
  U_DCT2D_ix65206z2093 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao6_s(7),
      ADR2 => romo2datao7_s(6),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z276
    );
  U_DCT2D_reg_databuf_reg_3_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_3_6_DYMUX,
      CE => U_DCT2D_databuf_reg_3_6_CEINV,
      CLK => U_DCT2D_databuf_reg_3_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_3_6_FFY_RST,
      O => U_DCT2D_databuf_reg_3_Q(7)
    );
  U_DCT2D_databuf_reg_3_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_3_6_FFY_RST
    );
  U_DCT2D_ix60669z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_3_6_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_4_6_Q,
      O => U_DCT2D_nx60669z1
    );
  U_DCT2D_reg_databuf_reg_3_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_3_6_DXMUX,
      CE => U_DCT2D_databuf_reg_3_6_CEINV,
      CLK => U_DCT2D_databuf_reg_3_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_3_6_FFX_RST,
      O => U_DCT2D_databuf_reg_3_Q(6)
    );
  U_DCT2D_databuf_reg_3_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_3_6_FFX_RST
    );
  U_DCT2D_ix63660z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_3_10_Q,
      ADR1 => U_DCT2D_latchbuf_reg_4_10_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx63660z1
    );
  U_DCT2D_reg_databuf_reg_3_9_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_3_8_DYMUX,
      CE => U_DCT2D_databuf_reg_3_8_CEINV,
      CLK => U_DCT2D_databuf_reg_3_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_3_8_FFY_RST,
      O => U_DCT2D_databuf_reg_3_Q(9)
    );
  U_DCT2D_databuf_reg_3_8_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_3_8_FFY_RST
    );
  U_DCT2D_ix65206z1364 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao2_s(4),
      ADR2 => VCC,
      ADR3 => rome2datao3_s(3),
      O => U_DCT2D_nx65206z37
    );
  U_DCT2D_reg_databuf_reg_5_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_5_10_DXMUX,
      CE => U_DCT2D_databuf_reg_5_10_CEINV,
      CLK => U_DCT2D_databuf_reg_5_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_5_10_FFX_RST,
      O => U_DCT2D_databuf_reg_5_Q(10)
    );
  U_DCT2D_databuf_reg_5_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_10_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_5_10_FFX_RST
    );
  U_DCT2D_databuf_reg_5_10_FFX_RSTAND_7616 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_5_10_FFX_RSTAND
    );
  U_DCT1D_ix55684z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_4_Q(1),
      ADR1 => U_DCT1D_latchbuf_reg_3_Q(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx55684z1
    );
  U_DCT1D_reg_databuf_reg_3_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_3_0_DYMUX,
      CE => U_DCT1D_databuf_reg_3_0_CEINV,
      CLK => U_DCT1D_databuf_reg_3_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_3_0_FFY_RST,
      O => U_DCT1D_databuf_reg_3_Q(1)
    );
  U_DCT1D_databuf_reg_3_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_3_0_FFY_RST
    );
  U_DCT1D_ix54687z1321 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_3_Q(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_4_Q(0),
      O => U_DCT1D_nx54687z1
    );
  U_DCT2D_ix65206z1410 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao0_s(4),
      ADR2 => rome2datao1_s(3),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z74
    );
  U_DCT1D_reg_databuf_reg_3_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_3_0_DXMUX,
      CE => U_DCT1D_databuf_reg_3_0_CEINV,
      CLK => U_DCT1D_databuf_reg_3_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_3_0_FFX_RST,
      O => U_DCT1D_databuf_reg_3_Q(0)
    );
  U_DCT1D_databuf_reg_3_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_3_0_FFX_RST
    );
  U_DCT1D_ix57678z1321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_3_Q(3),
      ADR2 => U_DCT1D_latchbuf_reg_4_Q(3),
      ADR3 => VCC,
      O => U_DCT1D_nx57678z1
    );
  U_DCT1D_reg_databuf_reg_5_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_5_4_DXMUX,
      CE => U_DCT1D_databuf_reg_5_4_CEINV,
      CLK => U_DCT1D_databuf_reg_5_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_5_4_FFX_RST,
      O => U_DCT1D_databuf_reg_5_Q(4)
    );
  U_DCT1D_databuf_reg_5_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_5_4_FFX_RST
    );
  U_DCT1D_ix51396z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_1_Q(7),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_6_Q(7),
      O => U_DCT1D_nx51396z1
    );
  U_DCT1D_reg_databuf_reg_5_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_5_6_DYMUX,
      CE => U_DCT1D_databuf_reg_5_6_CEINV,
      CLK => U_DCT1D_databuf_reg_5_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_5_6_FFY_RST,
      O => U_DCT1D_databuf_reg_5_Q(7)
    );
  U_DCT1D_databuf_reg_5_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_5_6_FFY_RST
    );
  U_DCT1D_ix50399z1324 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_1_Q(6),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_6_Q(6),
      O => U_DCT1D_nx50399z1
    );
  U_DCT1D_nx52393z1_rt_7617 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx52393z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx52393z1_rt
    );
  U_DCT1D_reg_databuf_reg_5_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_5_6_DXMUX,
      CE => U_DCT1D_databuf_reg_5_6_CEINV,
      CLK => U_DCT1D_databuf_reg_5_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_5_6_FFX_RST,
      O => U_DCT1D_databuf_reg_5_Q(6)
    );
  U_DCT1D_databuf_reg_5_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_5_6_FFX_RST
    );
  U_DCT2D_ix62663z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_3_8_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_4_8_Q,
      O => U_DCT2D_nx62663z1
    );
  U_DCT2D_nx14976z1_rt_7618 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT2D_nx14976z1,
      ADR3 => VCC,
      O => U_DCT2D_nx14976z1_rt
    );
  U_DCT2D_reg_databuf_reg_3_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_3_8_DXMUX,
      CE => U_DCT2D_databuf_reg_3_8_CEINV,
      CLK => U_DCT2D_databuf_reg_3_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_3_8_FFX_RST,
      O => U_DCT2D_databuf_reg_3_Q(8)
    );
  U_DCT2D_databuf_reg_3_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_3_8_FFX_RST
    );
  U_DCT2D_reg_databuf_reg_3_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_3_10_DXMUX,
      CE => U_DCT2D_databuf_reg_3_10_CEINV,
      CLK => U_DCT2D_databuf_reg_3_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_3_10_FFX_RST,
      O => U_DCT2D_databuf_reg_3_Q(10)
    );
  U_DCT2D_databuf_reg_3_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_10_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_3_10_FFX_RST
    );
  U_DCT2D_databuf_reg_3_10_FFX_RSTAND_7619 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_3_10_FFX_RSTAND
    );
  U_DCT2D_ix65206z1357 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao2_s(6),
      ADR1 => rome2datao3_s(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z31
    );
  U_DCT2D_ix65206z1367 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao2_s(3),
      ADR2 => VCC,
      ADR3 => rome2datao3_s(2),
      O => U_DCT2D_nx65206z40
    );
  U_DCT2D_ix59672z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_3_5_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_4_5_Q,
      O => U_DCT2D_nx59672z1
    );
  U_DCT2D_reg_databuf_reg_3_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_3_4_DYMUX,
      CE => U_DCT2D_databuf_reg_3_4_CEINV,
      CLK => U_DCT2D_databuf_reg_3_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_3_4_FFY_RST,
      O => U_DCT2D_databuf_reg_3_Q(5)
    );
  U_DCT2D_databuf_reg_3_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_3_4_FFY_RST
    );
  U_DCT2D_ix58675z1321 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_3_4_Q,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_4_4_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx58675z1
    );
  U_DCT2D_reg_databuf_reg_3_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_3_4_DXMUX,
      CE => U_DCT2D_databuf_reg_3_4_CEINV,
      CLK => U_DCT2D_databuf_reg_3_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_3_4_FFX_RST,
      O => U_DCT2D_databuf_reg_3_Q(4)
    );
  U_DCT2D_databuf_reg_3_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_3_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_3_4_FFX_RST
    );
  U_DCT2D_ix61666z1321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_3_7_Q,
      ADR2 => U_DCT2D_latchbuf_reg_4_7_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx61666z1
    );
  U_DCT2D_ix65206z1336 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao2_s(12),
      ADR1 => rome2datao3_s(11),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z13
    );
  U_DCT2D_ix65206z1346 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao2_s(9),
      ADR2 => VCC,
      ADR3 => rome2datao3_s(8),
      O => U_DCT2D_nx65206z22
    );
  U_DCT2D_ix65206z1329 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao2_s(13),
      ADR1 => rome2datao3_s(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z7
    );
  U_DCT2D_ix65206z1339 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao2_s(11),
      ADR2 => VCC,
      ADR3 => rome2datao3_s(10),
      O => U_DCT2D_nx65206z16
    );
  U_DCT1D_ix59700z1832 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1347(18),
      ADR1 => U_DCT1D_nx59700z384,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z383
    );
  U_DCT1D_ix59700z1822 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z253,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1347(20),
      O => U_DCT1D_nx59700z377
    );
  U_DCT2D_ix40279z1324 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_2_1_Q,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_5_1_Q,
      O => U_DCT2D_nx40279z1
    );
  U_DCT2D_reg_databuf_reg_6_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_6_0_DYMUX,
      CE => U_DCT2D_databuf_reg_6_0_CEINV,
      CLK => U_DCT2D_databuf_reg_6_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_6_0_FFY_RST,
      O => U_DCT2D_databuf_reg_6_Q(1)
    );
  U_DCT2D_databuf_reg_6_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_6_0_FFY_RST
    );
  U_DCT2D_ix65206z1785 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2datao6_s(12),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2datao7_s(11),
      O => U_DCT2D_nx65206z342
    );
  U_DCT2D_ix65206z1795 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2datao6_s(9),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2datao7_s(8),
      O => U_DCT2D_nx65206z351
    );
  U_DCT2D_ix65206z1778 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2datao6_s(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2datao7_s(13),
      O => U_DCT2D_nx65206z336
    );
  U_DCT2D_ix65206z1788 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao6_s(11),
      ADR2 => rome2datao7_s(10),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z345
    );
  U_DCT1D_ix59700z1855 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1347(14),
      ADR1 => U_DCT1D_nx59700z400,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z399
    );
  U_DCT1D_ix59700z1827 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z253,
      ADR1 => U_DCT1D_rtlc5n1347(19),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z380
    );
  U_DCT1D_ix59700z1843 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z392,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1347(16),
      O => U_DCT1D_nx59700z391
    );
  U_DCT2D_ix47258z1324 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_2_8_Q,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_5_8_Q,
      O => U_DCT2D_nx47258z1
    );
  U_DCT2D_nx8385z1_rt_7620 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_nx8385z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx8385z1_rt
    );
  U_DCT2D_reg_databuf_reg_6_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_6_8_DXMUX,
      CE => U_DCT2D_databuf_reg_6_8_CEINV,
      CLK => U_DCT2D_databuf_reg_6_8_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_6_8_FFX_RST,
      O => U_DCT2D_databuf_reg_6_Q(8)
    );
  U_DCT2D_databuf_reg_6_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_8_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_6_8_FFX_RST
    );
  U_DCT2D_reg_databuf_reg_6_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_6_10_DXMUX,
      CE => U_DCT2D_databuf_reg_6_10_CEINV,
      CLK => U_DCT2D_databuf_reg_6_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_6_10_FFX_RST,
      O => U_DCT2D_databuf_reg_6_Q(10)
    );
  U_DCT2D_databuf_reg_6_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_10_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_6_10_FFX_RST
    );
  U_DCT2D_databuf_reg_6_10_FFX_RSTAND_7621 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_databuf_reg_6_10_FFX_RSTAND
    );
  U_DCT1D_ix59983z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_7_Q(1),
      ADR1 => U_DCT1D_latchbuf_reg_0_Q(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59983z1
    );
  U_DCT1D_reg_databuf_reg_0_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_0_0_DYMUX,
      CE => U_DCT1D_databuf_reg_0_0_CEINV,
      CLK => U_DCT1D_databuf_reg_0_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_0_0_FFY_RST,
      O => U_DCT1D_databuf_reg_0_Q(1)
    );
  U_DCT1D_databuf_reg_0_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_0_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_0_0_FFY_RST
    );
  U_DCT2D_reg_databuf_reg_6_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_6_2_DXMUX,
      CE => U_DCT2D_databuf_reg_6_2_CEINV,
      CLK => U_DCT2D_databuf_reg_6_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_6_2_FFX_RST,
      O => U_DCT2D_databuf_reg_6_Q(2)
    );
  U_DCT2D_databuf_reg_6_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_6_2_FFX_RST
    );
  U_DCT2D_ix44267z1324 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_2_5_Q,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_5_5_Q,
      O => U_DCT2D_nx44267z1
    );
  U_DCT2D_reg_databuf_reg_6_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_6_4_DYMUX,
      CE => U_DCT2D_databuf_reg_6_4_CEINV,
      CLK => U_DCT2D_databuf_reg_6_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_6_4_FFY_RST,
      O => U_DCT2D_databuf_reg_6_Q(5)
    );
  U_DCT2D_databuf_reg_6_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_6_4_FFY_RST
    );
  U_DCT2D_ix43270z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_2_4_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_5_4_Q,
      O => U_DCT2D_nx43270z1
    );
  U_DCT2D_reg_databuf_reg_6_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_6_4_DXMUX,
      CE => U_DCT2D_databuf_reg_6_4_CEINV,
      CLK => U_DCT2D_databuf_reg_6_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_6_4_FFX_RST,
      O => U_DCT2D_databuf_reg_6_Q(4)
    );
  U_DCT2D_databuf_reg_6_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_6_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_6_4_FFX_RST
    );
  U_DCT2D_ix46261z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_2_7_Q,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_5_7_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx46261z1
    );
  ix53675z18787 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(1),
      ADR2 => rome2addro4_s(3),
      ADR3 => rome2addro4_s(2),
      O => nx53675z305
    );
  ix53675z25553 : X_LUT4
    generic map(
      INIT => X"50D4"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(1),
      ADR2 => rome2addro4_s(3),
      ADR3 => rome2addro4_s(2),
      O => nx53675z303
    );
  ix53675z12313 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => rome2addro4_s(3),
      ADR1 => rome2addro4_s(1),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(0),
      O => nx53675z311
    );
  ix53675z4958 : X_LUT4
    generic map(
      INIT => X"08CE"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(1),
      ADR2 => rome2addro4_s(3),
      ADR3 => rome2addro4_s(2),
      O => nx53675z306
    );
  ix53675z24569 : X_LUT4
    generic map(
      INIT => X"18A6"
    )
    port map (
      ADR0 => rome2addro4_s(3),
      ADR1 => rome2addro4_s(1),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(0),
      O => nx53675z309
    );
  ix53675z9054 : X_LUT4
    generic map(
      INIT => X"492C"
    )
    port map (
      ADR0 => rome2addro4_s(3),
      ADR1 => rome2addro4_s(1),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(0),
      O => nx53675z312
    );
  ix53675z18002 : X_LUT4
    generic map(
      INIT => X"088E"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(1),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(3),
      O => nx53675z68
    );
  ix53675z61546 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro4_s(3),
      ADR1 => rome2addro4_s(1),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(0),
      O => nx53675z308
    );
  ix53675z15627 : X_LUT4
    generic map(
      INIT => X"18C6"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(3),
      ADR3 => rome2addro9_s(1),
      O => nx53675z601
    );
  ix53675z31158 : X_LUT4
    generic map(
      INIT => X"50D4"
    )
    port map (
      ADR0 => rome2addro9_s(1),
      ADR1 => rome2addro9_s(3),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(0),
      O => nx53675z610
    );
  ix53675z12738 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => rome2addro9_s(3),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(0),
      O => nx53675z606
    );
  ix53675z8476 : X_LUT4
    generic map(
      INIT => X"294A"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(3),
      ADR3 => rome2addro9_s(1),
      O => nx53675z598
    );
  ix53675z35219 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => rome2addro9_s(3),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(0),
      O => nx53675z603
    );
  ix53675z4399 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => rome2addro9_s(3),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(0),
      O => nx53675z607
    );
  ix53675z19228 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => rome2addro9_s(1),
      ADR1 => rome2addro9_s(3),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(0),
      O => nx53675z612
    );
  ix53675z21898 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => rome2addro9_s(3),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(0),
      O => nx53675z604
    );
  ix53675z25997 : X_LUT4
    generic map(
      INIT => X"08CE"
    )
    port map (
      ADR0 => rome2addro9_s(1),
      ADR1 => rome2addro9_s(3),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(0),
      O => nx53675z613
    );
  ix53675z13202 : X_LUT4
    generic map(
      INIT => X"4D04"
    )
    port map (
      ADR0 => rome2addro9_s(1),
      ADR1 => rome2addro9_s(0),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(3),
      O => nx53675z618
    );
  ix53675z40685 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => rome2addro9_s(1),
      ADR1 => rome2addro9_s(3),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(0),
      O => nx53675z609
    );
  ix53675z18291 : X_LUT4
    generic map(
      INIT => X"20B2"
    )
    port map (
      ADR0 => rome2addro4_s(2),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(1),
      ADR3 => rome2addro4_s(0),
      O => nx53675z269
    );
  ix53675z8011 : X_LUT4
    generic map(
      INIT => X"24D2"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => rome2addro4_s(2),
      ADR2 => rome2addro4_s(0),
      ADR3 => rome2addro4_s(3),
      O => nx53675z273
    );
  ix53675z61212 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => rome2addro4_s(2),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(1),
      ADR3 => rome2addro4_s(0),
      O => nx53675z266
    );
  ix53675z14162 : X_LUT4
    generic map(
      INIT => X"2B0A"
    )
    port map (
      ADR0 => rome2addro4_s(2),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(1),
      ADR3 => rome2addro4_s(0),
      O => nx53675z270
    );
  ix53675z18747 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(2),
      ADR2 => rome2addro4_s(1),
      ADR3 => rome2addro4_s(3),
      O => nx53675z275
    );
  ix53675z3915 : X_LUT4
    generic map(
      INIT => X"7310"
    )
    port map (
      ADR0 => rome2addro4_s(2),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(1),
      ADR3 => rome2addro4_s(0),
      O => nx53675z267
    );
  ix53675z15162 : X_LUT4
    generic map(
      INIT => X"1C86"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(2),
      ADR2 => rome2addro4_s(1),
      ADR3 => rome2addro4_s(3),
      O => nx53675z276
    );
  ix53675z12273 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(1),
      O => nx53675z281
    );
  ix53675z7436 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => rome2addro4_s(2),
      ADR2 => rome2addro4_s(0),
      ADR3 => rome2addro4_s(3),
      O => nx53675z272
    );
  ix53675z34754 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(1),
      O => nx53675z278
    );
  ix53675z65640 : X_LUT4
    generic map(
      INIT => X"DD44"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro9_s(2),
      O => nx53675z1458
    );
  ix53675z4093 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => rome2addro6_s(3),
      ADR1 => rome2addro6_s(0),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => nx53675z391
    );
  ix53675z42405 : X_LUT4
    generic map(
      INIT => X"A45A"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(2),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(3),
      O => nx53675z1463
    );
  ix53675z23903 : X_LUT4
    generic map(
      INIT => X"1C30"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1455
    );
  ix53675z59086 : X_LUT4
    generic map(
      INIT => X"AD94"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(2),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(3),
      O => nx53675z1460
    );
  ix53675z45735 : X_LUT4
    generic map(
      INIT => X"C378"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(2),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(3),
      O => nx53675z1461
    );
  ix53675z53372 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(2),
      ADR2 => VCC,
      ADR3 => romo2addro9_s(3),
      O => nx53675z1464
    );
  ix53675z18469 : X_LUT4
    generic map(
      INIT => X"7110"
    )
    port map (
      ADR0 => rome2addro6_s(3),
      ADR1 => rome2addro6_s(0),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => nx53675z393
    );
  ix53675z14340 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => rome2addro6_s(3),
      ADR1 => rome2addro6_s(0),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => nx53675z394
    );
  U_DCT2D_ix65206z31421 : X_LUT4
    generic map(
      INIT => X"72D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1483(7),
      ADR2 => U_DCT2D_rtlc5n1494(7),
      ADR3 => U_DCT2D_rtlc5n1482(7),
      O => U_DCT2D_nx65206z499
    );
  U_DCT2D_ix65206z33587 : X_LUT4
    generic map(
      INIT => X"72D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => romo2datao6_s(0),
      ADR2 => rome2datao4_s(2),
      ADR3 => U_DCT2D_rtlc5n1482(6),
      O => U_DCT2D_nx65206z502
    );
  U_DCT2D_ix65206z31397 : X_LUT4
    generic map(
      INIT => X"72D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1483(11),
      ADR2 => U_DCT2D_rtlc5n1498(11),
      ADR3 => U_DCT2D_rtlc5n1482(11),
      O => U_DCT2D_nx65206z487
    );
  U_DCT2D_ix65206z31415 : X_LUT4
    generic map(
      INIT => X"72D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1483(8),
      ADR2 => U_DCT2D_rtlc5n1498(8),
      ADR3 => U_DCT2D_rtlc5n1482(8),
      O => U_DCT2D_nx65206z496
    );
  U_DCT1D_ix46411z1324 : X_LUT4
    generic map(
      INIT => X"C3C3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_1_Q(2),
      ADR2 => U_DCT1D_latchbuf_reg_6_Q(2),
      ADR3 => VCC,
      O => U_DCT1D_nx46411z1
    );
  U_DCT1D_reg_databuf_reg_5_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_5_2_DXMUX,
      CE => U_DCT1D_databuf_reg_5_2_CEINV,
      CLK => U_DCT1D_databuf_reg_5_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_5_2_FFX_RST,
      O => U_DCT1D_databuf_reg_5_Q(2)
    );
  U_DCT1D_databuf_reg_5_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_5_2_FFX_RST
    );
  U_DCT1D_ix49402z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_1_Q(5),
      ADR1 => U_DCT1D_latchbuf_reg_6_Q(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx49402z1
    );
  U_DCT1D_reg_databuf_reg_5_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_5_4_DYMUX,
      CE => U_DCT1D_databuf_reg_5_4_CEINV,
      CLK => U_DCT1D_databuf_reg_5_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_5_4_FFY_RST,
      O => U_DCT1D_databuf_reg_5_Q(5)
    );
  U_DCT1D_databuf_reg_5_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_5_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_5_4_FFY_RST
    );
  U_DCT1D_ix48405z1324 : X_LUT4
    generic map(
      INIT => X"C3C3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_1_Q(4),
      ADR2 => U_DCT1D_latchbuf_reg_6_Q(4),
      ADR3 => VCC,
      O => U_DCT1D_nx48405z1
    );
  U_DCT2D_reg_databuf_reg_5_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_5_4_DYMUX,
      CE => U_DCT2D_databuf_reg_5_4_CEINV,
      CLK => U_DCT2D_databuf_reg_5_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_5_4_FFY_RST,
      O => U_DCT2D_databuf_reg_5_Q(5)
    );
  U_DCT2D_databuf_reg_5_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_5_4_FFY_RST
    );
  U_DCT2D_ix48405z1324 : X_LUT4
    generic map(
      INIT => X"C3C3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_1_4_Q,
      ADR2 => U_DCT2D_latchbuf_reg_6_4_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx48405z1
    );
  U_DCT2D_reg_databuf_reg_5_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_5_4_DXMUX,
      CE => U_DCT2D_databuf_reg_5_4_CEINV,
      CLK => U_DCT2D_databuf_reg_5_4_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_5_4_FFX_RST,
      O => U_DCT2D_databuf_reg_5_Q(4)
    );
  U_DCT2D_databuf_reg_5_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_4_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_5_4_FFX_RST
    );
  U_DCT2D_ix51396z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_1_7_Q,
      ADR1 => U_DCT2D_latchbuf_reg_6_7_Q,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx51396z1
    );
  U_DCT2D_reg_databuf_reg_5_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_5_6_DYMUX,
      CE => U_DCT2D_databuf_reg_5_6_CEINV,
      CLK => U_DCT2D_databuf_reg_5_6_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_5_6_FFY_RST,
      O => U_DCT2D_databuf_reg_5_Q(7)
    );
  U_DCT2D_databuf_reg_5_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_6_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_5_6_FFY_RST
    );
  U_DCT2D_ix50399z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_1_6_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_6_6_Q,
      O => U_DCT2D_nx50399z1
    );
  U_DCT1D_ix59700z2093 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao4_s(7),
      ADR2 => VCC,
      ADR3 => romodatao5_s(6),
      O => U_DCT1D_nx59700z278
    );
  U_DCT1D_ix59700z1688 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao4_s(12),
      ADR1 => romodatao5_s(11),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z263
    );
  U_DCT1D_ix59700z1698 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao4_s(9),
      ADR1 => romodatao5_s(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z272
    );
  U_DCT1D_ix46261z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_2_Q(7),
      ADR1 => U_DCT1D_latchbuf_reg_5_Q(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx46261z1
    );
  U_DCT1D_reg_databuf_reg_6_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_6_6_DYMUX,
      CE => U_DCT1D_databuf_reg_6_6_CEINV,
      CLK => U_DCT1D_databuf_reg_6_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_6_6_FFY_RST,
      O => U_DCT1D_databuf_reg_6_Q(7)
    );
  U_DCT1D_databuf_reg_6_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_6_6_FFY_RST
    );
  U_DCT1D_ix59700z1512 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao2_s(2),
      ADR1 => romodatao3_s(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z159
    );
  U_DCT1D_ix45264z1324 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_2_Q(6),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_5_Q(6),
      O => U_DCT1D_nx45264z1
    );
  U_DCT1D_nx47258z1_rt_7622 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx47258z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx47258z1_rt
    );
  U_DCT1D_reg_databuf_reg_6_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_6_6_DXMUX,
      CE => U_DCT1D_databuf_reg_6_6_CEINV,
      CLK => U_DCT1D_databuf_reg_6_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_6_6_FFX_RST,
      O => U_DCT1D_databuf_reg_6_Q(6)
    );
  U_DCT1D_databuf_reg_6_6_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_6_6_FFX_RST
    );
  U_DCT1D_reg_databuf_reg_6_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_6_8_DXMUX,
      CE => U_DCT1D_databuf_reg_6_8_CEINV,
      CLK => U_DCT1D_databuf_reg_6_8_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_6_8_FFX_RST,
      O => U_DCT1D_databuf_reg_6_Q(8)
    );
  U_DCT1D_databuf_reg_6_8_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_8_FFX_RSTAND,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_6_8_FFX_RST
    );
  U_DCT1D_databuf_reg_6_8_FFX_RSTAND_7623 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_databuf_reg_6_8_FFX_RSTAND
    );
  U_DCT1D_reg_databuf_reg_3_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_3_4_DYMUX,
      CE => U_DCT1D_databuf_reg_3_4_CEINV,
      CLK => U_DCT1D_databuf_reg_3_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_3_4_FFY_RST,
      O => U_DCT1D_databuf_reg_3_Q(5)
    );
  U_DCT1D_databuf_reg_3_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_3_4_FFY_RST
    );
  U_DCT1D_ix58675z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_4_Q(4),
      ADR1 => U_DCT1D_latchbuf_reg_3_Q(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx58675z1
    );
  U_DCT1D_reg_databuf_reg_3_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_3_4_DXMUX,
      CE => U_DCT1D_databuf_reg_3_4_CEINV,
      CLK => U_DCT1D_databuf_reg_3_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_3_4_FFX_RST,
      O => U_DCT1D_databuf_reg_3_Q(4)
    );
  U_DCT1D_databuf_reg_3_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_3_4_FFX_RST
    );
  U_DCT1D_ix61666z1321 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_3_Q(7),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_4_Q(7),
      ADR3 => VCC,
      O => U_DCT1D_nx61666z1
    );
  U_DCT1D_reg_databuf_reg_3_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_3_6_DYMUX,
      CE => U_DCT1D_databuf_reg_3_6_CEINV,
      CLK => U_DCT1D_databuf_reg_3_6_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_3_6_FFY_RST,
      O => U_DCT1D_databuf_reg_3_Q(7)
    );
  U_DCT1D_databuf_reg_3_6_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_6_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_3_6_FFY_RST
    );
  U_DCT1D_ix60669z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_3_Q(6),
      ADR1 => U_DCT1D_latchbuf_reg_4_Q(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx60669z1
    );
  U_DCT1D_ix59700z1681 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romodatao4_s(13),
      ADR1 => VCC,
      ADR2 => romodatao5_s(13),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z257
    );
  U_DCT1D_ix59700z2065 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romodatao4_s(11),
      ADR1 => VCC,
      ADR2 => romodatao5_s(10),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z266
    );
  U_DCT1D_ix59700z1684 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao4_s(13),
      ADR1 => romodatao5_s(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z260
    );
  U_DCT2D_reg_databuf_reg_5_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_5_2_DYMUX,
      CE => U_DCT2D_databuf_reg_5_2_CEINV,
      CLK => U_DCT2D_databuf_reg_5_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_5_2_FFY_RST,
      O => U_DCT2D_databuf_reg_5_Q(3)
    );
  U_DCT2D_databuf_reg_5_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_5_2_FFY_RST
    );
  U_DCT2D_ix46411z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_1_2_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_6_2_Q,
      O => U_DCT2D_nx46411z1
    );
  U_DCT2D_reg_databuf_reg_5_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_databuf_reg_5_2_DXMUX,
      CE => U_DCT2D_databuf_reg_5_2_CEINV,
      CLK => U_DCT2D_databuf_reg_5_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_databuf_reg_5_2_FFX_RST,
      O => U_DCT2D_databuf_reg_5_Q(2)
    );
  U_DCT2D_databuf_reg_5_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_databuf_reg_5_2_SRINV,
      I1 => GSR,
      O => U_DCT2D_databuf_reg_5_2_FFX_RST
    );
  U_DCT2D_ix49402z1324 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_1_5_Q,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_6_5_Q,
      O => U_DCT2D_nx49402z1
    );
  U_DCT1D_ix59700z1477 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao2_s(12),
      ADR1 => romodatao3_s(11),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z129
    );
  U_DCT1D_ix59700z1657 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao2_s(9),
      ADR1 => romodatao3_s(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z138
    );
  U_DCT1D_ix59700z1470 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romodatao2_s(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romodatao3_s(13),
      O => U_DCT1D_nx59700z123
    );
  U_DCT1D_ix59700z1480 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao2_s(11),
      ADR2 => VCC,
      ADR3 => romodatao3_s(10),
      O => U_DCT1D_nx59700z132
    );
  U_DCT1D_reg_databuf_reg_3_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_3_2_DYMUX,
      CE => U_DCT1D_databuf_reg_3_2_CEINV,
      CLK => U_DCT1D_databuf_reg_3_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_3_2_FFY_RST,
      O => U_DCT1D_databuf_reg_3_Q(3)
    );
  U_DCT1D_databuf_reg_3_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_3_2_FFY_RST
    );
  U_DCT1D_ix56681z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_4_Q(2),
      ADR1 => U_DCT1D_latchbuf_reg_3_Q(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx56681z1
    );
  U_DCT1D_reg_databuf_reg_3_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_3_2_DXMUX,
      CE => U_DCT1D_databuf_reg_3_2_CEINV,
      CLK => U_DCT1D_databuf_reg_3_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_3_2_FFX_RST,
      O => U_DCT1D_databuf_reg_3_Q(2)
    );
  U_DCT1D_databuf_reg_3_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_3_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_3_2_FFX_RST
    );
  U_DCT1D_ix59672z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_3_Q(5),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_4_Q(5),
      O => U_DCT1D_nx59672z1
    );
  U_DCT1D_nx62663z1_rt_7624 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx62663z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx62663z1_rt
    );
  U_DCT2D_ix65206z1379 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao0_s(13),
      ADR2 => VCC,
      ADR3 => rome2datao1_s(12),
      O => U_DCT2D_nx65206z47
    );
  U_DCT2D_ix65206z1813 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao6_s(4),
      ADR2 => VCC,
      ADR3 => rome2datao7_s(3),
      O => U_DCT2D_nx65206z366
    );
  U_DCT2D_ix65206z1806 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rome2datao6_s(6),
      ADR1 => VCC,
      ADR2 => rome2datao7_s(5),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z360
    );
  U_DCT2D_ix65206z1816 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao6_s(3),
      ADR2 => VCC,
      ADR3 => rome2datao7_s(2),
      O => U_DCT2D_nx65206z369
    );
  U_DCT2D_ix65206z1781 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2datao6_s(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2datao7_s(12),
      O => U_DCT2D_nx65206z339
    );
  U_DCT1D_ix40279z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_5_Q(1),
      ADR1 => U_DCT1D_latchbuf_reg_2_Q(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx40279z1
    );
  U_DCT2D_ix65206z1396 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao1_s(7),
      ADR1 => rome2datao0_s(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z62
    );
  U_DCT2D_ix65206z1407 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao0_s(5),
      ADR2 => rome2datao1_s(4),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z71
    );
  U_DCT2D_ix65206z1389 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao0_s(10),
      ADR2 => VCC,
      ADR3 => rome2datao1_s(9),
      O => U_DCT2D_nx65206z56
    );
  U_DCT2D_ix65206z1400 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao0_s(7),
      ADR1 => rome2datao1_s(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z65
    );
  U_DCT2D_ix65206z1382 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao0_s(12),
      ADR1 => rome2datao1_s(11),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z50
    );
  U_DCT2D_ix65206z1393 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao0_s(9),
      ADR1 => rome2datao1_s(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z59
    );
  U_DCT2D_ix65206z1429 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao0_s(13),
      ADR1 => rome2datao1_s(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z44
    );
  U_DCT2D_ix65206z1386 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao0_s(11),
      ADR2 => rome2datao1_s(10),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z53
    );
  U_DCT1D_reg_databuf_reg_6_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_6_0_DYMUX,
      CE => U_DCT1D_databuf_reg_6_0_CEINV,
      CLK => U_DCT1D_databuf_reg_6_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_6_0_FFY_RST,
      O => U_DCT1D_databuf_reg_6_Q(1)
    );
  U_DCT1D_databuf_reg_6_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_6_0_FFY_RST
    );
  U_DCT1D_ix39282z1324 : X_LUT4
    generic map(
      INIT => X"C3C3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_2_Q(0),
      ADR2 => U_DCT1D_latchbuf_reg_5_Q(0),
      ADR3 => VCC,
      O => U_DCT1D_nx39282z1
    );
  U_DCT1D_reg_databuf_reg_6_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_6_0_DXMUX,
      CE => U_DCT1D_databuf_reg_6_0_CEINV,
      CLK => U_DCT1D_databuf_reg_6_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_6_0_FFX_RST,
      O => U_DCT1D_databuf_reg_6_Q(0)
    );
  U_DCT1D_databuf_reg_6_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_6_0_FFX_RST
    );
  U_DCT1D_ix42273z1324 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_2_Q(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_5_Q(3),
      O => U_DCT1D_nx42273z1
    );
  U_DCT1D_reg_databuf_reg_6_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_6_2_DYMUX,
      CE => U_DCT1D_databuf_reg_6_2_CEINV,
      CLK => U_DCT1D_databuf_reg_6_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_6_2_FFY_RST,
      O => U_DCT1D_databuf_reg_6_Q(3)
    );
  U_DCT1D_databuf_reg_6_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_6_2_FFY_RST
    );
  U_DCT1D_ix41276z1324 : X_LUT4
    generic map(
      INIT => X"C3C3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_2_Q(2),
      ADR2 => U_DCT1D_latchbuf_reg_5_Q(2),
      ADR3 => VCC,
      O => U_DCT1D_nx41276z1
    );
  U_DCT1D_ix59700z1491 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao2_s(8),
      ADR2 => romodatao3_s(7),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z141
    );
  U_DCT1D_ix59700z1502 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romodatao2_s(5),
      ADR1 => VCC,
      ADR2 => romodatao3_s(4),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z150
    );
  U_DCT1D_ix59700z1484 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao2_s(10),
      ADR2 => VCC,
      ADR3 => romodatao3_s(9),
      O => U_DCT1D_nx59700z135
    );
  U_DCT1D_ix59700z1495 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao2_s(7),
      ADR2 => VCC,
      ADR3 => romodatao3_s(6),
      O => U_DCT1D_nx59700z144
    );
  U_DCT2D_ix65206z1799 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao6_s(8),
      ADR2 => VCC,
      ADR3 => rome2datao7_s(7),
      O => U_DCT2D_nx65206z354
    );
  U_DCT2D_ix65206z1809 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao7_s(4),
      ADR1 => rome2datao6_s(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z363
    );
  U_DCT2D_ix65206z1792 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2datao6_s(10),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2datao7_s(9),
      O => U_DCT2D_nx65206z348
    );
  U_DCT2D_ix65206z1802 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao6_s(7),
      ADR1 => rome2datao7_s(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z357
    );
  U_DCT1D_reg_databuf_reg_6_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_6_2_DXMUX,
      CE => U_DCT1D_databuf_reg_6_2_CEINV,
      CLK => U_DCT1D_databuf_reg_6_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_6_2_FFX_RST,
      O => U_DCT1D_databuf_reg_6_Q(2)
    );
  U_DCT1D_databuf_reg_6_2_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_2_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_6_2_FFX_RST
    );
  U_DCT1D_ix44267z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latchbuf_reg_2_Q(5),
      ADR2 => VCC,
      ADR3 => U_DCT1D_latchbuf_reg_5_Q(5),
      O => U_DCT1D_nx44267z1
    );
  U_DCT1D_reg_databuf_reg_6_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_6_4_DYMUX,
      CE => U_DCT1D_databuf_reg_6_4_CEINV,
      CLK => U_DCT1D_databuf_reg_6_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_6_4_FFY_RST,
      O => U_DCT1D_databuf_reg_6_Q(5)
    );
  U_DCT1D_databuf_reg_6_4_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_6_4_FFY_RST
    );
  U_DCT1D_ix43270z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_5_Q(4),
      ADR1 => U_DCT1D_latchbuf_reg_2_Q(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx43270z1
    );
  U_DCT1D_reg_databuf_reg_6_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_databuf_reg_6_4_DXMUX,
      CE => U_DCT1D_databuf_reg_6_4_CEINV,
      CLK => U_DCT1D_databuf_reg_6_4_CLKINV,
      SET => GND,
      RST => U_DCT1D_databuf_reg_6_4_FFX_RST,
      O => U_DCT1D_databuf_reg_6_Q(4)
    );
  U_DCT1D_databuf_reg_6_4_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_databuf_reg_6_4_SRINV,
      I1 => GSR,
      O => U_DCT1D_databuf_reg_6_4_FFX_RST
    );
  U_DCT2D_ix65206z31403 : X_LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1483(10),
      ADR2 => U_DCT2D_rtlc5n1482(10),
      ADR3 => U_DCT2D_rtlc5n1498(10),
      O => U_DCT2D_nx65206z490
    );
  U_DCT2D_ix65206z31373 : X_LUT4
    generic map(
      INIT => X"72D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1483(15),
      ADR2 => U_DCT2D_rtlc5n1498(15),
      ADR3 => U_DCT2D_rtlc5n1482(15),
      O => U_DCT2D_nx65206z475
    );
  U_DCT2D_ix65206z31391 : X_LUT4
    generic map(
      INIT => X"72D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1483(12),
      ADR2 => U_DCT2D_rtlc5n1498(12),
      ADR3 => U_DCT2D_rtlc5n1482(12),
      O => U_DCT2D_nx65206z484
    );
  U_DCT1D_ix59700z1343 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao2_s(10),
      ADR2 => romedatao3_s(9),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z19
    );
  U_DCT1D_ix59700z1353 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romedatao3_s(6),
      ADR1 => romedatao2_s(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z28
    );
  U_DCT1D_ix59700z1336 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romedatao2_s(12),
      ADR1 => romedatao3_s(11),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z13
    );
  U_DCT1D_ix59700z1346 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao2_s(9),
      ADR2 => romedatao3_s(8),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z22
    );
  U_DCT2D_ix65206z2058 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_nx115_bus(13),
      ADR1 => U_DCT2D_nx65206z521,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z520
    );
  U_DCT2D_ix65206z2073 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z533,
      ADR1 => VCC,
      ADR2 => U_DCT2D_nx115_bus(10),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z532
    );
  U_DCT2D_ix65206z2050 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z3,
      ADR1 => VCC,
      ADR2 => U_DCT2D_nx115_bus(15),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z514
    );
  U_DCT2D_ix65206z2063 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z525,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_nx115_bus(12),
      O => U_DCT2D_nx65206z524
    );
  U_DCT1D_ix59700z1505 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao2_s(4),
      ADR2 => VCC,
      ADR3 => romodatao3_s(3),
      O => U_DCT1D_nx59700z153
    );
  U_DCT1D_ix59700z1516 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao2_s(1),
      ADR2 => VCC,
      ADR3 => romodatao3_s(0),
      O => U_DCT1D_nx59700z162
    );
  U_DCT1D_ix59700z1498 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao2_s(6),
      ADR1 => romodatao3_s(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z147
    );
  U_DCT1D_ix59700z1509 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao2_s(3),
      ADR2 => VCC,
      ADR3 => romodatao3_s(2),
      O => U_DCT1D_nx59700z156
    );
  U_DCT1D_ix59700z1629 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao2_s(13),
      ADR1 => romodatao3_s(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z126
    );
  U_DCT2D_ix65206z2234 : X_LUT4
    generic map(
      INIT => X"66CC"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_nx65206z567,
      ADR2 => VCC,
      ADR3 => U_DCT2D_rtlc5n1482(5),
      O => U_DCT2D_nx65206z566
    );
  U_DCT2D_ix65206z2112 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z561,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_nx115_bus(3),
      O => U_DCT2D_nx65206z560
    );
  U_DCT2D_ix65206z2238 : X_LUT4
    generic map(
      INIT => X"6A6A"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z570,
      ADR1 => romo2datao4_s(0),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z569
    );
  U_DCT1D_ix59700z1933 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z456,
      ADR2 => U_DCT1D_rtlc5n1359(14),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z455
    );
  U_DCT1D_ix59700z1918 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z444,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1359(17),
      O => U_DCT1D_nx59700z443
    );
  U_DCT1D_ix59700z1910 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1359(19),
      ADR1 => U_DCT1D_nx59700z3,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z437
    );
  U_DCT1D_ix59700z1923 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z448,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1359(16),
      O => U_DCT1D_nx59700z447
    );
  U_DCT2D_ix65206z2261 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1499(15),
      ADR1 => VCC,
      ADR2 => U_DCT2D_rtlc5n1501(15),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z675
    );
  U_DCT2D_ix65206z2278 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1499(12),
      ADR2 => U_DCT2D_rtlc5n1501(12),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z684
    );
  U_DCT2D_ix65206z2266 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1501(14),
      ADR1 => U_DCT2D_rtlc5n1499(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z678
    );
  U_DCT2D_ix65206z2251 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1499(17),
      ADR1 => U_DCT2D_rtlc5n1501(17),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z669
    );
  U_DCT2D_ix65206z2757 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z3,
      ADR1 => U_DCT2D_nx115_bus(18),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z505
    );
  U_DCT2D_ix65206z2291 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1484(9),
      ADR1 => U_DCT2D_rtlc5n1499(9),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z691
    );
  U_DCT2D_ix65206z2409 : X_LUT4
    generic map(
      INIT => X"6C6C"
    )
    port map (
      ADR0 => romo2datao8_s(0),
      ADR1 => U_DCT2D_rtlc5n1499(8),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z693
    );
  U_DCT2D_ix65206z2283 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1499(11),
      ADR2 => U_DCT2D_rtlc5n1501(11),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z687
    );
  U_DCT2D_ix65206z2287 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1499(10),
      ADR1 => U_DCT2D_rtlc5n1501(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z689
    );
  U_DCT2D_ix65206z3225 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1499(13),
      ADR1 => U_DCT2D_rtlc5n1501(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z681
    );
  U_DCT2D_nx65206z1_rt_7625 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_nx65206z1,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z1_rt
    );
  U_DCT2D_ix65206z3151 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1499(20),
      ADR2 => U_DCT2D_rtlc5n1501(20),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z660
    );
  U_DCT2D_ix65206z2224 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1501(22),
      ADR1 => U_DCT2D_rtlc5n1499(22),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z654
    );
  U_DCT1D_ix59700z2095 : X_LUT4
    generic map(
      INIT => X"66CC"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => U_DCT1D_nx59700z490,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1346(5),
      O => U_DCT1D_nx59700z489
    );
  U_DCT1D_ix59700z2099 : X_LUT4
    generic map(
      INIT => X"66AA"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z493,
      ADR1 => romodatao4_s(0),
      ADR2 => VCC,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z492
    );
  U_DCT1D_ix59700z1977 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z487,
      ADR2 => U_DCT1D_rtlc5n1359(6),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z486
    );
  U_DCT1D_ix59700z1961 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z476,
      ADR1 => U_DCT1D_rtlc5n1359(9),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z475
    );
  U_DCT1D_ix59700z1949 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1359(11),
      ADR1 => U_DCT1D_nx59700z468,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z467
    );
  U_DCT1D_ix59700z2615 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z480,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1359(8),
      O => U_DCT1D_nx59700z479
    );
  U_DCT1D_ix59700z1329 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romedatao2_s(13),
      ADR1 => VCC,
      ADR2 => romedatao3_s(13),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z7
    );
  U_DCT1D_ix59700z1339 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao2_s(11),
      ADR2 => VCC,
      ADR3 => romedatao3_s(10),
      O => U_DCT1D_nx59700z16
    );
  U_DCT1D_ix59700z1332 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romedatao2_s(13),
      ADR1 => romedatao3_s(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z10
    );
  U_DCT2D_ix65206z2765 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_nx65206z3,
      ADR2 => VCC,
      ADR3 => U_DCT2D_nx115_bus(17),
      O => U_DCT2D_nx65206z508
    );
  U_DCT2D_ix65206z2054 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z3,
      ADR1 => U_DCT2D_nx115_bus(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z517
    );
  U_DCT2D_ix65206z2046 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_nx65206z3,
      ADR2 => VCC,
      ADR3 => U_DCT2D_nx115_bus(16),
      O => U_DCT2D_nx65206z511
    );
  U_DCT2D_ix65206z50312 : X_LUT4
    generic map(
      INIT => X"D1E2"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1493(6),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1485(6),
      ADR3 => U_DCT2D_rtlc5n1492(6),
      O => U_DCT2D_nx65206z244
    );
  U_DCT2D_ix65206z50294 : X_LUT4
    generic map(
      INIT => X"DE12"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1493(9),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1492(9),
      ADR3 => U_DCT2D_rtlc5n1485(9),
      O => U_DCT2D_nx65206z235
    );
  U_DCT2D_ix65206z50282 : X_LUT4
    generic map(
      INIT => X"CC5A"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1492(11),
      ADR1 => U_DCT2D_rtlc5n1485(11),
      ADR2 => U_DCT2D_rtlc5n1493(11),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z229
    );
  U_DCT2D_ix65206z50300 : X_LUT4
    generic map(
      INIT => X"DE12"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1492(8),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1493(8),
      ADR3 => U_DCT2D_rtlc5n1485(8),
      O => U_DCT2D_nx65206z238
    );
  U_DCT1D_ix59700z1357 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romedatao3_s(5),
      ADR1 => romedatao2_s(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z31
    );
  U_DCT1D_ix59700z1367 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao2_s(3),
      ADR2 => VCC,
      ADR3 => romedatao3_s(2),
      O => U_DCT1D_nx59700z40
    );
  U_DCT1D_ix59700z1350 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao2_s(8),
      ADR2 => VCC,
      ADR3 => romedatao3_s(7),
      O => U_DCT1D_nx59700z25
    );
  U_DCT1D_ix59700z1360 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao2_s(5),
      ADR2 => VCC,
      ADR3 => romedatao3_s(4),
      O => U_DCT1D_nx59700z34
    );
  U_DCT1D_ix59700z2591 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z472,
      ADR2 => U_DCT1D_rtlc5n1359(10),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z471
    );
  U_DCT1D_ix59700z1938 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z460,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1359(13),
      O => U_DCT1D_nx59700z459
    );
  U_DCT1D_ix59700z1928 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1359(15),
      ADR1 => U_DCT1D_nx59700z452,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z451
    );
  U_DCT1D_ix59700z1943 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z464,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1359(12),
      O => U_DCT1D_nx59700z463
    );
  U_DCT2D_ix65206z2241 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1499(19),
      ADR2 => U_DCT2D_rtlc5n1501(19),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z663
    );
  U_DCT2D_ix65206z2256 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1499(16),
      ADR2 => U_DCT2D_rtlc5n1501(16),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z672
    );
  U_DCT2D_ix65206z2246 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1501(18),
      ADR1 => U_DCT2D_rtlc5n1499(18),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z666
    );
  U_DCT2D_ix65206z2229 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1501(21),
      ADR1 => U_DCT2D_rtlc5n1499(21),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z657
    );
  U_DCT2D_ix65206z1734 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao5_s(13),
      ADR1 => rome2datao4_s(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z299
    );
  U_DCT2D_ix65206z1744 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao4_s(11),
      ADR2 => rome2datao5_s(10),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z308
    );
  U_DCT2D_ix65206z2157 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao5_s(12),
      ADR1 => rome2datao4_s(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z302
    );
  U_DCT1D_ix59700z1455 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao1_s(3),
      ADR1 => romodatao0_s(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z111
    );
  U_DCT1D_ix59700z1466 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao0_s(1),
      ADR2 => VCC,
      ADR3 => romodatao1_s(0),
      O => U_DCT1D_nx59700z120
    );
  U_DCT1D_ix59700z1448 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao0_s(6),
      ADR2 => romodatao1_s(5),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z105
    );
  U_DCT1D_ix59700z1601 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao0_s(3),
      ADR1 => romodatao1_s(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z114
    );
  U_DCT1D_ix59700z45340 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => romedatao8_s(11),
      ADR1 => U_DCT1D_rtlc5n1350(19),
      ADR2 => romodatao8_s(11),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z498
    );
  U_DCT1D_reg_ramdatai_s_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramdatai_s_4_DYMUX,
      CE => ramdatai_s_4_CEINV,
      CLK => ramdatai_s_4_CLKINV,
      SET => GND,
      RST => ramdatai_s_4_FFY_RST,
      O => ramdatai_s(5)
    );
  ramdatai_s_4_FFY_RSTOR : X_OR2
    port map (
      I0 => ramdatai_s_4_SRINV,
      I1 => GSR,
      O => ramdatai_s_4_FFY_RST
    );
  U_DCT1D_ix59700z45353 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => romedatao8_s(8),
      ADR1 => U_DCT1D_rtlc5n1350(16),
      ADR2 => romodatao8_s(8),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z507
    );
  U_DCT1D_reg_ramdatai_s_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramdatai_s_4_DXMUX,
      CE => ramdatai_s_4_CEINV,
      CLK => ramdatai_s_4_CLKINV,
      SET => GND,
      RST => ramdatai_s_4_FFX_RST,
      O => ramdatai_s(4)
    );
  ramdatai_s_4_FFX_RSTOR : X_OR2
    port map (
      I0 => ramdatai_s_4_SRINV,
      I1 => GSR,
      O => ramdatai_s_4_FFX_RST
    );
  U_DCT2D_ix65206z31379 : X_LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1483(14),
      ADR2 => U_DCT2D_rtlc5n1482(14),
      ADR3 => U_DCT2D_rtlc5n1498(14),
      O => U_DCT2D_nx65206z478
    );
  U_DCT2D_ix65206z31350 : X_LUT4
    generic map(
      INIT => X"72D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1483(19),
      ADR2 => U_DCT2D_rtlc5n1498(19),
      ADR3 => U_DCT2D_rtlc5n1482(19),
      O => U_DCT2D_nx65206z463
    );
  U_DCT2D_ix65206z31367 : X_LUT4
    generic map(
      INIT => X"72D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1483(16),
      ADR2 => U_DCT2D_rtlc5n1498(16),
      ADR3 => U_DCT2D_rtlc5n1482(16),
      O => U_DCT2D_nx65206z472
    );
  U_DCT2D_ix65206z50318 : X_LUT4
    generic map(
      INIT => X"AA3C"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1485(5),
      ADR1 => U_DCT2D_rtlc5n1492(5),
      ADR2 => U_DCT2D_rtlc5n1493(5),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z247
    );
  U_DCT2D_ix65206z50306 : X_LUT4
    generic map(
      INIT => X"D1E2"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1492(7),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1485(7),
      ADR3 => U_DCT2D_rtlc5n1493(7),
      O => U_DCT2D_nx65206z241
    );
  U_DCT1D_ix59700z1723 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao4_s(2),
      ADR2 => romodatao5_s(1),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z293
    );
  U_DCT1D_ix59700z1716 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romodatao4_s(4),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romodatao5_s(3),
      O => U_DCT1D_nx59700z287
    );
  U_DCT1D_ix59700z1726 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao4_s(1),
      ADR1 => romodatao5_s(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z296
    );
  U_DCT1D_ix59700z1709 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao4_s(6),
      ADR2 => romodatao5_s(5),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z281
    );
  U_DCT1D_ix59700z55462 : X_LUT4
    generic map(
      INIT => X"AA3C"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1346(16),
      ADR1 => romedatao5_s(11),
      ADR2 => romedatao4_s(12),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z305
    );
  U_DCT1D_ix59700z55470 : X_LUT4
    generic map(
      INIT => X"F066"
    )
    port map (
      ADR0 => romedatao4_s(10),
      ADR1 => romedatao5_s(9),
      ADR2 => U_DCT1D_rtlc5n1346(14),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z311
    );
  U_DCT1D_ix59700z55482 : X_LUT4
    generic map(
      INIT => X"AA3C"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1346(11),
      ADR1 => romedatao4_s(7),
      ADR2 => romedatao5_s(6),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z320
    );
  U_DCT1D_ix59700z55474 : X_LUT4
    generic map(
      INIT => X"F066"
    )
    port map (
      ADR0 => romedatao4_s(9),
      ADR1 => romedatao5_s(8),
      ADR2 => U_DCT1D_rtlc5n1346(13),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z314
    );
  U_DCT1D_ix59700z2121 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romodatao4_s(3),
      ADR1 => VCC,
      ADR2 => romodatao5_s(2),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z290
    );
  U_DCT1D_ix59700z1702 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romodatao4_s(8),
      ADR1 => VCC,
      ADR2 => romodatao5_s(7),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z275
    );
  U_DCT1D_ix59700z1712 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao5_s(4),
      ADR1 => romodatao4_s(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z284
    );
  U_DCT1D_ix59700z1695 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao4_s(10),
      ADR2 => romodatao5_s(9),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z269
    );
  U_DCT1D_ix59700z55454 : X_LUT4
    generic map(
      INIT => X"F066"
    )
    port map (
      ADR0 => romedatao5_s(13),
      ADR1 => romedatao4_s(13),
      ADR2 => U_DCT1D_rtlc5n1346(18),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z299
    );
  U_DCT1D_ix59700z55466 : X_LUT4
    generic map(
      INIT => X"AA3C"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1346(15),
      ADR1 => romedatao4_s(11),
      ADR2 => romedatao5_s(10),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z308
    );
  U_DCT1D_ix59700z55458 : X_LUT4
    generic map(
      INIT => X"F066"
    )
    port map (
      ADR0 => romedatao5_s(12),
      ADR1 => romedatao4_s(13),
      ADR2 => U_DCT1D_rtlc5n1346(17),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z302
    );
  U_DCT2D_ix65206z31355 : X_LUT4
    generic map(
      INIT => X"7D28"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1483(18),
      ADR2 => U_DCT2D_rtlc5n1482(18),
      ADR3 => U_DCT2D_rtlc5n1498(18),
      O => U_DCT2D_nx65206z466
    );
  U_DCT2D_ix65206z31345 : X_LUT4
    generic map(
      INIT => X"72D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1483(20),
      ADR2 => U_DCT2D_rtlc5n1498(20),
      ADR3 => U_DCT2D_rtlc5n1482(19),
      O => U_DCT2D_nx65206z460
    );
  U_DCT1D_ix59700z45357 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => romedatao8_s(7),
      ADR1 => U_DCT1D_rtlc5n1350(15),
      ADR2 => romodatao8_s(7),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z510
    );
  U_DCT1D_ix59700z45378 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => romedatao8_s(2),
      ADR1 => U_DCT1D_rtlc5n1350(10),
      ADR2 => romodatao8_s(2),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z524
    );
  U_DCT1D_ix59700z45366 : X_LUT4
    generic map(
      INIT => X"A599"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1350(13),
      ADR1 => romedatao8_s(5),
      ADR2 => romodatao8_s(5),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z516
    );
  U_DCT1D_reg_ramdatai_s_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramdatai_s_0_DYMUX,
      CE => ramdatai_s_0_CEINV,
      CLK => ramdatai_s_0_CLKINV,
      SET => GND,
      RST => ramdatai_s_0_FFY_RST,
      O => ramdatai_s(1)
    );
  ramdatai_s_0_FFY_RSTOR : X_OR2
    port map (
      I0 => ramdatai_s_0_SRINV,
      I1 => GSR,
      O => ramdatai_s_0_FFY_RST
    );
  U_DCT1D_ix59700z45370 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => romedatao8_s(4),
      ADR1 => U_DCT1D_rtlc5n1350(12),
      ADR2 => romodatao8_s(4),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z519
    );
  U_DCT1D_ix59700z55494 : X_LUT4
    generic map(
      INIT => X"CC5A"
    )
    port map (
      ADR0 => romedatao5_s(3),
      ADR1 => U_DCT1D_rtlc5n1346(8),
      ADR2 => romedatao4_s(4),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z329
    );
  U_DCT1D_ix59700z55486 : X_LUT4
    generic map(
      INIT => X"CC5A"
    )
    port map (
      ADR0 => romedatao4_s(6),
      ADR1 => U_DCT1D_rtlc5n1346(10),
      ADR2 => romedatao5_s(5),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z323
    );
  U_DCT1D_ix59700z55478 : X_LUT4
    generic map(
      INIT => X"CC5A"
    )
    port map (
      ADR0 => romedatao5_s(7),
      ADR1 => U_DCT1D_rtlc5n1346(12),
      ADR2 => romedatao4_s(8),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z317
    );
  U_DCT1D_ix59700z55490 : X_LUT4
    generic map(
      INIT => X"F066"
    )
    port map (
      ADR0 => romedatao4_s(5),
      ADR1 => romedatao5_s(4),
      ADR2 => U_DCT1D_rtlc5n1346(9),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z326
    );
  U_DCT2D_ix65206z2221 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2datao4_s(4),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2datao5_s(3),
      O => U_DCT2D_nx65206z329
    );
  U_DCT2D_ix65206z1762 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao5_s(5),
      ADR1 => rome2datao4_s(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z323
    );
  U_DCT2D_ix65206z1773 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao5_s(2),
      ADR1 => rome2datao4_s(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z332
    );
  U_DCT2D_ix65206z1755 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao5_s(7),
      ADR1 => rome2datao4_s(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z317
    );
  U_DCT2D_ix65206z1765 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rome2datao4_s(5),
      ADR1 => VCC,
      ADR2 => rome2datao5_s(4),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z326
    );
  U_DCT2D_ix65206z1885 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1494(9),
      ADR2 => VCC,
      ADR3 => U_DCT2D_rtlc5n1495(9),
      O => U_DCT2D_nx65206z408
    );
  U_DCT2D_ix65206z1873 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1494(11),
      ADR1 => VCC,
      ADR2 => U_DCT2D_rtlc5n1495(11),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z402
    );
  U_DCT2D_ix65206z1891 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1494(8),
      ADR2 => VCC,
      ADR3 => rome2datao6_s(2),
      O => U_DCT2D_nx65206z411
    );
  U_DCT1D_reg_ramdatai_s_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramdatai_s_6_DYMUX,
      CE => ramdatai_s_6_CEINV,
      CLK => ramdatai_s_6_CLKINV,
      SET => GND,
      RST => ramdatai_s_6_FFY_RST,
      O => ramdatai_s(7)
    );
  ramdatai_s_6_FFY_RSTOR : X_OR2
    port map (
      I0 => ramdatai_s_6_SRINV,
      I1 => GSR,
      O => ramdatai_s_6_FFY_RST
    );
  U_DCT1D_ix59700z45344 : X_LUT4
    generic map(
      INIT => X"A599"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1350(18),
      ADR1 => romedatao8_s(10),
      ADR2 => romodatao8_s(10),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z501
    );
  U_DCT1D_reg_ramdatai_s_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramdatai_s_6_DXMUX,
      CE => ramdatai_s_6_CEINV,
      CLK => ramdatai_s_6_CLKINV,
      SET => GND,
      RST => ramdatai_s_6_FFX_RST,
      O => ramdatai_s(6)
    );
  ramdatai_s_6_FFX_RSTOR : X_OR2
    port map (
      I0 => ramdatai_s_6_SRINV,
      I1 => GSR,
      O => ramdatai_s_6_FFX_RST
    );
  U_DCT1D_reg_ramdatai_s_9_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramdatai_s_8_DYMUX,
      CE => ramdatai_s_8_CEINV,
      CLK => ramdatai_s_8_CLKINV,
      SET => GND,
      RST => ramdatai_s_8_FFY_RST,
      O => ramdatai_s(9)
    );
  ramdatai_s_8_FFY_RSTOR : X_OR2
    port map (
      I0 => ramdatai_s_8_SRINV,
      I1 => GSR,
      O => ramdatai_s_8_FFY_RST
    );
  U_DCT1D_ix59700z45335 : X_LUT4
    generic map(
      INIT => X"C399"
    )
    port map (
      ADR0 => romedatao8_s(12),
      ADR1 => U_DCT1D_rtlc5n1350(20),
      ADR2 => romodatao8_s(12),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z495
    );
  U_DCT1D_reg_ramdatai_s_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramdatai_s_8_DXMUX,
      CE => ramdatai_s_8_CEINV,
      CLK => ramdatai_s_8_CLKINV,
      SET => GND,
      RST => ramdatai_s_8_FFX_RST,
      O => ramdatai_s(8)
    );
  ramdatai_s_8_FFX_RSTOR : X_OR2
    port map (
      I0 => ramdatai_s_8_SRINV,
      I1 => GSR,
      O => ramdatai_s_8_FFX_RST
    );
  ix54672z24117 : X_LUT4
    generic map(
      INIT => X"00FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro1_s(2),
      ADR2 => romoaddro1_s(3),
      ADR3 => romoaddro1_s(0),
      O => nx54672z681
    );
  ix54672z23108 : X_LUT4
    generic map(
      INIT => X"02DC"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(2),
      ADR2 => romoaddro1_s(3),
      ADR3 => romoaddro1_s(0),
      O => nx54672z686
    );
  ix54672z51692 : X_LUT4
    generic map(
      INIT => X"DD44"
    )
    port map (
      ADR0 => romoaddro1_s(3),
      ADR1 => romoaddro1_s(2),
      ADR2 => VCC,
      ADR3 => romoaddro1_s(1),
      O => nx54672z690
    );
  ix54672z11067 : X_LUT4
    generic map(
      INIT => X"4242"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => VCC,
      O => nx54672z695
    );
  ix54672z6343 : X_LUT4
    generic map(
      INIT => X"3B3C"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(2),
      ADR2 => romoaddro1_s(3),
      ADR3 => romoaddro1_s(0),
      O => nx54672z687
    );
  ix54672z64552 : X_LUT4
    generic map(
      INIT => X"8E8E"
    )
    port map (
      ADR0 => romoaddro1_s(2),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(1),
      ADR3 => VCC,
      O => nx54672z696
    );
  ix54672z41317 : X_LUT4
    generic map(
      INIT => X"C338"
    )
    port map (
      ADR0 => romoaddro1_s(2),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(1),
      O => nx54672z701
    );
  ix54672z5174 : X_LUT4
    generic map(
      INIT => X"4254"
    )
    port map (
      ADR0 => romoaddro1_s(2),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(1),
      O => nx54672z692
    );
  ix54672z22815 : X_LUT4
    generic map(
      INIT => X"1838"
    )
    port map (
      ADR0 => romoaddro1_s(2),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(1),
      O => nx54672z693
    );
  ix54672z57998 : X_LUT4
    generic map(
      INIT => X"E81E"
    )
    port map (
      ADR0 => romoaddro1_s(2),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(1),
      O => nx54672z698
    );
  U_DCT2D_ix65206z50264 : X_LUT4
    generic map(
      INIT => X"D1E2"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1493(14),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1485(14),
      ADR3 => U_DCT2D_rtlc5n1492(14),
      O => U_DCT2D_nx65206z220
    );
  U_DCT2D_ix65206z50250 : X_LUT4
    generic map(
      INIT => X"8BB8"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1485(17),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1493(17),
      ADR3 => U_DCT2D_rtlc5n1492(15),
      O => U_DCT2D_nx65206z211
    );
  U_DCT2D_nx65206z4_rt_7626 : X_LUT4
    generic map(
      INIT => X"AAAA"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z4,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z4_rt
    );
  U_DCT2D_ix65206z50254 : X_LUT4
    generic map(
      INIT => X"BE14"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1492(15),
      ADR2 => U_DCT2D_rtlc5n1493(16),
      ADR3 => U_DCT2D_rtlc5n1485(16),
      O => U_DCT2D_nx65206z214
    );
  U_DCT1D_ix59700z1463 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao0_s(2),
      ADR1 => romodatao1_s(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z117
    );
  U_DCT2D_ix65206z1748 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao4_s(10),
      ADR1 => rome2datao5_s(9),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z311
    );
  U_DCT2D_ix65206z1758 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2datao4_s(7),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2datao5_s(6),
      O => U_DCT2D_nx65206z320
    );
  U_DCT2D_ix65206z1741 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao4_s(12),
      ADR2 => VCC,
      ADR3 => rome2datao5_s(11),
      O => U_DCT2D_nx65206z305
    );
  U_DCT2D_ix65206z1751 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao4_s(9),
      ADR1 => rome2datao5_s(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z314
    );
  U_DCT1D_ix59700z1441 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romodatao0_s(8),
      ADR1 => VCC,
      ADR2 => romodatao1_s(7),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z99
    );
  U_DCT1D_ix59700z1452 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao1_s(4),
      ADR1 => romodatao0_s(5),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z108
    );
  U_DCT1D_ix59700z1434 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao1_s(9),
      ADR1 => romodatao0_s(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z93
    );
  U_DCT1D_ix59700z1444 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao0_s(7),
      ADR1 => romodatao1_s(6),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z102
    );
  U_DCT1D_ix59700z23970 : X_LUT4
    generic map(
      INIT => X"36C6"
    )
    port map (
      ADR0 => romedatao7_s(8),
      ADR1 => U_DCT1D_nx59700z351,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => romodatao7_s(8),
      O => U_DCT1D_nx59700z350
    );
  U_DCT1D_ix59700z23964 : X_LUT4
    generic map(
      INIT => X"5A66"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z345,
      ADR1 => romedatao7_s(10),
      ADR2 => romodatao7_s(10),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z344
    );
  U_DCT2D_ix65206z1837 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1494(17),
      ADR2 => U_DCT2D_rtlc5n1495(17),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z384
    );
  U_DCT2D_ix65206z1855 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1495(14),
      ADR1 => U_DCT2D_rtlc5n1494(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z393
    );
  U_DCT2D_ix65206z1828 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1494(19),
      ADR1 => U_DCT2D_rtlc5n1495(19),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z378
    );
  U_DCT2D_ix65206z1843 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1494(16),
      ADR2 => U_DCT2D_rtlc5n1495(16),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z387
    );
  U_DCT2D_ix65206z1470 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romo2datao2_s(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romo2datao3_s(13),
      O => U_DCT2D_nx65206z123
    );
  U_DCT2D_ix65206z1480 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao3_s(10),
      ADR1 => romo2datao2_s(11),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z132
    );
  U_DCT2D_ix65206z1629 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao2_s(13),
      ADR1 => romo2datao3_s(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z126
    );
  U_DCT2D_ix65206z50288 : X_LUT4
    generic map(
      INIT => X"D1E2"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1493(10),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1485(10),
      ADR3 => U_DCT2D_rtlc5n1492(10),
      O => U_DCT2D_nx65206z232
    );
  U_DCT2D_ix65206z50270 : X_LUT4
    generic map(
      INIT => X"D1E2"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1493(13),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1485(13),
      ADR3 => U_DCT2D_rtlc5n1492(13),
      O => U_DCT2D_nx65206z223
    );
  U_DCT2D_ix65206z50259 : X_LUT4
    generic map(
      INIT => X"CC5A"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1492(15),
      ADR1 => U_DCT2D_rtlc5n1485(15),
      ADR2 => U_DCT2D_rtlc5n1493(15),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z217
    );
  U_DCT2D_ix65206z50276 : X_LUT4
    generic map(
      INIT => X"DE12"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1493(12),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1492(12),
      ADR3 => U_DCT2D_rtlc5n1485(12),
      O => U_DCT2D_nx65206z226
    );
  U_DCT1D_ix59700z1427 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao0_s(12),
      ADR2 => VCC,
      ADR3 => romodatao1_s(11),
      O => U_DCT1D_nx59700z87
    );
  U_DCT1D_ix59700z1437 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romodatao0_s(9),
      ADR1 => VCC,
      ADR2 => romodatao1_s(8),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z96
    );
  U_DCT1D_ix59700z1420 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romodatao0_s(13),
      ADR1 => VCC,
      ADR2 => romodatao1_s(13),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z81
    );
  U_DCT1D_ix59700z1430 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romodatao0_s(11),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romodatao1_s(10),
      O => U_DCT1D_nx59700z90
    );
  U_DCT1D_ix59700z1423 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao0_s(13),
      ADR1 => romodatao1_s(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z84
    );
  U_DCT2D_ix65206z1512 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao2_s(2),
      ADR2 => VCC,
      ADR3 => romo2datao3_s(1),
      O => U_DCT2D_nx65206z159
    );
  U_DCT2D_ix65206z1505 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao2_s(4),
      ADR1 => romo2datao3_s(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z153
    );
  U_DCT2D_ix65206z1516 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao2_s(1),
      ADR1 => romo2datao3_s(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z162
    );
  U_DCT2D_ix65206z2323 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1495(21),
      ADR1 => U_DCT2D_rtlc5n1494(19),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z372
    );
  U_DCT2D_ix65206z1832 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1495(18),
      ADR1 => U_DCT2D_rtlc5n1494(18),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z381
    );
  U_DCT2D_nx65206z296_rt_7627 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_nx65206z296,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z296_rt
    );
  U_DCT2D_ix65206z1824 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1494(19),
      ADR1 => VCC,
      ADR2 => U_DCT2D_rtlc5n1495(20),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z375
    );
  U_DCT1D_ix59700z1410 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao0_s(4),
      ADR2 => VCC,
      ADR3 => romedatao1_s(3),
      O => U_DCT1D_nx59700z74
    );
  ix53675z13834 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(2),
      O => nx53675z41
    );
  ix53675z18419 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(3),
      O => nx53675z46
    );
  ix53675z3587 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(2),
      O => nx53675z38
    );
  ix53675z25185 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(3),
      O => nx53675z44
    );
  ix53675z18499 : X_LUT4
    generic map(
      INIT => X"7118"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(2),
      ADR3 => rome2addro0_s(1),
      O => nx53675z58
    );
  ix53675z4590 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(3),
      O => nx53675z47
    );
  ix53675z11945 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => rome2addro0_s(1),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(0),
      ADR3 => rome2addro0_s(2),
      O => nx53675z52
    );
  ix53675z33860 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(3),
      O => nx53675z43
    );
  ix53675z61178 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro0_s(1),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(0),
      ADR3 => rome2addro0_s(2),
      O => nx53675z49
    );
  ix53675z8686 : X_LUT4
    generic map(
      INIT => X"2692"
    )
    port map (
      ADR0 => rome2addro0_s(1),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(0),
      ADR3 => rome2addro0_s(3),
      O => nx53675z53
    );
  U_DCT2D_ix65206z1484 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao2_s(10),
      ADR2 => VCC,
      ADR3 => romo2datao3_s(9),
      O => U_DCT2D_nx65206z135
    );
  U_DCT2D_ix65206z1495 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao2_s(7),
      ADR2 => VCC,
      ADR3 => romo2datao3_s(6),
      O => U_DCT2D_nx65206z144
    );
  U_DCT2D_ix65206z1477 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao2_s(12),
      ADR2 => VCC,
      ADR3 => romo2datao3_s(11),
      O => U_DCT2D_nx65206z129
    );
  U_DCT2D_ix65206z1657 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao2_s(9),
      ADR2 => romo2datao3_s(8),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z138
    );
  ix53675z24201 : X_LUT4
    generic map(
      INIT => X"1C86"
    )
    port map (
      ADR0 => rome2addro0_s(1),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(0),
      ADR3 => rome2addro0_s(2),
      O => nx53675z50
    );
  ix53675z4380 : X_LUT4
    generic map(
      INIT => X"2B22"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(3),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(1),
      O => nx53675z592
    );
  ix53675z33876 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(2),
      ADR3 => rome2addro0_s(1),
      O => nx53675z55
    );
  ix53675z27402 : X_LUT4
    generic map(
      INIT => X"6696"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(2),
      ADR3 => rome2addro0_s(1),
      O => nx53675z59
    );
  ix53675z18756 : X_LUT4
    generic map(
      INIT => X"7110"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(3),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(1),
      O => nx53675z594
    );
  ix53675z16899 : X_LUT4
    generic map(
      INIT => X"2DD2"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(2),
      ADR3 => rome2addro0_s(1),
      O => nx53675z56
    );
  ix53675z14627 : X_LUT4
    generic map(
      INIT => X"20F2"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(3),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(1),
      O => nx53675z595
    );
  ix53675z19212 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(3),
      ADR3 => rome2addro9_s(1),
      O => nx53675z600
    );
  ix53675z61677 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(3),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(1),
      O => nx53675z591
    );
  ix53675z7901 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(3),
      ADR3 => rome2addro9_s(1),
      O => nx53675z597
    );
  ix53675z25273 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z108
    );
  ix53675z26245 : X_LUT4
    generic map(
      INIT => X"4B24"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(2),
      O => nx53675z32
    );
  ix53675z12033 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => rome2addro1_s(1),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(3),
      ADR3 => rome2addro1_s(2),
      O => nx53675z116
    );
  ix53675z61266 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro1_s(1),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(3),
      ADR3 => rome2addro1_s(2),
      O => nx53675z113
    );
  ix53675z8774 : X_LUT4
    generic map(
      INIT => X"5924"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(3),
      ADR3 => rome2addro1_s(1),
      O => nx53675z117
    );
  ix53675z12369 : X_LUT4
    generic map(
      INIT => X"088E"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(2),
      O => nx53675z34
    );
  ix53675z24289 : X_LUT4
    generic map(
      INIT => X"3492"
    )
    port map (
      ADR0 => rome2addro1_s(1),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(3),
      ADR3 => rome2addro1_s(2),
      O => nx53675z114
    );
  ix53675z24180 : X_LUT4
    generic map(
      INIT => X"4694"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(2),
      O => nx53675z35
    );
  ix53675z11929 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(2),
      O => nx53675z40
    );
  ix53675z7370 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(2),
      O => nx53675z31
    );
  ix53675z61162 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(2),
      O => nx53675z37
    );
  U_DCT2D_ix65206z1926 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao4_s(6),
      ADR2 => romo2datao5_s(5),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z439
    );
  U_DCT2D_ix65206z1937 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao4_s(3),
      ADR1 => romo2datao5_s(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z448
    );
  U_DCT2D_ix65206z1919 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romo2datao4_s(8),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romo2datao5_s(7),
      O => U_DCT2D_nx65206z433
    );
  U_DCT2D_ix65206z1930 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao4_s(5),
      ADR2 => VCC,
      ADR3 => romo2datao5_s(4),
      O => U_DCT2D_nx65206z442
    );
  U_DCT1D_ix59700z1403 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao0_s(6),
      ADR2 => VCC,
      ADR3 => romedatao1_s(5),
      O => U_DCT1D_nx59700z68
    );
  U_DCT1D_ix59700z1414 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romedatao0_s(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romedatao1_s(2),
      O => U_DCT1D_nx59700z77
    );
  U_DCT1D_ix59700z1396 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao0_s(8),
      ADR2 => VCC,
      ADR3 => romedatao1_s(7),
      O => U_DCT1D_nx59700z62
    );
  U_DCT1D_ix59700z1407 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao0_s(5),
      ADR2 => romedatao1_s(4),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z71
    );
  U_DCT1D_ix59700z50259 : X_LUT4
    generic map(
      INIT => X"A3AC"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1348(15),
      ADR1 => U_DCT1D_rtlc5n1355(15),
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_rtlc5n1354(15),
      O => U_DCT1D_nx59700z217
    );
  U_DCT1D_ix59700z50276 : X_LUT4
    generic map(
      INIT => X"A3AC"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1348(12),
      ADR1 => U_DCT1D_rtlc5n1354(12),
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_rtlc5n1355(12),
      O => U_DCT1D_nx59700z226
    );
  U_DCT1D_ix59700z50250 : X_LUT4
    generic map(
      INIT => X"DE12"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1355(17),
      ADR1 => U_DCT1D_state_reg(0),
      ADR2 => U_DCT1D_rtlc5n1354(15),
      ADR3 => U_DCT1D_rtlc5n1348(17),
      O => U_DCT1D_nx59700z211
    );
  U_DCT1D_ix59700z50264 : X_LUT4
    generic map(
      INIT => X"DE12"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1354(14),
      ADR1 => U_DCT1D_state_reg(0),
      ADR2 => U_DCT1D_rtlc5n1355(14),
      ADR3 => U_DCT1D_rtlc5n1348(14),
      O => U_DCT1D_nx59700z220
    );
  U_DCT1D_ix59700z1429 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romedatao0_s(13),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romedatao1_s(13),
      O => U_DCT1D_nx59700z44
    );
  U_DCT1D_ix59700z1386 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romedatao0_s(11),
      ADR1 => romedatao1_s(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z53
    );
  U_DCT1D_ix59700z1379 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romedatao0_s(13),
      ADR1 => romedatao1_s(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z47
    );
  U_DCT2D_ix65206z1498 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao2_s(6),
      ADR2 => VCC,
      ADR3 => romo2datao3_s(5),
      O => U_DCT2D_nx65206z147
    );
  U_DCT2D_ix65206z1509 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao3_s(2),
      ADR1 => romo2datao2_s(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z156
    );
  U_DCT2D_ix65206z1491 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao2_s(8),
      ADR1 => romo2datao3_s(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z141
    );
  U_DCT2D_ix65206z1502 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao2_s(5),
      ADR2 => VCC,
      ADR3 => romo2datao3_s(4),
      O => U_DCT2D_nx65206z150
    );
  U_DCT1D_ix59700z50318 : X_LUT4
    generic map(
      INIT => X"DE12"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1355(5),
      ADR1 => U_DCT1D_state_reg(0),
      ADR2 => U_DCT1D_rtlc5n1354(5),
      ADR3 => U_DCT1D_rtlc5n1348(5),
      O => U_DCT1D_nx59700z247
    );
  U_DCT1D_ix59700z50306 : X_LUT4
    generic map(
      INIT => X"A3AC"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1348(7),
      ADR1 => U_DCT1D_rtlc5n1355(7),
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_rtlc5n1354(7),
      O => U_DCT1D_nx59700z241
    );
  U_DCT1D_ix59700z50294 : X_LUT4
    generic map(
      INIT => X"BE14"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => U_DCT1D_rtlc5n1355(9),
      ADR2 => U_DCT1D_rtlc5n1354(9),
      ADR3 => U_DCT1D_rtlc5n1348(9),
      O => U_DCT1D_nx59700z235
    );
  U_DCT1D_ix59700z50312 : X_LUT4
    generic map(
      INIT => X"DE12"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1354(6),
      ADR1 => U_DCT1D_state_reg(0),
      ADR2 => U_DCT1D_rtlc5n1355(6),
      ADR3 => U_DCT1D_rtlc5n1348(6),
      O => U_DCT1D_nx59700z244
    );
  U_DCT2D_ix65206z1861 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1494(13),
      ADR2 => U_DCT2D_rtlc5n1495(13),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z396
    );
  U_DCT2D_ix65206z1879 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1495(10),
      ADR1 => U_DCT2D_rtlc5n1494(10),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z405
    );
  U_DCT2D_ix65206z1849 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1494(15),
      ADR1 => U_DCT2D_rtlc5n1495(15),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z390
    );
  U_DCT2D_ix65206z1867 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1494(12),
      ADR2 => VCC,
      ADR3 => U_DCT2D_rtlc5n1495(12),
      O => U_DCT2D_nx65206z399
    );
  U_DCT1D_ix59700z1389 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romedatao0_s(10),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romedatao1_s(9),
      O => U_DCT1D_nx59700z56
    );
  U_DCT1D_ix59700z1400 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao0_s(7),
      ADR2 => VCC,
      ADR3 => romedatao1_s(6),
      O => U_DCT1D_nx59700z65
    );
  U_DCT1D_ix59700z1382 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao0_s(12),
      ADR2 => VCC,
      ADR3 => romedatao1_s(11),
      O => U_DCT1D_nx59700z50
    );
  U_DCT1D_ix59700z1393 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romedatao0_s(9),
      ADR1 => romedatao1_s(8),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z59
    );
  ix53675z26333 : X_LUT4
    generic map(
      INIT => X"294A"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(3),
      O => nx53675z96
    );
  ix53675z12017 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z104
    );
  ix53675z24268 : X_LUT4
    generic map(
      INIT => X"6318"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(3),
      O => nx53675z99
    );
  ix53675z3675 : X_LUT4
    generic map(
      INIT => X"44D4"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z102
    );
  ix53675z13922 : X_LUT4
    generic map(
      INIT => X"4F04"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z105
    );
  ix53675z18507 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z110
    );
  ix53675z61250 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z101
    );
  ix53675z33948 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z107
    );
  ix53675z4678 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z111
    );
  U_DCT1D_ix59700z23982 : X_LUT4
    generic map(
      INIT => X"3C66"
    )
    port map (
      ADR0 => romedatao7_s(4),
      ADR1 => U_DCT1D_nx59700z363,
      ADR2 => romodatao7_s(4),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z362
    );
  U_DCT1D_ix59700z23976 : X_LUT4
    generic map(
      INIT => X"3C66"
    )
    port map (
      ADR0 => romedatao7_s(6),
      ADR1 => U_DCT1D_nx59700z357,
      ADR2 => romodatao7_s(6),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z356
    );
  ix54672z14794 : X_LUT4
    generic map(
      INIT => X"2962"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(0),
      O => nx54672z17
    );
  ix54672z28429 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro0_s(0),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(1),
      ADR3 => romeaddro0_s(2),
      O => nx54672z63
    );
  ix54672z7643 : X_LUT4
    generic map(
      INIT => X"4B24"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(0),
      O => nx54672z14
    );
  ix54672z43584 : X_LUT4
    generic map(
      INIT => X"A1A0"
    )
    port map (
      ADR0 => romoaddro0_s(2),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(0),
      ADR3 => romoaddro0_s(3),
      O => nx54672z630
    );
  ix54672z13736 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romeaddro0_s(1),
      ADR3 => romeaddro0_s(2),
      O => nx54672z64
    );
  ix54672z41214 : X_LUT4
    generic map(
      INIT => X"9866"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(3),
      O => nx54672z624
    );
  ix54672z28426 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro0_s(0),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(1),
      ADR3 => romeaddro0_s(2),
      O => U1_ROME0_modgen_rom_ix2_nx_rm64_16_u
    );
  ix54672z1567 : X_LUT4
    generic map(
      INIT => X"2222"
    )
    port map (
      ADR0 => romeaddro0_s(0),
      ADR1 => romeaddro0_s(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z61
    );
  ix54672z57895 : X_LUT4
    generic map(
      INIT => X"D992"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(3),
      O => nx54672z621
    );
  ix54672z52181 : X_LUT4
    generic map(
      INIT => X"C33C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(3),
      O => nx54672z625
    );
  U_DCT1D_ix59700z1737 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1345(15),
      ADR1 => U_DCT1D_rtlc5n1344(15),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z171
    );
  U_DCT1D_ix59700z1542 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1344(12),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1345(12),
      O => U_DCT1D_nx59700z180
    );
  U_DCT1D_ix59700z1519 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_rtlc5n1344(15),
      ADR2 => U_DCT1D_rtlc5n1345(17),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z165
    );
  U_DCT1D_ix59700z1532 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1345(14),
      ADR1 => U_DCT1D_rtlc5n1344(14),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z174
    );
  U_DCT1D_nx59700z78_rt_7628 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT1D_nx59700z78,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z78_rt
    );
  ix53675z21065 : X_LUT4
    generic map(
      INIT => X"20BA"
    )
    port map (
      ADR0 => rome2addro0_s(1),
      ADR1 => rome2addro0_s(0),
      ADR2 => rome2addro0_s(3),
      ADR3 => rome2addro0_s(2),
      O => nx53675z20
    );
  ix53675z11905 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => rome2addro0_s(1),
      ADR1 => rome2addro0_s(0),
      ADR2 => rome2addro0_s(3),
      ADR3 => rome2addro0_s(2),
      O => nx53675z22
    );
  ix53675z18395 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => rome2addro0_s(2),
      ADR1 => rome2addro0_s(1),
      ADR2 => rome2addro0_s(3),
      ADR3 => rome2addro0_s(0),
      O => nx53675z28
    );
  ix53675z3566 : X_LUT4
    generic map(
      INIT => X"0C8E"
    )
    port map (
      ADR0 => rome2addro0_s(1),
      ADR1 => rome2addro0_s(0),
      ADR2 => rome2addro0_s(3),
      ADR3 => rome2addro0_s(2),
      O => nx53675z23
    );
  ix53675z30325 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => rome2addro0_s(2),
      ADR1 => rome2addro0_s(1),
      ADR2 => rome2addro0_s(3),
      ADR3 => rome2addro0_s(0),
      O => nx53675z26
    );
  ix53675z25164 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => rome2addro0_s(2),
      ADR1 => rome2addro0_s(1),
      ADR2 => rome2addro0_s(3),
      ADR3 => rome2addro0_s(0),
      O => nx53675z29
    );
  ix53675z18748 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => rome2addro9_s(3),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(0),
      O => nx53675z588
    );
  ix53675z39852 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => rome2addro0_s(2),
      ADR1 => rome2addro0_s(1),
      ADR2 => rome2addro0_s(3),
      ADR3 => rome2addro0_s(0),
      O => nx53675z25
    );
  U_DCT1D_ix59700z23959 : X_LUT4
    generic map(
      INIT => X"5A66"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z335,
      ADR1 => romedatao7_s(12),
      ADR2 => romodatao7_s(12),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z339
    );
  U_DCT1D_ix59700z1589 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1345(3),
      ADR1 => U_DCT1D_rtlc5n1344(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z207
    );
  U_DCT1D_ix59700z1593 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romodatao2_s(0),
      ADR1 => U_DCT1D_rtlc5n1344(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z209
    );
  U_DCT1D_ix59700z1578 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_rtlc5n1344(5),
      ADR2 => U_DCT1D_rtlc5n1345(5),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z201
    );
  U_DCT1D_ix59700z1568 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1345(7),
      ADR1 => U_DCT1D_rtlc5n1344(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z195
    );
  U_DCT2D_ix65206z1912 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao4_s(10),
      ADR2 => VCC,
      ADR3 => romo2datao5_s(9),
      O => U_DCT2D_nx65206z427
    );
  U_DCT2D_ix65206z1923 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao4_s(7),
      ADR2 => VCC,
      ADR3 => romo2datao5_s(6),
      O => U_DCT2D_nx65206z436
    );
  U_DCT2D_ix65206z1905 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao5_s(11),
      ADR1 => romo2datao4_s(12),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z421
    );
  U_DCT2D_ix65206z1916 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao4_s(9),
      ADR2 => VCC,
      ADR3 => romo2datao5_s(8),
      O => U_DCT2D_nx65206z430
    );
  ix53675z14720 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(0),
      ADR3 => rome2addro10_s(3),
      O => nx53675z660
    );
  ix53675z4473 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(0),
      ADR3 => rome2addro10_s(3),
      O => nx53675z657
    );
  ix53675z26427 : X_LUT4
    generic map(
      INIT => X"6138"
    )
    port map (
      ADR0 => rome2addro2_s(0),
      ADR1 => rome2addro2_s(1),
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(3),
      O => nx53675z161
    );
  ix53675z7994 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(2),
      O => nx53675z662
    );
  ix53675z15720 : X_LUT4
    generic map(
      INIT => X"4B24"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(2),
      O => nx53675z666
    );
  ix53675z12551 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => rome2addro2_s(0),
      ADR1 => rome2addro2_s(1),
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(3),
      O => nx53675z163
    );
  ix53675z8569 : X_LUT4
    generic map(
      INIT => X"4694"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(2),
      O => nx53675z663
    );
  ix53675z24362 : X_LUT4
    generic map(
      INIT => X"5924"
    )
    port map (
      ADR0 => rome2addro2_s(0),
      ADR1 => rome2addro2_s(1),
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(3),
      O => nx53675z164
    );
  ix53675z12457 : X_LUT4
    generic map(
      INIT => X"4D04"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(3),
      O => nx53675z98
    );
  ix53675z11927 : X_LUT4
    generic map(
      INIT => X"05A0"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1299
    );
  ix53675z52552 : X_LUT4
    generic map(
      INIT => X"F550"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro7_s(2),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1294
    );
  ix53675z58858 : X_LUT4
    generic map(
      INIT => X"E836"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(2),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1302
    );
  ix53675z7203 : X_LUT4
    generic map(
      INIT => X"7656"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(3),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1291
    );
  ix53675z65412 : X_LUT4
    generic map(
      INIT => X"DD44"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro7_s(2),
      O => nx53675z1300
    );
  ix53675z42177 : X_LUT4
    generic map(
      INIT => X"9964"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(2),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1305
    );
  ix53675z6034 : X_LUT4
    generic map(
      INIT => X"02D4"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(3),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1296
    );
  ix53675z23675 : X_LUT4
    generic map(
      INIT => X"1C30"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(3),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1297
    );
  U_DCT1D_ix59700z1523 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_rtlc5n1344(15),
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1345(16),
      O => U_DCT1D_nx59700z168
    );
  U_DCT2D_ix65206z1940 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao4_s(2),
      ADR2 => VCC,
      ADR3 => romo2datao5_s(1),
      O => U_DCT2D_nx65206z451
    );
  U_DCT2D_ix65206z1933 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao5_s(3),
      ADR1 => romo2datao4_s(4),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z445
    );
  U_DCT2D_ix65206z1944 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao4_s(1),
      ADR2 => VCC,
      ADR3 => romo2datao5_s(0),
      O => U_DCT2D_nx65206z454
    );
  U_DCT2D_ix65206z1898 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao4_s(13),
      ADR1 => romo2datao5_s(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z415
    );
  U_DCT2D_ix65206z1909 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao4_s(11),
      ADR2 => romo2datao5_s(10),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z424
    );
  U_DCT2D_ix65206z1902 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2datao4_s(13),
      ADR1 => VCC,
      ADR2 => romo2datao5_s(12),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z418
    );
  ix53675z3769 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(1),
      ADR3 => rome2addro2_s(0),
      O => nx53675z167
    );
  ix53675z34786 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(3),
      O => nx53675z692
    );
  ix53675z5516 : X_LUT4
    generic map(
      INIT => X"50D4"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(3),
      O => nx53675z696
    );
  ix53675z12111 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(1),
      ADR3 => rome2addro2_s(0),
      O => nx53675z169
    );
  ix53675z26111 : X_LUT4
    generic map(
      INIT => X"7310"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(3),
      O => nx53675z693
    );
  ix53675z14016 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(1),
      ADR3 => rome2addro2_s(0),
      O => nx53675z170
    );
  ix53675z18601 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(0),
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(1),
      O => nx53675z175
    );
  ix53675z61344 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(1),
      ADR3 => rome2addro2_s(0),
      O => nx53675z166
    );
  ix53675z34042 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(0),
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(1),
      O => nx53675z172
    );
  ix53675z25034 : X_LUT4
    generic map(
      INIT => X"6518"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(3),
      O => nx53675z634
    );
  ix53675z34693 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(3),
      ADR3 => rome2addro9_s(1),
      O => nx53675z627
    );
  ix53675z5423 : X_LUT4
    generic map(
      INIT => X"3B02"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(3),
      ADR3 => rome2addro9_s(1),
      O => nx53675z631
    );
  ix53675z12778 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(3),
      O => nx53675z636
    );
  ix53675z26018 : X_LUT4
    generic map(
      INIT => X"7150"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(3),
      ADR3 => rome2addro9_s(1),
      O => nx53675z628
    );
  ix53675z9519 : X_LUT4
    generic map(
      INIT => X"3492"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(3),
      O => nx53675z637
    );
  ix53675z19332 : X_LUT4
    generic map(
      INIT => X"24B2"
    )
    port map (
      ADR0 => rome2addro9_s(1),
      ADR1 => rome2addro9_s(3),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(0),
      O => nx53675z642
    );
  ix53675z62011 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(3),
      O => nx53675z633
    );
  ix53675z34709 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro9_s(1),
      ADR1 => rome2addro9_s(3),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(0),
      O => nx53675z639
    );
  ix53675z48101 : X_LUT4
    generic map(
      INIT => X"BF0A"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(3),
      ADR2 => romo2addro0_s(1),
      ADR3 => romo2addro0_s(0),
      O => nx53675z725
    );
  ix53675z54822 : X_LUT4
    generic map(
      INIT => X"F3F2"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(3),
      ADR2 => romo2addro0_s(1),
      ADR3 => romo2addro0_s(0),
      O => nx53675z722
    );
  ix53675z29293 : X_LUT4
    generic map(
      INIT => X"5A50"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => VCC,
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(3),
      O => nx53675z1293
    );
  ix53675z10255 : X_LUT4
    generic map(
      INIT => X"6668"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(2),
      ADR2 => romo2addro0_s(0),
      ADR3 => romo2addro0_s(1),
      O => nx53675z727
    );
  ix53675z40909 : X_LUT4
    generic map(
      INIT => X"D23C"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(2),
      ADR2 => romo2addro0_s(0),
      ADR3 => romo2addro0_s(1),
      O => nx53675z731
    );
  ix53675z58972 : X_LUT4
    generic map(
      INIT => X"99AA"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro0_s(0),
      O => nx53675z736
    );
  ix53675z54630 : X_LUT4
    generic map(
      INIT => X"AB54"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(2),
      ADR2 => romo2addro0_s(0),
      ADR3 => romo2addro0_s(1),
      O => nx53675z728
    );
  ix53675z14663 : X_LUT4
    generic map(
      INIT => X"2244"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro0_s(2),
      O => nx53675z737
    );
  ix53675z42707 : X_LUT4
    generic map(
      INIT => X"C3F2"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(0),
      ADR2 => romo2addro0_s(1),
      ADR3 => romo2addro0_s(2),
      O => nx53675z733
    );
  ix53675z24200 : X_LUT4
    generic map(
      INIT => X"3322"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro0_s(2),
      O => nx53675z734
    );
  ix53675z14619 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => rome2addro9_s(3),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(0),
      O => nx53675z589
    );
  ix53675z4372 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => rome2addro9_s(3),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(0),
      O => nx53675z586
    );
  ix53675z17566 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z584
    );
  ix53675z24074 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2addro8_s(3),
      ADR2 => rome2addro8_s(0),
      ADR3 => VCC,
      O => U2_ROME8_modgen_rom_ix2_nx_rm64_16_l
    );
  ix53675z18849 : X_LUT4
    generic map(
      INIT => X"088E"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(0),
      ADR3 => rome2addro10_s(3),
      O => nx53675z659
    );
  ix53675z19305 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(2),
      O => nx53675z665
    );
  ix54672z23005 : X_LUT4
    generic map(
      INIT => X"5158"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(3),
      O => nx54672z609
    );
  ix54672z51589 : X_LUT4
    generic map(
      INIT => X"C0FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(3),
      O => nx54672z613
    );
  ix54672z10964 : X_LUT4
    generic map(
      INIT => X"0A50"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(3),
      O => nx54672z618
    );
  ix54672z6240 : X_LUT4
    generic map(
      INIT => X"0FDA"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(3),
      O => nx54672z610
    );
  ix54672z64449 : X_LUT4
    generic map(
      INIT => X"AF0A"
    )
    port map (
      ADR0 => romoaddro0_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(3),
      O => nx54672z619
    );
  ix54672z3778 : X_LUT4
    generic map(
      INIT => X"3366"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro0_s(2),
      O => nx54672z660
    );
  ix54672z5071 : X_LUT4
    generic map(
      INIT => X"4524"
    )
    port map (
      ADR0 => romoaddro0_s(2),
      ADR1 => romoaddro0_s(0),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(3),
      O => nx54672z615
    );
  ix54672z22712 : X_LUT4
    generic map(
      INIT => X"224C"
    )
    port map (
      ADR0 => romoaddro0_s(2),
      ADR1 => romoaddro0_s(0),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(3),
      O => nx54672z616
    );
  ix54672z54529 : X_LUT4
    generic map(
      INIT => X"C3F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro0_s(3),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(2),
      O => nx54672z657
    );
  ix54672z13968 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(2),
      ADR3 => romeaddro2_s(1),
      O => nx54672z134
    );
  ix54672z3721 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(2),
      ADR3 => romeaddro2_s(1),
      O => nx54672z131
    );
  ix54672z3634 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(2),
      ADR2 => romeaddro1_s(3),
      ADR3 => romeaddro1_s(0),
      O => nx54672z72
    );
  ix54672z18011 : X_LUT4
    generic map(
      INIT => X"088E"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(2),
      ADR2 => romeaddro1_s(3),
      ADR3 => romeaddro1_s(0),
      O => nx54672z74
    );
  ix54672z13882 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(2),
      ADR2 => romeaddro1_s(3),
      ADR3 => romeaddro1_s(0),
      O => nx54672z75
    );
  ix54672z22958 : X_LUT4
    generic map(
      INIT => X"5700"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z744
    );
  ix54672z60931 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(2),
      ADR2 => romeaddro1_s(3),
      ADR3 => romeaddro1_s(0),
      O => nx54672z71
    );
  ix54672z13918 : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => VCC,
      ADR2 => romeaddro2_s(1),
      ADR3 => VCC,
      O => nx54672z193
    );
  ix54672z22966 : X_LUT4
    generic map(
      INIT => X"02AA"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(1),
      ADR3 => romoaddro2_s(0),
      O => nx54672z750
    );
  ix54672z1749 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romeaddro2_s(0),
      ADR2 => VCC,
      ADR3 => romeaddro2_s(3),
      O => nx54672z190
    );
  ix54672z25542 : X_LUT4
    generic map(
      INIT => X"57A8"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z756
    );
  ix54672z54850 : X_LUT4
    generic map(
      INIT => X"F3F2"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(1),
      ADR3 => romoaddro2_s(0),
      O => nx54672z748
    );
  ix54672z48129 : X_LUT4
    generic map(
      INIT => X"BF0A"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(1),
      ADR3 => romoaddro2_s(0),
      O => nx54672z751
    );
  ix54672z10283 : X_LUT4
    generic map(
      INIT => X"1EE0"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z753
    );
  ix54672z54658 : X_LUT4
    generic map(
      INIT => X"C3C6"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z754
    );
  ix54672z40937 : X_LUT4
    generic map(
      INIT => X"996A"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z757
    );
  ix54672z18097 : X_LUT4
    generic map(
      INIT => X"7110"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(2),
      ADR3 => romeaddro2_s(1),
      O => nx54672z133
    );
  ix54672z17081 : X_LUT4
    generic map(
      INIT => X"5A96"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(3),
      O => nx54672z185
    );
  ix54672z61360 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(3),
      O => nx54672z178
    );
  ix54672z8868 : X_LUT4
    generic map(
      INIT => X"42B4"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(2),
      O => nx54672z182
    );
  ix54672z18681 : X_LUT4
    generic map(
      INIT => X"24B2"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(3),
      O => nx54672z187
    );
  ix54672z24383 : X_LUT4
    generic map(
      INIT => X"2692"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(2),
      O => nx54672z179
    );
  ix54672z27584 : X_LUT4
    generic map(
      INIT => X"39C6"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(3),
      O => nx54672z188
    );
  ix54672z28611 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(3),
      O => nx54672z192
    );
  ix54672z34058 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(3),
      O => nx54672z184
    );
  ix54672z28608 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(3),
      O => U1_ROME2_modgen_rom_ix2_nx_rm64_16_u
    );
  ix54672z2220 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro0_s(0),
      O => nx54672z652
    );
  ix54672z18477 : X_LUT4
    generic map(
      INIT => X"20B2"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z399
    );
  ix54672z17453 : X_LUT4
    generic map(
      INIT => X"6696"
    )
    port map (
      ADR0 => romeaddro6_s(2),
      ADR1 => romeaddro6_s(1),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(3),
      O => nx54672z445
    );
  ix54672z61398 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z396
    );
  ix54672z14348 : X_LUT4
    generic map(
      INIT => X"50D4"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z400
    );
  ix54672z19053 : X_LUT4
    generic map(
      INIT => X"188E"
    )
    port map (
      ADR0 => romeaddro6_s(2),
      ADR1 => romeaddro6_s(1),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(3),
      O => nx54672z447
    );
  ix54672z4101 : X_LUT4
    generic map(
      INIT => X"08CE"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z397
    );
  ix54672z27956 : X_LUT4
    generic map(
      INIT => X"2DD2"
    )
    port map (
      ADR0 => romeaddro6_s(2),
      ADR1 => romeaddro6_s(1),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(3),
      O => nx54672z448
    );
  ix54672z28983 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro6_s(0),
      ADR1 => romeaddro6_s(3),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(1),
      O => nx54672z452
    );
  ix54672z34430 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro6_s(2),
      ADR1 => romeaddro6_s(1),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(3),
      O => nx54672z444
    );
  ix54672z28980 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro6_s(0),
      ADR1 => romeaddro6_s(3),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(1),
      O => U1_ROME6_modgen_rom_ix2_nx_rm64_16_u
    );
  ix53675z54917 : X_LUT4
    generic map(
      INIT => X"BBBA"
    )
    port map (
      ADR0 => romo2addro1_s(1),
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(2),
      ADR3 => romo2addro1_s(0),
      O => nx53675z793
    );
  ix53675z8203 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => rome2addro9_s(1),
      ADR1 => rome2addro9_s(0),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(3),
      O => nx53675z615
    );
  ix53675z25013 : X_LUT4
    generic map(
      INIT => X"3942"
    )
    port map (
      ADR0 => rome2addro9_s(1),
      ADR1 => rome2addro9_s(0),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(3),
      O => nx53675z619
    );
  ix53675z23033 : X_LUT4
    generic map(
      INIT => X"10F0"
    )
    port map (
      ADR0 => romo2addro1_s(1),
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(2),
      ADR3 => romo2addro1_s(0),
      O => nx53675z795
    );
  ix53675z27078 : X_LUT4
    generic map(
      INIT => X"6158"
    )
    port map (
      ADR0 => rome2addro9_s(1),
      ADR1 => rome2addro9_s(0),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(3),
      O => nx53675z616
    );
  ix53675z48196 : X_LUT4
    generic map(
      INIT => X"F750"
    )
    port map (
      ADR0 => romo2addro1_s(1),
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(2),
      ADR3 => romo2addro1_s(0),
      O => nx53675z796
    );
  ix53675z25514 : X_LUT4
    generic map(
      INIT => X"3C6C"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(2),
      ADR2 => romo2addro0_s(0),
      ADR3 => romo2addro0_s(1),
      O => nx53675z730
    );
  ix53675z22938 : X_LUT4
    generic map(
      INIT => X"02AA"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(3),
      ADR2 => romo2addro0_s(1),
      ADR3 => romo2addro0_s(0),
      O => nx53675z724
    );
  ix53675z26090 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(2),
      O => nx53675z678
    );
  ix53675z4513 : X_LUT4
    generic map(
      INIT => X"08AE"
    )
    port map (
      ADR0 => rome2addro10_s(0),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(2),
      ADR3 => rome2addro10_s(3),
      O => nx53675z687
    );
  ix53675z13295 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => rome2addro10_s(0),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(2),
      ADR3 => rome2addro10_s(3),
      O => nx53675z683
    );
  ix53675z31251 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(2),
      O => nx53675z675
    );
  ix53675z8296 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => rome2addro10_s(0),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(2),
      ADR3 => rome2addro10_s(3),
      O => nx53675z680
    );
  ix53675z25106 : X_LUT4
    generic map(
      INIT => X"5924"
    )
    port map (
      ADR0 => rome2addro10_s(0),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(2),
      ADR3 => rome2addro10_s(3),
      O => nx53675z684
    );
  ix53675z12855 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => rome2addro10_s(0),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(2),
      ADR3 => rome2addro10_s(3),
      O => nx53675z689
    );
  ix53675z27171 : X_LUT4
    generic map(
      INIT => X"6138"
    )
    port map (
      ADR0 => rome2addro10_s(0),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(2),
      ADR3 => rome2addro10_s(3),
      O => nx53675z681
    );
  ix53675z14760 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => rome2addro10_s(0),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(2),
      ADR3 => rome2addro10_s(3),
      O => nx53675z690
    );
  ix53675z19345 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(3),
      O => nx53675z695
    );
  ix53675z62088 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro10_s(0),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(2),
      ADR3 => rome2addro10_s(3),
      O => nx53675z686
    );
  ix53675z16915 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2addro1_s(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2addro1_s(2),
      O => nx53675z129
    );
  ix53675z23422 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(3),
      O => U2_ROME1_modgen_rom_ix2_nx_rm64_16_l
    );
  ix53675z3547 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => rome2addro0_s(3),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(0),
      O => nx53675z8
    );
  ix53675z17923 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => rome2addro0_s(3),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(0),
      O => nx53675z10
    );
  ix53675z13794 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => rome2addro0_s(3),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(0),
      O => nx53675z11
    );
  ix53675z18379 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(2),
      ADR3 => rome2addro0_s(1),
      O => nx53675z16
    );
  ix53675z60844 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => rome2addro0_s(3),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(0),
      O => nx53675z7
    );
  ix53675z7068 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(2),
      ADR3 => rome2addro0_s(1),
      O => nx53675z13
    );
  ix53675z21991 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(2),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(0),
      O => nx53675z669
    );
  ix53675z43597 : X_LUT4
    generic map(
      INIT => X"CF32"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(0),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(1),
      O => nx53675z1363
    );
  ix53675z15553 : X_LUT4
    generic map(
      INIT => X"2424"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(3),
      ADR3 => VCC,
      O => nx53675z1367
    );
  ix53675z12831 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(2),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(0),
      O => nx53675z671
    );
  ix53675z25090 : X_LUT4
    generic map(
      INIT => X"00FA"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1364
    );
  ix53675z4492 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(2),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(0),
      O => nx53675z672
    );
  ix53675z19321 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(2),
      O => nx53675z677
    );
  ix53675z35312 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(2),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(0),
      O => nx53675z668
    );
  ix53675z40778 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(2),
      O => nx53675z674
    );
  ix53675z4000 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => rome2addro5_s(2),
      ADR1 => rome2addro5_s(0),
      ADR2 => rome2addro5_s(3),
      ADR3 => rome2addro5_s(1),
      O => nx53675z326
    );
  ix53675z18376 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => rome2addro5_s(2),
      ADR1 => rome2addro5_s(0),
      ADR2 => rome2addro5_s(3),
      ADR3 => rome2addro5_s(1),
      O => nx53675z328
    );
  ix53675z14247 : X_LUT4
    generic map(
      INIT => X"08AE"
    )
    port map (
      ADR0 => rome2addro5_s(2),
      ADR1 => rome2addro5_s(0),
      ADR2 => rome2addro5_s(3),
      ADR3 => rome2addro5_s(1),
      O => nx53675z329
    );
  ix53675z3729 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(1),
      ADR3 => rome2addro2_s(0),
      O => nx53675z137
    );
  ix53675z18105 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(1),
      ADR3 => rome2addro2_s(0),
      O => nx53675z139
    );
  ix53675z13976 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(1),
      ADR3 => rome2addro2_s(0),
      O => nx53675z140
    );
  ix53675z7250 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(1),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(2),
      O => nx53675z142
    );
  ix53675z18561 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(1),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(2),
      O => nx53675z145
    );
  ix53675z61026 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(1),
      ADR3 => rome2addro2_s(0),
      O => nx53675z136
    );
  ix53675z4772 : X_LUT4
    generic map(
      INIT => X"4F04"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(0),
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(1),
      O => nx53675z176
    );
  ix53675z17081 : X_LUT4
    generic map(
      INIT => X"4BB4"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(0),
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(1),
      O => nx53675z185
    );
  ix53675z12127 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(1),
      ADR3 => rome2addro2_s(0),
      O => nx53675z181
    );
  ix53675z25367 : X_LUT4
    generic map(
      INIT => X"2B22"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(0),
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(1),
      O => nx53675z173
    );
  ix53675z61360 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(1),
      ADR3 => rome2addro2_s(0),
      O => nx53675z178
    );
  ix53675z8868 : X_LUT4
    generic map(
      INIT => X"6138"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(1),
      ADR3 => rome2addro2_s(0),
      O => nx53675z182
    );
  ix53675z28608 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro2_s(1),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(3),
      O => U2_ROME2_modgen_rom_ix2_nx_rm64_16_u
    );
  ix53675z18681 : X_LUT4
    generic map(
      INIT => X"7118"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(0),
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(1),
      O => nx53675z187
    );
  ix53675z24383 : X_LUT4
    generic map(
      INIT => X"249A"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(1),
      ADR3 => rome2addro2_s(0),
      O => nx53675z179
    );
  ix53675z27584 : X_LUT4
    generic map(
      INIT => X"6696"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(0),
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(1),
      O => nx53675z188
    );
  ix53675z34058 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(0),
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(1),
      O => nx53675z184
    );
  ix53675z28611 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro2_s(1),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(3),
      O => nx53675z192
    );
  ix53675z13873 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(1),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(3),
      O => nx53675z69
    );
  ix53675z3626 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(1),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(3),
      O => nx53675z66
    );
  ix53675z7731 : X_LUT4
    generic map(
      INIT => X"42B4"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(1),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(3),
      O => nx53675z78
    );
  ix53675z18467 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(1),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(3),
      O => nx53675z80
    );
  ix53675z18587 : X_LUT4
    generic map(
      INIT => X"2B42"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(3),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(1),
      O => nx53675z122
    );
  ix53675z14882 : X_LUT4
    generic map(
      INIT => X"2692"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(1),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(3),
      O => nx53675z81
    );
  ix53675z11993 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z86
    );
  ix53675z7156 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(1),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(3),
      O => nx53675z77
    );
  ix53675z34474 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z83
    );
  ix53675z3654 : X_LUT4
    generic map(
      INIT => X"44D4"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z87
    );
  ix53675z3721 : X_LUT4
    generic map(
      INIT => X"20F2"
    )
    port map (
      ADR0 => rome2addro2_s(1),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(3),
      O => nx53675z131
    );
  ix53675z13918 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => rome2addro2_s(1),
      ADR1 => rome2addro2_s(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z193
    );
  ix53675z18097 : X_LUT4
    generic map(
      INIT => X"088E"
    )
    port map (
      ADR0 => rome2addro2_s(1),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(3),
      O => nx53675z133
    );
  ix53675z1749 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rome2addro2_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2addro2_s(3),
      O => nx53675z190
    );
  ix53675z13968 : X_LUT4
    generic map(
      INIT => X"44D4"
    )
    port map (
      ADR0 => rome2addro2_s(1),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(3),
      O => nx53675z134
    );
  ix53675z18011 : X_LUT4
    generic map(
      INIT => X"7110"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z74
    );
  ix53675z60931 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z71
    );
  ix53675z21153 : X_LUT4
    generic map(
      INIT => X"20F2"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z84
    );
  ix53675z33964 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(3),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(1),
      O => nx53675z119
    );
  ix53675z27490 : X_LUT4
    generic map(
      INIT => X"3C96"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(3),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(1),
      O => nx53675z123
    );
  ix53675z28517 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(1),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(3),
      O => nx53675z127
    );
  ix53675z16987 : X_LUT4
    generic map(
      INIT => X"659A"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(3),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(1),
      O => nx53675z120
    );
  ix53675z13824 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2addro1_s(1),
      ADR2 => VCC,
      ADR3 => rome2addro1_s(2),
      O => nx53675z128
    );
  ix53675z28514 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(1),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(3),
      O => U2_ROME1_modgen_rom_ix2_nx_rm64_16_u
    );
  ix53675z1655 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2addro1_s(0),
      ADR2 => VCC,
      ADR3 => rome2addro1_s(3),
      O => nx53675z125
    );
  ix53675z4865 : X_LUT4
    generic map(
      INIT => X"7130"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z241
    );
  ix53675z18774 : X_LUT4
    generic map(
      INIT => X"42D4"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z252
    );
  ix53675z25460 : X_LUT4
    generic map(
      INIT => X"20BA"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z238
    );
  ix53675z34151 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z249
    );
  ix53675z27677 : X_LUT4
    generic map(
      INIT => X"59A6"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z253
    );
  ix53675z17174 : X_LUT4
    generic map(
      INIT => X"693C"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z250
    );
  ix53675z17101 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rome2addro3_s(2),
      ADR3 => rome2addro3_s(1),
      O => nx53675z259
    );
  ix53675z13882 : X_LUT4
    generic map(
      INIT => X"4F04"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z75
    );
  ix53675z23934 : X_LUT4
    generic map(
      INIT => X"1F00"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1427
    );
  ix53675z3634 : X_LUT4
    generic map(
      INIT => X"44D4"
    )
    port map (
      ADR0 => rome2addro1_s(3),
      ADR1 => rome2addro1_s(0),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z72
    );
  ix53675z55818 : X_LUT4
    generic map(
      INIT => X"BBBA"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1425
    );
  ix53675z49097 : X_LUT4
    generic map(
      INIT => X"F570"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1428
    );
  ix53675z18841 : X_LUT4
    generic map(
      INIT => X"20B2"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(3),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(0),
      O => nx53675z653
    );
  ix53675z4465 : X_LUT4
    generic map(
      INIT => X"7310"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(3),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(0),
      O => nx53675z651
    );
  ix53675z14712 : X_LUT4
    generic map(
      INIT => X"2B0A"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(3),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(0),
      O => nx53675z654
    );
  ix53675z55940 : X_LUT4
    generic map(
      INIT => X"AFAE"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1510
    );
  ix53675z23264 : X_LUT4
    generic map(
      INIT => X"444C"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(1),
      ADR3 => romo2addro3_s(3),
      O => nx53675z959
    );
  ix53675z49219 : X_LUT4
    generic map(
      INIT => X"DF44"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1513
    );
  ix53675z60013 : X_LUT4
    generic map(
      INIT => X"C800"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(1),
      ADR3 => romo2addro3_s(3),
      O => nx53675z956
    );
  ix53675z48427 : X_LUT4
    generic map(
      INIT => X"8EAE"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(1),
      ADR3 => romo2addro3_s(3),
      O => nx53675z960
    );
  ix53675z3002 : X_LUT4
    generic map(
      INIT => X"00FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro3_s(0),
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(3),
      O => nx53675z1019
    );
  ix53675z55148 : X_LUT4
    generic map(
      INIT => X"F0FE"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(1),
      ADR3 => romo2addro3_s(3),
      O => nx53675z957
    );
  ix53675z2797 : X_LUT4
    generic map(
      INIT => X"0050"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => VCC,
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(3),
      O => nx53675z1016
    );
  ix53675z2495 : X_LUT4
    generic map(
      INIT => X"FEFE"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => romo2addro3_s(0),
      ADR2 => romo2addro3_s(2),
      ADR3 => VCC,
      O => nx53675z1020
    );
  ix53675z14794 : X_LUT4
    generic map(
      INIT => X"24D2"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(2),
      ADR3 => rome2addro0_s(1),
      O => nx53675z17
    );
  ix53675z4420 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => rome2addro9_s(3),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(0),
      O => nx53675z622
    );
  ix53675z28429 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(3),
      O => nx53675z63
    );
  ix53675z7643 : X_LUT4
    generic map(
      INIT => X"2962"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(3),
      ADR2 => rome2addro0_s(2),
      ADR3 => rome2addro0_s(1),
      O => nx53675z14
    );
  ix53675z28426 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(1),
      ADR3 => rome2addro0_s(3),
      O => U2_ROME0_modgen_rom_ix2_nx_rm64_16_u
    );
  ix53675z13736 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => rome2addro0_s(1),
      ADR1 => rome2addro0_s(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z64
    );
  ix53675z12762 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => rome2addro9_s(3),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(0),
      O => nx53675z624
    );
  ix53675z1567 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rome2addro0_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2addro0_s(3),
      O => nx53675z61
    );
  ix53675z14667 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => rome2addro9_s(3),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(0),
      O => nx53675z625
    );
  ix53675z19252 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(3),
      ADR3 => rome2addro9_s(1),
      O => nx53675z630
    );
  ix53675z61995 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro9_s(3),
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => rome2addro9_s(0),
      O => nx53675z621
    );
  ix53675z28235 : X_LUT4
    generic map(
      INIT => X"639C"
    )
    port map (
      ADR0 => rome2addro9_s(1),
      ADR1 => rome2addro9_s(3),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(0),
      O => nx53675z643
    );
  ix53675z3539 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => rome2addro0_s(1),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(3),
      ADR3 => rome2addro0_s(0),
      O => nx53675z2
    );
  ix53675z29262 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(1),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(3),
      O => nx53675z647
    );
  ix53675z17732 : X_LUT4
    generic map(
      INIT => X"695A"
    )
    port map (
      ADR0 => rome2addro9_s(1),
      ADR1 => rome2addro9_s(3),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(0),
      O => nx53675z640
    );
  ix53675z29259 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => rome2addro9_s(1),
      ADR2 => rome2addro9_s(2),
      ADR3 => rome2addro9_s(3),
      O => U2_ROME9_modgen_rom_ix2_nx_rm64_16_u
    );
  ix53675z14569 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2addro9_s(1),
      ADR2 => rome2addro9_s(2),
      ADR3 => VCC,
      O => nx53675z648
    );
  ix53675z17915 : X_LUT4
    generic map(
      INIT => X"088E"
    )
    port map (
      ADR0 => rome2addro0_s(1),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(3),
      ADR3 => rome2addro0_s(0),
      O => nx53675z4
    );
  ix53675z2400 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rome2addro9_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2addro9_s(3),
      O => nx53675z645
    );
  ix53675z13786 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => rome2addro0_s(1),
      ADR1 => rome2addro0_s(2),
      ADR2 => rome2addro0_s(3),
      ADR3 => rome2addro0_s(0),
      O => nx53675z5
    );
  ix53675z23144 : X_LUT4
    generic map(
      INIT => X"1F00"
    )
    port map (
      ADR0 => romo2addro2_s(3),
      ADR1 => romo2addro2_s(1),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(2),
      O => nx53675z874
    );
  ix53675z55028 : X_LUT4
    generic map(
      INIT => X"DDDC"
    )
    port map (
      ADR0 => romo2addro2_s(3),
      ADR1 => romo2addro2_s(1),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(2),
      O => nx53675z872
    );
  ix53675z48307 : X_LUT4
    generic map(
      INIT => X"F370"
    )
    port map (
      ADR0 => romo2addro2_s(3),
      ADR1 => romo2addro2_s(1),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(2),
      O => nx53675z875
    );
  ix53675z59790 : X_LUT4
    generic map(
      INIT => X"C080"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(2),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(1),
      O => nx53675z798
    );
  ix53675z2891 : X_LUT4
    generic map(
      INIT => X"0F0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(2),
      O => nx53675z940
    );
  ix53675z2384 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romo2addro2_s(1),
      ADR1 => romo2addro2_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(2),
      O => nx53675z941
    );
  ix53675z2686 : X_LUT4
    generic map(
      INIT => X"000A"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z937
    );
  ix53675z2621 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z938
    );
  ix53675z23041 : X_LUT4
    generic map(
      INIT => X"444C"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(2),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(1),
      O => nx53675z801
    );
  ix53675z54733 : X_LUT4
    generic map(
      INIT => X"F10E"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(2),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(1),
      O => nx53675z805
    );
  ix53675z48204 : X_LUT4
    generic map(
      INIT => X"8AEE"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(2),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(1),
      O => nx53675z802
    );
  ix53675z25617 : X_LUT4
    generic map(
      INIT => X"666C"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(2),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(1),
      O => nx53675z807
    );
  ix53675z54925 : X_LUT4
    generic map(
      INIT => X"FF0E"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(2),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(1),
      O => nx53675z799
    );
  ix53675z41012 : X_LUT4
    generic map(
      INIT => X"9A66"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(2),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(1),
      O => nx53675z808
    );
  ix53675z59075 : X_LUT4
    generic map(
      INIT => X"C6C6"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(1),
      ADR3 => VCC,
      O => nx53675z813
    );
  ix53675z10358 : X_LUT4
    generic map(
      INIT => X"3C68"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(2),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(1),
      O => nx53675z804
    );
  ix53675z42810 : X_LUT4
    generic map(
      INIT => X"F05E"
    )
    port map (
      ADR0 => romo2addro1_s(2),
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(1),
      ADR3 => romo2addro1_s(0),
      O => nx53675z810
    );
  ix53675z14766 : X_LUT4
    generic map(
      INIT => X"1818"
    )
    port map (
      ADR0 => romo2addro1_s(2),
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(1),
      ADR3 => VCC,
      O => nx53675z814
    );
  ix53675z55452 : X_LUT4
    generic map(
      INIT => X"CC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro7_s(3),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1327
    );
  ix53675z3454 : X_LUT4
    generic map(
      INIT => X"00FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro7_s(2),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(3),
      O => nx53675z1335
    );
  ix53675z2947 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro7_s(2),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1336
    );
  ix53675z3249 : X_LUT4
    generic map(
      INIT => X"0044"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(2),
      ADR2 => VCC,
      ADR3 => romo2addro7_s(3),
      O => nx53675z1332
    );
  ix53675z3184 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro7_s(3),
      O => nx53675z1333
    );
  ix53675z4743 : X_LUT4
    generic map(
      INIT => X"5656"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(2),
      ADR3 => VCC,
      O => nx53675z1341
    );
  ix53675z10924 : X_LUT4
    generic map(
      INIT => X"1E1E"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(2),
      ADR3 => VCC,
      O => nx53675z1342
    );
  ix53675z57391 : X_LUT4
    generic map(
      INIT => X"AF50"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro7_s(2),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1338
    );
  ix53675z25073 : X_LUT4
    generic map(
      INIT => X"0F5A"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1339
    );
  ix53675z64635 : X_LUT4
    generic map(
      INIT => X"AF0A"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro0_s(1),
      ADR3 => romo2addro0_s(2),
      O => nx53675z749
    );
  ix53675z41400 : X_LUT4
    generic map(
      INIT => X"A54A"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(2),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(1),
      O => nx53675z754
    );
  ix53675z22898 : X_LUT4
    generic map(
      INIT => X"4622"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(3),
      ADR2 => romo2addro0_s(1),
      ADR3 => romo2addro0_s(2),
      O => nx53675z746
    );
  ix53675z44730 : X_LUT4
    generic map(
      INIT => X"969A"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(2),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(1),
      O => nx53675z752
    );
  ix53675z52367 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(1),
      O => nx53675z755
    );
  ix53675z43770 : X_LUT4
    generic map(
      INIT => X"AA10"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(1),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(0),
      O => nx53675z760
    );
  ix53675z58081 : X_LUT4
    generic map(
      INIT => X"E856"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(2),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(1),
      O => nx53675z751
    );
  ix53675z22619 : X_LUT4
    generic map(
      INIT => X"50D4"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(1),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(0),
      O => nx53675z757
    );
  ix53675z38280 : X_LUT4
    generic map(
      INIT => X"C242"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(1),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(0),
      O => nx53675z758
    );
  ix53675z61923 : X_LUT4
    generic map(
      INIT => X"EC80"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(1),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(0),
      O => nx53675z761
    );
  ix53675z21180 : X_LUT4
    generic map(
      INIT => X"459A"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(1),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(0),
      O => nx53675z766
    );
  ix53675z28760 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro1_s(1),
      ADR3 => VCC,
      O => nx53675z870
    );
  ix53675z15803 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro1_s(1),
      ADR3 => VCC,
      O => U2_ROMO1_modgen_rom_ix0_nx_rm64_16_l
    );
  ix53675z28516 : X_LUT4
    generic map(
      INIT => X"22CC"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro0_s(1),
      O => nx53675z742
    );
  ix53675z51775 : X_LUT4
    generic map(
      INIT => X"F550"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro0_s(2),
      ADR3 => romo2addro0_s(1),
      O => nx53675z743
    );
  ix53675z11150 : X_LUT4
    generic map(
      INIT => X"0A50"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro0_s(1),
      ADR3 => romo2addro0_s(0),
      O => nx53675z748
    );
  ix53675z23191 : X_LUT4
    generic map(
      INIT => X"3432"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(0),
      ADR2 => romo2addro0_s(2),
      ADR3 => romo2addro0_s(1),
      O => nx53675z739
    );
  ix53675z6426 : X_LUT4
    generic map(
      INIT => X"5E1E"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(0),
      ADR2 => romo2addro0_s(2),
      ADR3 => romo2addro0_s(1),
      O => nx53675z740
    );
  ix53675z5257 : X_LUT4
    generic map(
      INIT => X"108E"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(3),
      ADR2 => romo2addro0_s(1),
      ADR3 => romo2addro0_s(2),
      O => nx53675z745
    );
  ix53675z3822 : X_LUT4
    generic map(
      INIT => X"08AE"
    )
    port map (
      ADR0 => rome2addro3_s(0),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(2),
      ADR3 => rome2addro3_s(3),
      O => nx53675z202
    );
  ix53675z19475 : X_LUT4
    generic map(
      INIT => X"1A86"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(1),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(0),
      O => nx53675z763
    );
  ix53675z36809 : X_LUT4
    generic map(
      INIT => X"934C"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(1),
      ADR2 => romo2addro0_s(2),
      ADR3 => romo2addro0_s(0),
      O => nx53675z767
    );
  ix53675z18198 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => rome2addro3_s(0),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(2),
      ADR3 => rome2addro3_s(3),
      O => nx53675z204
    );
  ix53675z27932 : X_LUT4
    generic map(
      INIT => X"3E96"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(1),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(0),
      O => nx53675z764
    );
  ix53675z18694 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z240
    );
  ix53675z14069 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => rome2addro3_s(0),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(2),
      ADR3 => rome2addro3_s(3),
      O => nx53675z205
    );
  ix53675z34135 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z237
    );
  ix53675z24303 : X_LUT4
    generic map(
      INIT => X"5454"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(2),
      ADR3 => VCC,
      O => nx53675z811
    );
  ix53675z28619 : X_LUT4
    generic map(
      INIT => X"3C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro1_s(0),
      ADR2 => romo2addro1_s(1),
      ADR3 => romo2addro1_s(3),
      O => nx53675z819
    );
  ix53675z23294 : X_LUT4
    generic map(
      INIT => X"02DC"
    )
    port map (
      ADR0 => romo2addro1_s(1),
      ADR1 => romo2addro1_s(2),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(0),
      O => nx53675z816
    );
  ix53675z51878 : X_LUT4
    generic map(
      INIT => X"C0FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro1_s(2),
      ADR2 => romo2addro1_s(1),
      ADR3 => romo2addro1_s(3),
      O => nx53675z820
    );
  ix53675z6622 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro1_s(2),
      ADR3 => VCC,
      O => U2_ROMO1_modgen_rom_ix0_nx_rm64_16_u
    );
  ix53675z11253 : X_LUT4
    generic map(
      INIT => X"03C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(0),
      ADR3 => romo2addro1_s(1),
      O => nx53675z825
    );
  ix53675z6529 : X_LUT4
    generic map(
      INIT => X"3B3C"
    )
    port map (
      ADR0 => romo2addro1_s(1),
      ADR1 => romo2addro1_s(2),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(0),
      O => nx53675z817
    );
  ix53675z64738 : X_LUT4
    generic map(
      INIT => X"C0FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(2),
      ADR3 => romo2addro1_s(1),
      O => nx53675z826
    );
  ix53675z5360 : X_LUT4
    generic map(
      INIT => X"2432"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => romo2addro1_s(2),
      ADR2 => romo2addro1_s(0),
      ADR3 => romo2addro1_s(1),
      O => nx53675z822
    );
  ix53675z23001 : X_LUT4
    generic map(
      INIT => X"1C30"
    )
    port map (
      ADR0 => romo2addro1_s(1),
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(0),
      ADR3 => romo2addro1_s(2),
      O => nx53675z823
    );
  ix53675z25675 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro1_s(2),
      ADR3 => VCC,
      O => nx53675z869
    );
  ix53675z15668 : X_LUT4
    generic map(
      INIT => X"0A50"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro9_s(1),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1446
    );
  ix53675z29521 : X_LUT4
    generic map(
      INIT => X"44AA"
    )
    port map (
      ADR0 => romo2addro9_s(0),
      ADR1 => romo2addro9_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro9_s(1),
      O => nx53675z1451
    );
  ix53675z25205 : X_LUT4
    generic map(
      INIT => X"3322"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => romo2addro9_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro9_s(2),
      O => nx53675z1443
    );
  ix53675z52780 : X_LUT4
    generic map(
      INIT => X"BB22"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro9_s(2),
      O => nx53675z1452
    );
  ix53675z12155 : X_LUT4
    generic map(
      INIT => X"1188"
    )
    port map (
      ADR0 => romo2addro9_s(0),
      ADR1 => romo2addro9_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro9_s(1),
      O => nx53675z1457
    );
  ix53675z24196 : X_LUT4
    generic map(
      INIT => X"0F24"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1448
    );
  ix53675z7431 : X_LUT4
    generic map(
      INIT => X"23FC"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1449
    );
  ix53675z6262 : X_LUT4
    generic map(
      INIT => X"02D4"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1454
    );
  ix53675z14976 : X_LUT4
    generic map(
      INIT => X"6318"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(1),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(2),
      O => nx53675z146
    );
  ix53675z12087 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro2_s(1),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(3),
      O => nx53675z151
    );
  ix53675z7825 : X_LUT4
    generic map(
      INIT => X"5294"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(1),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(2),
      O => nx53675z143
    );
  ix53675z21247 : X_LUT4
    generic map(
      INIT => X"2B22"
    )
    port map (
      ADR0 => rome2addro2_s(1),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(3),
      O => nx53675z149
    );
  ix53675z3748 : X_LUT4
    generic map(
      INIT => X"20F2"
    )
    port map (
      ADR0 => rome2addro2_s(1),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(3),
      O => nx53675z152
    );
  ix53675z18577 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(1),
      O => nx53675z157
    );
  ix53675z34568 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => rome2addro2_s(1),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(3),
      O => nx53675z148
    );
  ix53675z40034 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(1),
      O => nx53675z154
    );
  ix53675z30507 : X_LUT4
    generic map(
      INIT => X"08CE"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(1),
      O => nx53675z155
    );
  ix53675z25346 : X_LUT4
    generic map(
      INIT => X"2B0A"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => rome2addro2_s(2),
      ADR2 => rome2addro2_s(0),
      ADR3 => rome2addro2_s(1),
      O => nx53675z158
    );
  ix53675z45620 : X_LUT4
    generic map(
      INIT => X"B54A"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1382
    );
  ix53675z53257 : X_LUT4
    generic map(
      INIT => X"9696"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => VCC,
      O => nx53675z1385
    );
  ix53675z28822 : X_LUT4
    generic map(
      INIT => X"5E96"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(2),
      ADR2 => romo2addro8_s(1),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1394
    );
  ix53675z44660 : X_LUT4
    generic map(
      INIT => X"F002"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1390
    );
  ix53675z23509 : X_LUT4
    generic map(
      INIT => X"0A8E"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1387
    );
  ix53675z62813 : X_LUT4
    generic map(
      INIT => X"EC80"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1391
    );
  ix53675z20253 : X_LUT4
    generic map(
      INIT => X"6518"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(1),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1314
    );
  ix53675z22070 : X_LUT4
    generic map(
      INIT => X"31C6"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(2),
      ADR2 => romo2addro8_s(1),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1396
    );
  ix53675z39170 : X_LUT4
    generic map(
      INIT => X"9818"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1388
    );
  ix53675z37699 : X_LUT4
    generic map(
      INIT => X"8770"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(2),
      ADR2 => romo2addro8_s(1),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1397
    );
  ix53675z20365 : X_LUT4
    generic map(
      INIT => X"4694"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(2),
      ADR2 => romo2addro8_s(1),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1393
    );
  ix53675z21958 : X_LUT4
    generic map(
      INIT => X"31C6"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(1),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1317
    );
  ix53675z26346 : X_LUT4
    generic map(
      INIT => X"666A"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(3),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1321
    );
  ix53675z37587 : X_LUT4
    generic map(
      INIT => X"943C"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(1),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1318
    );
  ix53675z41024 : X_LUT4
    generic map(
      INIT => X"8F70"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(3),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1323
    );
  ix53675z28710 : X_LUT4
    generic map(
      INIT => X"6D5A"
    )
    port map (
      ADR0 => romo2addro7_s(3),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(1),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1315
    );
  ix53675z11349 : X_LUT4
    generic map(
      INIT => X"5A78"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(3),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1324
    );
  ix53675z26396 : X_LUT4
    generic map(
      INIT => X"3CC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro7_s(2),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(3),
      O => nx53675z1329
    );
  ix53675z30167 : X_LUT4
    generic map(
      INIT => X"639C"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(3),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1320
    );
  ix53675z7225 : X_LUT4
    generic map(
      INIT => X"3388"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(2),
      ADR2 => VCC,
      ADR3 => romo2addro7_s(3),
      O => nx53675z1326
    );
  ix53675z42261 : X_LUT4
    generic map(
      INIT => X"F00C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro7_s(2),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1330
    );
  U_DCT1D_reg_latchbuf_reg_1_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_5_DXMUX,
      CE => U_DCT1D_latchbuf_reg_1_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_1_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_1_5_FFX_RST,
      O => U_DCT1D_latchbuf_reg_1_Q(5)
    );
  U_DCT1D_latchbuf_reg_1_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_1_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_1_5_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_1_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_7_DYMUX,
      CE => U_DCT1D_latchbuf_reg_1_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_1_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_1_7_FFY_RST,
      O => U_DCT1D_latchbuf_reg_1_Q(6)
    );
  U_DCT1D_latchbuf_reg_1_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_1_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_1_7_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_1_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_7_DXMUX,
      CE => U_DCT1D_latchbuf_reg_1_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_1_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_1_7_FFX_RST,
      O => U_DCT1D_latchbuf_reg_1_Q(7)
    );
  U_DCT1D_latchbuf_reg_1_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_1_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_1_7_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_2_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_1_DYMUX,
      CE => U_DCT1D_latchbuf_reg_2_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_2_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_2_1_FFY_RST,
      O => U_DCT1D_latchbuf_reg_2_Q(0)
    );
  U_DCT1D_latchbuf_reg_2_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_2_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_2_1_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_2_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_1_DXMUX,
      CE => U_DCT1D_latchbuf_reg_2_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_2_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_2_1_FFX_RST,
      O => U_DCT1D_latchbuf_reg_2_Q(1)
    );
  U_DCT1D_latchbuf_reg_2_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_2_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_2_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_2_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_3_DYMUX,
      CE => U_DCT1D_latchbuf_reg_2_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_2_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_2_3_FFY_RST,
      O => U_DCT1D_latchbuf_reg_2_Q(2)
    );
  U_DCT1D_latchbuf_reg_2_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_2_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_2_3_FFY_RST
    );
  ix53675z43260 : X_LUT4
    generic map(
      INIT => X"B5B4"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => romo2addro5_s(2),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1126
    );
  ix53675z15216 : X_LUT4
    generic map(
      INIT => X"0A50"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1130
    );
  ix53675z29069 : X_LUT4
    generic map(
      INIT => X"5A0A"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1135
    );
  ix53675z24753 : X_LUT4
    generic map(
      INIT => X"0F0A"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro5_s(0),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1127
    );
  ix53675z52328 : X_LUT4
    generic map(
      INIT => X"A0FA"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1136
    );
  ix53675z11703 : X_LUT4
    generic map(
      INIT => X"0A50"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(0),
      O => nx53675z1141
    );
  ix53675z23744 : X_LUT4
    generic map(
      INIT => X"0B4A"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(0),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1132
    );
  ix53675z6979 : X_LUT4
    generic map(
      INIT => X"55DA"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(0),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1133
    );
  ix53675z5810 : X_LUT4
    generic map(
      INIT => X"108E"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => romo2addro5_s(0),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1138
    );
  ix53675z12406 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => rome2addro5_s(1),
      ADR1 => rome2addro5_s(3),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z376
    );
  ix53675z18960 : X_LUT4
    generic map(
      INIT => X"42D4"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(1),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z382
    );
  ix53675z24662 : X_LUT4
    generic map(
      INIT => X"18C6"
    )
    port map (
      ADR0 => rome2addro5_s(1),
      ADR1 => rome2addro5_s(3),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z374
    );
  ix53675z9147 : X_LUT4
    generic map(
      INIT => X"294A"
    )
    port map (
      ADR0 => rome2addro5_s(1),
      ADR1 => rome2addro5_s(3),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z377
    );
  ix53675z17360 : X_LUT4
    generic map(
      INIT => X"693C"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(1),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z380
    );
  ix53675z27863 : X_LUT4
    generic map(
      INIT => X"659A"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(1),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z383
    );
  ix53675z26351 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1343
    );
  ix53675z34337 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(1),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z379
    );
  ix53675z7298 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romo2addro7_s(3),
      O => U2_ROMO7_modgen_rom_ix0_nx_rm64_16_u
    );
  ix53675z24081 : X_LUT4
    generic map(
      INIT => X"04BA"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(3),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1369
    );
  ix53675z52665 : X_LUT4
    generic map(
      INIT => X"88EE"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro8_s(3),
      O => nx53675z1373
    );
  ix53675z12040 : X_LUT4
    generic map(
      INIT => X"0A50"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro8_s(1),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1378
    );
  ix53675z7316 : X_LUT4
    generic map(
      INIT => X"5D5A"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(3),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1370
    );
  ix53675z65525 : X_LUT4
    generic map(
      INIT => X"A0FA"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(1),
      O => nx53675z1379
    );
  ix53675z42290 : X_LUT4
    generic map(
      INIT => X"9964"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1384
    );
  ix53675z6147 : X_LUT4
    generic map(
      INIT => X"2342"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(2),
      ADR2 => romo2addro8_s(1),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1375
    );
  ix53675z23788 : X_LUT4
    generic map(
      INIT => X"1588"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(2),
      ADR2 => romo2addro8_s(1),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1376
    );
  ix53675z58971 : X_LUT4
    generic map(
      INIT => X"C9B2"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1381
    );
  ix53675z23609 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2addro3_s(0),
      ADR2 => VCC,
      ADR3 => rome2addro3_s(3),
      O => U2_ROME3_modgen_rom_ix2_nx_rm64_16_l
    );
  ix53675z25944 : X_LUT4
    generic map(
      INIT => X"3CC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(3),
      O => nx53675z1013
    );
  ix53675z3814 : X_LUT4
    generic map(
      INIT => X"08AE"
    )
    port map (
      ADR0 => rome2addro3_s(0),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(2),
      ADR3 => rome2addro3_s(3),
      O => nx53675z196
    );
  ix53675z41809 : X_LUT4
    generic map(
      INIT => X"AA44"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => romo2addro3_s(2),
      ADR2 => VCC,
      ADR3 => romo2addro3_s(0),
      O => nx53675z1014
    );
  ix53675z55000 : X_LUT4
    generic map(
      INIT => X"AA50"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => VCC,
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(3),
      O => nx53675z1011
    );
  ix53675z18190 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => rome2addro3_s(0),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(2),
      ADR3 => rome2addro3_s(3),
      O => nx53675z198
    );
  ix53675z14061 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => rome2addro3_s(0),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(2),
      ADR3 => rome2addro3_s(3),
      O => nx53675z199
    );
  ix53675z29406 : X_LUT4
    generic map(
      INIT => X"6644"
    )
    port map (
      ADR0 => romo2addro8_s(1),
      ADR1 => romo2addro8_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro8_s(3),
      O => nx53675z1372
    );
  ix53675z24455 : X_LUT4
    generic map(
      INIT => X"492C"
    )
    port map (
      ADR0 => rome2addro3_s(2),
      ADR1 => rome2addro3_s(3),
      ADR2 => rome2addro3_s(0),
      ADR3 => rome2addro3_s(1),
      O => nx53675z229
    );
  ix53675z25952 : X_LUT4
    generic map(
      INIT => X"3C6C"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1044
    );
  ix53675z26520 : X_LUT4
    generic map(
      INIT => X"18A6"
    )
    port map (
      ADR0 => rome2addro3_s(2),
      ADR1 => rome2addro3_s(3),
      ADR2 => rome2addro3_s(0),
      ADR3 => rome2addro3_s(1),
      O => nx53675z226
    );
  ix53675z55068 : X_LUT4
    generic map(
      INIT => X"AA56"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1042
    );
  ix53675z41347 : X_LUT4
    generic map(
      INIT => X"96A6"
    )
    port map (
      ADR0 => romo2addro4_s(0),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(1),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1045
    );
  ix53675z4290 : X_LUT4
    generic map(
      INIT => X"333C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro3_s(3),
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(0),
      O => nx53675z1025
    );
  ix53675z10693 : X_LUT4
    generic map(
      INIT => X"36C8"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1041
    );
  ix53675z55041 : X_LUT4
    generic map(
      INIT => X"CF30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro3_s(3),
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(1),
      O => nx53675z1022
    );
  ix53675z10471 : X_LUT4
    generic map(
      INIT => X"0F5A"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(1),
      O => nx53675z1026
    );
  ix53675z28371 : X_LUT4
    generic map(
      INIT => X"59E6"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1078
    );
  ix53675z29664 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2addro9_s(0),
      ADR1 => romo2addro9_s(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1502
    );
  ix53675z16707 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => romo2addro9_s(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROMO9_modgen_rom_ix0_nx_rm64_16_l
    );
  ix53675z23149 : X_LUT4
    generic map(
      INIT => X"3C16"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1080
    );
  ix53675z23256 : X_LUT4
    generic map(
      INIT => X"0A2A"
    )
    port map (
      ADR0 => romo2addro3_s(2),
      ADR1 => romo2addro3_s(1),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(3),
      O => nx53675z953
    );
  ix53675z37249 : X_LUT4
    generic map(
      INIT => X"8770"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1081
    );
  ix53675z48419 : X_LUT4
    generic map(
      INIT => X"B2F2"
    )
    port map (
      ADR0 => romo2addro3_s(2),
      ADR1 => romo2addro3_s(1),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(3),
      O => nx53675z954
    );
  ix53675z2732 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => romo2addro3_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro3_s(3),
      O => nx53675z1017
    );
  ix53675z23152 : X_LUT4
    generic map(
      INIT => X"0A2A"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(3),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(1),
      O => nx53675z880
    );
  ix53675z54844 : X_LUT4
    generic map(
      INIT => X"AA56"
    )
    port map (
      ADR0 => romo2addro2_s(1),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(2),
      ADR3 => romo2addro2_s(3),
      O => nx53675z884
    );
  ix53675z59901 : X_LUT4
    generic map(
      INIT => X"8880"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(3),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(1),
      O => nx53675z877
    );
  ix53675z48315 : X_LUT4
    generic map(
      INIT => X"B0FA"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(3),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(1),
      O => nx53675z881
    );
  ix53675z25728 : X_LUT4
    generic map(
      INIT => X"3C78"
    )
    port map (
      ADR0 => romo2addro2_s(1),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(2),
      ADR3 => romo2addro2_s(3),
      O => nx53675z886
    );
  ix53675z55036 : X_LUT4
    generic map(
      INIT => X"FF32"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(3),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(1),
      O => nx53675z878
    );
  ix53675z41123 : X_LUT4
    generic map(
      INIT => X"969C"
    )
    port map (
      ADR0 => romo2addro2_s(1),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(2),
      ADR3 => romo2addro2_s(3),
      O => nx53675z887
    );
  ix53675z59186 : X_LUT4
    generic map(
      INIT => X"F05A"
    )
    port map (
      ADR0 => romo2addro2_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z892
    );
  ix53675z10469 : X_LUT4
    generic map(
      INIT => X"1EE0"
    )
    port map (
      ADR0 => romo2addro2_s(1),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(2),
      ADR3 => romo2addro2_s(3),
      O => nx53675z883
    );
  ix53675z42921 : X_LUT4
    generic map(
      INIT => X"BB54"
    )
    port map (
      ADR0 => romo2addro2_s(0),
      ADR1 => romo2addro2_s(2),
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z889
    );
  ix53675z25127 : X_LUT4
    generic map(
      INIT => X"4B24"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(0),
      ADR3 => rome2addro10_s(3),
      O => nx53675z699
    );
  ix53675z29436 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1344
    );
  ix53675z16479 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romo2addro7_s(3),
      O => U2_ROMO7_modgen_rom_ix0_nx_rm64_16_l
    );
  ix53675z12871 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(0),
      ADR3 => rome2addro10_s(3),
      O => nx53675z701
    );
  ix53675z29355 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(2),
      O => nx53675z712
    );
  ix53675z9612 : X_LUT4
    generic map(
      INIT => X"4694"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(0),
      ADR3 => rome2addro10_s(3),
      O => nx53675z702
    );
  ix53675z19425 : X_LUT4
    generic map(
      INIT => X"42D4"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(2),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(0),
      O => nx53675z707
    );
  ix53675z62104 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(1),
      ADR2 => rome2addro10_s(0),
      ADR3 => rome2addro10_s(3),
      O => nx53675z698
    );
  ix53675z34802 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(2),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(0),
      O => nx53675z704
    );
  ix53675z28328 : X_LUT4
    generic map(
      INIT => X"59A6"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(2),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(0),
      O => nx53675z708
    );
  ix53675z14877 : X_LUT4
    generic map(
      INIT => X"03C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro2_s(2),
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z893
    );
  ix53675z28730 : X_LUT4
    generic map(
      INIT => X"22CC"
    )
    port map (
      ADR0 => romo2addro2_s(3),
      ADR1 => romo2addro2_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(1),
      O => nx53675z898
    );
  ix53675z24414 : X_LUT4
    generic map(
      INIT => X"5454"
    )
    port map (
      ADR0 => romo2addro2_s(0),
      ADR1 => romo2addro2_s(2),
      ADR2 => romo2addro2_s(3),
      ADR3 => VCC,
      O => nx53675z890
    );
  ix53675z51989 : X_LUT4
    generic map(
      INIT => X"DD44"
    )
    port map (
      ADR0 => romo2addro2_s(3),
      ADR1 => romo2addro2_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(2),
      O => nx53675z899
    );
  ix53675z11364 : X_LUT4
    generic map(
      INIT => X"4242"
    )
    port map (
      ADR0 => romo2addro2_s(1),
      ADR1 => romo2addro2_s(3),
      ADR2 => romo2addro2_s(0),
      ADR3 => VCC,
      O => nx53675z904
    );
  ix53675z23405 : X_LUT4
    generic map(
      INIT => X"0F42"
    )
    port map (
      ADR0 => romo2addro2_s(3),
      ADR1 => romo2addro2_s(1),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(2),
      O => nx53675z895
    );
  ix53675z6640 : X_LUT4
    generic map(
      INIT => X"45FA"
    )
    port map (
      ADR0 => romo2addro2_s(3),
      ADR1 => romo2addro2_s(1),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(2),
      O => nx53675z896
    );
  ix53675z5471 : X_LUT4
    generic map(
      INIT => X"02D4"
    )
    port map (
      ADR0 => romo2addro2_s(1),
      ADR1 => romo2addro2_s(3),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(2),
      O => nx53675z901
    );
  ix53675z64849 : X_LUT4
    generic map(
      INIT => X"DD44"
    )
    port map (
      ADR0 => romo2addro2_s(1),
      ADR1 => romo2addro2_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(2),
      O => nx53675z905
    );
  ix53675z17194 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(1),
      O => nx53675z324
    );
  ix53675z23702 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => rome2addro4_s(3),
      ADR1 => VCC,
      ADR2 => rome2addro4_s(0),
      ADR3 => VCC,
      O => U2_ROME4_modgen_rom_ix2_nx_rm64_16_l
    );
  ix53675z30413 : X_LUT4
    generic map(
      INIT => X"4F04"
    )
    port map (
      ADR0 => rome2addro1_s(0),
      ADR1 => rome2addro1_s(3),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z90
    );
  ix53675z18483 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(1),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(3),
      O => nx53675z92
    );
  ix53675z25252 : X_LUT4
    generic map(
      INIT => X"4F04"
    )
    port map (
      ADR0 => rome2addro1_s(2),
      ADR1 => rome2addro1_s(1),
      ADR2 => rome2addro1_s(0),
      ADR3 => rome2addro1_s(3),
      O => nx53675z93
    );
  ix53675z39940 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => rome2addro1_s(0),
      ADR1 => rome2addro1_s(3),
      ADR2 => rome2addro1_s(1),
      ADR3 => rome2addro1_s(2),
      O => nx53675z89
    );
  ix53675z24056 : X_LUT4
    generic map(
      INIT => X"04CC"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1512
    );
  ix53675z17825 : X_LUT4
    generic map(
      INIT => X"693C"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(2),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(0),
      O => nx53675z705
    );
  ix53675z29352 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(0),
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(2),
      O => U2_ROME10_modgen_rom_ix2_nx_rm64_16_u
    );
  ix53675z14662 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rome2addro10_s(1),
      ADR3 => rome2addro10_s(2),
      O => nx53675z713
    );
  ix53675z2493 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => rome2addro10_s(3),
      ADR1 => rome2addro10_s(0),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z710
    );
  ix53675z17752 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2addro10_s(2),
      ADR1 => rome2addro10_s(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z714
    );
  ix53675z24260 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2addro10_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2addro10_s(3),
      O => U2_ROME10_modgen_rom_ix2_nx_rm64_16_l
    );
  ix53675z48645 : X_LUT4
    generic map(
      INIT => X"CF4C"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => romo2addro5_s(0),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1112
    );
  ix53675z44323 : X_LUT4
    generic map(
      INIT => X"AA10"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(3),
      ADR3 => romo2addro5_s(0),
      O => nx53675z1153
    );
  ix53675z38833 : X_LUT4
    generic map(
      INIT => X"C242"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(3),
      ADR3 => romo2addro5_s(0),
      O => nx53675z1151
    );
  ix53675z28485 : X_LUT4
    generic map(
      INIT => X"6B3C"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => romo2addro5_s(3),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1157
    );
  ix53675z62476 : X_LUT4
    generic map(
      INIT => X"EC80"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(3),
      ADR3 => romo2addro5_s(0),
      O => nx53675z1154
    );
  ix53675z29942 : X_LUT4
    generic map(
      INIT => X"639C"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(3),
      ADR3 => romo2addro5_s(0),
      O => nx53675z1162
    );
  ix53675z21733 : X_LUT4
    generic map(
      INIT => X"51A6"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => romo2addro5_s(3),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1159
    );
  ix53675z23172 : X_LUT4
    generic map(
      INIT => X"50D4"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(3),
      ADR3 => romo2addro5_s(0),
      O => nx53675z1150
    );
  ix53675z37362 : X_LUT4
    generic map(
      INIT => X"925A"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => romo2addro5_s(3),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1160
    );
  ix53675z20028 : X_LUT4
    generic map(
      INIT => X"6318"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => romo2addro5_s(3),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1156
    );
  ix53675z40799 : X_LUT4
    generic map(
      INIT => X"9C3C"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(3),
      ADR3 => romo2addro5_s(0),
      O => nx53675z1165
    );
  U_DCT2D_reg_romoaddro5_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro5_s_1_DYMUX,
      CE => romo2addro5_s_1_CEINV,
      CLK => romo2addro5_s_1_CLKINV,
      SET => GND,
      RST => romo2addro5_s_1_FFY_RST,
      O => romo2addro5_s(0)
    );
  romo2addro5_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro5_s_1_SRINV,
      I1 => GSR,
      O => romo2addro5_s_1_FFY_RST
    );
  U_DCT2D_reg_romoaddro5_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro5_s_1_DXMUX,
      CE => romo2addro5_s_1_CEINV,
      CLK => romo2addro5_s_1_CLKINV,
      SET => GND,
      RST => romo2addro5_s_1_FFX_RST,
      O => romo2addro5_s(1)
    );
  romo2addro5_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro5_s_1_SRINV,
      I1 => GSR,
      O => romo2addro5_s_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_5_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_3_DYMUX,
      CE => U_DCT1D_latchbuf_reg_5_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_5_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_5_3_FFY_RST,
      O => U_DCT1D_latchbuf_reg_5_Q(2)
    );
  U_DCT1D_latchbuf_reg_5_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_5_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_5_3_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_5_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_3_DXMUX,
      CE => U_DCT1D_latchbuf_reg_5_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_5_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_5_3_FFX_RST,
      O => U_DCT1D_latchbuf_reg_5_Q(3)
    );
  U_DCT1D_latchbuf_reg_5_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_5_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_5_3_FFX_RST
    );
  U_DCT2D_reg_romoaddro5_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro5_s_3_DYMUX,
      CE => romo2addro5_s_3_CEINV,
      CLK => romo2addro5_s_3_CLKINV,
      SET => GND,
      RST => romo2addro5_s_3_FFY_RST,
      O => romo2addro5_s(2)
    );
  romo2addro5_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro5_s_3_SRINV,
      I1 => GSR,
      O => romo2addro5_s_3_FFY_RST
    );
  U_DCT2D_reg_romoaddro5_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro5_s_3_DXMUX,
      CE => romo2addro5_s_3_CEINV,
      CLK => romo2addro5_s_3_CLKINV,
      SET => GND,
      RST => romo2addro5_s_3_FFX_RST,
      O => romo2addro5_s(3)
    );
  romo2addro5_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro5_s_3_SRINV,
      I1 => GSR,
      O => romo2addro5_s_3_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_5_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_5_DYMUX,
      CE => U_DCT1D_latchbuf_reg_5_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_5_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_5_5_FFY_RST,
      O => U_DCT1D_latchbuf_reg_5_Q(4)
    );
  U_DCT1D_latchbuf_reg_5_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_5_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_5_5_FFY_RST
    );
  ix53675z3934 : X_LUT4
    generic map(
      INIT => X"2B22"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(1),
      O => nx53675z282
    );
  ix53675z18867 : X_LUT4
    generic map(
      INIT => X"188E"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => rome2addro4_s(2),
      ADR2 => rome2addro4_s(0),
      ADR3 => rome2addro4_s(3),
      O => nx53675z317
    );
  ix53675z21433 : X_LUT4
    generic map(
      INIT => X"4F04"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(1),
      O => nx53675z279
    );
  ix53675z34244 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => rome2addro4_s(2),
      ADR2 => rome2addro4_s(0),
      ADR3 => rome2addro4_s(3),
      O => nx53675z314
    );
  ix53675z27770 : X_LUT4
    generic map(
      INIT => X"4BB4"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => rome2addro4_s(2),
      ADR2 => rome2addro4_s(0),
      ADR3 => rome2addro4_s(3),
      O => nx53675z318
    );
  ix53675z28797 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => rome2addro4_s(0),
      ADR2 => rome2addro4_s(3),
      ADR3 => rome2addro4_s(2),
      O => nx53675z322
    );
  ix53675z17267 : X_LUT4
    generic map(
      INIT => X"6696"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => rome2addro4_s(2),
      ADR2 => rome2addro4_s(0),
      ADR3 => rome2addro4_s(3),
      O => nx53675z315
    );
  ix53675z14104 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => VCC,
      ADR2 => rome2addro4_s(2),
      ADR3 => VCC,
      O => nx53675z323
    );
  ix53675z28794 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => rome2addro4_s(0),
      ADR2 => rome2addro4_s(3),
      ADR3 => rome2addro4_s(2),
      O => U2_ROME4_modgen_rom_ix2_nx_rm64_16_u
    );
  ix53675z1935 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2addro4_s(0),
      ADR2 => rome2addro4_s(3),
      ADR3 => VCC,
      O => nx53675z320
    );
  ix53675z17008 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rome2addro2_s(2),
      ADR3 => rome2addro2_s(1),
      O => nx53675z194
    );
  ix53675z23516 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2addro2_s(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2addro2_s(0),
      O => U2_ROME2_modgen_rom_ix2_nx_rm64_16_l
    );
  ix53675z55635 : X_LUT4
    generic map(
      INIT => X"F10E"
    )
    port map (
      ADR0 => romo2addro9_s(2),
      ADR1 => romo2addro9_s(0),
      ADR2 => romo2addro9_s(3),
      ADR3 => romo2addro9_s(1),
      O => nx53675z1437
    );
  ix53675z26519 : X_LUT4
    generic map(
      INIT => X"666A"
    )
    port map (
      ADR0 => romo2addro9_s(2),
      ADR1 => romo2addro9_s(0),
      ADR2 => romo2addro9_s(3),
      ADR3 => romo2addro9_s(1),
      O => nx53675z1439
    );
  ix53675z43712 : X_LUT4
    generic map(
      INIT => X"99BA"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(0),
      ADR2 => romo2addro9_s(3),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1442
    );
  ix53675z41914 : X_LUT4
    generic map(
      INIT => X"9C66"
    )
    port map (
      ADR0 => romo2addro9_s(2),
      ADR1 => romo2addro9_s(0),
      ADR2 => romo2addro9_s(3),
      ADR3 => romo2addro9_s(1),
      O => nx53675z1440
    );
  ix53675z11260 : X_LUT4
    generic map(
      INIT => X"5A68"
    )
    port map (
      ADR0 => romo2addro9_s(2),
      ADR1 => romo2addro9_s(0),
      ADR2 => romo2addro9_s(3),
      ADR3 => romo2addro9_s(1),
      O => nx53675z1436
    );
  ix53675z59977 : X_LUT4
    generic map(
      INIT => X"A5AA"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro9_s(1),
      ADR3 => romo2addro9_s(0),
      O => nx53675z1445
    );
  ix53675z23112 : X_LUT4
    generic map(
      INIT => X"1C30"
    )
    port map (
      ADR0 => romo2addro2_s(1),
      ADR1 => romo2addro2_s(3),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(2),
      O => nx53675z902
    );
  ix53675z17659 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2addro9_s(2),
      ADR2 => rome2addro9_s(1),
      ADR3 => VCC,
      O => nx53675z649
    );
  ix53675z24167 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2addro9_s(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2addro9_s(0),
      O => U2_ROME9_modgen_rom_ix2_nx_rm64_16_l
    );
  ix53675z24048 : X_LUT4
    generic map(
      INIT => X"04CC"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1506
    );
  ix53675z49211 : X_LUT4
    generic map(
      INIT => X"DF44"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1507
    );
  ix53675z55140 : X_LUT4
    generic map(
      INIT => X"CCFE"
    )
    port map (
      ADR0 => romo2addro3_s(2),
      ADR1 => romo2addro3_s(1),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(3),
      O => nx53675z951
    );
  ix53675z4179 : X_LUT4
    generic map(
      INIT => X"555A"
    )
    port map (
      ADR0 => romo2addro2_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro2_s(2),
      ADR3 => romo2addro2_s(0),
      O => nx53675z946
    );
  ix53675z10360 : X_LUT4
    generic map(
      INIT => X"5566"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(0),
      O => nx53675z947
    );
  ix53675z54930 : X_LUT4
    generic map(
      INIT => X"9C9C"
    )
    port map (
      ADR0 => romo2addro2_s(3),
      ADR1 => romo2addro2_s(1),
      ADR2 => romo2addro2_s(2),
      ADR3 => VCC,
      O => nx53675z943
    );
  ix53675z24509 : X_LUT4
    generic map(
      INIT => X"11EE"
    )
    port map (
      ADR0 => romo2addro2_s(3),
      ADR1 => romo2addro2_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(0),
      O => nx53675z944
    );
  ix53675z25787 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romo2addro2_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romo2addro2_s(2),
      O => nx53675z948
    );
  ix53675z28872 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romo2addro2_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romo2addro2_s(1),
      O => nx53675z949
    );
  ix53675z6734 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro2_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(2),
      O => U2_ROMO2_modgen_rom_ix0_nx_rm64_16_u
    );
  ix53675z55834 : X_LUT4
    generic map(
      INIT => X"F50A"
    )
    port map (
      ADR0 => romo2addro10_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1575
    );
  ix53675z11264 : X_LUT4
    generic map(
      INIT => X"555A"
    )
    port map (
      ADR0 => romo2addro10_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro10_s(0),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1579
    );
  ix53675z25413 : X_LUT4
    generic map(
      INIT => X"333C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro10_s(0),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1576
    );
  ix53675z26691 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro10_s(0),
      ADR2 => romo2addro10_s(2),
      ADR3 => VCC,
      O => nx53675z1580
    );
  ix53675z29776 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro10_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro10_s(1),
      O => nx53675z1581
    );
  ix53675z7638 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romo2addro10_s(2),
      ADR3 => romo2addro10_s(3),
      O => U2_ROMO10_modgen_rom_ix0_nx_rm64_16_u
    );
  ix53675z16819 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(1),
      O => U2_ROMO10_modgen_rom_ix0_nx_rm64_16_l
    );
  ix53675z26579 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2addro9_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro9_s(0),
      ADR3 => VCC,
      O => nx53675z1501
    );
  ix53675z7526 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romo2addro9_s(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romo2addro9_s(3),
      O => U2_ROMO9_modgen_rom_ix0_nx_rm64_16_u
    );
  ix53675z29098 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romo2addro4_s(0),
      O => nx53675z1107
    );
  ix53675z4287 : X_LUT4
    generic map(
      INIT => X"0C8E"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z527
    );
  ix53675z16141 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romo2addro4_s(3),
      O => U2_ROMO4_modgen_rom_ix0_nx_rm64_16_l
    );
  ix53675z18663 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z529
    );
  ix53675z14534 : X_LUT4
    generic map(
      INIT => X"3B02"
    )
    port map (
      ADR0 => rome2addro8_s(0),
      ADR1 => rome2addro8_s(1),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z530
    );
  ix53675z19119 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(3),
      ADR2 => rome2addro8_s(0),
      ADR3 => rome2addro8_s(1),
      O => nx53675z535
    );
  ix53675z61584 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z526
    );
  ix53675z7808 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(3),
      ADR2 => rome2addro8_s(0),
      ADR3 => rome2addro8_s(1),
      O => nx53675z532
    );
  ix53675z8383 : X_LUT4
    generic map(
      INIT => X"6138"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(3),
      ADR2 => rome2addro8_s(0),
      ADR3 => rome2addro8_s(1),
      O => nx53675z533
    );
  ix53675z15534 : X_LUT4
    generic map(
      INIT => X"249A"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(3),
      ADR2 => rome2addro8_s(0),
      ADR3 => rome2addro8_s(1),
      O => nx53675z536
    );
  ix53675z12645 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => rome2addro8_s(3),
      ADR1 => rome2addro8_s(1),
      ADR2 => rome2addro8_s(0),
      ADR3 => rome2addro8_s(2),
      O => nx53675z541
    );
  ix53675z62588 : X_LUT4
    generic map(
      INIT => X"E8A0"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(2),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1233
    );
  ix53675z21845 : X_LUT4
    generic map(
      INIT => X"495A"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(0),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1238
    );
  ix53675z38945 : X_LUT4
    generic map(
      INIT => X"B00C"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(2),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1230
    );
  ix53675z28597 : X_LUT4
    generic map(
      INIT => X"39E6"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(0),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1236
    );
  ix53675z26283 : X_LUT4
    generic map(
      INIT => X"6868"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(3),
      ADR2 => romo2addro6_s(0),
      ADR3 => VCC,
      O => nx53675z1250
    );
  ix53675z37474 : X_LUT4
    generic map(
      INIT => X"943C"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(0),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1239
    );
  ix53675z40911 : X_LUT4
    generic map(
      INIT => X"9C3C"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(3),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1244
    );
  ix53675z20140 : X_LUT4
    generic map(
      INIT => X"18A6"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(0),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1235
    );
  ix53675z30054 : X_LUT4
    generic map(
      INIT => X"6696"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(3),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1241
    );
  ix53675z11236 : X_LUT4
    generic map(
      INIT => X"1EF0"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(3),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1245
    );
  ix53675z15915 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro2_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(1),
      O => U2_ROMO2_modgen_rom_ix0_nx_rm64_16_l
    );
  ix53675z41503 : X_LUT4
    generic map(
      INIT => X"C338"
    )
    port map (
      ADR0 => romo2addro1_s(2),
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(0),
      ADR3 => romo2addro1_s(1),
      O => nx53675z831
    );
  ix53675z38383 : X_LUT4
    generic map(
      INIT => X"C422"
    )
    port map (
      ADR0 => romo2addro1_s(2),
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(0),
      ADR3 => romo2addro1_s(3),
      O => nx53675z835
    );
  ix53675z58184 : X_LUT4
    generic map(
      INIT => X"E81E"
    )
    port map (
      ADR0 => romo2addro1_s(2),
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(0),
      ADR3 => romo2addro1_s(1),
      O => nx53675z828
    );
  ix53675z44833 : X_LUT4
    generic map(
      INIT => X"96B4"
    )
    port map (
      ADR0 => romo2addro1_s(2),
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(0),
      ADR3 => romo2addro1_s(1),
      O => nx53675z829
    );
  ix53675z52470 : X_LUT4
    generic map(
      INIT => X"9696"
    )
    port map (
      ADR0 => romo2addro1_s(1),
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(2),
      ADR3 => VCC,
      O => nx53675z832
    );
  ix53675z43873 : X_LUT4
    generic map(
      INIT => X"A1A0"
    )
    port map (
      ADR0 => romo2addro1_s(2),
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(0),
      ADR3 => romo2addro1_s(3),
      O => nx53675z837
    );
  ix53675z62026 : X_LUT4
    generic map(
      INIT => X"E8C0"
    )
    port map (
      ADR0 => romo2addro1_s(2),
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(0),
      ADR3 => romo2addro1_s(3),
      O => nx53675z838
    );
  ix53675z21283 : X_LUT4
    generic map(
      INIT => X"31C6"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => romo2addro1_s(0),
      ADR2 => romo2addro1_s(1),
      ADR3 => romo2addro1_s(2),
      O => nx53675z843
    );
  ix53675z22722 : X_LUT4
    generic map(
      INIT => X"5D04"
    )
    port map (
      ADR0 => romo2addro1_s(2),
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(0),
      ADR3 => romo2addro1_s(3),
      O => nx53675z834
    );
  ix53675z19578 : X_LUT4
    generic map(
      INIT => X"6518"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => romo2addro1_s(0),
      ADR2 => romo2addro1_s(1),
      ADR3 => romo2addro1_s(2),
      O => nx53675z840
    );
  ix53675z2406 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro0_s(1),
      O => nx53675z782
    );
  ix53675z3964 : X_LUT4
    generic map(
      INIT => X"0F5A"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(0),
      O => nx53675z790
    );
  ix53675z21340 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => rome2addro3_s(2),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(0),
      ADR3 => rome2addro3_s(3),
      O => nx53675z214
    );
  ix53675z54715 : X_LUT4
    generic map(
      INIT => X"F50A"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(1),
      O => nx53675z787
    );
  ix53675z10145 : X_LUT4
    generic map(
      INIT => X"0F5A"
    )
    port map (
      ADR0 => romo2addro0_s(1),
      ADR1 => VCC,
      ADR2 => romo2addro0_s(2),
      ADR3 => romo2addro0_s(0),
      O => nx53675z791
    );
  ix53675z24294 : X_LUT4
    generic map(
      INIT => X"05FA"
    )
    port map (
      ADR0 => romo2addro0_s(1),
      ADR1 => VCC,
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(0),
      O => nx53675z788
    );
  ix53675z12180 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro3_s(2),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(0),
      ADR3 => rome2addro3_s(3),
      O => nx53675z216
    );
  ix53675z3841 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => rome2addro3_s(2),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(0),
      ADR3 => rome2addro3_s(3),
      O => nx53675z217
    );
  ix53675z12644 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => rome2addro3_s(2),
      ADR1 => rome2addro3_s(3),
      ADR2 => rome2addro3_s(0),
      ADR3 => rome2addro3_s(1),
      O => nx53675z228
    );
  ix53675z34661 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => rome2addro3_s(2),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(0),
      ADR3 => rome2addro3_s(3),
      O => nx53675z213
    );
  ix53675z7645 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => rome2addro3_s(2),
      ADR1 => rome2addro3_s(3),
      ADR2 => rome2addro3_s(0),
      ADR3 => rome2addro3_s(1),
      O => nx53675z225
    );
  ix53675z24620 : X_LUT4
    generic map(
      INIT => X"3366"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro3_s(1),
      O => nx53675z1023
    );
  ix53675z22930 : X_LUT4
    generic map(
      INIT => X"222A"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(0),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(1),
      O => nx53675z718
    );
  ix53675z48093 : X_LUT4
    generic map(
      INIT => X"C4FC"
    )
    port map (
      ADR0 => romo2addro0_s(3),
      ADR1 => romo2addro0_s(0),
      ADR2 => romo2addro0_s(2),
      ADR3 => romo2addro0_s(1),
      O => nx53675z719
    );
  ix53675z54814 : X_LUT4
    generic map(
      INIT => X"FF0E"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(0),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(1),
      O => nx53675z716
    );
  ix53675z55712 : X_LUT4
    generic map(
      INIT => X"CCFE"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(0),
      ADR3 => romo2addro8_s(3),
      O => nx53675z1352
    );
  ix53675z23828 : X_LUT4
    generic map(
      INIT => X"0A2A"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(0),
      ADR3 => romo2addro8_s(3),
      O => nx53675z1354
    );
  ix53675z48991 : X_LUT4
    generic map(
      INIT => X"B2F2"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(0),
      ADR3 => romo2addro8_s(3),
      O => nx53675z1355
    );
  ix53675z60577 : X_LUT4
    generic map(
      INIT => X"A800"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(0),
      ADR3 => romo2addro8_s(3),
      O => nx53675z1351
    );
  ix53675z41136 : X_LUT4
    generic map(
      INIT => X"93CC"
    )
    port map (
      ADR0 => romo2addro8_s(0),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(3),
      O => nx53675z1402
    );
  ix53675z30279 : X_LUT4
    generic map(
      INIT => X"6966"
    )
    port map (
      ADR0 => romo2addro8_s(0),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(3),
      O => nx53675z1399
    );
  ix53675z55932 : X_LUT4
    generic map(
      INIT => X"AFAE"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1504
    );
  ix53675z60091 : X_LUT4
    generic map(
      INIT => X"9C9C"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(0),
      ADR3 => VCC,
      O => nx53675z1524
    );
  ix53675z15782 : X_LUT4
    generic map(
      INIT => X"500A"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => VCC,
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(2),
      O => nx53675z1525
    );
  ix53675z3795 : X_LUT4
    generic map(
      INIT => X"3330"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(0),
      ADR3 => romo2addro10_s(2),
      O => nx53675z1572
    );
  ix53675z43826 : X_LUT4
    generic map(
      INIT => X"99BA"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(0),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(2),
      O => nx53675z1521
    );
  ix53675z25319 : X_LUT4
    generic map(
      INIT => X"0F0A"
    )
    port map (
      ADR0 => romo2addro10_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro10_s(0),
      ADR3 => romo2addro10_s(2),
      O => nx53675z1522
    );
  ix53675z3288 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => VCC,
      ADR2 => romo2addro10_s(0),
      ADR3 => romo2addro10_s(2),
      O => nx53675z1573
    );
  ix53675z3590 : X_LUT4
    generic map(
      INIT => X"1100"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro10_s(2),
      O => nx53675z1569
    );
  ix53675z3525 : X_LUT4
    generic map(
      INIT => X"FEFE"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(0),
      ADR3 => VCC,
      O => nx53675z1570
    );
  ix53675z5083 : X_LUT4
    generic map(
      INIT => X"05FA"
    )
    port map (
      ADR0 => romo2addro10_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro10_s(0),
      ADR3 => romo2addro10_s(3),
      O => nx53675z1578
    );
  ix53675z30786 : X_LUT4
    generic map(
      INIT => X"20F2"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(0),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(1),
      O => nx53675z350
    );
  ix53675z4027 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => rome2addro5_s(1),
      ADR1 => rome2addro5_s(2),
      ADR2 => rome2addro5_s(3),
      ADR3 => rome2addro5_s(0),
      O => nx53675z347
    );
  ix53675z18856 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(0),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(1),
      O => nx53675z352
    );
  ix53675z21526 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => rome2addro5_s(1),
      ADR1 => rome2addro5_s(2),
      ADR2 => rome2addro5_s(3),
      ADR3 => rome2addro5_s(0),
      O => nx53675z344
    );
  ix53675z25625 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => rome2addro5_s(3),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(1),
      O => nx53675z353
    );
  ix53675z28890 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => rome2addro5_s(2),
      ADR2 => rome2addro5_s(1),
      ADR3 => rome2addro5_s(3),
      O => nx53675z387
    );
  ix53675z40313 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(0),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(1),
      O => nx53675z349
    );
  ix53675z28887 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => rome2addro5_s(2),
      ADR2 => rome2addro5_s(1),
      ADR3 => rome2addro5_s(3),
      O => U2_ROME5_modgen_rom_ix2_nx_rm64_16_u
    );
  ix53675z14197 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => rome2addro5_s(1),
      ADR1 => rome2addro5_s(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z388
    );
  ix53675z36912 : X_LUT4
    generic map(
      INIT => X"943C"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => romo2addro1_s(0),
      ADR2 => romo2addro1_s(1),
      ADR3 => romo2addro1_s(2),
      O => nx53675z844
    );
  ix53675z40349 : X_LUT4
    generic map(
      INIT => X"9C3C"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(2),
      O => nx53675z849
    );
  ix53675z28035 : X_LUT4
    generic map(
      INIT => X"6D5A"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => romo2addro1_s(0),
      ADR2 => romo2addro1_s(1),
      ADR3 => romo2addro1_s(2),
      O => nx53675z841
    );
  ix53675z25671 : X_LUT4
    generic map(
      INIT => X"57A8"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(2),
      O => nx53675z847
    );
  ix53675z10674 : X_LUT4
    generic map(
      INIT => X"1EF0"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(2),
      O => nx53675z850
    );
  ix53675z25721 : X_LUT4
    generic map(
      INIT => X"3CC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(2),
      ADR3 => romo2addro1_s(0),
      O => nx53675z855
    );
  ix53675z29492 : X_LUT4
    generic map(
      INIT => X"6696"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(3),
      ADR3 => romo2addro1_s(2),
      O => nx53675z846
    );
  ix53675z6550 : X_LUT4
    generic map(
      INIT => X"4A4A"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(2),
      ADR3 => VCC,
      O => nx53675z852
    );
  ix53675z41586 : X_LUT4
    generic map(
      INIT => X"CC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(2),
      ADR3 => romo2addro1_s(0),
      O => nx53675z856
    );
  ix53675z10571 : X_LUT4
    generic map(
      INIT => X"1EF0"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(1),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(2),
      O => nx53675z773
    );
  ix53675z25618 : X_LUT4
    generic map(
      INIT => X"6688"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(2),
      ADR2 => VCC,
      ADR3 => romo2addro0_s(3),
      O => nx53675z778
    );
  ix53675z25568 : X_LUT4
    generic map(
      INIT => X"57A8"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(1),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(2),
      O => nx53675z770
    );
  ix53675z6447 : X_LUT4
    generic map(
      INIT => X"5588"
    )
    port map (
      ADR0 => romo2addro0_s(2),
      ADR1 => romo2addro0_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro0_s(3),
      O => nx53675z775
    );
  ix53675z41483 : X_LUT4
    generic map(
      INIT => X"AA50"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro0_s(2),
      ADR3 => romo2addro0_s(1),
      O => nx53675z779
    );
  ix53675z54674 : X_LUT4
    generic map(
      INIT => X"CC22"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro0_s(3),
      O => nx53675z776
    );
  ix53675z2676 : X_LUT4
    generic map(
      INIT => X"3322"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro0_s(2),
      O => nx53675z784
    );
  ix53675z2471 : X_LUT4
    generic map(
      INIT => X"1100"
    )
    port map (
      ADR0 => romo2addro0_s(1),
      ADR1 => romo2addro0_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro0_s(2),
      O => nx53675z781
    );
  ix53675z2169 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(2),
      ADR2 => VCC,
      ADR3 => romo2addro0_s(1),
      O => nx53675z785
    );
  ix53675z14290 : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => rome2addro6_s(2),
      ADR1 => VCC,
      ADR2 => rome2addro6_s(1),
      ADR3 => VCC,
      O => nx53675z453
    );
  ix53675z2121 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2addro6_s(3),
      O => nx53675z450
    );
  ix53675z17380 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2addro6_s(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2addro6_s(1),
      O => nx53675z454
    );
  ix53675z23888 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROME6_modgen_rom_ix2_nx_rm64_16_l
    );
  ix53675z40246 : X_LUT4
    generic map(
      INIT => X"9C3C"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(1),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(2),
      O => nx53675z772
    );
  ix53675z29389 : X_LUT4
    generic map(
      INIT => X"6696"
    )
    port map (
      ADR0 => romo2addro0_s(0),
      ADR1 => romo2addro0_s(1),
      ADR2 => romo2addro0_s(3),
      ADR3 => romo2addro0_s(2),
      O => nx53675z769
    );
  ix53675z54777 : X_LUT4
    generic map(
      INIT => X"9988"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => romo2addro1_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro1_s(0),
      O => nx53675z853
    );
  ix53675z18477 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(1),
      ADR3 => rome2addro6_s(3),
      O => nx53675z399
    );
  ix53675z17453 : X_LUT4
    generic map(
      INIT => X"2DD2"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => nx53675z445
    );
  ix53675z61398 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(1),
      ADR3 => rome2addro6_s(3),
      O => nx53675z396
    );
  ix53675z14348 : X_LUT4
    generic map(
      INIT => X"0C8E"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(1),
      ADR3 => rome2addro6_s(3),
      O => nx53675z400
    );
  ix53675z19053 : X_LUT4
    generic map(
      INIT => X"7118"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => nx53675z447
    );
  ix53675z4101 : X_LUT4
    generic map(
      INIT => X"20BA"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(1),
      ADR3 => rome2addro6_s(3),
      O => nx53675z397
    );
  ix53675z27956 : X_LUT4
    generic map(
      INIT => X"6696"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => nx53675z448
    );
  ix53675z28980 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => U2_ROME6_modgen_rom_ix2_nx_rm64_16_u
    );
  ix53675z28983 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => nx53675z452
    );
  ix53675z34430 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => nx53675z444
    );
  ix53675z49106 : X_LUT4
    generic map(
      INIT => X"F570"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1434
    );
  ix53675z23490 : X_LUT4
    generic map(
      INIT => X"0A2A"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(0),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1117
    );
  ix53675z57863 : X_LUT4
    generic map(
      INIT => X"BBBA"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1431
    );
  ix53675z60239 : X_LUT4
    generic map(
      INIT => X"A800"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(0),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1114
    );
  ix53675z48653 : X_LUT4
    generic map(
      INIT => X"B2F2"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(0),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1118
    );
  ix53675z3116 : X_LUT4
    generic map(
      INIT => X"5550"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(2),
      O => nx53675z1098
    );
  ix53675z55374 : X_LUT4
    generic map(
      INIT => X"DDDC"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(0),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1115
    );
  ix53675z2609 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romo2addro4_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1099
    );
  ix53675z2911 : X_LUT4
    generic map(
      INIT => X"0500"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(1),
      ADR3 => romo2addro4_s(2),
      O => nx53675z1095
    );
  ix53675z2846 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1096
    );
  ix53675z28142 : X_LUT4
    generic map(
      INIT => X"3C96"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(1),
      O => nx53675z578
    );
  ix53675z12592 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(1),
      O => nx53675z506
    );
  ix53675z17639 : X_LUT4
    generic map(
      INIT => X"59A6"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(1),
      O => nx53675z575
    );
  ix53675z24848 : X_LUT4
    generic map(
      INIT => X"492C"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(1),
      O => nx53675z504
    );
  ix53675z23603 : X_LUT4
    generic map(
      INIT => X"222A"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(0),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1196
    );
  ix53675z9333 : X_LUT4
    generic map(
      INIT => X"6518"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(1),
      O => nx53675z507
    );
  ix53675z19146 : X_LUT4
    generic map(
      INIT => X"2B42"
    )
    port map (
      ADR0 => rome2addro7_s(1),
      ADR1 => rome2addro7_s(0),
      ADR2 => rome2addro7_s(3),
      ADR3 => rome2addro7_s(2),
      O => nx53675z512
    );
  ix53675z61825 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(1),
      O => nx53675z503
    );
  ix53675z34523 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro7_s(1),
      ADR1 => rome2addro7_s(0),
      ADR2 => rome2addro7_s(3),
      ADR3 => rome2addro7_s(2),
      O => nx53675z509
    );
  ix53675z28049 : X_LUT4
    generic map(
      INIT => X"693C"
    )
    port map (
      ADR0 => rome2addro7_s(1),
      ADR1 => rome2addro7_s(0),
      ADR2 => rome2addro7_s(3),
      ADR3 => rome2addro7_s(2),
      O => nx53675z513
    );
  ix53675z15441 : X_LUT4
    generic map(
      INIT => X"2692"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(3),
      O => nx53675z471
    );
  ix53675z29076 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(1),
      O => nx53675z517
    );
  ix53675z8290 : X_LUT4
    generic map(
      INIT => X"42B4"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(3),
      O => nx53675z468
    );
  ix53675z14383 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2addro7_s(2),
      ADR2 => VCC,
      ADR3 => rome2addro7_s(1),
      O => nx53675z518
    );
  ix53675z29073 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(1),
      O => U2_ROME7_modgen_rom_ix2_nx_rm64_16_u
    );
  ix53675z2214 : X_LUT4
    generic map(
      INIT => X"2222"
    )
    port map (
      ADR0 => rome2addro7_s(0),
      ADR1 => rome2addro7_s(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z515
    );
  ix53675z2028 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2addro5_s(3),
      O => nx53675z385
    );
  ix53675z17287 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2addro5_s(2),
      ADR2 => VCC,
      ADR3 => rome2addro5_s(1),
      O => nx53675z389
    );
  ix53675z23795 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => rome2addro5_s(3),
      O => U2_ROME5_modgen_rom_ix2_nx_rm64_16_l
    );
  ix53675z23820 : X_LUT4
    generic map(
      INIT => X"222A"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(0),
      ADR2 => romo2addro8_s(1),
      ADR3 => romo2addro8_s(3),
      O => nx53675z1348
    );
  ix53675z48983 : X_LUT4
    generic map(
      INIT => X"8ECE"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(0),
      ADR2 => romo2addro8_s(1),
      ADR3 => romo2addro8_s(3),
      O => nx53675z1349
    );
  ix53675z25532 : X_LUT4
    generic map(
      INIT => X"08CE"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(0),
      O => nx53675z288
    );
  ix53675z30693 : X_LUT4
    generic map(
      INIT => X"50D4"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(0),
      O => nx53675z285
    );
  ix53675z3955 : X_LUT4
    generic map(
      INIT => X"2B22"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(1),
      O => nx53675z297
    );
  ix53675z12737 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => rome2addro4_s(3),
      ADR1 => rome2addro4_s(2),
      ADR2 => rome2addro4_s(1),
      ADR3 => rome2addro4_s(0),
      O => nx53675z293
    );
  ix53675z7738 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => rome2addro4_s(3),
      ADR1 => rome2addro4_s(0),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(1),
      O => nx53675z290
    );
  ix53675z24548 : X_LUT4
    generic map(
      INIT => X"2962"
    )
    port map (
      ADR0 => rome2addro4_s(3),
      ADR1 => rome2addro4_s(0),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(1),
      O => nx53675z294
    );
  ix53675z12297 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(1),
      O => nx53675z299
    );
  ix53675z26613 : X_LUT4
    generic map(
      INIT => X"24D2"
    )
    port map (
      ADR0 => rome2addro4_s(3),
      ADR1 => rome2addro4_s(0),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(1),
      O => nx53675z291
    );
  ix53675z14202 : X_LUT4
    generic map(
      INIT => X"20F2"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(1),
      O => nx53675z300
    );
  ix53675z61530 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(1),
      O => nx53675z296
    );
  ix53675z18654 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z210
    );
  ix53675z7343 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z207
    );
  ix54672z4194 : X_LUT4
    generic map(
      INIT => X"2B22"
    )
    port map (
      ADR0 => romeaddro7_s(0),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(2),
      ADR3 => romeaddro7_s(1),
      O => nx54672z462
    );
  ix54672z10599 : X_LUT4
    generic map(
      INIT => X"666C"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(1),
      O => nx54672z799
    );
  ix54672z18570 : X_LUT4
    generic map(
      INIT => X"7110"
    )
    port map (
      ADR0 => romeaddro7_s(0),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(2),
      ADR3 => romeaddro7_s(1),
      O => nx54672z464
    );
  ix54672z25596 : X_LUT4
    generic map(
      INIT => X"5A6A"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(1),
      O => nx54672z796
    );
  ix54672z19026 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(0),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(2),
      O => nx54672z470
    );
  ix54672z14441 : X_LUT4
    generic map(
      INIT => X"20F2"
    )
    port map (
      ADR0 => romeaddro7_s(0),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(2),
      ADR3 => romeaddro7_s(1),
      O => nx54672z465
    );
  ix54672z7715 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(0),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(2),
      O => nx54672z467
    );
  ix54672z15441 : X_LUT4
    generic map(
      INIT => X"5924"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(0),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(2),
      O => nx54672z471
    );
  ix53675z55704 : X_LUT4
    generic map(
      INIT => X"F0FE"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(0),
      ADR2 => romo2addro8_s(1),
      ADR3 => romo2addro8_s(3),
      O => nx53675z1346
    );
  ix53675z4857 : X_LUT4
    generic map(
      INIT => X"0F5A"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro8_s(3),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1420
    );
  ix53675z4194 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => rome2addro7_s(0),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z462
    );
  ix53675z11038 : X_LUT4
    generic map(
      INIT => X"5566"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro8_s(0),
      O => nx53675z1421
    );
  ix53675z59629 : X_LUT4
    generic map(
      INIT => X"C6C6"
    )
    port map (
      ADR0 => romo2addro8_s(2),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(3),
      ADR3 => VCC,
      O => nx53675z1417
    );
  ix53675z25187 : X_LUT4
    generic map(
      INIT => X"03FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(3),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1418
    );
  ix53675z18570 : X_LUT4
    generic map(
      INIT => X"7110"
    )
    port map (
      ADR0 => rome2addro7_s(0),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z464
    );
  ix53675z7715 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(3),
      O => nx53675z467
    );
  ix53675z14441 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => rome2addro7_s(0),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z465
    );
  ix53675z19026 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(3),
      O => nx53675z470
    );
  ix53675z3296 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro8_s(0),
      O => nx53675z1412
    );
  ix53675z18384 : X_LUT4
    generic map(
      INIT => X"7110"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(0),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(1),
      O => nx53675z334
    );
  ix53675z4008 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(0),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(1),
      O => nx53675z332
    );
  ix53675z8104 : X_LUT4
    generic map(
      INIT => X"2962"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => rome2addro5_s(3),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(1),
      O => nx53675z338
    );
  ix53675z14255 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(0),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(1),
      O => nx53675z335
    );
  ix53675z34847 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => rome2addro5_s(1),
      ADR1 => rome2addro5_s(2),
      ADR2 => rome2addro5_s(3),
      ADR3 => rome2addro5_s(0),
      O => nx53675z343
    );
  ix53675z18840 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => rome2addro5_s(3),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(1),
      O => nx53675z340
    );
  ix53675z61305 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(0),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(1),
      O => nx53675z331
    );
  ix53675z15255 : X_LUT4
    generic map(
      INIT => X"24D2"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => rome2addro5_s(3),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(1),
      O => nx53675z341
    );
  ix53675z7529 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => rome2addro5_s(3),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(1),
      O => nx53675z337
    );
  ix53675z12366 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro5_s(1),
      ADR1 => rome2addro5_s(2),
      ADR2 => rome2addro5_s(3),
      ADR3 => rome2addro5_s(0),
      O => nx53675z346
    );
  ix53675z3412 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro9_s(1),
      ADR3 => romo2addro9_s(0),
      O => nx53675z1491
    );
  ix53675z23376 : X_LUT4
    generic map(
      INIT => X"3070"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(0),
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1038
    );
  ix53675z55260 : X_LUT4
    generic map(
      INIT => X"AAFE"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(0),
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1036
    );
  ix53675z48539 : X_LUT4
    generic map(
      INIT => X"D4DC"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(0),
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1039
    );
  ix53675z5583 : X_LUT4
    generic map(
      INIT => X"2342"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(1),
      ADR3 => romo2addro3_s(3),
      O => nx53675z980
    );
  ix53675z59298 : X_LUT4
    generic map(
      INIT => X"DD22"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => romo2addro3_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro3_s(3),
      O => nx53675z971
    );
  ix53675z60125 : X_LUT4
    generic map(
      INIT => X"E000"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(0),
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1035
    );
  ix53675z14989 : X_LUT4
    generic map(
      INIT => X"05A0"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(1),
      O => nx53675z972
    );
  ix53675z43033 : X_LUT4
    generic map(
      INIT => X"AF54"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => romo2addro3_s(3),
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(1),
      O => nx53675z968
    );
  ix53675z24526 : X_LUT4
    generic map(
      INIT => X"5550"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(3),
      O => nx53675z969
    );
  ix53675z11476 : X_LUT4
    generic map(
      INIT => X"0C30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro3_s(0),
      ADR2 => romo2addro3_s(1),
      ADR3 => romo2addro3_s(3),
      O => nx53675z983
    );
  ix53675z3862 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => rome2addro3_s(2),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(0),
      ADR3 => rome2addro3_s(3),
      O => nx53675z232
    );
  ix53675z15069 : X_LUT4
    generic map(
      INIT => X"492C"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z211
    );
  ix53675z12204 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro3_s(2),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(0),
      ADR3 => rome2addro3_s(3),
      O => nx53675z234
    );
  ix53675z7918 : X_LUT4
    generic map(
      INIT => X"6518"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z208
    );
  ix53675z14109 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => rome2addro3_s(2),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(0),
      ADR3 => rome2addro3_s(3),
      O => nx53675z235
    );
  ix53675z3682 : X_LUT4
    generic map(
      INIT => X"5544"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => romo2addro9_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro9_s(2),
      O => nx53675z1493
    );
  ix53675z61437 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro3_s(2),
      ADR1 => rome2addro3_s(1),
      ADR2 => rome2addro3_s(0),
      ADR3 => rome2addro3_s(3),
      O => nx53675z231
    );
  ix53675z3477 : X_LUT4
    generic map(
      INIT => X"0500"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro9_s(1),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1490
    );
  ix53675z3175 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romo2addro9_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro9_s(1),
      ADR3 => romo2addro9_s(0),
      O => nx53675z1494
    );
  ix53675z11461 : X_LUT4
    generic map(
      INIT => X"1FE0"
    )
    port map (
      ADR0 => romo2addro8_s(0),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(3),
      O => nx53675z1403
    );
  ix53675z26508 : X_LUT4
    generic map(
      INIT => X"5AA0"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1408
    );
  ix53675z26458 : X_LUT4
    generic map(
      INIT => X"5A78"
    )
    port map (
      ADR0 => romo2addro8_s(0),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(3),
      O => nx53675z1400
    );
  ix53675z42373 : X_LUT4
    generic map(
      INIT => X"AA50"
    )
    port map (
      ADR0 => romo2addro8_s(1),
      ADR1 => VCC,
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1409
    );
  ix53675z7337 : X_LUT4
    generic map(
      INIT => X"0FA0"
    )
    port map (
      ADR0 => romo2addro8_s(1),
      ADR1 => VCC,
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(3),
      O => nx53675z1405
    );
  ix53675z55564 : X_LUT4
    generic map(
      INIT => X"AA44"
    )
    port map (
      ADR0 => romo2addro8_s(1),
      ADR1 => romo2addro8_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro8_s(3),
      O => nx53675z1406
    );
  ix53675z5571 : X_LUT4
    generic map(
      INIT => X"5550"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1414
    );
  ix53675z3361 : X_LUT4
    generic map(
      INIT => X"1010"
    )
    port map (
      ADR0 => romo2addro8_s(3),
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => VCC,
      O => nx53675z1411
    );
  ix53675z3060 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro8_s(1),
      ADR2 => romo2addro8_s(2),
      ADR3 => romo2addro8_s(0),
      O => nx53675z1415
    );
  ix53675z26008 : X_LUT4
    generic map(
      INIT => X"56AA"
    )
    port map (
      ADR0 => romo2addro4_s(2),
      ADR1 => romo2addro4_s(1),
      ADR2 => romo2addro4_s(3),
      ADR3 => romo2addro4_s(0),
      O => nx53675z1084
    );
  ix53675z29550 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2addro8_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro8_s(1),
      ADR3 => VCC,
      O => nx53675z1423
    );
  ix53675z16593 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro8_s(3),
      ADR2 => romo2addro8_s(1),
      ADR3 => VCC,
      O => U2_ROMO8_modgen_rom_ix0_nx_rm64_16_l
    );
  ix53675z40686 : X_LUT4
    generic map(
      INIT => X"9C3C"
    )
    port map (
      ADR0 => romo2addro4_s(2),
      ADR1 => romo2addro4_s(1),
      ADR2 => romo2addro4_s(3),
      ADR3 => romo2addro4_s(0),
      O => nx53675z1086
    );
  ix53675z11011 : X_LUT4
    generic map(
      INIT => X"5A78"
    )
    port map (
      ADR0 => romo2addro4_s(2),
      ADR1 => romo2addro4_s(1),
      ADR2 => romo2addro4_s(3),
      ADR3 => romo2addro4_s(0),
      O => nx53675z1087
    );
  ix53675z18763 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(0),
      O => nx53675z287
    );
  ix53675z29829 : X_LUT4
    generic map(
      INIT => X"639C"
    )
    port map (
      ADR0 => romo2addro4_s(2),
      ADR1 => romo2addro4_s(1),
      ADR2 => romo2addro4_s(3),
      ADR3 => romo2addro4_s(0),
      O => nx53675z1083
    );
  ix53675z40220 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => rome2addro4_s(1),
      ADR1 => rome2addro4_s(3),
      ADR2 => rome2addro4_s(2),
      ADR3 => rome2addro4_s(0),
      O => nx53675z284
    );
  ix53675z28937 : X_LUT4
    generic map(
      INIT => X"6D5A"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => romo2addro9_s(0),
      ADR2 => romo2addro9_s(1),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1473
    );
  ix53675z30394 : X_LUT4
    generic map(
      INIT => X"5A96"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1478
    );
  ix53675z11576 : X_LUT4
    generic map(
      INIT => X"36CC"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1482
    );
  ix53675z7412 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro8_s(3),
      ADR2 => romo2addro8_s(2),
      ADR3 => VCC,
      O => U2_ROMO8_modgen_rom_ix0_nx_rm64_16_u
    );
  ix53675z26624 : X_LUT4
    generic map(
      INIT => X"6688"
    )
    port map (
      ADR0 => romo2addro9_s(0),
      ADR1 => romo2addro9_s(2),
      ADR2 => VCC,
      ADR3 => romo2addro9_s(3),
      O => nx53675z1487
    );
  ix53675z26573 : X_LUT4
    generic map(
      INIT => X"1FE0"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1479
    );
  ix53675z42489 : X_LUT4
    generic map(
      INIT => X"AA44"
    )
    port map (
      ADR0 => romo2addro9_s(0),
      ADR1 => romo2addro9_s(2),
      ADR2 => VCC,
      ADR3 => romo2addro9_s(1),
      O => nx53675z1488
    );
  ix53675z7452 : X_LUT4
    generic map(
      INIT => X"6644"
    )
    port map (
      ADR0 => romo2addro9_s(2),
      ADR1 => romo2addro9_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro9_s(1),
      O => nx53675z1484
    );
  ix53675z57789 : X_LUT4
    generic map(
      INIT => X"CC22"
    )
    port map (
      ADR0 => romo2addro9_s(0),
      ADR1 => romo2addro9_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro9_s(1),
      O => nx53675z1485
    );
  ix53675z26465 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2addro8_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro8_s(2),
      ADR3 => VCC,
      O => nx53675z1422
    );
  ix53675z17473 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rome2addro7_s(2),
      ADR3 => rome2addro7_s(1),
      O => nx53675z519
    );
  ix53675z23981 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(3),
      O => U2_ROME7_modgen_rom_ix2_nx_rm64_16_l
    );
  ix53675z39285 : X_LUT4
    generic map(
      INIT => X"C422"
    )
    port map (
      ADR0 => romo2addro9_s(2),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(1),
      O => nx53675z1467
    );
  ix53675z44775 : X_LUT4
    generic map(
      INIT => X"A0A4"
    )
    port map (
      ADR0 => romo2addro9_s(2),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(1),
      O => nx53675z1469
    );
  ix53675z41251 : X_LUT4
    generic map(
      INIT => X"A666"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1481
    );
  ix53675z62928 : X_LUT4
    generic map(
      INIT => X"F880"
    )
    port map (
      ADR0 => romo2addro9_s(2),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(1),
      O => nx53675z1470
    );
  ix53675z22185 : X_LUT4
    generic map(
      INIT => X"31C6"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => romo2addro9_s(0),
      ADR2 => romo2addro9_s(1),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1475
    );
  ix53675z23624 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => romo2addro9_s(2),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(1),
      O => nx53675z1466
    );
  ix53675z20480 : X_LUT4
    generic map(
      INIT => X"6518"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => romo2addro9_s(0),
      ADR2 => romo2addro9_s(1),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1472
    );
  ix53675z37814 : X_LUT4
    generic map(
      INIT => X"943C"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => romo2addro9_s(0),
      ADR2 => romo2addro9_s(1),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1476
    );
  ix53675z44944 : X_LUT4
    generic map(
      INIT => X"96B4"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(3),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(1),
      O => nx53675z908
    );
  ix53675z52581 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(1),
      O => nx53675z911
    );
  ix53675z28146 : X_LUT4
    generic map(
      INIT => X"2DDA"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z920
    );
  ix53675z43984 : X_LUT4
    generic map(
      INIT => X"8988"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(1),
      ADR3 => romo2addro2_s(3),
      O => nx53675z916
    );
  ix53675z22833 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(1),
      ADR3 => romo2addro2_s(3),
      O => nx53675z913
    );
  ix53675z62137 : X_LUT4
    generic map(
      INIT => X"E8C0"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(1),
      ADR3 => romo2addro2_s(3),
      O => nx53675z917
    );
  ix53675z21394 : X_LUT4
    generic map(
      INIT => X"6616"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z922
    );
  ix53675z38494 : X_LUT4
    generic map(
      INIT => X"D00A"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(1),
      ADR3 => romo2addro2_s(3),
      O => nx53675z914
    );
  ix53675z37023 : X_LUT4
    generic map(
      INIT => X"934C"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z923
    );
  ix53675z40460 : X_LUT4
    generic map(
      INIT => X"8F70"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z928
    );
  ix53675z19689 : X_LUT4
    generic map(
      INIT => X"294A"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z919
    );
  ix53675z65754 : X_LUT4
    generic map(
      INIT => X"C0FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(2),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1537
    );
  ix53675z42519 : X_LUT4
    generic map(
      INIT => X"A558"
    )
    port map (
      ADR0 => romo2addro10_s(3),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(1),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1542
    );
  ix53675z24017 : X_LUT4
    generic map(
      INIT => X"4262"
    )
    port map (
      ADR0 => romo2addro10_s(0),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(2),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1534
    );
  ix53675z39399 : X_LUT4
    generic map(
      INIT => X"8C30"
    )
    port map (
      ADR0 => romo2addro10_s(0),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(2),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1546
    );
  ix53675z45849 : X_LUT4
    generic map(
      INIT => X"9D62"
    )
    port map (
      ADR0 => romo2addro10_s(3),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(1),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1540
    );
  ix53675z53486 : X_LUT4
    generic map(
      INIT => X"9696"
    )
    port map (
      ADR0 => romo2addro10_s(3),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(1),
      ADR3 => VCC,
      O => nx53675z1543
    );
  ix53675z44889 : X_LUT4
    generic map(
      INIT => X"C0C2"
    )
    port map (
      ADR0 => romo2addro10_s(3),
      ADR1 => romo2addro10_s(0),
      ADR2 => romo2addro10_s(2),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1548
    );
  ix53675z59200 : X_LUT4
    generic map(
      INIT => X"E18E"
    )
    port map (
      ADR0 => romo2addro10_s(3),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(1),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1539
    );
  ix53675z63042 : X_LUT4
    generic map(
      INIT => X"EC80"
    )
    port map (
      ADR0 => romo2addro10_s(3),
      ADR1 => romo2addro10_s(0),
      ADR2 => romo2addro10_s(2),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1549
    );
  ix53675z22299 : X_LUT4
    generic map(
      INIT => X"6616"
    )
    port map (
      ADR0 => romo2addro10_s(2),
      ADR1 => romo2addro10_s(0),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1554
    );
  ix53675z23738 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => romo2addro10_s(0),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(2),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1545
    );
  ix53675z26799 : X_LUT4
    generic map(
      INIT => X"1C86"
    )
    port map (
      ADR0 => rome2addro6_s(3),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(1),
      ADR3 => rome2addro6_s(0),
      O => nx53675z421
    );
  ix53675z25718 : X_LUT4
    generic map(
      INIT => X"44D4"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(1),
      ADR3 => rome2addro6_s(2),
      O => nx53675z418
    );
  ix53675z12923 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => rome2addro6_s(3),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(1),
      ADR3 => rome2addro6_s(0),
      O => nx53675z423
    );
  ix53675z30879 : X_LUT4
    generic map(
      INIT => X"4F04"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(1),
      ADR3 => rome2addro6_s(2),
      O => nx53675z415
    );
  ix53675z26058 : X_LUT4
    generic map(
      INIT => X"6868"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => VCC,
      O => nx53675z1092
    );
  ix53675z24734 : X_LUT4
    generic map(
      INIT => X"249A"
    )
    port map (
      ADR0 => rome2addro6_s(3),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(1),
      ADR3 => rome2addro6_s(0),
      O => nx53675z424
    );
  ix53675z12483 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(3),
      ADR3 => rome2addro6_s(0),
      O => nx53675z429
    );
  ix53675z7924 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => rome2addro6_s(3),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(1),
      ADR3 => rome2addro6_s(0),
      O => nx53675z420
    );
  ix53675z61716 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(3),
      ADR3 => rome2addro6_s(0),
      O => nx53675z426
    );
  ix53675z14388 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(3),
      ADR3 => rome2addro6_s(0),
      O => nx53675z430
    );
  ix53675z64961 : X_LUT4
    generic map(
      INIT => X"CF0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(1),
      ADR3 => romo2addro3_s(3),
      O => nx53675z984
    );
  ix53675z25898 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => romo2addro3_s(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1027
    );
  ix53675z23224 : X_LUT4
    generic map(
      INIT => X"442A"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(1),
      ADR3 => romo2addro3_s(3),
      O => nx53675z981
    );
  ix53675z30441 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romo2addro3_s(0),
      O => nx53675z1028
    );
  ix53675z6845 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(3),
      ADR3 => VCC,
      O => U2_ROMO3_modgen_rom_ix0_nx_rm64_16_u
    );
  ix53675z16026 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => VCC,
      ADR2 => romo2addro3_s(3),
      ADR3 => VCC,
      O => U2_ROMO3_modgen_rom_ix0_nx_rm64_16_l
    );
  ix53675z41614 : X_LUT4
    generic map(
      INIT => X"C338"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(3),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(1),
      O => nx53675z910
    );
  ix53675z58295 : X_LUT4
    generic map(
      INIT => X"E81E"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(3),
      ADR2 => romo2addro2_s(0),
      ADR3 => romo2addro2_s(1),
      O => nx53675z907
    );
  ix53675z4186 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => rome2addro7_s(0),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z456
    );
  ix53675z18933 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(0),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(3),
      O => nx53675z405
    );
  ix53675z8197 : X_LUT4
    generic map(
      INIT => X"18C6"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(0),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(3),
      O => nx53675z403
    );
  ix53675z21619 : X_LUT4
    generic map(
      INIT => X"2B22"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(0),
      ADR3 => rome2addro6_s(3),
      O => nx53675z409
    );
  ix53675z15348 : X_LUT4
    generic map(
      INIT => X"5294"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(0),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(3),
      O => nx53675z406
    );
  ix53675z12459 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(0),
      ADR3 => rome2addro6_s(3),
      O => nx53675z411
    );
  ix53675z7622 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(0),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(3),
      O => nx53675z402
    );
  ix53675z4120 : X_LUT4
    generic map(
      INIT => X"20F2"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(0),
      ADR3 => rome2addro6_s(3),
      O => nx53675z412
    );
  ix53675z34940 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(0),
      ADR3 => rome2addro6_s(3),
      O => nx53675z408
    );
  ix53675z18949 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(1),
      ADR3 => rome2addro6_s(2),
      O => nx53675z417
    );
  ix53675z40406 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(1),
      ADR3 => rome2addro6_s(2),
      O => nx53675z414
    );
  ix53675z29603 : X_LUT4
    generic map(
      INIT => X"639C"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z925
    );
  ix53675z10785 : X_LUT4
    generic map(
      INIT => X"5A78"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z929
    );
  ix53675z29635 : X_LUT4
    generic map(
      INIT => X"0CF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(0),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1530
    );
  ix53675z25782 : X_LUT4
    generic map(
      INIT => X"666A"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => romo2addro2_s(3),
      ADR3 => romo2addro2_s(1),
      O => nx53675z926
    );
  ix53675z52894 : X_LUT4
    generic map(
      INIT => X"BB22"
    )
    port map (
      ADR0 => romo2addro10_s(2),
      ADR1 => romo2addro10_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro10_s(1),
      O => nx53675z1531
    );
  ix53675z12269 : X_LUT4
    generic map(
      INIT => X"1188"
    )
    port map (
      ADR0 => romo2addro10_s(0),
      ADR1 => romo2addro10_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro10_s(1),
      O => nx53675z1536
    );
  ix53675z24310 : X_LUT4
    generic map(
      INIT => X"1A0E"
    )
    port map (
      ADR0 => romo2addro10_s(2),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(0),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1527
    );
  ix53675z7545 : X_LUT4
    generic map(
      INIT => X"7656"
    )
    port map (
      ADR0 => romo2addro10_s(2),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(0),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1528
    );
  ix53675z6376 : X_LUT4
    generic map(
      INIT => X"180E"
    )
    port map (
      ADR0 => romo2addro10_s(0),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(2),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1533
    );
  ix53675z26706 : X_LUT4
    generic map(
      INIT => X"492C"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => rome2addro5_s(2),
      ADR2 => rome2addro5_s(1),
      ADR3 => rome2addro5_s(3),
      O => nx53675z356
    );
  ix53675z25646 : X_LUT4
    generic map(
      INIT => X"08AE"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(1),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z368
    );
  ix53675z61623 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(1),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z361
    );
  ix53675z14295 : X_LUT4
    generic map(
      INIT => X"7130"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(1),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z365
    );
  ix53675z18880 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(1),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z370
    );
  ix53675z4048 : X_LUT4
    generic map(
      INIT => X"5D04"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(1),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z362
    );
  ix53675z5051 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(1),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z371
    );
  ix53675z35033 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(3),
      ADR3 => rome2addro7_s(0),
      O => nx53675z473
    );
  ix53675z12552 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(3),
      ADR3 => rome2addro7_s(0),
      O => nx53675z476
    );
  ix53675z34321 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(1),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z367
    );
  ix53675z2272 : X_LUT4
    generic map(
      INIT => X"FEFE"
    )
    port map (
      ADR0 => romo2addro1_s(0),
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(2),
      ADR3 => VCC,
      O => nx53675z862
    );
  ix53675z2509 : X_LUT4
    generic map(
      INIT => X"FEFE"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(0),
      ADR3 => VCC,
      O => nx53675z859
    );
  ix53675z4067 : X_LUT4
    generic map(
      INIT => X"5656"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => romo2addro1_s(0),
      ADR2 => romo2addro1_s(2),
      ADR3 => VCC,
      O => nx53675z867
    );
  ix53675z10248 : X_LUT4
    generic map(
      INIT => X"0F3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro1_s(0),
      ADR2 => romo2addro1_s(2),
      ADR3 => romo2addro1_s(1),
      O => nx53675z868
    );
  ix53675z54818 : X_LUT4
    generic map(
      INIT => X"CF30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro1_s(3),
      ADR2 => romo2addro1_s(2),
      ADR3 => romo2addro1_s(1),
      O => nx53675z864
    );
  ix53675z24397 : X_LUT4
    generic map(
      INIT => X"3366"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => romo2addro1_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro1_s(1),
      O => nx53675z865
    );
  ix53675z18562 : X_LUT4
    generic map(
      INIT => X"7110"
    )
    port map (
      ADR0 => rome2addro7_s(0),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z458
    );
  ix53675z14433 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => rome2addro7_s(0),
      ADR1 => rome2addro7_s(3),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z459
    );
  ix53675z4141 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(3),
      ADR3 => rome2addro6_s(0),
      O => nx53675z427
    );
  ix53675z6887 : X_LUT4
    generic map(
      INIT => X"44AA"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro4_s(2),
      O => nx53675z1089
    );
  ix53675z41923 : X_LUT4
    generic map(
      INIT => X"F00A"
    )
    port map (
      ADR0 => romo2addro4_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1093
    );
  ix53675z55114 : X_LUT4
    generic map(
      INIT => X"AA50"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1090
    );
  ix53675z4405 : X_LUT4
    generic map(
      INIT => X"05FA"
    )
    port map (
      ADR0 => romo2addro4_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1104
    );
  ix53675z10586 : X_LUT4
    generic map(
      INIT => X"11EE"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro4_s(2),
      O => nx53675z1105
    );
  ix53675z55155 : X_LUT4
    generic map(
      INIT => X"AA5A"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1101
    );
  ix53675z26295 : X_LUT4
    generic map(
      INIT => X"3366"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro4_s(3),
      O => nx53675z1102
    );
  ix53675z11815 : X_LUT4
    generic map(
      INIT => X"0A50"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1220
    );
  ix53675z31065 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z545
    );
  ix53675z35126 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => rome2addro8_s(3),
      ADR1 => rome2addro8_s(1),
      ADR2 => rome2addro8_s(0),
      ADR3 => rome2addro8_s(2),
      O => nx53675z538
    );
  ix53675z4306 : X_LUT4
    generic map(
      INIT => X"50D4"
    )
    port map (
      ADR0 => rome2addro8_s(3),
      ADR1 => rome2addro8_s(1),
      ADR2 => rome2addro8_s(0),
      ADR3 => rome2addro8_s(2),
      O => nx53675z542
    );
  ix53675z19135 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z547
    );
  ix53675z21805 : X_LUT4
    generic map(
      INIT => X"08CE"
    )
    port map (
      ADR0 => rome2addro8_s(3),
      ADR1 => rome2addro8_s(1),
      ADR2 => rome2addro8_s(0),
      ADR3 => rome2addro8_s(2),
      O => nx53675z539
    );
  ix53675z25904 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z548
    );
  ix53675z18283 : X_LUT4
    generic map(
      INIT => X"4D04"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(1),
      ADR2 => rome2addro4_s(3),
      ADR3 => rome2addro4_s(2),
      O => nx53675z263
    );
  ix53675z40592 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z544
    );
  ix53675z65188 : X_LUT4
    generic map(
      INIT => X"AF0A"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1142
    );
  ix53675z3229 : X_LUT4
    generic map(
      INIT => X"3322"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => romo2addro5_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro5_s(2),
      O => nx53675z1177
    );
  ix53675z23451 : X_LUT4
    generic map(
      INIT => X"2644"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => romo2addro5_s(0),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1139
    );
  ix53675z3024 : X_LUT4
    generic map(
      INIT => X"0300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro5_s(3),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1174
    );
  ix53675z2722 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1178
    );
  ix53675z2959 : X_LUT4
    generic map(
      INIT => X"FEFE"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => romo2addro5_s(3),
      ADR2 => romo2addro5_s(1),
      ADR3 => VCC,
      O => nx53675z1175
    );
  ix53675z4517 : X_LUT4
    generic map(
      INIT => X"0F5A"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro5_s(3),
      ADR3 => romo2addro5_s(0),
      O => nx53675z1183
    );
  ix53675z10698 : X_LUT4
    generic map(
      INIT => X"5566"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro5_s(0),
      O => nx53675z1184
    );
  ix53675z55268 : X_LUT4
    generic map(
      INIT => X"C6C6"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(3),
      ADR3 => VCC,
      O => nx53675z1180
    );
  ix53675z24847 : X_LUT4
    generic map(
      INIT => X"11EE"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => romo2addro5_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro5_s(0),
      O => nx53675z1181
    );
  ix53675z26233 : X_LUT4
    generic map(
      INIT => X"57A8"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(3),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1242
    );
  ix53675z7112 : X_LUT4
    generic map(
      INIT => X"6464"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(3),
      ADR2 => romo2addro6_s(1),
      ADR3 => VCC,
      O => nx53675z1247
    );
  ix53675z42148 : X_LUT4
    generic map(
      INIT => X"A4A4"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(2),
      ADR2 => romo2addro6_s(1),
      ADR3 => VCC,
      O => nx53675z1251
    );
  ix53675z55339 : X_LUT4
    generic map(
      INIT => X"C2C2"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(3),
      ADR2 => romo2addro6_s(1),
      ADR3 => VCC,
      O => nx53675z1248
    );
  ix53675z3341 : X_LUT4
    generic map(
      INIT => X"3322"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro6_s(0),
      O => nx53675z1256
    );
  ix53675z2834 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(0),
      O => nx53675z1257
    );
  ix53675z3136 : X_LUT4
    generic map(
      INIT => X"0202"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(3),
      ADR2 => romo2addro6_s(1),
      ADR3 => VCC,
      O => nx53675z1253
    );
  ix53675z3071 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro6_s(3),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(0),
      O => nx53675z1254
    );
  ix53675z59525 : X_LUT4
    generic map(
      INIT => X"F50A"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1129
    );
  ix53675z55252 : X_LUT4
    generic map(
      INIT => X"FF54"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1030
    );
  ix53675z20594 : X_LUT4
    generic map(
      INIT => X"294A"
    )
    port map (
      ADR0 => romo2addro10_s(2),
      ADR1 => romo2addro10_s(0),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1551
    );
  ix53675z37928 : X_LUT4
    generic map(
      INIT => X"934C"
    )
    port map (
      ADR0 => romo2addro10_s(2),
      ADR1 => romo2addro10_s(0),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1555
    );
  ix53675z23368 : X_LUT4
    generic map(
      INIT => X"0C4C"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1032
    );
  ix53675z29051 : X_LUT4
    generic map(
      INIT => X"2DDA"
    )
    port map (
      ADR0 => romo2addro10_s(2),
      ADR1 => romo2addro10_s(0),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(1),
      O => nx53675z1552
    );
  ix53675z48531 : X_LUT4
    generic map(
      INIT => X"D0FC"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1033
    );
  ix53675z2779 : X_LUT4
    generic map(
      INIT => X"5550"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro1_s(0),
      ADR3 => romo2addro1_s(2),
      O => nx53675z861
    );
  ix53675z2574 : X_LUT4
    generic map(
      INIT => X"1010"
    )
    port map (
      ADR0 => romo2addro1_s(3),
      ADR1 => romo2addro1_s(1),
      ADR2 => romo2addro1_s(2),
      ADR3 => VCC,
      O => nx53675z858
    );
  ix53675z42065 : X_LUT4
    generic map(
      INIT => X"9694"
    )
    port map (
      ADR0 => romo2addro6_s(3),
      ADR1 => romo2addro6_s(0),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1226
    );
  ix53675z65300 : X_LUT4
    generic map(
      INIT => X"AF0A"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1221
    );
  ix53675z23563 : X_LUT4
    generic map(
      INIT => X"502A"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(2),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1218
    );
  ix53675z45395 : X_LUT4
    generic map(
      INIT => X"9C66"
    )
    port map (
      ADR0 => romo2addro6_s(3),
      ADR1 => romo2addro6_s(0),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1224
    );
  ix53675z53032 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => romo2addro6_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1227
    );
  ix53675z23482 : X_LUT4
    generic map(
      INIT => X"3700"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => romo2addro5_s(0),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1111
    );
  ix53675z58746 : X_LUT4
    generic map(
      INIT => X"E386"
    )
    port map (
      ADR0 => romo2addro6_s(3),
      ADR1 => romo2addro6_s(0),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1223
    );
  ix53675z55366 : X_LUT4
    generic map(
      INIT => X"F5F4"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => romo2addro5_s(0),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1109
    );
  ix53675z55478 : X_LUT4
    generic map(
      INIT => X"F5F4"
    )
    port map (
      ADR0 => romo2addro6_s(3),
      ADR1 => romo2addro6_s(0),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1188
    );
  ix53675z57847 : X_LUT4
    generic map(
      INIT => X"A5F0"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro9_s(1),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1496
    );
  ix53675z11152 : X_LUT4
    generic map(
      INIT => X"03FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro9_s(0),
      ADR2 => romo2addro9_s(1),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1500
    );
  ix53675z25301 : X_LUT4
    generic map(
      INIT => X"05FA"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro9_s(1),
      ADR3 => romo2addro9_s(0),
      O => nx53675z1497
    );
  ix53675z23594 : X_LUT4
    generic map(
      INIT => X"3700"
    )
    port map (
      ADR0 => romo2addro6_s(3),
      ADR1 => romo2addro6_s(0),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1190
    );
  ix53675z48757 : X_LUT4
    generic map(
      INIT => X"CF4C"
    )
    port map (
      ADR0 => romo2addro6_s(3),
      ADR1 => romo2addro6_s(0),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1191
    );
  ix53675z44435 : X_LUT4
    generic map(
      INIT => X"8988"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(2),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1232
    );
  ix53675z23284 : X_LUT4
    generic map(
      INIT => X"7310"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(2),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1229
    );
  ix53675z14154 : X_LUT4
    generic map(
      INIT => X"3B02"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(1),
      ADR2 => rome2addro4_s(3),
      ADR3 => rome2addro4_s(2),
      O => nx53675z264
    );
  ix53675z3907 : X_LUT4
    generic map(
      INIT => X"0A8E"
    )
    port map (
      ADR0 => rome2addro4_s(0),
      ADR1 => rome2addro4_s(1),
      ADR2 => rome2addro4_s(3),
      ADR3 => rome2addro4_s(2),
      O => nx53675z261
    );
  ix53675z4279 : X_LUT4
    generic map(
      INIT => X"0C8E"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z521
    );
  ix53675z18655 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z523
    );
  ix53675z14526 : X_LUT4
    generic map(
      INIT => X"5D04"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z524
    );
  ix53675z12390 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => rome2addro5_s(3),
      ADR1 => rome2addro5_s(1),
      ADR2 => rome2addro5_s(2),
      ADR3 => rome2addro5_s(0),
      O => nx53675z364
    );
  ix53675z12830 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => rome2addro5_s(2),
      ADR2 => rome2addro5_s(1),
      ADR3 => rome2addro5_s(3),
      O => nx53675z358
    );
  ix53675z7831 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => rome2addro5_s(2),
      ADR2 => rome2addro5_s(1),
      ADR3 => rome2addro5_s(3),
      O => nx53675z355
    );
  ix53675z24641 : X_LUT4
    generic map(
      INIT => X"6518"
    )
    port map (
      ADR0 => rome2addro5_s(0),
      ADR1 => rome2addro5_s(2),
      ADR2 => rome2addro5_s(1),
      ADR3 => rome2addro5_s(3),
      O => nx53675z359
    );
  ix53675z14011 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(2),
      O => nx53675z258
    );
  ix53675z59411 : X_LUT4
    generic map(
      INIT => X"AA5A"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1050
    );
  ix53675z1842 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => rome2addro3_s(3),
      ADR3 => rome2addro3_s(0),
      O => nx53675z255
    );
  ix53675z43145 : X_LUT4
    generic map(
      INIT => X"CF32"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(0),
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1047
    );
  ix53675z15102 : X_LUT4
    generic map(
      INIT => X"05A0"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1051
    );
  ix53675z44096 : X_LUT4
    generic map(
      INIT => X"C1C0"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => romo2addro3_s(0),
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(3),
      O => nx53675z995
    );
  ix53675z24638 : X_LUT4
    generic map(
      INIT => X"00FA"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(0),
      O => nx53675z1048
    );
  ix53675z22945 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => romo2addro3_s(0),
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(3),
      O => nx53675z992
    );
  ix53675z38606 : X_LUT4
    generic map(
      INIT => X"8A50"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => romo2addro3_s(0),
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(3),
      O => nx53675z993
    );
  ix53675z62249 : X_LUT4
    generic map(
      INIT => X"E888"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => romo2addro3_s(0),
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(3),
      O => nx53675z996
    );
  ix53675z40572 : X_LUT4
    generic map(
      INIT => X"D52A"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(1),
      O => nx53675z1007
    );
  ix53675z11124 : X_LUT4
    generic map(
      INIT => X"5A78"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(3),
      ADR3 => romo2addro5_s(0),
      O => nx53675z1166
    );
  ix53675z26171 : X_LUT4
    generic map(
      INIT => X"6688"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => romo2addro5_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro5_s(2),
      O => nx53675z1171
    );
  ix53675z26121 : X_LUT4
    generic map(
      INIT => X"56AA"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(3),
      ADR3 => romo2addro5_s(0),
      O => nx53675z1163
    );
  ix53675z42036 : X_LUT4
    generic map(
      INIT => X"A5A0"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1172
    );
  ix53675z7000 : X_LUT4
    generic map(
      INIT => X"33C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro5_s(2),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1168
    );
  ix53675z55227 : X_LUT4
    generic map(
      INIT => X"F00A"
    )
    port map (
      ADR0 => romo2addro5_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1169
    );
  ix53675z26013 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(0),
      O => nx53675z1106
    );
  ix53675z6960 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(3),
      O => U2_ROMO4_modgen_rom_ix0_nx_rm64_16_u
    );
  ix53675z25832 : X_LUT4
    generic map(
      INIT => X"0A8E"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(2),
      O => nx53675z498
    );
  ix53675z61809 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(0),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z491
    );
  ix53675z14481 : X_LUT4
    generic map(
      INIT => X"4F04"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(0),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z495
    );
  ix53675z19066 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(2),
      O => nx53675z500
    );
  ix53675z4234 : X_LUT4
    generic map(
      INIT => X"44D4"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(0),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z492
    );
  ix53675z5237 : X_LUT4
    generic map(
      INIT => X"40DC"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(2),
      O => nx53675z501
    );
  ix53675z23943 : X_LUT4
    generic map(
      INIT => X"1F00"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1433
    );
  ix53675z34507 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(0),
      ADR3 => rome2addro7_s(2),
      O => nx53675z497
    );
  ix53675z60691 : X_LUT4
    generic map(
      INIT => X"C800"
    )
    port map (
      ADR0 => romo2addro9_s(1),
      ADR1 => romo2addro9_s(3),
      ADR2 => romo2addro9_s(0),
      ADR3 => romo2addro9_s(2),
      O => nx53675z1430
    );
  ix53675z18670 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(0),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(2),
      O => nx53675z222
    );
  ix53675z24476 : X_LUT4
    generic map(
      INIT => X"249A"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z244
    );
  ix53675z40127 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(0),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(2),
      O => nx53675z219
    );
  ix53675z25439 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(0),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(2),
      O => nx53675z223
    );
  ix53675z12220 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z246
    );
  ix53675z30600 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(0),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(2),
      O => nx53675z220
    );
  ix53675z8961 : X_LUT4
    generic map(
      INIT => X"6138"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z247
    );
  ix53675z28704 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro3_s(1),
      ADR1 => rome2addro3_s(0),
      ADR2 => rome2addro3_s(3),
      ADR3 => rome2addro3_s(2),
      O => nx53675z257
    );
  ix53675z61453 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(2),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(0),
      O => nx53675z243
    );
  ix53675z28701 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro3_s(3),
      ADR1 => rome2addro3_s(0),
      ADR2 => rome2addro3_s(1),
      ADR3 => rome2addro3_s(2),
      O => U2_ROME3_modgen_rom_ix2_nx_rm64_16_u
    );
  ix53675z26687 : X_LUT4
    generic map(
      INIT => X"1FE0"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(0),
      ADR3 => romo2addro10_s(2),
      O => nx53675z1558
    );
  ix53675z29715 : X_LUT4
    generic map(
      INIT => X"2DD2"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(1),
      O => nx53675z1004
    );
  ix53675z10897 : X_LUT4
    generic map(
      INIT => X"666A"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(1),
      O => nx53675z1008
    );
  ix53675z41365 : X_LUT4
    generic map(
      INIT => X"A666"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(0),
      ADR3 => romo2addro10_s(2),
      O => nx53675z1560
    );
  ix53675z25894 : X_LUT4
    generic map(
      INIT => X"3C6C"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(1),
      O => nx53675z1005
    );
  ix53675z11690 : X_LUT4
    generic map(
      INIT => X"36CC"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(0),
      ADR3 => romo2addro10_s(2),
      O => nx53675z1561
    );
  ix53675z26737 : X_LUT4
    generic map(
      INIT => X"6688"
    )
    port map (
      ADR0 => romo2addro10_s(3),
      ADR1 => romo2addro10_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro10_s(2),
      O => nx53675z1566
    );
  ix53675z30508 : X_LUT4
    generic map(
      INIT => X"5A96"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(0),
      ADR3 => romo2addro10_s(2),
      O => nx53675z1557
    );
  ix53675z7566 : X_LUT4
    generic map(
      INIT => X"22CC"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro10_s(2),
      O => nx53675z1563
    );
  ix53675z4213 : X_LUT4
    generic map(
      INIT => X"4F04"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(3),
      ADR3 => rome2addro7_s(0),
      O => nx53675z477
    );
  ix53675z19042 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(0),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z482
    );
  ix53675z21712 : X_LUT4
    generic map(
      INIT => X"44D4"
    )
    port map (
      ADR0 => rome2addro7_s(2),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(3),
      ADR3 => rome2addro7_s(0),
      O => nx53675z474
    );
  ix53675z30972 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(0),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z480
    );
  ix53675z25811 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(0),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z483
    );
  ix53675z13016 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(2),
      ADR3 => rome2addro7_s(0),
      O => nx53675z488
    );
  ix53675z40499 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(0),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z479
    );
  ix53675z8017 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(2),
      ADR3 => rome2addro7_s(0),
      O => nx53675z485
    );
  ix53675z26892 : X_LUT4
    generic map(
      INIT => X"3492"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(2),
      ADR3 => rome2addro7_s(0),
      O => nx53675z486
    );
  ix53675z24827 : X_LUT4
    generic map(
      INIT => X"18A6"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(1),
      ADR2 => rome2addro7_s(2),
      ADR3 => rome2addro7_s(0),
      O => nx53675z489
    );
  ix53675z12576 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => rome2addro7_s(3),
      ADR1 => rome2addro7_s(0),
      ADR2 => rome2addro7_s(1),
      ADR3 => rome2addro7_s(2),
      O => nx53675z494
    );
  ix54672z54628 : X_LUT4
    generic map(
      INIT => X"F5F4"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(2),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(0),
      O => nx54672z586
    );
  ix54672z39852 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(0),
      O => nx54672z25
    );
  ix54672z25164 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(0),
      O => nx54672z29
    );
  ix54672z22744 : X_LUT4
    generic map(
      INIT => X"04CC"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(2),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(0),
      O => nx54672z588
    );
  ix54672z30325 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(0),
      O => nx54672z26
    );
  ix54672z47907 : X_LUT4
    generic map(
      INIT => X"DF0C"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(2),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(0),
      O => nx54672z589
    );
  ix53675z2307 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => VCC,
      O => nx53675z580
    );
  ix53675z7185 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROMO6_modgen_rom_ix0_nx_rm64_16_u
    );
  ix53675z57907 : X_LUT4
    generic map(
      INIT => X"A5A6"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1516
    );
  ix53675z29323 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1265
    );
  ix53675z16366 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2addro6_s(3),
      ADR1 => romo2addro6_s(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROMO6_modgen_rom_ix0_nx_rm64_16_l
    );
  ix53675z26633 : X_LUT4
    generic map(
      INIT => X"36CC"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1518
    );
  ix53675z42028 : X_LUT4
    generic map(
      INIT => X"9B64"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1519
    );
  ix53675z11373 : X_LUT4
    generic map(
      INIT => X"3C68"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(2),
      ADR2 => romo2addro10_s(3),
      ADR3 => romo2addro10_s(0),
      O => nx53675z1515
    );
  ix53675z23707 : X_LUT4
    generic map(
      INIT => X"1F00"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(3),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1269
    );
  ix53675z23337 : X_LUT4
    generic map(
      INIT => X"224C"
    )
    port map (
      ADR0 => romo2addro4_s(2),
      ADR1 => romo2addro4_s(0),
      ADR2 => romo2addro4_s(1),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1060
    );
  ix53675z38719 : X_LUT4
    generic map(
      INIT => X"A244"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1072
    );
  ix53675z58520 : X_LUT4
    generic map(
      INIT => X"B994"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(0),
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1065
    );
  ix53675z45169 : X_LUT4
    generic map(
      INIT => X"C36C"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(0),
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1066
    );
  ix53675z52806 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1069
    );
  ix53675z44209 : X_LUT4
    generic map(
      INIT => X"C0C2"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1074
    );
  ix53675z62362 : X_LUT4
    generic map(
      INIT => X"F880"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1075
    );
  ix53675z34414 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(3),
      ADR3 => rome2addro6_s(0),
      O => nx53675z432
    );
  ix53675z18973 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(3),
      ADR3 => rome2addro6_s(0),
      O => nx53675z435
    );
  ix53675z23058 : X_LUT4
    generic map(
      INIT => X"2B22"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(2),
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1071
    );
  ix53675z42602 : X_LUT4
    generic map(
      INIT => X"9988"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro10_s(2),
      O => nx53675z1567
    );
  ix53675z55793 : X_LUT4
    generic map(
      INIT => X"9898"
    )
    port map (
      ADR0 => romo2addro10_s(1),
      ADR1 => romo2addro10_s(3),
      ADR2 => romo2addro10_s(0),
      ADR3 => VCC,
      O => nx53675z1564
    );
  ix53675z28955 : X_LUT4
    generic map(
      INIT => X"0AF0"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(0),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1056
    );
  ix53675z52214 : X_LUT4
    generic map(
      INIT => X"F550"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1057
    );
  ix53675z11589 : X_LUT4
    generic map(
      INIT => X"4422"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro4_s(3),
      O => nx53675z1062
    );
  ix53675z23630 : X_LUT4
    generic map(
      INIT => X"3432"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(0),
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1053
    );
  ix53675z6865 : X_LUT4
    generic map(
      INIT => X"5E1E"
    )
    port map (
      ADR0 => romo2addro4_s(3),
      ADR1 => romo2addro4_s(0),
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(1),
      O => nx53675z1054
    );
  ix53675z5696 : X_LUT4
    generic map(
      INIT => X"4524"
    )
    port map (
      ADR0 => romo2addro4_s(2),
      ADR1 => romo2addro4_s(0),
      ADR2 => romo2addro4_s(1),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1059
    );
  ix53675z41839 : X_LUT4
    generic map(
      INIT => X"9866"
    )
    port map (
      ADR0 => romo2addro4_s(1),
      ADR1 => romo2addro4_s(0),
      ADR2 => romo2addro4_s(2),
      ADR3 => romo2addro4_s(3),
      O => nx53675z1068
    );
  ix53675z65074 : X_LUT4
    generic map(
      INIT => X"BB22"
    )
    port map (
      ADR0 => romo2addro4_s(2),
      ADR1 => romo2addro4_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro4_s(3),
      O => nx53675z1063
    );
  ix53675z26125 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romo2addro5_s(0),
      O => nx53675z1185
    );
  ix53675z7072 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro5_s(3),
      ADR3 => VCC,
      O => U2_ROMO5_modgen_rom_ix0_nx_rm64_16_u
    );
  ix53675z54956 : X_LUT4
    generic map(
      INIT => X"A5B4"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(1),
      ADR3 => romo2addro3_s(0),
      O => nx53675z963
    );
  ix53675z29210 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro5_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro5_s(0),
      O => nx53675z1186
    );
  ix53675z16253 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(3),
      ADR3 => VCC,
      O => U2_ROMO5_modgen_rom_ix0_nx_rm64_16_l
    );
  ix53675z25840 : X_LUT4
    generic map(
      INIT => X"36CC"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(1),
      ADR3 => romo2addro3_s(0),
      O => nx53675z965
    );
  ix53675z41235 : X_LUT4
    generic map(
      INIT => X"D32C"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(1),
      ADR3 => romo2addro3_s(0),
      O => nx53675z966
    );
  ix53675z27153 : X_LUT4
    generic map(
      INIT => X"6688"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(3),
      O => nx53675z934
    );
  ix53675z10581 : X_LUT4
    generic map(
      INIT => X"6668"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(1),
      ADR3 => romo2addro3_s(0),
      O => nx53675z962
    );
  ix53675z6661 : X_LUT4
    generic map(
      INIT => X"5588"
    )
    port map (
      ADR0 => romo2addro2_s(2),
      ADR1 => romo2addro2_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(3),
      O => nx53675z931
    );
  ix53675z5144 : X_LUT4
    generic map(
      INIT => X"2B22"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(3),
      ADR3 => rome2addro6_s(0),
      O => nx53675z436
    );
  ix53675z12499 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => nx53675z441
    );
  ix53675z25739 : X_LUT4
    generic map(
      INIT => X"20F2"
    )
    port map (
      ADR0 => rome2addro6_s(1),
      ADR1 => rome2addro6_s(2),
      ADR2 => rome2addro6_s(3),
      ADR3 => rome2addro6_s(0),
      O => nx53675z433
    );
  ix53675z24755 : X_LUT4
    generic map(
      INIT => X"4964"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => nx53675z439
    );
  ix53675z9240 : X_LUT4
    generic map(
      INIT => X"2D42"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => nx53675z442
    );
  ix53675z26067 : X_LUT4
    generic map(
      INIT => X"666A"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(0),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1123
    );
  ix53675z61732 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro6_s(0),
      ADR1 => rome2addro6_s(3),
      ADR2 => rome2addro6_s(2),
      ADR3 => rome2addro6_s(1),
      O => nx53675z438
    );
  ix53675z10807 : X_LUT4
    generic map(
      INIT => X"56A8"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(0),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1120
    );
  ix53675z56775 : X_LUT4
    generic map(
      INIT => X"F01E"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(0),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1121
    );
  ix53675z41462 : X_LUT4
    generic map(
      INIT => X"96C6"
    )
    port map (
      ADR0 => romo2addro5_s(2),
      ADR1 => romo2addro5_s(0),
      ADR2 => romo2addro5_s(1),
      ADR3 => romo2addro5_s(3),
      O => nx53675z1124
    );
  ix53675z4971 : X_LUT4
    generic map(
      INIT => X"5566"
    )
    port map (
      ADR0 => romo2addro9_s(3),
      ADR1 => romo2addro9_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro9_s(2),
      O => nx53675z1499
    );
  ix53675z41698 : X_LUT4
    generic map(
      INIT => X"9988"
    )
    port map (
      ADR0 => romo2addro2_s(1),
      ADR1 => romo2addro2_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(2),
      O => nx53675z935
    );
  ix53675z26985 : X_LUT4
    generic map(
      INIT => X"249A"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(1),
      O => nx53675z551
    );
  ix53675z54888 : X_LUT4
    generic map(
      INIT => X"AA44"
    )
    port map (
      ADR0 => romo2addro2_s(1),
      ADR1 => romo2addro2_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro2_s(3),
      O => nx53675z932
    );
  ix53675z13109 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(1),
      O => nx53675z553
    );
  ix53675z24920 : X_LUT4
    generic map(
      INIT => X"6138"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(1),
      O => nx53675z554
    );
  ix53675z12669 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => rome2addro8_s(0),
      ADR1 => rome2addro8_s(1),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z559
    );
  ix53675z8110 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(1),
      O => nx53675z550
    );
  ix53675z61902 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro8_s(0),
      ADR1 => rome2addro8_s(1),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z556
    );
  ix53675z14574 : X_LUT4
    generic map(
      INIT => X"3B02"
    )
    port map (
      ADR0 => rome2addro8_s(0),
      ADR1 => rome2addro8_s(1),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z560
    );
  ix53675z17546 : X_LUT4
    generic map(
      INIT => X"59A6"
    )
    port map (
      ADR0 => rome2addro7_s(1),
      ADR1 => rome2addro7_s(0),
      ADR2 => rome2addro7_s(3),
      ADR3 => rome2addro7_s(2),
      O => nx53675z510
    );
  ix53675z55599 : X_LUT4
    generic map(
      INIT => X"CCFE"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(1),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(3),
      O => nx53675z1273
    );
  ix53675z60351 : X_LUT4
    generic map(
      INIT => X"A800"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(0),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1193
    );
  ix53675z48766 : X_LUT4
    generic map(
      INIT => X"8ECE"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(0),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1197
    );
  ix53675z23715 : X_LUT4
    generic map(
      INIT => X"0A2A"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(1),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(3),
      O => nx53675z1275
    );
  ix53675z57183 : X_LUT4
    generic map(
      INIT => X"F0FE"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(0),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(3),
      O => nx53675z1194
    );
  ix53675z48878 : X_LUT4
    generic map(
      INIT => X"B2F2"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(1),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(3),
      O => nx53675z1276
    );
  ix53675z26291 : X_LUT4
    generic map(
      INIT => X"37C8"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(3),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1281
    );
  ix53675z60464 : X_LUT4
    generic map(
      INIT => X"A800"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(1),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(3),
      O => nx53675z1272
    );
  ix53675z11032 : X_LUT4
    generic map(
      INIT => X"1EE0"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(3),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1278
    );
  ix53675z45283 : X_LUT4
    generic map(
      INIT => X"B45A"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(0),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1145
    );
  ix53675z52920 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => romo2addro5_s(1),
      ADR2 => VCC,
      ADR3 => romo2addro5_s(2),
      O => nx53675z1148
    );
  ix53675z28842 : X_LUT4
    generic map(
      INIT => X"0AF0"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(1),
      O => nx53675z977
    );
  ix53675z52101 : X_LUT4
    generic map(
      INIT => X"F550"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => VCC,
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(1),
      O => nx53675z978
    );
  ix53675z29169 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro8_s(0),
      ADR1 => rome2addro8_s(1),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z582
    );
  ix53675z23517 : X_LUT4
    generic map(
      INIT => X"5158"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => romo2addro3_s(1),
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(3),
      O => nx53675z974
    );
  ix53675z6752 : X_LUT4
    generic map(
      INIT => X"0FDA"
    )
    port map (
      ADR0 => romo2addro3_s(0),
      ADR1 => romo2addro3_s(1),
      ADR2 => romo2addro3_s(2),
      ADR3 => romo2addro3_s(3),
      O => nx53675z975
    );
  ix53675z29166 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => rome2addro8_s(0),
      ADR1 => rome2addro8_s(1),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => U2_ROME8_modgen_rom_ix2_nx_rm64_16_u
    );
  ix53675z26238 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => VCC,
      ADR2 => romo2addro6_s(2),
      ADR3 => VCC,
      O => nx53675z1264
    );
  ix53675z14476 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2addro8_s(1),
      ADR2 => VCC,
      ADR3 => rome2addro8_s(2),
      O => nx53675z583
    );
  ix53675z41686 : X_LUT4
    generic map(
      INIT => X"996C"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(3),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1282
    );
  ix53675z29181 : X_LUT4
    generic map(
      INIT => X"33C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(3),
      ADR3 => romo2addro6_s(0),
      O => nx53675z1214
    );
  ix53675z26179 : X_LUT4
    generic map(
      INIT => X"1FE0"
    )
    port map (
      ADR0 => romo2addro6_s(3),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(0),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1202
    );
  ix53675z55407 : X_LUT4
    generic map(
      INIT => X"A5A6"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(3),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1279
    );
  ix53675z10920 : X_LUT4
    generic map(
      INIT => X"56A8"
    )
    port map (
      ADR0 => romo2addro6_s(3),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(0),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1199
    );
  ix53675z41574 : X_LUT4
    generic map(
      INIT => X"C378"
    )
    port map (
      ADR0 => romo2addro6_s(3),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(0),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1203
    );
  ix53675z59637 : X_LUT4
    generic map(
      INIT => X"C6C6"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(3),
      ADR2 => romo2addro6_s(1),
      ADR3 => VCC,
      O => nx53675z1208
    );
  ix53675z55295 : X_LUT4
    generic map(
      INIT => X"999C"
    )
    port map (
      ADR0 => romo2addro6_s(3),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(0),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1200
    );
  ix53675z15328 : X_LUT4
    generic map(
      INIT => X"1818"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(3),
      ADR2 => romo2addro6_s(1),
      ADR3 => VCC,
      O => nx53675z1209
    );
  ix53675z43372 : X_LUT4
    generic map(
      INIT => X"A5F4"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(3),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(2),
      O => nx53675z1205
    );
  ix53675z24865 : X_LUT4
    generic map(
      INIT => X"5454"
    )
    port map (
      ADR0 => romo2addro6_s(0),
      ADR1 => romo2addro6_s(3),
      ADR2 => romo2addro6_s(2),
      ADR3 => VCC,
      O => nx53675z1206
    );
  ix54672z26333 : X_LUT4
    generic map(
      INIT => X"5924"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z96
    );
  ix54672z54632 : X_LUT4
    generic map(
      INIT => X"F30C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro1_s(2),
      ADR2 => romoaddro1_s(3),
      ADR3 => romoaddro1_s(1),
      O => nx54672z734
    );
  ix54672z10062 : X_LUT4
    generic map(
      INIT => X"333C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro1_s(2),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(1),
      O => nx54672z738
    );
  ix54672z24211 : X_LUT4
    generic map(
      INIT => X"333C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(3),
      ADR3 => romoaddro1_s(1),
      O => nx54672z735
    );
  ix54672z12457 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z98
    );
  ix54672z12017 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z104
    );
  ix54672z24268 : X_LUT4
    generic map(
      INIT => X"1C86"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z99
    );
  ix54672z61250 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z101
    );
  ix53675z45056 : X_LUT4
    generic map(
      INIT => X"C378"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(3),
      O => nx53675z987
    );
  ix53675z52693 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => romo2addro3_s(2),
      ADR2 => VCC,
      ADR3 => romo2addro3_s(3),
      O => nx53675z990
    );
  ix53675z21506 : X_LUT4
    generic map(
      INIT => X"3C16"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(1),
      O => nx53675z1001
    );
  ix53675z19801 : X_LUT4
    generic map(
      INIT => X"4964"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(1),
      O => nx53675z998
    );
  ix53675z37135 : X_LUT4
    generic map(
      INIT => X"8770"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(1),
      O => nx53675z1002
    );
  ix54672z11905 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(0),
      ADR3 => romeaddro0_s(3),
      O => nx54672z22
    );
  ix53675z28258 : X_LUT4
    generic map(
      INIT => X"59E6"
    )
    port map (
      ADR0 => romo2addro3_s(3),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(1),
      O => nx53675z999
    );
  ix54672z18395 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(0),
      O => nx54672z28
    );
  ix54672z21065 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(0),
      ADR3 => romeaddro0_s(3),
      O => nx54672z20
    );
  ix54672z3566 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(0),
      ADR3 => romeaddro0_s(3),
      O => nx54672z23
    );
  ix53675z48870 : X_LUT4
    generic map(
      INIT => X"F570"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(3),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1270
    );
  ix53675z55591 : X_LUT4
    generic map(
      INIT => X"BBBA"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(3),
      ADR2 => romo2addro7_s(0),
      ADR3 => romo2addro7_s(2),
      O => nx53675z1267
    );
  ix53675z59749 : X_LUT4
    generic map(
      INIT => X"BB44"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro7_s(3),
      O => nx53675z1287
    );
  ix53675z15440 : X_LUT4
    generic map(
      INIT => X"05A0"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro7_s(3),
      ADR3 => romo2addro7_s(1),
      O => nx53675z1288
    );
  ix53675z41726 : X_LUT4
    generic map(
      INIT => X"A45A"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(3),
      O => nx53675z989
    );
  ix53675z43484 : X_LUT4
    generic map(
      INIT => X"9B9A"
    )
    port map (
      ADR0 => romo2addro7_s(1),
      ADR1 => romo2addro7_s(0),
      ADR2 => romo2addro7_s(2),
      ADR3 => romo2addro7_s(3),
      O => nx53675z1284
    );
  ix53675z24977 : X_LUT4
    generic map(
      INIT => X"3322"
    )
    port map (
      ADR0 => romo2addro7_s(2),
      ADR1 => romo2addro7_s(0),
      ADR2 => VCC,
      ADR3 => romo2addro7_s(3),
      O => nx53675z1285
    );
  ix53675z58407 : X_LUT4
    generic map(
      INIT => X"AD94"
    )
    port map (
      ADR0 => romo2addro3_s(1),
      ADR1 => romo2addro3_s(2),
      ADR2 => romo2addro3_s(0),
      ADR3 => romo2addro3_s(3),
      O => nx53675z986
    );
  ix54672z47915 : X_LUT4
    generic map(
      INIT => X"B2BA"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(3),
      O => nx54672z595
    );
  ix54672z28330 : X_LUT4
    generic map(
      INIT => X"6622"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro0_s(3),
      O => nx54672z612
    );
  ix54672z25328 : X_LUT4
    generic map(
      INIT => X"36CC"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(2),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(0),
      O => nx54672z600
    );
  ix54672z54636 : X_LUT4
    generic map(
      INIT => X"CCFE"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(3),
      O => nx54672z592
    );
  ix54672z10069 : X_LUT4
    generic map(
      INIT => X"6668"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(2),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(0),
      O => nx54672z597
    );
  ix54672z40723 : X_LUT4
    generic map(
      INIT => X"9D62"
    )
    port map (
      ADR0 => romoaddro0_s(2),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(3),
      ADR3 => romoaddro0_s(0),
      O => nx54672z601
    );
  ix54672z58786 : X_LUT4
    generic map(
      INIT => X"A5AA"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(0),
      O => nx54672z606
    );
  ix54672z54444 : X_LUT4
    generic map(
      INIT => X"A5B4"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(2),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(0),
      O => nx54672z598
    );
  ix54672z14477 : X_LUT4
    generic map(
      INIT => X"0A50"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(2),
      O => nx54672z607
    );
  ix54672z42521 : X_LUT4
    generic map(
      INIT => X"C3F2"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(0),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(2),
      O => nx54672z603
    );
  ix54672z24014 : X_LUT4
    generic map(
      INIT => X"3322"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro0_s(2),
      O => nx54672z604
    );
  ix53675z4327 : X_LUT4
    generic map(
      INIT => X"0A8E"
    )
    port map (
      ADR0 => rome2addro8_s(0),
      ADR1 => rome2addro8_s(1),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(2),
      O => nx53675z557
    );
  ix53675z24941 : X_LUT4
    generic map(
      INIT => X"1C86"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(3),
      ADR2 => rome2addro8_s(0),
      ADR3 => rome2addro8_s(2),
      O => nx53675z569
    );
  ix53675z19159 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(1),
      ADR3 => rome2addro8_s(3),
      O => nx53675z565
    );
  ix53675z34600 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(1),
      ADR3 => rome2addro8_s(3),
      O => nx53675z562
    );
  ix53675z5330 : X_LUT4
    generic map(
      INIT => X"50D4"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(1),
      ADR3 => rome2addro8_s(3),
      O => nx53675z566
    );
  ix53675z12685 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(3),
      ADR2 => rome2addro8_s(0),
      ADR3 => rome2addro8_s(2),
      O => nx53675z571
    );
  ix53675z25925 : X_LUT4
    generic map(
      INIT => X"7310"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(1),
      ADR3 => rome2addro8_s(3),
      O => nx53675z563
    );
  ix53675z9426 : X_LUT4
    generic map(
      INIT => X"249A"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(3),
      ADR2 => rome2addro8_s(0),
      ADR3 => rome2addro8_s(2),
      O => nx53675z572
    );
  ix53675z19239 : X_LUT4
    generic map(
      INIT => X"2B42"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(1),
      O => nx53675z577
    );
  ix53675z61918 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => rome2addro8_s(1),
      ADR1 => rome2addro8_s(3),
      ADR2 => rome2addro8_s(0),
      ADR3 => rome2addro8_s(2),
      O => nx53675z568
    );
  ix53675z34616 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => rome2addro8_s(2),
      ADR1 => rome2addro8_s(0),
      ADR2 => rome2addro8_s(3),
      ADR3 => rome2addro8_s(1),
      O => nx53675z574
    );
  ix54672z9959 : X_LUT4
    generic map(
      INIT => X"05FA"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(2),
      O => nx54672z661
    );
  ix54672z24108 : X_LUT4
    generic map(
      INIT => X"555A"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(3),
      O => nx54672z658
    );
  ix54672z12111 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(3),
      O => nx54672z169
    );
  ix54672z3769 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(3),
      O => nx54672z167
    );
  ix54672z14016 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(3),
      O => nx54672z170
    );
  ix54672z18601 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(2),
      O => nx54672z175
    );
  ix54672z61344 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(3),
      O => nx54672z166
    );
  ix54672z34042 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(2),
      O => nx54672z172
    );
  ix54672z25367 : X_LUT4
    generic map(
      INIT => X"0A8E"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(2),
      O => nx54672z173
    );
  ix54672z4772 : X_LUT4
    generic map(
      INIT => X"40DC"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(2),
      O => nx54672z176
    );
  ix54672z12127 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(2),
      O => nx54672z181
    );
  ix54672z48018 : X_LUT4
    generic map(
      INIT => X"B0FA"
    )
    port map (
      ADR0 => romoaddro1_s(2),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(1),
      O => nx54672z672
    );
  ix54672z10172 : X_LUT4
    generic map(
      INIT => X"1EE0"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(3),
      O => nx54672z674
    );
  ix54672z40826 : X_LUT4
    generic map(
      INIT => X"969C"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(3),
      O => nx54672z678
    );
  ix54672z2593 : X_LUT4
    generic map(
      INIT => X"00FA"
    )
    port map (
      ADR0 => romoaddro1_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(3),
      O => nx54672z731
    );
  ix54672z54547 : X_LUT4
    generic map(
      INIT => X"AA56"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(3),
      O => nx54672z675
    );
  ix54672z2086 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romoaddro1_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(1),
      O => nx54672z732
    );
  ix54672z2388 : X_LUT4
    generic map(
      INIT => X"0050"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(3),
      O => nx54672z728
    );
  ix54672z2323 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(3),
      O => nx54672z729
    );
  ix54672z3881 : X_LUT4
    generic map(
      INIT => X"1E1E"
    )
    port map (
      ADR0 => romoaddro1_s(0),
      ADR1 => romoaddro1_s(2),
      ADR2 => romoaddro1_s(3),
      ADR3 => VCC,
      O => nx54672z737
    );
  ix53675z23856 : X_LUT4
    generic map(
      INIT => X"02DC"
    )
    port map (
      ADR0 => romo2addro6_s(1),
      ADR1 => romo2addro6_s(2),
      ADR2 => romo2addro6_s(3),
      ADR3 => romo2addro6_s(0),
      O => nx53675z1211
    );
  ix53675z52440 : X_LUT4
    generic map(
      INIT => X"8E8E"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(1),
      ADR2 => romo2addro6_s(3),
      ADR3 => VCC,
      O => nx53675z1215
    );
  ix53675z4630 : X_LUT4
    generic map(
      INIT => X"3366"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(3),
      ADR2 => VCC,
      ADR3 => romo2addro6_s(0),
      O => nx53675z1262
    );
  ix53675z7091 : X_LUT4
    generic map(
      INIT => X"3B3C"
    )
    port map (
      ADR0 => romo2addro6_s(1),
      ADR1 => romo2addro6_s(2),
      ADR2 => romo2addro6_s(3),
      ADR3 => romo2addro6_s(0),
      O => nx53675z1212
    );
  ix53675z10811 : X_LUT4
    generic map(
      INIT => X"555A"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => VCC,
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(0),
      O => nx53675z1263
    );
  ix53675z57165 : X_LUT4
    generic map(
      INIT => X"D2D2"
    )
    port map (
      ADR0 => romo2addro6_s(2),
      ADR1 => romo2addro6_s(3),
      ADR2 => romo2addro6_s(1),
      ADR3 => VCC,
      O => nx53675z1259
    );
  ix53675z24960 : X_LUT4
    generic map(
      INIT => X"03FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2addro6_s(3),
      ADR2 => romo2addro6_s(1),
      ADR3 => romo2addro6_s(0),
      O => nx53675z1260
    );
  ix53675z41953 : X_LUT4
    generic map(
      INIT => X"9694"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(0),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1147
    );
  ix53675z58634 : X_LUT4
    generic map(
      INIT => X"CB92"
    )
    port map (
      ADR0 => romo2addro5_s(3),
      ADR1 => romo2addro5_s(1),
      ADR2 => romo2addro5_s(0),
      ADR3 => romo2addro5_s(2),
      O => nx53675z1144
    );
  ix54672z24323 : X_LUT4
    generic map(
      INIT => X"0F5A"
    )
    port map (
      ADR0 => romoaddro2_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(3),
      O => nx54672z814
    );
  ix54672z25601 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro2_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro2_s(2),
      O => nx54672z818
    );
  ix54672z28686 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro2_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro2_s(1),
      O => nx54672z819
    );
  ix54672z6548 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romoaddro2_s(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romoaddro2_s(2),
      O => U1_ROMO2_modgen_rom_ix0_nx_rm64_16_u
    );
  ix54672z15729 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romoaddro2_s(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romoaddro2_s(1),
      O => U1_ROMO2_modgen_rom_ix0_nx_rm64_16_l
    );
  ix54672z58889 : X_LUT4
    generic map(
      INIT => X"F03C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(3),
      ADR3 => romoaddro1_s(1),
      O => nx54672z683
    );
  ix54672z42624 : X_LUT4
    generic map(
      INIT => X"CF32"
    )
    port map (
      ADR0 => romoaddro1_s(3),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(1),
      O => nx54672z680
    );
  ix54672z28433 : X_LUT4
    generic map(
      INIT => X"55A0"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro1_s(3),
      ADR3 => romoaddro1_s(0),
      O => nx54672z689
    );
  ix54672z14580 : X_LUT4
    generic map(
      INIT => X"03C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro1_s(2),
      ADR2 => romoaddro1_s(3),
      ADR3 => romoaddro1_s(1),
      O => nx54672z684
    );
  ix54672z48121 : X_LUT4
    generic map(
      INIT => X"BB2A"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z745
    );
  ix54672z54842 : X_LUT4
    generic map(
      INIT => X"CFCE"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z742
    );
  ix54672z2705 : X_LUT4
    generic map(
      INIT => X"0F0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro2_s(0),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z810
    );
  ix54672z2198 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romoaddro2_s(1),
      ADR1 => romoaddro2_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro2_s(2),
      O => nx54672z811
    );
  ix54672z2500 : X_LUT4
    generic map(
      INIT => X"0500"
    )
    port map (
      ADR0 => romoaddro2_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z807
    );
  ix54672z2435 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro2_s(0),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(1),
      O => nx54672z808
    );
  ix54672z3993 : X_LUT4
    generic map(
      INIT => X"05FA"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(3),
      O => nx54672z816
    );
  ix54672z54744 : X_LUT4
    generic map(
      INIT => X"99AA"
    )
    port map (
      ADR0 => romoaddro2_s(1),
      ADR1 => romoaddro2_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro2_s(2),
      O => nx54672z813
    );
  ix54672z10174 : X_LUT4
    generic map(
      INIT => X"05FA"
    )
    port map (
      ADR0 => romoaddro2_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(2),
      O => nx54672z817
    );
  ix54672z27677 : X_LUT4
    generic map(
      INIT => X"3C96"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z253
    );
  ix54672z17174 : X_LUT4
    generic map(
      INIT => X"659A"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z250
    );
  ix54672z17101 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romeaddro3_s(1),
      O => nx54672z259
    );
  ix54672z23609 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => VCC,
      O => U1_ROME3_modgen_rom_ix2_nx_rm64_16_l
    );
  ix54672z18190 : X_LUT4
    generic map(
      INIT => X"7110"
    )
    port map (
      ADR0 => romeaddro3_s(3),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(1),
      ADR3 => romeaddro3_s(2),
      O => nx54672z198
    );
  ix54672z17566 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romeaddro8_s(1),
      ADR1 => romeaddro8_s(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z584
    );
  ix54672z24074 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U1_ROME8_modgen_rom_ix2_nx_rm64_16_l
    );
  ix54672z26427 : X_LUT4
    generic map(
      INIT => X"3942"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(2),
      O => nx54672z161
    );
  ix54672z12551 : X_LUT4
    generic map(
      INIT => X"20B2"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(2),
      O => nx54672z163
    );
  ix54672z22855 : X_LUT4
    generic map(
      INIT => X"0A2A"
    )
    port map (
      ADR0 => romoaddro1_s(2),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(1),
      O => nx54672z671
    );
  ix54672z24362 : X_LUT4
    generic map(
      INIT => X"1A86"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(2),
      O => nx54672z164
    );
  ix54672z25431 : X_LUT4
    generic map(
      INIT => X"3C78"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(3),
      O => nx54672z677
    );
  ix54672z54739 : X_LUT4
    generic map(
      INIT => X"FF32"
    )
    port map (
      ADR0 => romoaddro1_s(2),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(1),
      O => nx54672z669
    );
  ix54672z54731 : X_LUT4
    generic map(
      INIT => X"BBBA"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(2),
      O => nx54672z663
    );
  ix54672z29360 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romoaddro8_s(1),
      O => nx54672z1293
    );
  ix54672z16402 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romoaddro8_s(1),
      O => U1_ROMO8_modgen_rom_ix0_nx_rm64_16_l
    );
  ix54672z22847 : X_LUT4
    generic map(
      INIT => X"1F00"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(2),
      O => nx54672z665
    );
  ix54672z48010 : X_LUT4
    generic map(
      INIT => X"F570"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(2),
      O => nx54672z666
    );
  ix54672z22752 : X_LUT4
    generic map(
      INIT => X"5070"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(3),
      O => nx54672z594
    );
  ix54672z59501 : X_LUT4
    generic map(
      INIT => X"E000"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(3),
      O => nx54672z591
    );
  ix54672z13922 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z105
    );
  ix54672z24289 : X_LUT4
    generic map(
      INIT => X"1C86"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z114
    );
  ix54672z18507 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(0),
      ADR2 => romeaddro1_s(3),
      ADR3 => romeaddro1_s(1),
      O => nx54672z110
    );
  ix54672z3675 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z102
    );
  ix54672z33948 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(0),
      ADR2 => romeaddro1_s(3),
      ADR3 => romeaddro1_s(1),
      O => nx54672z107
    );
  ix54672z4678 : X_LUT4
    generic map(
      INIT => X"5D04"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(0),
      ADR2 => romeaddro1_s(3),
      ADR3 => romeaddro1_s(1),
      O => nx54672z111
    );
  ix54672z7370 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => romeaddro0_s(1),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(0),
      ADR3 => romeaddro0_s(2),
      O => nx54672z31
    );
  ix54672z12033 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z116
    );
  ix54672z25273 : X_LUT4
    generic map(
      INIT => X"7130"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(0),
      ADR2 => romeaddro1_s(3),
      ADR3 => romeaddro1_s(1),
      O => nx54672z108
    );
  ix54672z8774 : X_LUT4
    generic map(
      INIT => X"249A"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z117
    );
  ix54672z61266 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z113
    );
  ix54672z12369 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => romeaddro0_s(1),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(0),
      ADR3 => romeaddro0_s(2),
      O => nx54672z34
    );
  ix54672z3587 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => romeaddro0_s(0),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(1),
      ADR3 => romeaddro0_s(2),
      O => nx54672z38
    );
  ix54672z24180 : X_LUT4
    generic map(
      INIT => X"1C86"
    )
    port map (
      ADR0 => romeaddro0_s(1),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(0),
      ADR3 => romeaddro0_s(2),
      O => nx54672z35
    );
  ix54672z11929 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => romeaddro0_s(0),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(1),
      ADR3 => romeaddro0_s(2),
      O => nx54672z40
    );
  ix54672z26245 : X_LUT4
    generic map(
      INIT => X"5924"
    )
    port map (
      ADR0 => romeaddro0_s(1),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(0),
      ADR3 => romeaddro0_s(2),
      O => nx54672z32
    );
  ix54672z13834 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => romeaddro0_s(0),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(1),
      ADR3 => romeaddro0_s(2),
      O => nx54672z41
    );
  ix54672z18419 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(0),
      O => nx54672z46
    );
  ix54672z61162 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro0_s(0),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(1),
      ADR3 => romeaddro0_s(2),
      O => nx54672z37
    );
  ix54672z33860 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(0),
      O => nx54672z43
    );
  ix54672z4590 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(0),
      O => nx54672z47
    );
  ix54672z25185 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(0),
      O => nx54672z44
    );
  ix54672z16899 : X_LUT4
    generic map(
      INIT => X"39C6"
    )
    port map (
      ADR0 => romeaddro0_s(0),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(2),
      O => nx54672z56
    );
  ix54672z11945 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(1),
      ADR3 => romeaddro0_s(0),
      O => nx54672z52
    );
  ix54672z61178 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(1),
      ADR3 => romeaddro0_s(0),
      O => nx54672z49
    );
  ix54672z8686 : X_LUT4
    generic map(
      INIT => X"6158"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(1),
      ADR3 => romeaddro0_s(0),
      O => nx54672z53
    );
  ix54672z18499 : X_LUT4
    generic map(
      INIT => X"4D24"
    )
    port map (
      ADR0 => romeaddro0_s(0),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(2),
      O => nx54672z58
    );
  ix54672z24201 : X_LUT4
    generic map(
      INIT => X"429C"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(1),
      ADR3 => romeaddro0_s(0),
      O => nx54672z50
    );
  ix54672z27402 : X_LUT4
    generic map(
      INIT => X"695A"
    )
    port map (
      ADR0 => romeaddro0_s(0),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(2),
      O => nx54672z59
    );
  ix54672z26275 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romoaddro8_s(2),
      O => nx54672z1292
    );
  ix54672z33876 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro0_s(0),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(2),
      O => nx54672z55
    );
  ix54672z6454 : X_LUT4
    generic map(
      INIT => X"31EE"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(1),
      ADR3 => romoaddro2_s(2),
      O => nx54672z766
    );
  ix54672z5285 : X_LUT4
    generic map(
      INIT => X"4254"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(1),
      O => nx54672z771
    );
  ix54672z64663 : X_LUT4
    generic map(
      INIT => X"88EE"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro2_s(1),
      O => nx54672z775
    );
  ix54672z41428 : X_LUT4
    generic map(
      INIT => X"9686"
    )
    port map (
      ADR0 => romoaddro2_s(1),
      ADR1 => romoaddro2_s(0),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z780
    );
  ix54672z22926 : X_LUT4
    generic map(
      INIT => X"1838"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(1),
      O => nx54672z772
    );
  ix54672z44758 : X_LUT4
    generic map(
      INIT => X"C63C"
    )
    port map (
      ADR0 => romoaddro2_s(1),
      ADR1 => romoaddro2_s(0),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z778
    );
  ix54672z52395 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => romoaddro2_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z781
    );
  ix54672z43798 : X_LUT4
    generic map(
      INIT => X"F002"
    )
    port map (
      ADR0 => romoaddro2_s(3),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(2),
      O => nx54672z786
    );
  ix54672z58109 : X_LUT4
    generic map(
      INIT => X"B994"
    )
    port map (
      ADR0 => romoaddro2_s(1),
      ADR1 => romoaddro2_s(0),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z777
    );
  ix54672z22647 : X_LUT4
    generic map(
      INIT => X"08AE"
    )
    port map (
      ADR0 => romoaddro2_s(3),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(2),
      O => nx54672z783
    );
  ix54672z44647 : X_LUT4
    generic map(
      INIT => X"96B4"
    )
    port map (
      ADR0 => romoaddro1_s(2),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(1),
      O => nx54672z699
    );
  ix54672z52284 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => romoaddro1_s(2),
      ADR1 => romoaddro1_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro1_s(1),
      O => nx54672z702
    );
  ix54672z43687 : X_LUT4
    generic map(
      INIT => X"CC10"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(3),
      ADR3 => romoaddro1_s(2),
      O => nx54672z707
    );
  ix54672z38197 : X_LUT4
    generic map(
      INIT => X"85A0"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(3),
      ADR3 => romoaddro1_s(2),
      O => nx54672z705
    );
  ix54672z61840 : X_LUT4
    generic map(
      INIT => X"E888"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(3),
      ADR3 => romoaddro1_s(2),
      O => nx54672z708
    );
  ix54672z25489 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro1_s(2),
      ADR2 => romoaddro1_s(0),
      ADR3 => VCC,
      O => nx54672z739
    );
  ix54672z22536 : X_LUT4
    generic map(
      INIT => X"20F2"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(3),
      ADR3 => romoaddro1_s(2),
      O => nx54672z704
    );
  ix54672z6436 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro1_s(2),
      ADR2 => VCC,
      ADR3 => romoaddro1_s(3),
      O => U1_ROMO1_modgen_rom_ix0_nx_rm64_16_u
    );
  ix54672z28574 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romoaddro1_s(0),
      ADR3 => romoaddro1_s(1),
      O => nx54672z740
    );
  ix54672z15617 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro1_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro1_s(3),
      O => U1_ROMO1_modgen_rom_ix0_nx_rm64_16_l
    );
  ix54672z18787 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(3),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(1),
      O => nx54672z305
    );
  ix54672z25553 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(3),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(1),
      O => nx54672z303
    );
  ix54672z12313 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro4_s(3),
      ADR1 => romeaddro4_s(1),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(0),
      O => nx54672z311
    );
  ix54672z4958 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(3),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(1),
      O => nx54672z306
    );
  ix54672z24569 : X_LUT4
    generic map(
      INIT => X"18A6"
    )
    port map (
      ADR0 => romeaddro4_s(3),
      ADR1 => romeaddro4_s(1),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(0),
      O => nx54672z309
    );
  ix54672z9054 : X_LUT4
    generic map(
      INIT => X"492C"
    )
    port map (
      ADR0 => romeaddro4_s(3),
      ADR1 => romeaddro4_s(1),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(0),
      O => nx54672z312
    );
  ix54672z61546 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro4_s(3),
      ADR1 => romeaddro4_s(1),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(0),
      O => nx54672z308
    );
  ix54672z18002 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z68
    );
  ix54672z21153 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(1),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(3),
      O => nx54672z84
    );
  ix54672z18587 : X_LUT4
    generic map(
      INIT => X"2B42"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(0),
      ADR2 => romeaddro1_s(3),
      ADR3 => romeaddro1_s(1),
      O => nx54672z122
    );
  ix54672z33964 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(0),
      ADR2 => romeaddro1_s(3),
      ADR3 => romeaddro1_s(1),
      O => nx54672z119
    );
  ix54672z27490 : X_LUT4
    generic map(
      INIT => X"3C96"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(0),
      ADR2 => romeaddro1_s(3),
      ADR3 => romeaddro1_s(1),
      O => nx54672z123
    );
  ix54672z28517 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(1),
      ADR3 => romeaddro1_s(0),
      O => nx54672z127
    );
  ix54672z16987 : X_LUT4
    generic map(
      INIT => X"59A6"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(0),
      ADR2 => romeaddro1_s(3),
      ADR3 => romeaddro1_s(1),
      O => nx54672z120
    );
  ix54672z13824 : X_LUT4
    generic map(
      INIT => X"0A0A"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => VCC,
      ADR2 => romeaddro1_s(1),
      ADR3 => VCC,
      O => nx54672z128
    );
  ix54672z28514 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(1),
      ADR3 => romeaddro1_s(0),
      O => U1_ROME1_modgen_rom_ix2_nx_rm64_16_u
    );
  ix54672z1655 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romeaddro1_s(3),
      ADR2 => VCC,
      ADR3 => romeaddro1_s(0),
      O => nx54672z125
    );
  ix54672z40034 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(2),
      O => nx54672z154
    );
  ix54672z25346 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(2),
      O => nx54672z158
    );
  ix54672z30507 : X_LUT4
    generic map(
      INIT => X"2F02"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(2),
      O => nx54672z155
    );
  ix54672z17008 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romeaddro2_s(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romeaddro2_s(2),
      O => nx54672z194
    );
  ix54672z23516 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romeaddro2_s(0),
      ADR2 => VCC,
      ADR3 => romeaddro2_s(3),
      O => U1_ROME2_modgen_rom_ix2_nx_rm64_16_l
    );
  ix54672z44022 : X_LUT4
    generic map(
      INIT => X"F004"
    )
    port map (
      ADR0 => romoaddro4_s(1),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(0),
      ADR3 => romoaddro4_s(2),
      O => nx54672z944
    );
  ix54672z13873 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z69
    );
  ix54672z3626 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(2),
      O => nx54672z66
    );
  ix54672z7731 : X_LUT4
    generic map(
      INIT => X"2962"
    )
    port map (
      ADR0 => romeaddro1_s(0),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(2),
      ADR3 => romeaddro1_s(1),
      O => nx54672z78
    );
  ix54672z18467 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => romeaddro1_s(0),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(2),
      ADR3 => romeaddro1_s(1),
      O => nx54672z80
    );
  ix54672z14882 : X_LUT4
    generic map(
      INIT => X"24D2"
    )
    port map (
      ADR0 => romeaddro1_s(0),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(2),
      ADR3 => romeaddro1_s(1),
      O => nx54672z81
    );
  ix54672z11993 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(1),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(3),
      O => nx54672z86
    );
  ix54672z7156 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => romeaddro1_s(0),
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(2),
      ADR3 => romeaddro1_s(1),
      O => nx54672z77
    );
  ix54672z34474 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(1),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(3),
      O => nx54672z83
    );
  ix54672z3654 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(1),
      ADR2 => romeaddro1_s(0),
      ADR3 => romeaddro1_s(3),
      O => nx54672z87
    );
  ix54672z16915 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romeaddro1_s(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romeaddro1_s(2),
      O => nx54672z129
    );
  ix54672z23422 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romeaddro1_s(3),
      ADR2 => romeaddro1_s(0),
      ADR3 => VCC,
      O => U1_ROME1_modgen_rom_ix2_nx_rm64_16_l
    );
  ix54672z3547 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => romeaddro0_s(1),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(0),
      ADR3 => romeaddro0_s(2),
      O => nx54672z8
    );
  ix54672z17923 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => romeaddro0_s(1),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(0),
      ADR3 => romeaddro0_s(2),
      O => nx54672z10
    );
  ix54672z13794 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => romeaddro0_s(1),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(0),
      ADR3 => romeaddro0_s(2),
      O => nx54672z11
    );
  ix54672z18379 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(0),
      O => nx54672z16
    );
  ix54672z60844 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => romeaddro0_s(1),
      ADR1 => romeaddro0_s(3),
      ADR2 => romeaddro0_s(0),
      ADR3 => romeaddro0_s(2),
      O => nx54672z7
    );
  ix54672z7068 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(1),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(0),
      O => nx54672z13
    );
  ix54672z44544 : X_LUT4
    generic map(
      INIT => X"A56A"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(3),
      O => nx54672z622
    );
  ix54672z27746 : X_LUT4
    generic map(
      INIT => X"5E96"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(2),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(0),
      O => nx54672z634
    );
  ix54672z22433 : X_LUT4
    generic map(
      INIT => X"5D04"
    )
    port map (
      ADR0 => romoaddro0_s(2),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(0),
      ADR3 => romoaddro0_s(3),
      O => nx54672z627
    );
  ix54672z61737 : X_LUT4
    generic map(
      INIT => X"E8C0"
    )
    port map (
      ADR0 => romoaddro0_s(2),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(0),
      ADR3 => romoaddro0_s(3),
      O => nx54672z631
    );
  ix54672z20994 : X_LUT4
    generic map(
      INIT => X"31C6"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(2),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(0),
      O => nx54672z636
    );
  ix54672z38094 : X_LUT4
    generic map(
      INIT => X"C422"
    )
    port map (
      ADR0 => romoaddro0_s(2),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(0),
      ADR3 => romoaddro0_s(3),
      O => nx54672z628
    );
  ix54672z36623 : X_LUT4
    generic map(
      INIT => X"8770"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(2),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(0),
      O => nx54672z637
    );
  ix54672z40060 : X_LUT4
    generic map(
      INIT => X"C666"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(0),
      O => nx54672z642
    );
  ix54672z19289 : X_LUT4
    generic map(
      INIT => X"4694"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(2),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(0),
      O => nx54672z633
    );
  ix54672z29203 : X_LUT4
    generic map(
      INIT => X"39C6"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(0),
      O => nx54672z639
    );
  ix54672z3539 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(0),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(1),
      O => nx54672z2
    );
  ix54672z18198 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z204
    );
  ix54672z3822 : X_LUT4
    generic map(
      INIT => X"7130"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z202
    );
  ix54672z18694 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z240
    );
  ix54672z14069 : X_LUT4
    generic map(
      INIT => X"20BA"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z205
    );
  ix54672z25460 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z238
    );
  ix54672z4865 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z241
    );
  ix54672z18774 : X_LUT4
    generic map(
      INIT => X"2B42"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z252
    );
  ix54672z34135 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z237
    );
  ix54672z34151 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z249
    );
  ix54672z13976 : X_LUT4
    generic map(
      INIT => X"44D4"
    )
    port map (
      ADR0 => romeaddro2_s(1),
      ADR1 => romeaddro2_s(2),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(3),
      O => nx54672z140
    );
  ix54672z18561 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(2),
      ADR3 => romeaddro2_s(1),
      O => nx54672z145
    );
  ix54672z3729 : X_LUT4
    generic map(
      INIT => X"20F2"
    )
    port map (
      ADR0 => romeaddro2_s(1),
      ADR1 => romeaddro2_s(2),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(3),
      O => nx54672z137
    );
  ix54672z7825 : X_LUT4
    generic map(
      INIT => X"4964"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(2),
      ADR3 => romeaddro2_s(1),
      O => nx54672z143
    );
  ix54672z14976 : X_LUT4
    generic map(
      INIT => X"42B4"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(2),
      ADR3 => romeaddro2_s(1),
      O => nx54672z146
    );
  ix54672z12087 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(3),
      O => nx54672z151
    );
  ix54672z7250 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(2),
      ADR3 => romeaddro2_s(1),
      O => nx54672z142
    );
  ix54672z34568 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(3),
      O => nx54672z148
    );
  ix54672z21247 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(3),
      O => nx54672z149
    );
  ix54672z3748 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => romeaddro2_s(2),
      ADR1 => romeaddro2_s(1),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(3),
      O => nx54672z152
    );
  ix54672z18577 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => romeaddro2_s(3),
      ADR1 => romeaddro2_s(0),
      ADR2 => romeaddro2_s(1),
      ADR3 => romeaddro2_s(2),
      O => nx54672z157
    );
  ix54672z14061 : X_LUT4
    generic map(
      INIT => X"4F04"
    )
    port map (
      ADR0 => romeaddro3_s(3),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(1),
      ADR3 => romeaddro3_s(2),
      O => nx54672z199
    );
  ix54672z3814 : X_LUT4
    generic map(
      INIT => X"44D4"
    )
    port map (
      ADR0 => romeaddro3_s(3),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(1),
      ADR3 => romeaddro3_s(2),
      O => nx54672z196
    );
  ix54672z24662 : X_LUT4
    generic map(
      INIT => X"6518"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => romeaddro5_s(2),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(3),
      O => nx54672z374
    );
  ix54672z12406 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => romeaddro5_s(2),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(3),
      O => nx54672z376
    );
  ix54672z18960 : X_LUT4
    generic map(
      INIT => X"188E"
    )
    port map (
      ADR0 => romeaddro5_s(2),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(3),
      ADR3 => romeaddro5_s(0),
      O => nx54672z382
    );
  ix54672z9147 : X_LUT4
    generic map(
      INIT => X"3492"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => romeaddro5_s(2),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(3),
      O => nx54672z377
    );
  ix54672z34337 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro5_s(2),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(3),
      ADR3 => romeaddro5_s(0),
      O => nx54672z379
    );
  ix54672z17360 : X_LUT4
    generic map(
      INIT => X"6966"
    )
    port map (
      ADR0 => romeaddro5_s(2),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(3),
      ADR3 => romeaddro5_s(0),
      O => nx54672z380
    );
  ix54672z27863 : X_LUT4
    generic map(
      INIT => X"2DD2"
    )
    port map (
      ADR0 => romeaddro5_s(2),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(3),
      ADR3 => romeaddro5_s(0),
      O => nx54672z383
    );
  ix54672z11513 : X_LUT4
    generic map(
      INIT => X"0A50"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro5_s(1),
      ADR3 => romoaddro5_s(0),
      O => nx54672z1011
    );
  ix54672z10385 : X_LUT4
    generic map(
      INIT => X"5A6A"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(0),
      O => nx54672z643
    );
  ix54672z25432 : X_LUT4
    generic map(
      INIT => X"6688"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(2),
      ADR2 => VCC,
      ADR3 => romoaddro0_s(3),
      O => nx54672z648
    );
  ix54672z25382 : X_LUT4
    generic map(
      INIT => X"1EF0"
    )
    port map (
      ADR0 => romoaddro0_s(3),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(2),
      ADR3 => romoaddro0_s(0),
      O => nx54672z640
    );
  ix54672z41297 : X_LUT4
    generic map(
      INIT => X"A4A4"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => romoaddro0_s(2),
      ADR2 => romoaddro0_s(1),
      ADR3 => VCC,
      O => nx54672z649
    );
  ix54672z6261 : X_LUT4
    generic map(
      INIT => X"33C0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro0_s(2),
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(3),
      O => nx54672z645
    );
  ix54672z54488 : X_LUT4
    generic map(
      INIT => X"F00A"
    )
    port map (
      ADR0 => romoaddro0_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro0_s(1),
      ADR3 => romoaddro0_s(3),
      O => nx54672z646
    );
  ix54672z17915 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(0),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(1),
      O => nx54672z4
    );
  ix54672z13786 : X_LUT4
    generic map(
      INIT => X"08AE"
    )
    port map (
      ADR0 => romeaddro0_s(2),
      ADR1 => romeaddro0_s(0),
      ADR2 => romeaddro0_s(3),
      ADR3 => romeaddro0_s(1),
      O => nx54672z5
    );
  ix54672z18376 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(2),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(0),
      O => nx54672z328
    );
  ix54672z64998 : X_LUT4
    generic map(
      INIT => X"AF0A"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro5_s(1),
      ADR3 => romoaddro5_s(2),
      O => nx54672z1012
    );
  ix54672z4000 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(2),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(0),
      O => nx54672z326
    );
  ix54672z23261 : X_LUT4
    generic map(
      INIT => X"1588"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(1),
      ADR3 => romoaddro5_s(0),
      O => nx54672z1009
    );
  ix54672z14247 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(2),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(0),
      O => nx54672z329
    );
  ix54672z18105 : X_LUT4
    generic map(
      INIT => X"088E"
    )
    port map (
      ADR0 => romeaddro2_s(1),
      ADR1 => romeaddro2_s(2),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(3),
      O => nx54672z139
    );
  ix54672z61026 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => romeaddro2_s(1),
      ADR1 => romeaddro2_s(2),
      ADR2 => romeaddro2_s(0),
      ADR3 => romeaddro2_s(3),
      O => nx54672z136
    );
  ix54672z15840 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romoaddro3_s(1),
      O => U1_ROMO3_modgen_rom_ix0_nx_rm64_16_l
    );
  ix54672z59000 : X_LUT4
    generic map(
      INIT => X"A5F0"
    )
    port map (
      ADR0 => romoaddro2_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(0),
      O => nx54672z762
    );
  ix54672z14691 : X_LUT4
    generic map(
      INIT => X"500A"
    )
    port map (
      ADR0 => romoaddro2_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(2),
      O => nx54672z763
    );
  ix54672z28544 : X_LUT4
    generic map(
      INIT => X"44AA"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro2_s(1),
      O => nx54672z768
    );
  ix54672z42735 : X_LUT4
    generic map(
      INIT => X"F05E"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(1),
      ADR3 => romoaddro2_s(0),
      O => nx54672z759
    );
  ix54672z24228 : X_LUT4
    generic map(
      INIT => X"00FA"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(0),
      O => nx54672z760
    );
  ix54672z23219 : X_LUT4
    generic map(
      INIT => X"5524"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(1),
      ADR3 => romoaddro2_s(2),
      O => nx54672z765
    );
  ix54672z11178 : X_LUT4
    generic map(
      INIT => X"1188"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro2_s(1),
      O => nx54672z774
    );
  ix54672z51803 : X_LUT4
    generic map(
      INIT => X"BB22"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro2_s(1),
      O => nx54672z769
    );
  ix54672z25820 : X_LUT4
    generic map(
      INIT => X"57A8"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(2),
      O => nx54672z954
    );
  ix54672z59112 : X_LUT4
    generic map(
      INIT => X"BB44"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro3_s(3),
      O => nx54672z841
    );
  ix54672z23078 : X_LUT4
    generic map(
      INIT => X"04CC"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(1),
      ADR3 => romoaddro3_s(0),
      O => nx54672z829
    );
  ix54672z29529 : X_LUT4
    generic map(
      INIT => X"6966"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(3),
      O => nx54672z874
    );
  ix54672z54962 : X_LUT4
    generic map(
      INIT => X"F5F4"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(1),
      ADR3 => romoaddro3_s(0),
      O => nx54672z827
    );
  ix54672z48241 : X_LUT4
    generic map(
      INIT => X"DF0C"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(1),
      ADR3 => romoaddro3_s(0),
      O => nx54672z830
    );
  ix54672z14803 : X_LUT4
    generic map(
      INIT => X"4422"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => VCC,
      ADR3 => romoaddro3_s(3),
      O => nx54672z842
    );
  ix54672z42847 : X_LUT4
    generic map(
      INIT => X"9B9A"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(3),
      O => nx54672z838
    );
  ix54672z24340 : X_LUT4
    generic map(
      INIT => X"3330"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(3),
      O => nx54672z839
    );
  ix54672z40386 : X_LUT4
    generic map(
      INIT => X"95AA"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(3),
      O => nx54672z877
    );
  ix54672z14162 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(1),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(3),
      O => nx54672z270
    );
  ix54672z3915 : X_LUT4
    generic map(
      INIT => X"08AE"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(1),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(3),
      O => nx54672z267
    );
  ix54672z21433 : X_LUT4
    generic map(
      INIT => X"7130"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(3),
      O => nx54672z279
    );
  ix54672z18747 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => romeaddro4_s(3),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(0),
      O => nx54672z275
    );
  ix54672z7436 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => romeaddro4_s(3),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(0),
      O => nx54672z272
    );
  ix54672z15162 : X_LUT4
    generic map(
      INIT => X"492C"
    )
    port map (
      ADR0 => romeaddro4_s(3),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(0),
      O => nx54672z276
    );
  ix54672z12273 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(3),
      O => nx54672z281
    );
  ix54672z8011 : X_LUT4
    generic map(
      INIT => X"6518"
    )
    port map (
      ADR0 => romeaddro4_s(3),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(0),
      O => nx54672z273
    );
  ix54672z3934 : X_LUT4
    generic map(
      INIT => X"20BA"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(3),
      O => nx54672z282
    );
  ix54672z34754 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(3),
      O => nx54672z278
    );
  ix54672z18867 : X_LUT4
    generic map(
      INIT => X"188E"
    )
    port map (
      ADR0 => romeaddro4_s(1),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(3),
      ADR3 => romeaddro4_s(0),
      O => nx54672z317
    );
  ix54672z34244 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro4_s(1),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(3),
      ADR3 => romeaddro4_s(0),
      O => nx54672z314
    );
  ix54672z21432 : X_LUT4
    generic map(
      INIT => X"6616"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(2),
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(1),
      O => nx54672z950
    );
  ix54672z38532 : X_LUT4
    generic map(
      INIT => X"9188"
    )
    port map (
      ADR0 => romoaddro4_s(1),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(0),
      ADR3 => romoaddro4_s(2),
      O => nx54672z942
    );
  ix54672z62175 : X_LUT4
    generic map(
      INIT => X"E8A0"
    )
    port map (
      ADR0 => romoaddro4_s(1),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(0),
      ADR3 => romoaddro4_s(2),
      O => nx54672z945
    );
  ix54672z28184 : X_LUT4
    generic map(
      INIT => X"4BBC"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(2),
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(1),
      O => nx54672z948
    );
  ix54672z37061 : X_LUT4
    generic map(
      INIT => X"952A"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(2),
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(1),
      O => nx54672z951
    );
  ix54672z40498 : X_LUT4
    generic map(
      INIT => X"B43C"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(2),
      O => nx54672z956
    );
  ix54672z19727 : X_LUT4
    generic map(
      INIT => X"492C"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(2),
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(1),
      O => nx54672z947
    );
  ix54672z29641 : X_LUT4
    generic map(
      INIT => X"5A96"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(2),
      O => nx54672z953
    );
  ix54672z10823 : X_LUT4
    generic map(
      INIT => X"36CC"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(2),
      O => nx54672z957
    );
  ix54672z54954 : X_LUT4
    generic map(
      INIT => X"AFAE"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(3),
      ADR3 => romoaddro3_s(0),
      O => nx54672z821
    );
  ix54672z21097 : X_LUT4
    generic map(
      INIT => X"293C"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(3),
      O => nx54672z713
    );
  ix54672z27849 : X_LUT4
    generic map(
      INIT => X"65DA"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(3),
      O => nx54672z711
    );
  ix54672z25485 : X_LUT4
    generic map(
      INIT => X"5A78"
    )
    port map (
      ADR0 => romoaddro1_s(0),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(1),
      O => nx54672z717
    );
  ix54672z36726 : X_LUT4
    generic map(
      INIT => X"8666"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(3),
      O => nx54672z714
    );
  ix54672z40163 : X_LUT4
    generic map(
      INIT => X"B34C"
    )
    port map (
      ADR0 => romoaddro1_s(0),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(1),
      O => nx54672z719
    );
  ix54672z19392 : X_LUT4
    generic map(
      INIT => X"24D2"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(3),
      O => nx54672z710
    );
  ix54672z10488 : X_LUT4
    generic map(
      INIT => X"3C6C"
    )
    port map (
      ADR0 => romoaddro1_s(0),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(1),
      O => nx54672z720
    );
  ix54672z25535 : X_LUT4
    generic map(
      INIT => X"6868"
    )
    port map (
      ADR0 => romoaddro1_s(3),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(2),
      ADR3 => VCC,
      O => nx54672z725
    );
  ix54672z29306 : X_LUT4
    generic map(
      INIT => X"59A6"
    )
    port map (
      ADR0 => romoaddro1_s(0),
      ADR1 => romoaddro1_s(3),
      ADR2 => romoaddro1_s(2),
      ADR3 => romoaddro1_s(1),
      O => nx54672z716
    );
  ix54672z6364 : X_LUT4
    generic map(
      INIT => X"6262"
    )
    port map (
      ADR0 => romoaddro1_s(3),
      ADR1 => romoaddro1_s(2),
      ADR2 => romoaddro1_s(1),
      ADR3 => VCC,
      O => nx54672z722
    );
  ix54672z10711 : X_LUT4
    generic map(
      INIT => X"1FE0"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(3),
      O => nx54672z878
    );
  ix54672z2816 : X_LUT4
    generic map(
      INIT => X"00FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(0),
      ADR3 => romoaddro3_s(3),
      O => nx54672z889
    );
  ix54672z25708 : X_LUT4
    generic map(
      INIT => X"3C78"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(3),
      O => nx54672z875
    );
  ix54672z2309 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(0),
      ADR3 => romoaddro3_s(1),
      O => nx54672z890
    );
  ix54672z2611 : X_LUT4
    generic map(
      INIT => X"0044"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => VCC,
      ADR3 => romoaddro3_s(3),
      O => nx54672z886
    );
  ix54672z2546 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro3_s(0),
      ADR3 => romoaddro3_s(3),
      O => nx54672z887
    );
  ix54672z25712 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romoaddro3_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro3_s(2),
      ADR3 => VCC,
      O => nx54672z897
    );
  ix54672z6659 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro3_s(2),
      ADR3 => VCC,
      O => U1_ROMO3_modgen_rom_ix0_nx_rm64_16_u
    );
  ix54672z30069 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romoaddro3_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romoaddro3_s(1),
      O => nx54672z898
    );
  ix54672z61951 : X_LUT4
    generic map(
      INIT => X"E8C0"
    )
    port map (
      ADR0 => romoaddro2_s(3),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(2),
      O => nx54672z787
    );
  ix54672z23182 : X_LUT4
    generic map(
      INIT => X"02AA"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(0),
      O => nx54672z902
    );
  ix54672z38308 : X_LUT4
    generic map(
      INIT => X"9188"
    )
    port map (
      ADR0 => romoaddro2_s(3),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(2),
      O => nx54672z784
    );
  ix54672z55066 : X_LUT4
    generic map(
      INIT => X"F3F2"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(0),
      O => nx54672z900
    );
  ix54672z48345 : X_LUT4
    generic map(
      INIT => X"BF0A"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(0),
      O => nx54672z903
    );
  ix54672z23070 : X_LUT4
    generic map(
      INIT => X"04CC"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(3),
      ADR3 => romoaddro3_s(0),
      O => nx54672z823
    );
  ix54672z48233 : X_LUT4
    generic map(
      INIT => X"DF44"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(3),
      ADR3 => romoaddro3_s(0),
      O => nx54672z824
    );
  ix54672z41400 : X_LUT4
    generic map(
      INIT => X"9898"
    )
    port map (
      ADR0 => romoaddro1_s(1),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(2),
      ADR3 => VCC,
      O => nx54672z726
    );
  ix54672z4093 : X_LUT4
    generic map(
      INIT => X"08CE"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z391
    );
  ix54672z54591 : X_LUT4
    generic map(
      INIT => X"A4A4"
    )
    port map (
      ADR0 => romoaddro1_s(3),
      ADR1 => romoaddro1_s(0),
      ADR2 => romoaddro1_s(1),
      ADR3 => VCC,
      O => nx54672z723
    );
  ix54672z18469 : X_LUT4
    generic map(
      INIT => X"20B2"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z393
    );
  ix54672z14340 : X_LUT4
    generic map(
      INIT => X"50D4"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z394
    );
  ix54672z18291 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(1),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(3),
      O => nx54672z269
    );
  ix54672z61212 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(1),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(3),
      O => nx54672z266
    );
  ix54672z4186 : X_LUT4
    generic map(
      INIT => X"7130"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z456
    );
  ix54672z18933 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z405
    );
  ix54672z8197 : X_LUT4
    generic map(
      INIT => X"18C6"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z403
    );
  ix54672z21619 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => romeaddro6_s(0),
      ADR1 => romeaddro6_s(1),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z409
    );
  ix54672z15348 : X_LUT4
    generic map(
      INIT => X"5294"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z406
    );
  ix54672z12459 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro6_s(0),
      ADR1 => romeaddro6_s(1),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z411
    );
  ix54672z7622 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z402
    );
  ix54672z4120 : X_LUT4
    generic map(
      INIT => X"08AE"
    )
    port map (
      ADR0 => romeaddro6_s(0),
      ADR1 => romeaddro6_s(1),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z412
    );
  ix54672z18949 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(1),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(2),
      O => nx54672z417
    );
  ix54672z34940 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => romeaddro6_s(0),
      ADR1 => romeaddro6_s(1),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(3),
      O => nx54672z408
    );
  ix54672z40406 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(1),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(2),
      O => nx54672z414
    );
  ix54672z14290 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(1),
      O => nx54672z453
    );
  ix54672z2121 : X_LUT4
    generic map(
      INIT => X"2222"
    )
    port map (
      ADR0 => romeaddro6_s(0),
      ADR1 => romeaddro6_s(3),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z450
    );
  ix54672z17380 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romeaddro6_s(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romeaddro6_s(1),
      O => nx54672z454
    );
  ix54672z23888 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(3),
      O => U1_ROME6_modgen_rom_ix2_nx_rm64_16_l
    );
  ix54672z12180 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z216
    );
  ix54672z34661 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z213
    );
  ix54672z3841 : X_LUT4
    generic map(
      INIT => X"7130"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z217
    );
  ix54672z4008 : X_LUT4
    generic map(
      INIT => X"3B02"
    )
    port map (
      ADR0 => romeaddro5_s(1),
      ADR1 => romeaddro5_s(3),
      ADR2 => romeaddro5_s(2),
      ADR3 => romeaddro5_s(0),
      O => nx54672z332
    );
  ix54672z12644 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => romeaddro3_s(1),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(3),
      ADR3 => romeaddro3_s(2),
      O => nx54672z228
    );
  ix54672z21340 : X_LUT4
    generic map(
      INIT => X"5D04"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z214
    );
  ix54672z7645 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => romeaddro3_s(1),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(3),
      ADR3 => romeaddro3_s(2),
      O => nx54672z225
    );
  ix54672z24455 : X_LUT4
    generic map(
      INIT => X"3492"
    )
    port map (
      ADR0 => romeaddro3_s(1),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(3),
      ADR3 => romeaddro3_s(2),
      O => nx54672z229
    );
  ix54672z18384 : X_LUT4
    generic map(
      INIT => X"20B2"
    )
    port map (
      ADR0 => romeaddro5_s(1),
      ADR1 => romeaddro5_s(3),
      ADR2 => romeaddro5_s(2),
      ADR3 => romeaddro5_s(0),
      O => nx54672z334
    );
  ix54672z26520 : X_LUT4
    generic map(
      INIT => X"6518"
    )
    port map (
      ADR0 => romeaddro3_s(1),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(3),
      ADR3 => romeaddro3_s(2),
      O => nx54672z226
    );
  ix54672z14255 : X_LUT4
    generic map(
      INIT => X"7150"
    )
    port map (
      ADR0 => romeaddro5_s(1),
      ADR1 => romeaddro5_s(3),
      ADR2 => romeaddro5_s(2),
      ADR3 => romeaddro5_s(0),
      O => nx54672z335
    );
  ix54672z18840 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => romeaddro5_s(1),
      ADR1 => romeaddro5_s(2),
      ADR2 => romeaddro5_s(0),
      ADR3 => romeaddro5_s(3),
      O => nx54672z340
    );
  ix54672z61305 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => romeaddro5_s(1),
      ADR1 => romeaddro5_s(3),
      ADR2 => romeaddro5_s(2),
      ADR3 => romeaddro5_s(0),
      O => nx54672z331
    );
  ix54672z27770 : X_LUT4
    generic map(
      INIT => X"4BB4"
    )
    port map (
      ADR0 => romeaddro4_s(1),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(3),
      ADR3 => romeaddro4_s(0),
      O => nx54672z318
    );
  ix54672z28797 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(3),
      O => nx54672z322
    );
  ix54672z17267 : X_LUT4
    generic map(
      INIT => X"6966"
    )
    port map (
      ADR0 => romeaddro4_s(1),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(3),
      ADR3 => romeaddro4_s(0),
      O => nx54672z315
    );
  ix54672z14104 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => VCC,
      O => nx54672z323
    );
  ix54672z28794 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(3),
      O => U1_ROME4_modgen_rom_ix2_nx_rm64_16_u
    );
  ix54672z1935 : X_LUT4
    generic map(
      INIT => X"00CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romeaddro4_s(0),
      ADR2 => VCC,
      ADR3 => romeaddro4_s(3),
      O => nx54672z320
    );
  ix54672z17194 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romeaddro4_s(2),
      ADR2 => VCC,
      ADR3 => romeaddro4_s(1),
      O => nx54672z324
    );
  ix54672z23702 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romeaddro4_s(3),
      O => U1_ROME4_modgen_rom_ix2_nx_rm64_16_l
    );
  ix54672z30413 : X_LUT4
    generic map(
      INIT => X"2B0A"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(0),
      ADR2 => romeaddro1_s(1),
      ADR3 => romeaddro1_s(3),
      O => nx54672z90
    );
  ix54672z18483 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(0),
      ADR2 => romeaddro1_s(1),
      ADR3 => romeaddro1_s(3),
      O => nx54672z92
    );
  ix54672z25252 : X_LUT4
    generic map(
      INIT => X"7310"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(0),
      ADR2 => romeaddro1_s(1),
      ADR3 => romeaddro1_s(3),
      O => nx54672z93
    );
  ix54672z2490 : X_LUT4
    generic map(
      INIT => X"0F0A"
    )
    port map (
      ADR0 => romoaddro0_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro0_s(3),
      ADR3 => romoaddro0_s(0),
      O => nx54672z654
    );
  ix54672z39940 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => romeaddro1_s(2),
      ADR1 => romeaddro1_s(0),
      ADR2 => romeaddro1_s(1),
      ADR3 => romeaddro1_s(3),
      O => nx54672z89
    );
  ix54672z2285 : X_LUT4
    generic map(
      INIT => X"0202"
    )
    port map (
      ADR0 => romoaddro0_s(2),
      ADR1 => romoaddro0_s(1),
      ADR2 => romoaddro0_s(3),
      ADR3 => VCC,
      O => nx54672z651
    );
  ix54672z1983 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romoaddro0_s(2),
      ADR1 => romoaddro0_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro0_s(0),
      O => nx54672z655
    );
  ix54672z25625 : X_LUT4
    generic map(
      INIT => X"08AE"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(2),
      ADR3 => romeaddro5_s(0),
      O => nx54672z353
    );
  ix54672z28890 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro5_s(1),
      ADR1 => romeaddro5_s(2),
      ADR2 => romeaddro5_s(3),
      ADR3 => romeaddro5_s(0),
      O => nx54672z387
    );
  ix54672z30786 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(2),
      ADR3 => romeaddro5_s(0),
      O => nx54672z350
    );
  ix54672z28887 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro5_s(2),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(0),
      ADR3 => romeaddro5_s(3),
      O => U1_ROME5_modgen_rom_ix2_nx_rm64_16_u
    );
  ix54672z14197 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(2),
      ADR3 => VCC,
      O => nx54672z388
    );
  ix54672z2028 : X_LUT4
    generic map(
      INIT => X"00AA"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romeaddro5_s(3),
      O => nx54672z385
    );
  ix54672z17287 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romeaddro5_s(2),
      ADR3 => romeaddro5_s(1),
      O => nx54672z389
    );
  ix54672z15069 : X_LUT4
    generic map(
      INIT => X"5924"
    )
    port map (
      ADR0 => romeaddro3_s(1),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(3),
      ADR3 => romeaddro3_s(2),
      O => nx54672z211
    );
  ix54672z12204 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z234
    );
  ix54672z7918 : X_LUT4
    generic map(
      INIT => X"1C86"
    )
    port map (
      ADR0 => romeaddro3_s(1),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(3),
      ADR3 => romeaddro3_s(2),
      O => nx54672z208
    );
  ix54672z3862 : X_LUT4
    generic map(
      INIT => X"7130"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z232
    );
  ix54672z14109 : X_LUT4
    generic map(
      INIT => X"20BA"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z235
    );
  ix54672z18562 : X_LUT4
    generic map(
      INIT => X"2B02"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z458
    );
  ix54672z61437 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z231
    );
  ix54672z14433 : X_LUT4
    generic map(
      INIT => X"20BA"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z459
    );
  ix54672z21526 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(2),
      ADR3 => romeaddro5_s(3),
      O => nx54672z344
    );
  ix54672z7529 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(2),
      ADR2 => romeaddro5_s(0),
      ADR3 => romeaddro5_s(1),
      O => nx54672z337
    );
  ix54672z15255 : X_LUT4
    generic map(
      INIT => X"429C"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(2),
      ADR2 => romeaddro5_s(0),
      ADR3 => romeaddro5_s(1),
      O => nx54672z341
    );
  ix54672z12366 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(2),
      ADR3 => romeaddro5_s(3),
      O => nx54672z346
    );
  ix54672z8104 : X_LUT4
    generic map(
      INIT => X"6158"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(2),
      ADR2 => romeaddro5_s(0),
      ADR3 => romeaddro5_s(1),
      O => nx54672z338
    );
  ix54672z4027 : X_LUT4
    generic map(
      INIT => X"08AE"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(2),
      ADR3 => romeaddro5_s(3),
      O => nx54672z347
    );
  ix54672z18856 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(0),
      ADR3 => romeaddro5_s(2),
      O => nx54672z352
    );
  ix54672z34847 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(2),
      ADR3 => romeaddro5_s(3),
      O => nx54672z343
    );
  ix54672z40313 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(2),
      ADR3 => romeaddro5_s(0),
      O => nx54672z349
    );
  ix54672z45205 : X_LUT4
    generic map(
      INIT => X"A578"
    )
    port map (
      ADR0 => romoaddro6_s(2),
      ADR1 => romoaddro6_s(1),
      ADR2 => romoaddro6_s(0),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1094
    );
  ix54672z52842 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => romoaddro6_s(2),
      ADR1 => romoaddro6_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro6_s(3),
      O => nx54672z1097
    );
  ix54672z41763 : X_LUT4
    generic map(
      INIT => X"9866"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(3),
      O => nx54672z1017
    );
  ix54672z45093 : X_LUT4
    generic map(
      INIT => X"A56A"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(3),
      O => nx54672z1015
    );
  ix54672z52730 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => romoaddro5_s(2),
      ADR1 => romoaddro5_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro5_s(3),
      O => nx54672z1018
    );
  ix54672z44133 : X_LUT4
    generic map(
      INIT => X"CC02"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(1),
      ADR3 => romoaddro5_s(0),
      O => nx54672z1023
    );
  ix54672z58444 : X_LUT4
    generic map(
      INIT => X"D992"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(3),
      O => nx54672z1014
    );
  ix54672z22982 : X_LUT4
    generic map(
      INIT => X"22B2"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(1),
      ADR3 => romoaddro5_s(0),
      O => nx54672z1020
    );
  ix54672z62286 : X_LUT4
    generic map(
      INIT => X"F880"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(1),
      ADR3 => romoaddro5_s(0),
      O => nx54672z1024
    );
  ix54672z64775 : X_LUT4
    generic map(
      INIT => X"DD44"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => VCC,
      ADR3 => romoaddro3_s(3),
      O => nx54672z854
    );
  ix54672z43910 : X_LUT4
    generic map(
      INIT => X"C1C0"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(0),
      ADR3 => romoaddro3_s(3),
      O => nx54672z865
    );
  ix54672z27960 : X_LUT4
    generic map(
      INIT => X"3E96"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(0),
      O => nx54672z790
    );
  ix54672z23038 : X_LUT4
    generic map(
      INIT => X"0C70"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(0),
      ADR3 => romoaddro3_s(3),
      O => nx54672z851
    );
  ix54672z22759 : X_LUT4
    generic map(
      INIT => X"3B02"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(0),
      ADR3 => romoaddro3_s(3),
      O => nx54672z862
    );
  ix54672z62063 : X_LUT4
    generic map(
      INIT => X"E8A0"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(0),
      ADR3 => romoaddro3_s(3),
      O => nx54672z866
    );
  ix54672z29417 : X_LUT4
    generic map(
      INIT => X"4BB4"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(1),
      O => nx54672z795
    );
  ix54672z21208 : X_LUT4
    generic map(
      INIT => X"459A"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(0),
      O => nx54672z792
    );
  ix54672z38420 : X_LUT4
    generic map(
      INIT => X"A244"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(0),
      ADR3 => romoaddro3_s(3),
      O => nx54672z863
    );
  ix54672z36837 : X_LUT4
    generic map(
      INIT => X"934C"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(0),
      O => nx54672z793
    );
  ix54672z19503 : X_LUT4
    generic map(
      INIT => X"1A86"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(3),
      ADR3 => romoaddro2_s(0),
      O => nx54672z789
    );
  ix54672z40274 : X_LUT4
    generic map(
      INIT => X"B34C"
    )
    port map (
      ADR0 => romoaddro2_s(2),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(0),
      ADR3 => romoaddro2_s(1),
      O => nx54672z798
    );
  ix54672z48353 : X_LUT4
    generic map(
      INIT => X"DD4C"
    )
    port map (
      ADR0 => romoaddro4_s(1),
      ADR1 => romoaddro4_s(0),
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(2),
      O => nx54672z909
    );
  ix54672z59224 : X_LUT4
    generic map(
      INIT => X"A6A6"
    )
    port map (
      ADR0 => romoaddro4_s(3),
      ADR1 => romoaddro4_s(0),
      ADR2 => romoaddro4_s(1),
      ADR3 => VCC,
      O => nx54672z920
    );
  ix54672z55074 : X_LUT4
    generic map(
      INIT => X"AFAE"
    )
    port map (
      ADR0 => romoaddro4_s(1),
      ADR1 => romoaddro4_s(0),
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(2),
      O => nx54672z906
    );
  ix54672z25870 : X_LUT4
    generic map(
      INIT => X"6688"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro4_s(2),
      O => nx54672z962
    );
  ix54672z42959 : X_LUT4
    generic map(
      INIT => X"C3F2"
    )
    port map (
      ADR0 => romoaddro4_s(3),
      ADR1 => romoaddro4_s(0),
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(2),
      O => nx54672z917
    );
  ix54672z14915 : X_LUT4
    generic map(
      INIT => X"2244"
    )
    port map (
      ADR0 => romoaddro4_s(3),
      ADR1 => romoaddro4_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro4_s(2),
      O => nx54672z921
    );
  ix54672z28768 : X_LUT4
    generic map(
      INIT => X"6622"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro4_s(3),
      O => nx54672z926
    );
  ix54672z24452 : X_LUT4
    generic map(
      INIT => X"3322"
    )
    port map (
      ADR0 => romoaddro4_s(3),
      ADR1 => romoaddro4_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro4_s(2),
      O => nx54672z918
    );
  ix54672z52027 : X_LUT4
    generic map(
      INIT => X"CF0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro4_s(1),
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(2),
      O => nx54672z927
    );
  ix54672z23443 : X_LUT4
    generic map(
      INIT => X"0D2C"
    )
    port map (
      ADR0 => romoaddro4_s(1),
      ADR1 => romoaddro4_s(2),
      ADR2 => romoaddro4_s(0),
      ADR3 => romoaddro4_s(3),
      O => nx54672z923
    );
  ix54672z6678 : X_LUT4
    generic map(
      INIT => X"33BC"
    )
    port map (
      ADR0 => romoaddro4_s(1),
      ADR1 => romoaddro4_s(2),
      ADR2 => romoaddro4_s(0),
      ADR3 => romoaddro4_s(3),
      O => nx54672z924
    );
  ix54672z23795 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romeaddro5_s(3),
      ADR2 => VCC,
      ADR3 => romeaddro5_s(0),
      O => U1_ROME5_modgen_rom_ix2_nx_rm64_16_l
    );
  ix54672z58556 : X_LUT4
    generic map(
      INIT => X"CB92"
    )
    port map (
      ADR0 => romoaddro6_s(2),
      ADR1 => romoaddro6_s(1),
      ADR2 => romoaddro6_s(0),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1093
    );
  ix54672z28991 : X_LUT4
    generic map(
      INIT => X"5A0A"
    )
    port map (
      ADR0 => romoaddro6_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1084
    );
  ix54672z11625 : X_LUT4
    generic map(
      INIT => X"2244"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro6_s(0),
      O => nx54672z1090
    );
  ix54672z52250 : X_LUT4
    generic map(
      INIT => X"D4D4"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(1),
      ADR3 => VCC,
      O => nx54672z1085
    );
  ix54672z6901 : X_LUT4
    generic map(
      INIT => X"33E6"
    )
    port map (
      ADR0 => romoaddro6_s(0),
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1082
    );
  ix54672z65110 : X_LUT4
    generic map(
      INIT => X"8E8E"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(1),
      ADR3 => VCC,
      O => nx54672z1091
    );
  ix54672z5732 : X_LUT4
    generic map(
      INIT => X"3118"
    )
    port map (
      ADR0 => romoaddro6_s(1),
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(3),
      ADR3 => romoaddro6_s(0),
      O => nx54672z1087
    );
  ix54672z23373 : X_LUT4
    generic map(
      INIT => X"07C0"
    )
    port map (
      ADR0 => romoaddro6_s(1),
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(3),
      ADR3 => romoaddro6_s(0),
      O => nx54672z1088
    );
  ix54672z41875 : X_LUT4
    generic map(
      INIT => X"C23C"
    )
    port map (
      ADR0 => romoaddro6_s(2),
      ADR1 => romoaddro6_s(1),
      ADR2 => romoaddro6_s(0),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1096
    );
  ix54672z38643 : X_LUT4
    generic map(
      INIT => X"A424"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(1),
      ADR3 => romoaddro5_s(0),
      O => nx54672z1021
    );
  ix54672z25931 : X_LUT4
    generic map(
      INIT => X"666C"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(1),
      ADR3 => romoaddro5_s(3),
      O => nx54672z1033
    );
  ix54672z21543 : X_LUT4
    generic map(
      INIT => X"0DD2"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(0),
      O => nx54672z1029
    );
  ix54672z19838 : X_LUT4
    generic map(
      INIT => X"5294"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(0),
      O => nx54672z1026
    );
  ix54672z37172 : X_LUT4
    generic map(
      INIT => X"934C"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(0),
      O => nx54672z1030
    );
  ix54672z40609 : X_LUT4
    generic map(
      INIT => X"87F0"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(1),
      ADR3 => romoaddro5_s(3),
      O => nx54672z1035
    );
  ix54672z28295 : X_LUT4
    generic map(
      INIT => X"7696"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(0),
      O => nx54672z1027
    );
  ix54672z10934 : X_LUT4
    generic map(
      INIT => X"37C8"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(1),
      ADR3 => romoaddro5_s(3),
      O => nx54672z1036
    );
  ix54672z29752 : X_LUT4
    generic map(
      INIT => X"695A"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(1),
      ADR3 => romoaddro5_s(3),
      O => nx54672z1032
    );
  ix54672z25981 : X_LUT4
    generic map(
      INIT => X"6868"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(0),
      ADR2 => romoaddro5_s(2),
      ADR3 => VCC,
      O => nx54672z1041
    );
  ix54672z6810 : X_LUT4
    generic map(
      INIT => X"5A0A"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(1),
      O => nx54672z1038
    );
  ix54672z41049 : X_LUT4
    generic map(
      INIT => X"9B64"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(3),
      ADR3 => romoaddro3_s(0),
      O => nx54672z836
    );
  ix54672z26781 : X_LUT4
    generic map(
      INIT => X"6868"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(3),
      ADR2 => romoaddro2_s(2),
      ADR3 => VCC,
      O => nx54672z804
    );
  ix54672z54770 : X_LUT4
    generic map(
      INIT => X"A5A6"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(3),
      ADR3 => romoaddro3_s(0),
      O => nx54672z833
    );
  ix54672z41512 : X_LUT4
    generic map(
      INIT => X"9898"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(2),
      ADR3 => VCC,
      O => nx54672z805
    );
  ix54672z6475 : X_LUT4
    generic map(
      INIT => X"4A4A"
    )
    port map (
      ADR0 => romoaddro2_s(3),
      ADR1 => romoaddro2_s(1),
      ADR2 => romoaddro2_s(2),
      ADR3 => VCC,
      O => nx54672z801
    );
  ix54672z54702 : X_LUT4
    generic map(
      INIT => X"CC22"
    )
    port map (
      ADR0 => romoaddro2_s(0),
      ADR1 => romoaddro2_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro2_s(1),
      O => nx54672z802
    );
  ix54672z18763 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(3),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(1),
      O => nx54672z287
    );
  ix54672z40220 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(3),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(1),
      O => nx54672z284
    );
  ix54672z25532 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(3),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(1),
      O => nx54672z288
    );
  ix54672z55177 : X_LUT4
    generic map(
      INIT => X"AFAE"
    )
    port map (
      ADR0 => romoaddro5_s(1),
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(3),
      ADR3 => romoaddro5_s(0),
      O => nx54672z979
    );
  ix54672z41846 : X_LUT4
    generic map(
      INIT => X"F00A"
    )
    port map (
      ADR0 => romoaddro5_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro5_s(0),
      ADR3 => romoaddro5_s(1),
      O => nx54672z1042
    );
  ix54672z55037 : X_LUT4
    generic map(
      INIT => X"AA50"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro5_s(0),
      ADR3 => romoaddro5_s(1),
      O => nx54672z1039
    );
  ix54672z23293 : X_LUT4
    generic map(
      INIT => X"04CC"
    )
    port map (
      ADR0 => romoaddro5_s(1),
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(3),
      ADR3 => romoaddro5_s(0),
      O => nx54672z981
    );
  ix54672z48456 : X_LUT4
    generic map(
      INIT => X"BF22"
    )
    port map (
      ADR0 => romoaddro5_s(2),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(3),
      ADR3 => romoaddro5_s(0),
      O => nx54672z982
    );
  ix54672z23190 : X_LUT4
    generic map(
      INIT => X"3700"
    )
    port map (
      ADR0 => romoaddro4_s(1),
      ADR1 => romoaddro4_s(0),
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(2),
      O => nx54672z908
    );
  ix54672z59939 : X_LUT4
    generic map(
      INIT => X"E000"
    )
    port map (
      ADR0 => romoaddro4_s(1),
      ADR1 => romoaddro4_s(0),
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(2),
      O => nx54672z905
    );
  ix54672z11046 : X_LUT4
    generic map(
      INIT => X"3C78"
    )
    port map (
      ADR0 => romoaddro6_s(0),
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(3),
      ADR3 => romoaddro6_s(1),
      O => nx54672z1115
    );
  ix54672z26093 : X_LUT4
    generic map(
      INIT => X"6868"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(2),
      ADR3 => VCC,
      O => nx54672z1120
    );
  ix54672z26043 : X_LUT4
    generic map(
      INIT => X"666C"
    )
    port map (
      ADR0 => romoaddro6_s(0),
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(3),
      ADR3 => romoaddro6_s(1),
      O => nx54672z1112
    );
  ix54672z6922 : X_LUT4
    generic map(
      INIT => X"55A0"
    )
    port map (
      ADR0 => romoaddro6_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1117
    );
  ix54672z41958 : X_LUT4
    generic map(
      INIT => X"C2C2"
    )
    port map (
      ADR0 => romoaddro6_s(2),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(1),
      ADR3 => VCC,
      O => nx54672z1121
    );
  ix54672z55149 : X_LUT4
    generic map(
      INIT => X"A4A4"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(1),
      ADR3 => VCC,
      O => nx54672z1118
    );
  ix54672z3151 : X_LUT4
    generic map(
      INIT => X"5544"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(2),
      ADR2 => VCC,
      ADR3 => romoaddro6_s(0),
      O => nx54672z1126
    );
  ix54672z2644 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(0),
      O => nx54672z1127
    );
  ix54672z2946 : X_LUT4
    generic map(
      INIT => X"0404"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(1),
      ADR3 => VCC,
      O => nx54672z1123
    );
  ix54672z6699 : X_LUT4
    generic map(
      INIT => X"30CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(2),
      O => nx54672z959
    );
  ix54672z41735 : X_LUT4
    generic map(
      INIT => X"A5A0"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(2),
      O => nx54672z963
    );
  ix54672z54926 : X_LUT4
    generic map(
      INIT => X"F00A"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(3),
      O => nx54672z960
    );
  ix54672z2928 : X_LUT4
    generic map(
      INIT => X"0F0A"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(0),
      O => nx54672z968
    );
  ix54672z2421 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro4_s(0),
      O => nx54672z969
    );
  ix54672z2723 : X_LUT4
    generic map(
      INIT => X"0202"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(1),
      ADR2 => romoaddro4_s(3),
      ADR3 => VCC,
      O => nx54672z965
    );
  ix54672z2658 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romoaddro4_s(3),
      ADR1 => romoaddro4_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro4_s(0),
      O => nx54672z966
    );
  ix54672z4216 : X_LUT4
    generic map(
      INIT => X"0F5A"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(0),
      O => nx54672z974
    );
  ix54672z54967 : X_LUT4
    generic map(
      INIT => X"F50A"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(1),
      O => nx54672z971
    );
  ix54672z10397 : X_LUT4
    generic map(
      INIT => X"555A"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(0),
      O => nx54672z975
    );
  ix54672z24546 : X_LUT4
    generic map(
      INIT => X"05FA"
    )
    port map (
      ADR0 => romoaddro4_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(0),
      O => nx54672z972
    );
  ix54672z25824 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro4_s(2),
      ADR3 => VCC,
      O => nx54672z976
    );
  ix54672z28909 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z977
    );
  ix54672z6771 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romoaddro4_s(2),
      ADR3 => romoaddro4_s(3),
      O => U1_ROMO4_modgen_rom_ix0_nx_rm64_16_u
    );
  ix54672z15952 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro4_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro4_s(3),
      O => U1_ROMO4_modgen_rom_ix0_nx_rm64_16_l
    );
  ix54672z11290 : X_LUT4
    generic map(
      INIT => X"4422"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro3_s(3),
      O => nx54672z853
    );
  ix54672z5397 : X_LUT4
    generic map(
      INIT => X"3118"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(0),
      ADR3 => romoaddro3_s(3),
      O => nx54672z850
    );
  ix54672z30693 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(3),
      ADR2 => romeaddro4_s(2),
      ADR3 => romeaddro4_s(1),
      O => nx54672z285
    );
  ix54672z3955 : X_LUT4
    generic map(
      INIT => X"4F04"
    )
    port map (
      ADR0 => romeaddro4_s(2),
      ADR1 => romeaddro4_s(1),
      ADR2 => romeaddro4_s(3),
      ADR3 => romeaddro4_s(0),
      O => nx54672z297
    );
  ix54672z12737 : X_LUT4
    generic map(
      INIT => X"088E"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(3),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(2),
      O => nx54672z293
    );
  ix54672z7738 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(3),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(2),
      O => nx54672z290
    );
  ix54672z24548 : X_LUT4
    generic map(
      INIT => X"4694"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(3),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(2),
      O => nx54672z294
    );
  ix54672z12297 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => romeaddro4_s(2),
      ADR1 => romeaddro4_s(1),
      ADR2 => romeaddro4_s(3),
      ADR3 => romeaddro4_s(0),
      O => nx54672z299
    );
  ix54672z26613 : X_LUT4
    generic map(
      INIT => X"4B24"
    )
    port map (
      ADR0 => romeaddro4_s(0),
      ADR1 => romeaddro4_s(3),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(2),
      O => nx54672z291
    );
  ix54672z14202 : X_LUT4
    generic map(
      INIT => X"2B22"
    )
    port map (
      ADR0 => romeaddro4_s(2),
      ADR1 => romeaddro4_s(1),
      ADR2 => romeaddro4_s(3),
      ADR3 => romeaddro4_s(0),
      O => nx54672z300
    );
  ix54672z18654 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro3_s(1),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(3),
      ADR3 => romeaddro3_s(2),
      O => nx54672z210
    );
  ix54672z61530 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro4_s(2),
      ADR1 => romeaddro4_s(1),
      ADR2 => romeaddro4_s(3),
      ADR3 => romeaddro4_s(0),
      O => nx54672z296
    );
  ix54672z7343 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => romeaddro3_s(1),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(3),
      ADR3 => romeaddro3_s(2),
      O => nx54672z207
    );
  ix54672z55289 : X_LUT4
    generic map(
      INIT => X"CCFE"
    )
    port map (
      ADR0 => romoaddro6_s(0),
      ADR1 => romoaddro6_s(1),
      ADR2 => romoaddro6_s(2),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1058
    );
  ix54672z41610 : X_LUT4
    generic map(
      INIT => X"C378"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => romoaddro8_s(1),
      ADR2 => romoaddro8_s(0),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1231
    );
  ix54672z23405 : X_LUT4
    generic map(
      INIT => X"5070"
    )
    port map (
      ADR0 => romoaddro6_s(0),
      ADR1 => romoaddro6_s(1),
      ADR2 => romoaddro6_s(2),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1060
    );
  ix54672z57071 : X_LUT4
    generic map(
      INIT => X"999C"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => romoaddro8_s(1),
      ADR2 => romoaddro8_s(0),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1228
    );
  ix54672z48568 : X_LUT4
    generic map(
      INIT => X"B2BA"
    )
    port map (
      ADR0 => romoaddro6_s(0),
      ADR1 => romoaddro6_s(1),
      ADR2 => romoaddro6_s(2),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1061
    );
  ix54672z25936 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romoaddro5_s(2),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romoaddro5_s(0),
      O => nx54672z1055
    );
  ix54672z6883 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro5_s(2),
      ADR3 => VCC,
      O => U1_ROMO5_modgen_rom_ix0_nx_rm64_16_u
    );
  ix54672z29021 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro5_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro5_s(0),
      O => nx54672z1056
    );
  ix54672z55219 : X_LUT4
    generic map(
      INIT => X"F01E"
    )
    port map (
      ADR0 => romoaddro7_s(2),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1149
    );
  ix54672z26103 : X_LUT4
    generic map(
      INIT => X"666A"
    )
    port map (
      ADR0 => romoaddro7_s(2),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1151
    );
  ix54672z59561 : X_LUT4
    generic map(
      INIT => X"B4B4"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(3),
      ADR3 => VCC,
      O => nx54672z1157
    );
  ix54672z41498 : X_LUT4
    generic map(
      INIT => X"96C6"
    )
    port map (
      ADR0 => romoaddro7_s(2),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1152
    );
  ix54672z10395 : X_LUT4
    generic map(
      INIT => X"3C68"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(3),
      ADR3 => romoaddro3_s(0),
      O => nx54672z832
    );
  ix54672z15252 : X_LUT4
    generic map(
      INIT => X"500A"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro7_s(3),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1158
    );
  ix54672z25654 : X_LUT4
    generic map(
      INIT => X"36CC"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(3),
      ADR3 => romoaddro3_s(0),
      O => nx54672z835
    );
  ix54672z43296 : X_LUT4
    generic map(
      INIT => X"99BA"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(3),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1154
    );
  ix54672z24789 : X_LUT4
    generic map(
      INIT => X"5550"
    )
    port map (
      ADR0 => romoaddro7_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro7_s(3),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1155
    );
  ix54672z8383 : X_LUT4
    generic map(
      INIT => X"5294"
    )
    port map (
      ADR0 => romeaddro8_s(3),
      ADR1 => romeaddro8_s(1),
      ADR2 => romeaddro8_s(0),
      ADR3 => romeaddro8_s(2),
      O => nx54672z533
    );
  ix54672z61584 : X_LUT4
    generic map(
      INIT => X"E880"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(1),
      ADR3 => romeaddro8_s(3),
      O => nx54672z526
    );
  ix54672z14534 : X_LUT4
    generic map(
      INIT => X"0A8E"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(1),
      ADR3 => romeaddro8_s(3),
      O => nx54672z530
    );
  ix54672z19119 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => romeaddro8_s(3),
      ADR1 => romeaddro8_s(1),
      ADR2 => romeaddro8_s(0),
      ADR3 => romeaddro8_s(2),
      O => nx54672z535
    );
  ix54672z4287 : X_LUT4
    generic map(
      INIT => X"40DC"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(1),
      ADR3 => romeaddro8_s(3),
      O => nx54672z527
    );
  ix54672z15534 : X_LUT4
    generic map(
      INIT => X"6318"
    )
    port map (
      ADR0 => romeaddro8_s(3),
      ADR1 => romeaddro8_s(1),
      ADR2 => romeaddro8_s(0),
      ADR3 => romeaddro8_s(2),
      O => nx54672z536
    );
  ix54672z12645 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(1),
      ADR3 => romeaddro8_s(3),
      O => nx54672z541
    );
  ix54672z7808 : X_LUT4
    generic map(
      INIT => X"1668"
    )
    port map (
      ADR0 => romeaddro8_s(3),
      ADR1 => romeaddro8_s(1),
      ADR2 => romeaddro8_s(0),
      ADR3 => romeaddro8_s(2),
      O => nx54672z532
    );
  ix54672z35126 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(1),
      ADR3 => romeaddro8_s(3),
      O => nx54672z538
    );
  ix54672z28407 : X_LUT4
    generic map(
      INIT => X"65DA"
    )
    port map (
      ADR0 => romoaddro6_s(1),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(2),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1106
    );
  ix54672z23094 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => romoaddro6_s(2),
      ADR1 => romoaddro6_s(3),
      ADR2 => romoaddro6_s(0),
      ADR3 => romoaddro6_s(1),
      O => nx54672z1099
    );
  ix54672z62398 : X_LUT4
    generic map(
      INIT => X"F880"
    )
    port map (
      ADR0 => romoaddro6_s(2),
      ADR1 => romoaddro6_s(3),
      ADR2 => romoaddro6_s(0),
      ADR3 => romoaddro6_s(1),
      O => nx54672z1103
    );
  ix54672z21655 : X_LUT4
    generic map(
      INIT => X"293C"
    )
    port map (
      ADR0 => romoaddro6_s(1),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(2),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1108
    );
  ix54672z38755 : X_LUT4
    generic map(
      INIT => X"C422"
    )
    port map (
      ADR0 => romoaddro6_s(2),
      ADR1 => romoaddro6_s(3),
      ADR2 => romoaddro6_s(0),
      ADR3 => romoaddro6_s(1),
      O => nx54672z1100
    );
  ix54672z37284 : X_LUT4
    generic map(
      INIT => X"8666"
    )
    port map (
      ADR0 => romoaddro6_s(1),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(2),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1109
    );
  ix54672z40721 : X_LUT4
    generic map(
      INIT => X"8F70"
    )
    port map (
      ADR0 => romoaddro6_s(0),
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(3),
      ADR3 => romoaddro6_s(1),
      O => nx54672z1114
    );
  ix54672z19950 : X_LUT4
    generic map(
      INIT => X"24D2"
    )
    port map (
      ADR0 => romoaddro6_s(1),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(2),
      ADR3 => romoaddro6_s(3),
      O => nx54672z1105
    );
  ix54672z29864 : X_LUT4
    generic map(
      INIT => X"659A"
    )
    port map (
      ADR0 => romoaddro6_s(0),
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(3),
      ADR3 => romoaddro6_s(1),
      O => nx54672z1111
    );
  ix54672z9333 : X_LUT4
    generic map(
      INIT => X"294A"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(2),
      ADR3 => romeaddro7_s(0),
      O => nx54672z507
    );
  ix54672z19146 : X_LUT4
    generic map(
      INIT => X"2B42"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(0),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(2),
      O => nx54672z512
    );
  ix54672z24848 : X_LUT4
    generic map(
      INIT => X"18C6"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(2),
      ADR3 => romeaddro7_s(0),
      O => nx54672z504
    );
  ix54672z34523 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(0),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(2),
      O => nx54672z509
    );
  ix54672z28049 : X_LUT4
    generic map(
      INIT => X"693C"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(0),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(2),
      O => nx54672z513
    );
  ix54672z11851 : X_LUT4
    generic map(
      INIT => X"0A50"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(0),
      O => nx54672z1248
    );
  ix54672z17546 : X_LUT4
    generic map(
      INIT => X"59A6"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(0),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(2),
      O => nx54672z510
    );
  ix54672z65336 : X_LUT4
    generic map(
      INIT => X"AF0A"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1249
    );
  ix54672z5958 : X_LUT4
    generic map(
      INIT => X"3118"
    )
    port map (
      ADR0 => romoaddro8_s(1),
      ADR1 => romoaddro8_s(2),
      ADR2 => romoaddro8_s(3),
      ADR3 => romoaddro8_s(0),
      O => nx54672z1245
    );
  ix54672z23599 : X_LUT4
    generic map(
      INIT => X"07C0"
    )
    port map (
      ADR0 => romoaddro8_s(1),
      ADR1 => romoaddro8_s(2),
      ADR2 => romoaddro8_s(3),
      ADR3 => romoaddro8_s(0),
      O => nx54672z1246
    );
  ix54672z42101 : X_LUT4
    generic map(
      INIT => X"9964"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => romoaddro8_s(0),
      ADR2 => romoaddro8_s(2),
      ADR3 => romoaddro8_s(1),
      O => nx54672z1254
    );
  ix54672z14295 : X_LUT4
    generic map(
      INIT => X"7310"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(0),
      ADR3 => romeaddro5_s(2),
      O => nx54672z365
    );
  ix54672z18880 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => romeaddro5_s(2),
      ADR1 => romeaddro5_s(0),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(3),
      O => nx54672z370
    );
  ix54672z4048 : X_LUT4
    generic map(
      INIT => X"50D4"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(0),
      ADR3 => romeaddro5_s(2),
      O => nx54672z362
    );
  ix54672z25646 : X_LUT4
    generic map(
      INIT => X"7310"
    )
    port map (
      ADR0 => romeaddro5_s(2),
      ADR1 => romeaddro5_s(0),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(3),
      O => nx54672z368
    );
  ix54672z5051 : X_LUT4
    generic map(
      INIT => X"50D4"
    )
    port map (
      ADR0 => romeaddro5_s(2),
      ADR1 => romeaddro5_s(0),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(3),
      O => nx54672z371
    );
  ix54672z23413 : X_LUT4
    generic map(
      INIT => X"1F00"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(1),
      ADR2 => romoaddro6_s(0),
      ADR3 => romoaddro6_s(2),
      O => nx54672z1066
    );
  ix54672z34321 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro5_s(2),
      ADR1 => romeaddro5_s(0),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(3),
      O => nx54672z367
    );
  ix54672z60162 : X_LUT4
    generic map(
      INIT => X"A800"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(1),
      ADR2 => romoaddro6_s(0),
      ADR3 => romoaddro6_s(2),
      O => nx54672z1063
    );
  ix54672z55297 : X_LUT4
    generic map(
      INIT => X"DDDC"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(1),
      ADR2 => romoaddro6_s(0),
      ADR3 => romoaddro6_s(2),
      O => nx54672z1064
    );
  ix54672z48576 : X_LUT4
    generic map(
      INIT => X"F370"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(1),
      ADR2 => romoaddro6_s(0),
      ADR3 => romoaddro6_s(2),
      O => nx54672z1067
    );
  ix54672z44245 : X_LUT4
    generic map(
      INIT => X"A0A4"
    )
    port map (
      ADR0 => romoaddro6_s(2),
      ADR1 => romoaddro6_s(3),
      ADR2 => romoaddro6_s(0),
      ADR3 => romoaddro6_s(1),
      O => nx54672z1102
    );
  ix54672z15026 : X_LUT4
    generic map(
      INIT => X"2244"
    )
    port map (
      ADR0 => romoaddro5_s(2),
      ADR1 => romoaddro5_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro5_s(3),
      O => nx54672z1000
    );
  ix54672z28879 : X_LUT4
    generic map(
      INIT => X"6622"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => romoaddro5_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro5_s(3),
      O => nx54672z1005
    );
  ix54672z24563 : X_LUT4
    generic map(
      INIT => X"3322"
    )
    port map (
      ADR0 => romoaddro5_s(2),
      ADR1 => romoaddro5_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro5_s(3),
      O => nx54672z997
    );
  ix54672z52138 : X_LUT4
    generic map(
      INIT => X"88EE"
    )
    port map (
      ADR0 => romoaddro5_s(2),
      ADR1 => romoaddro5_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro5_s(3),
      O => nx54672z1006
    );
  ix54672z3039 : X_LUT4
    generic map(
      INIT => X"0F0A"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro5_s(3),
      ADR3 => romoaddro5_s(2),
      O => nx54672z1047
    );
  ix54672z23554 : X_LUT4
    generic map(
      INIT => X"5158"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(3),
      O => nx54672z1002
    );
  ix54672z6789 : X_LUT4
    generic map(
      INIT => X"0FDA"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(3),
      O => nx54672z1003
    );
  ix54672z2834 : X_LUT4
    generic map(
      INIT => X"000A"
    )
    port map (
      ADR0 => romoaddro5_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro5_s(3),
      ADR3 => romoaddro5_s(1),
      O => nx54672z1044
    );
  ix54672z2532 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(1),
      O => nx54672z1048
    );
  ix54672z18655 : X_LUT4
    generic map(
      INIT => X"20B2"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(3),
      ADR2 => romeaddro8_s(1),
      ADR3 => romeaddro8_s(0),
      O => nx54672z523
    );
  ix54672z4279 : X_LUT4
    generic map(
      INIT => X"7310"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(3),
      ADR2 => romeaddro8_s(1),
      ADR3 => romeaddro8_s(0),
      O => nx54672z521
    );
  ix54672z14526 : X_LUT4
    generic map(
      INIT => X"2B0A"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(3),
      ADR2 => romeaddro8_s(1),
      ADR3 => romeaddro8_s(0),
      O => nx54672z524
    );
  ix54672z26706 : X_LUT4
    generic map(
      INIT => X"4B24"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => romeaddro5_s(3),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(2),
      O => nx54672z356
    );
  ix54672z12830 : X_LUT4
    generic map(
      INIT => X"088E"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => romeaddro5_s(3),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(2),
      O => nx54672z358
    );
  ix54672z24641 : X_LUT4
    generic map(
      INIT => X"4694"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => romeaddro5_s(3),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(2),
      O => nx54672z359
    );
  ix54672z61623 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(0),
      ADR3 => romeaddro5_s(2),
      O => nx54672z361
    );
  ix54672z12390 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => romeaddro5_s(3),
      ADR1 => romeaddro5_s(1),
      ADR2 => romeaddro5_s(0),
      ADR3 => romeaddro5_s(2),
      O => nx54672z364
    );
  ix54672z7831 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => romeaddro5_s(0),
      ADR1 => romeaddro5_s(3),
      ADR2 => romeaddro5_s(1),
      ADR3 => romeaddro5_s(2),
      O => nx54672z355
    );
  ix54672z25718 : X_LUT4
    generic map(
      INIT => X"0A8E"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(1),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(2),
      O => nx54672z418
    );
  ix54672z12923 : X_LUT4
    generic map(
      INIT => X"20B2"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(2),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(1),
      O => nx54672z423
    );
  ix54672z30879 : X_LUT4
    generic map(
      INIT => X"3B02"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(1),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(2),
      O => nx54672z415
    );
  ix54672z26799 : X_LUT4
    generic map(
      INIT => X"18C6"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(2),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(1),
      O => nx54672z421
    );
  ix54672z24734 : X_LUT4
    generic map(
      INIT => X"294A"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(2),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(1),
      O => nx54672z424
    );
  ix54672z12483 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(1),
      O => nx54672z429
    );
  ix54672z7924 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(2),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(1),
      O => nx54672z420
    );
  ix54672z61716 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(1),
      O => nx54672z426
    );
  ix54672z4141 : X_LUT4
    generic map(
      INIT => X"4D44"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(1),
      O => nx54672z427
    );
  ix54672z14388 : X_LUT4
    generic map(
      INIT => X"40F4"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(1),
      O => nx54672z430
    );
  ix54672z18663 : X_LUT4
    generic map(
      INIT => X"20B2"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(1),
      ADR3 => romeaddro8_s(3),
      O => nx54672z529
    );
  ix54672z2881 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(0),
      O => nx54672z1124
    );
  ix54672z23301 : X_LUT4
    generic map(
      INIT => X"02AA"
    )
    port map (
      ADR0 => romoaddro5_s(2),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(3),
      ADR3 => romoaddro5_s(0),
      O => nx54672z987
    );
  ix54672z54993 : X_LUT4
    generic map(
      INIT => X"999C"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(0),
      O => nx54672z991
    );
  ix54672z60050 : X_LUT4
    generic map(
      INIT => X"A080"
    )
    port map (
      ADR0 => romoaddro5_s(2),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(3),
      ADR3 => romoaddro5_s(0),
      O => nx54672z984
    );
  ix54672z48464 : X_LUT4
    generic map(
      INIT => X"BF22"
    )
    port map (
      ADR0 => romoaddro5_s(2),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(3),
      ADR3 => romoaddro5_s(0),
      O => nx54672z988
    );
  ix54672z25877 : X_LUT4
    generic map(
      INIT => X"1EF0"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(0),
      O => nx54672z993
    );
  ix54672z55185 : X_LUT4
    generic map(
      INIT => X"CFCE"
    )
    port map (
      ADR0 => romoaddro5_s(2),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(3),
      ADR3 => romoaddro5_s(0),
      O => nx54672z985
    );
  ix54672z41272 : X_LUT4
    generic map(
      INIT => X"C738"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(0),
      O => nx54672z994
    );
  ix54672z59335 : X_LUT4
    generic map(
      INIT => X"DD22"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => romoaddro5_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro5_s(3),
      O => nx54672z999
    );
  ix54672z10618 : X_LUT4
    generic map(
      INIT => X"5A68"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(0),
      O => nx54672z990
    );
  ix54672z43070 : X_LUT4
    generic map(
      INIT => X"9D9C"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => romoaddro5_s(1),
      ADR2 => romoaddro5_s(2),
      ADR3 => romoaddro5_s(3),
      O => nx54672z996
    );
  ix54672z4306 : X_LUT4
    generic map(
      INIT => X"40DC"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(1),
      ADR3 => romeaddro8_s(3),
      O => nx54672z542
    );
  ix54672z3907 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => romeaddro4_s(3),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(0),
      O => nx54672z261
    );
  ix54672z19135 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(2),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z547
    );
  ix54672z21805 : X_LUT4
    generic map(
      INIT => X"7150"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(1),
      ADR3 => romeaddro8_s(3),
      O => nx54672z539
    );
  ix54672z40592 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(2),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z544
    );
  ix54672z25904 : X_LUT4
    generic map(
      INIT => X"7150"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(2),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z548
    );
  ix54672z18283 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => romeaddro4_s(3),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(0),
      O => nx54672z263
    );
  ix54672z31065 : X_LUT4
    generic map(
      INIT => X"40DC"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(2),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z545
    );
  ix54672z14154 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => romeaddro4_s(3),
      ADR1 => romeaddro4_s(2),
      ADR2 => romeaddro4_s(1),
      ADR3 => romeaddro4_s(0),
      O => nx54672z264
    );
  ix54672z2769 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romoaddro5_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro5_s(3),
      ADR3 => romoaddro5_s(1),
      O => nx54672z1045
    );
  ix54672z5813 : X_LUT4
    generic map(
      INIT => X"03FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro5_s(2),
      ADR2 => romoaddro5_s(0),
      ADR3 => romoaddro5_s(3),
      O => nx54672z1053
    );
  ix54672z55522 : X_LUT4
    generic map(
      INIT => X"CFCE"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => romoaddro8_s(1),
      ADR2 => romoaddro8_s(3),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1222
    );
  ix54672z55078 : X_LUT4
    generic map(
      INIT => X"AA66"
    )
    port map (
      ADR0 => romoaddro5_s(1),
      ADR1 => romoaddro5_s(2),
      ADR2 => VCC,
      ADR3 => romoaddro5_s(3),
      O => nx54672z1050
    );
  ix54672z10509 : X_LUT4
    generic map(
      INIT => X"11EE"
    )
    port map (
      ADR0 => romoaddro5_s(1),
      ADR1 => romoaddro5_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro5_s(2),
      O => nx54672z1054
    );
  ix54672z24657 : X_LUT4
    generic map(
      INIT => X"3366"
    )
    port map (
      ADR0 => romoaddro5_s(1),
      ADR1 => romoaddro5_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro5_s(3),
      O => nx54672z1051
    );
  ix54672z23638 : X_LUT4
    generic map(
      INIT => X"5700"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => romoaddro8_s(1),
      ADR2 => romoaddro8_s(3),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1224
    );
  ix54672z48801 : X_LUT4
    generic map(
      INIT => X"BB2A"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => romoaddro8_s(1),
      ADR2 => romoaddro8_s(3),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1225
    );
  ix54672z60387 : X_LUT4
    generic map(
      INIT => X"E000"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => romoaddro8_s(1),
      ADR2 => romoaddro8_s(3),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1221
    );
  ix54672z26215 : X_LUT4
    generic map(
      INIT => X"1FE0"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => romoaddro8_s(1),
      ADR2 => romoaddro8_s(0),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1230
    );
  ix54672z10955 : X_LUT4
    generic map(
      INIT => X"56A8"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => romoaddro8_s(1),
      ADR2 => romoaddro8_s(0),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1227
    );
  ix54672z44982 : X_LUT4
    generic map(
      INIT => X"A758"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(1),
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(0),
      O => nx54672z936
    );
  ix54672z30972 : X_LUT4
    generic map(
      INIT => X"08AE"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z480
    );
  ix54672z35033 : X_LUT4
    generic map(
      INIT => X"8116"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z473
    );
  ix54672z4213 : X_LUT4
    generic map(
      INIT => X"7130"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z477
    );
  ix54672z19042 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z482
    );
  ix54672z21712 : X_LUT4
    generic map(
      INIT => X"5D04"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z474
    );
  ix54672z25811 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z483
    );
  ix54672z13016 : X_LUT4
    generic map(
      INIT => X"40D4"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(0),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(2),
      O => nx54672z488
    );
  ix54672z40499 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z479
    );
  ix54672z8017 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(0),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(2),
      O => nx54672z485
    );
  ix54672z5144 : X_LUT4
    generic map(
      INIT => X"4F04"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(1),
      O => nx54672z436
    );
  ix54672z26985 : X_LUT4
    generic map(
      INIT => X"5294"
    )
    port map (
      ADR0 => romeaddro8_s(1),
      ADR1 => romeaddro8_s(3),
      ADR2 => romeaddro8_s(2),
      ADR3 => romeaddro8_s(0),
      O => nx54672z551
    );
  ix54672z12499 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(2),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(3),
      O => nx54672z441
    );
  ix54672z25739 : X_LUT4
    generic map(
      INIT => X"2B22"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(1),
      O => nx54672z433
    );
  ix54672z61732 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(2),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(3),
      O => nx54672z438
    );
  ix54672z9240 : X_LUT4
    generic map(
      INIT => X"2692"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(2),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(3),
      O => nx54672z442
    );
  ix54672z13109 : X_LUT4
    generic map(
      INIT => X"4D04"
    )
    port map (
      ADR0 => romeaddro8_s(1),
      ADR1 => romeaddro8_s(3),
      ADR2 => romeaddro8_s(2),
      ADR3 => romeaddro8_s(0),
      O => nx54672z553
    );
  ix54672z24755 : X_LUT4
    generic map(
      INIT => X"2D42"
    )
    port map (
      ADR0 => romeaddro6_s(1),
      ADR1 => romeaddro6_s(2),
      ADR2 => romeaddro6_s(0),
      ADR3 => romeaddro6_s(3),
      O => nx54672z439
    );
  ix54672z24920 : X_LUT4
    generic map(
      INIT => X"18C6"
    )
    port map (
      ADR0 => romeaddro8_s(1),
      ADR1 => romeaddro8_s(3),
      ADR2 => romeaddro8_s(2),
      ADR3 => romeaddro8_s(0),
      O => nx54672z554
    );
  ix54672z8110 : X_LUT4
    generic map(
      INIT => X"177E"
    )
    port map (
      ADR0 => romeaddro8_s(1),
      ADR1 => romeaddro8_s(3),
      ADR2 => romeaddro8_s(2),
      ADR3 => romeaddro8_s(0),
      O => nx54672z550
    );
  ix54672z12669 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => romeaddro8_s(1),
      ADR1 => romeaddro8_s(3),
      ADR2 => romeaddro8_s(0),
      ADR3 => romeaddro8_s(2),
      O => nx54672z559
    );
  ix54672z61453 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro3_s(0),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(2),
      ADR3 => romeaddro3_s(1),
      O => nx54672z243
    );
  ix54672z8961 : X_LUT4
    generic map(
      INIT => X"2D42"
    )
    port map (
      ADR0 => romeaddro3_s(0),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(2),
      ADR3 => romeaddro3_s(1),
      O => nx54672z247
    );
  ix54672z28704 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => nx54672z257
    );
  ix54672z24476 : X_LUT4
    generic map(
      INIT => X"4964"
    )
    port map (
      ADR0 => romeaddro3_s(0),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(2),
      ADR3 => romeaddro3_s(1),
      O => nx54672z244
    );
  ix54672z14011 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romeaddro3_s(2),
      ADR3 => romeaddro3_s(1),
      O => nx54672z258
    );
  ix54672z18973 : X_LUT4
    generic map(
      INIT => X"6118"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(1),
      O => nx54672z435
    );
  ix54672z28701 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro3_s(2),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => romeaddro3_s(1),
      O => U1_ROME3_modgen_rom_ix2_nx_rm64_16_u
    );
  ix54672z1842 : X_LUT4
    generic map(
      INIT => X"3030"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(0),
      ADR3 => VCC,
      O => nx54672z255
    );
  ix54672z34414 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro6_s(3),
      ADR1 => romeaddro6_s(0),
      ADR2 => romeaddro6_s(2),
      ADR3 => romeaddro6_s(1),
      O => nx54672z432
    );
  ix54672z16064 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => romoaddro5_s(3),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => romoaddro5_s(1),
      O => U1_ROMO5_modgen_rom_ix0_nx_rm64_16_l
    );
  ix54672z11402 : X_LUT4
    generic map(
      INIT => X"4422"
    )
    port map (
      ADR0 => romoaddro4_s(1),
      ADR1 => romoaddro4_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro4_s(0),
      O => nx54672z932
    );
  ix54672z12552 : X_LUT4
    generic map(
      INIT => X"4294"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z476
    );
  ix54672z64887 : X_LUT4
    generic map(
      INIT => X"DD44"
    )
    port map (
      ADR0 => romoaddro4_s(1),
      ADR1 => romoaddro4_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro4_s(2),
      O => nx54672z933
    );
  ix54672z41652 : X_LUT4
    generic map(
      INIT => X"C32C"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(1),
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(0),
      O => nx54672z938
    );
  ix54672z5509 : X_LUT4
    generic map(
      INIT => X"108E"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(2),
      O => nx54672z929
    );
  ix54672z23150 : X_LUT4
    generic map(
      INIT => X"4622"
    )
    port map (
      ADR0 => romoaddro4_s(0),
      ADR1 => romoaddro4_s(3),
      ADR2 => romoaddro4_s(1),
      ADR3 => romoaddro4_s(2),
      O => nx54672z930
    );
  ix54672z58333 : X_LUT4
    generic map(
      INIT => X"C9B2"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(1),
      ADR2 => romoaddro4_s(3),
      ADR3 => romoaddro4_s(0),
      O => nx54672z935
    );
  ix54672z52619 : X_LUT4
    generic map(
      INIT => X"9696"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(1),
      ADR2 => romoaddro4_s(3),
      ADR3 => VCC,
      O => nx54672z939
    );
  odv1_OUTPUT_OTCLK1INV_7629 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => odv1_OUTPUT_OTCLK1INV
    );
  odv1_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramwe_repl0,
      O => odv1_O
    );
  odv1_OUTPUT_OFF_OCEINV_7630 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_NOT_rtlcs2,
      O => odv1_OUTPUT_OFF_OCEINV
    );
  odv1_OUTPUT_OFF_O1INV_7631 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => odv1_OUTPUT_OFF_O1INV
    );
  U_DCT1D_reg_ramwe_s_repl0 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => odv1_OUTPUT_OFF_O1INV,
      CE => odv1_OUTPUT_OFF_OCEINV,
      CLK => odv1_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => odv1_OUTPUT_OFF_OFF1_RST,
      O => ramwe_repl0
    );
  odv1_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => odv1_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => odv1_OUTPUT_OFF_OFF1_RST
    );
  odv1_OUTPUT_OFF_OFF1_RSTAND_7632 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => odv1_OUTPUT_OFF_OFF1_RSTAND
    );
  dcti_0_IFF_IFF1_RSTOR : X_OR2
    port map (
      I0 => dcti_0_IFF_ISR_USED,
      I1 => GSR,
      O => dcti_0_IFF_IFF1_RST
    );
  U_DCT1D_reg_latchbuf_reg_7_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcti_0_IFF_IFFDMUX,
      CE => dcti_0_IFF_ICEINV,
      CLK => dcti_0_IFF_ICLK1INV,
      SET => GND,
      RST => dcti_0_IFF_IFF1_RST,
      O => U_DCT1D_latchbuf_reg_7_Q(0)
    );
  dcti_0_IFF_IFFDMUX_7633 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti_0_INBUF,
      O => dcti_0_IFF_IFFDMUX
    );
  dcti_0_IFF_ISR_USED_7634 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcti_0_IFF_ISR_USED
    );
  dcti_0_IFF_ICLK1INV_7635 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcti_0_IFF_ICLK1INV
    );
  dcti_0_IFF_ICEINV_7636 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => dcti_0_IFF_ICEINV
    );
  dcti_1_IFF_IFFDMUX_7637 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti_1_INBUF,
      O => dcti_1_IFF_IFFDMUX
    );
  dcti_1_IFF_ICLK1INV_7638 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcti_1_IFF_ICLK1INV
    );
  dcti_1_IFF_ICEINV_7639 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => dcti_1_IFF_ICEINV
    );
  U_DCT1D_reg_latchbuf_reg_7_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcti_1_IFF_IFFDMUX,
      CE => dcti_1_IFF_ICEINV,
      CLK => dcti_1_IFF_ICLK1INV,
      SET => GND,
      RST => dcti_1_IFF_IFF1_RST,
      O => U_DCT1D_latchbuf_reg_7_Q(1)
    );
  dcti_1_IFF_IFF1_RSTOR : X_OR2
    port map (
      I0 => dcti_1_IFF_IFF1_RSTAND,
      I1 => GSR,
      O => dcti_1_IFF_IFF1_RST
    );
  dcti_1_IFF_IFF1_RSTAND_7640 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcti_1_IFF_IFF1_RSTAND
    );
  ix54672z24827 : X_LUT4
    generic map(
      INIT => X"3492"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(0),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(2),
      O => nx54672z489
    );
  ix54672z25832 : X_LUT4
    generic map(
      INIT => X"4D0C"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z498
    );
  ix54672z12576 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => romeaddro7_s(0),
      ADR1 => romeaddro7_s(2),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(1),
      O => nx54672z494
    );
  ix54672z26892 : X_LUT4
    generic map(
      INIT => X"6518"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(0),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(2),
      O => nx54672z486
    );
  ix54672z61809 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro7_s(0),
      ADR1 => romeaddro7_s(2),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(1),
      O => nx54672z491
    );
  ix54672z14481 : X_LUT4
    generic map(
      INIT => X"08CE"
    )
    port map (
      ADR0 => romeaddro7_s(0),
      ADR1 => romeaddro7_s(2),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(1),
      O => nx54672z495
    );
  ix54672z19066 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z500
    );
  ix54672z4234 : X_LUT4
    generic map(
      INIT => X"2B0A"
    )
    port map (
      ADR0 => romeaddro7_s(0),
      ADR1 => romeaddro7_s(2),
      ADR2 => romeaddro7_s(3),
      ADR3 => romeaddro7_s(1),
      O => nx54672z492
    );
  ix54672z5237 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z501
    );
  ix54672z34507 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro7_s(2),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(0),
      ADR3 => romeaddro7_s(1),
      O => nx54672z497
    );
  ix54672z59673 : X_LUT4
    generic map(
      INIT => X"DD22"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => romoaddro8_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro8_s(3),
      O => nx54672z1236
    );
  ix54672z43408 : X_LUT4
    generic map(
      INIT => X"9D9C"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => romoaddro8_s(1),
      ADR2 => romoaddro8_s(2),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1233
    );
  ix54672z15364 : X_LUT4
    generic map(
      INIT => X"2244"
    )
    port map (
      ADR0 => romoaddro8_s(2),
      ADR1 => romoaddro8_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro8_s(3),
      O => nx54672z1237
    );
  ix54672z29217 : X_LUT4
    generic map(
      INIT => X"6644"
    )
    port map (
      ADR0 => romoaddro8_s(1),
      ADR1 => romoaddro8_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro8_s(3),
      O => nx54672z1242
    );
  ix54672z24901 : X_LUT4
    generic map(
      INIT => X"5550"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro8_s(2),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1234
    );
  ix54672z52476 : X_LUT4
    generic map(
      INIT => X"A0FA"
    )
    port map (
      ADR0 => romoaddro8_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1243
    );
  ix54672z29105 : X_LUT4
    generic map(
      INIT => X"3C30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1163
    );
  ix54672z23892 : X_LUT4
    generic map(
      INIT => X"2362"
    )
    port map (
      ADR0 => romoaddro8_s(2),
      ADR1 => romoaddro8_s(0),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1239
    );
  ix54672z7127 : X_LUT4
    generic map(
      INIT => X"55E6"
    )
    port map (
      ADR0 => romoaddro8_s(2),
      ADR1 => romoaddro8_s(0),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1240
    );
  ix54672z23780 : X_LUT4
    generic map(
      INIT => X"5158"
    )
    port map (
      ADR0 => romoaddro7_s(0),
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(2),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1160
    );
  ix54672z52364 : X_LUT4
    generic map(
      INIT => X"C0FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(2),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1164
    );
  ix54672z11739 : X_LUT4
    generic map(
      INIT => X"1818"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => VCC,
      O => nx54672z1169
    );
  ix54672z7015 : X_LUT4
    generic map(
      INIT => X"0FDA"
    )
    port map (
      ADR0 => romoaddro7_s(0),
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(2),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1161
    );
  ix54672z44359 : X_LUT4
    generic map(
      INIT => X"CC10"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => romoaddro7_s(2),
      ADR2 => romoaddro7_s(3),
      ADR3 => romoaddro7_s(0),
      O => nx54672z1181
    );
  ix54672z65224 : X_LUT4
    generic map(
      INIT => X"AF0A"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1170
    );
  ix54672z41989 : X_LUT4
    generic map(
      INIT => X"C23C"
    )
    port map (
      ADR0 => romoaddro7_s(2),
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1175
    );
  ix54672z5846 : X_LUT4
    generic map(
      INIT => X"108E"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1166
    );
  ix54672z23487 : X_LUT4
    generic map(
      INIT => X"2644"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1167
    );
  ix54672z58670 : X_LUT4
    generic map(
      INIT => X"CB92"
    )
    port map (
      ADR0 => romoaddro7_s(2),
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1172
    );
  ix54672z52956 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => romoaddro7_s(2),
      ADR1 => romoaddro7_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro7_s(3),
      O => nx54672z1176
    );
  U_DCT2D_reg_latchbuf_reg_4_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_3_DXMUX,
      CE => U_DCT2D_latchbuf_reg_4_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_4_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_4_3_FFX_RST,
      O => U_DCT2D_latchbuf_reg_4_3_Q
    );
  U_DCT2D_latchbuf_reg_4_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_4_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_4_3_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_4_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_5_DYMUX,
      CE => U_DCT2D_latchbuf_reg_4_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_4_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_4_5_FFY_RST,
      O => U_DCT2D_latchbuf_reg_4_4_Q
    );
  U_DCT2D_latchbuf_reg_4_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_4_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_4_5_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_4_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_5_DXMUX,
      CE => U_DCT2D_latchbuf_reg_4_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_4_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_4_5_FFX_RST,
      O => U_DCT2D_latchbuf_reg_4_5_Q
    );
  U_DCT2D_latchbuf_reg_4_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_4_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_4_5_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_4_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_7_DYMUX,
      CE => U_DCT2D_latchbuf_reg_4_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_4_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_4_7_FFY_RST,
      O => U_DCT2D_latchbuf_reg_4_6_Q
    );
  U_DCT2D_latchbuf_reg_4_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_4_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_4_7_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_4_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_7_DXMUX,
      CE => U_DCT2D_latchbuf_reg_4_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_4_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_4_7_FFX_RST,
      O => U_DCT2D_latchbuf_reg_4_7_Q
    );
  U_DCT2D_latchbuf_reg_4_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_4_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_4_7_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_4_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_10_DYMUX,
      CE => U_DCT2D_latchbuf_reg_4_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_4_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_4_10_FFY_RST,
      O => U_DCT2D_latchbuf_reg_4_8_Q
    );
  U_DCT2D_latchbuf_reg_4_10_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_4_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_4_10_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_4_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_10_DXMUX,
      CE => U_DCT2D_latchbuf_reg_4_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_4_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_4_10_FFX_RST,
      O => U_DCT2D_latchbuf_reg_4_10_Q
    );
  U_DCT2D_latchbuf_reg_4_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_4_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_4_10_FFX_RST
    );
  ix54672z51915 : X_LUT4
    generic map(
      INIT => X"F550"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(1),
      O => nx54672z848
    );
  ix54672z21320 : X_LUT4
    generic map(
      INIT => X"239C"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(3),
      ADR3 => romoaddro3_s(2),
      O => nx54672z871
    );
  ix54672z6566 : X_LUT4
    generic map(
      INIT => X"5E1E"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(1),
      O => nx54672z845
    );
  ix54672z30600 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => romeaddro3_s(1),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(3),
      ADR3 => romeaddro3_s(2),
      O => nx54672z220
    );
  ix54672z28072 : X_LUT4
    generic map(
      INIT => X"5E96"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(3),
      ADR3 => romoaddro3_s(0),
      O => nx54672z869
    );
  ix54672z36949 : X_LUT4
    generic map(
      INIT => X"8666"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(3),
      ADR3 => romoaddro3_s(2),
      O => nx54672z872
    );
  ix54672z18670 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro3_s(1),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(3),
      ADR3 => romeaddro3_s(2),
      O => nx54672z222
    );
  ix54672z19615 : X_LUT4
    generic map(
      INIT => X"1C86"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(3),
      ADR3 => romoaddro3_s(0),
      O => nx54672z868
    );
  ix54672z25439 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => romeaddro3_s(1),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(3),
      ADR3 => romeaddro3_s(2),
      O => nx54672z223
    );
  ix54672z12220 : X_LUT4
    generic map(
      INIT => X"1886"
    )
    port map (
      ADR0 => romeaddro3_s(0),
      ADR1 => romeaddro3_s(3),
      ADR2 => romeaddro3_s(2),
      ADR3 => romeaddro3_s(1),
      O => nx54672z246
    );
  ix54672z40127 : X_LUT4
    generic map(
      INIT => X"9668"
    )
    port map (
      ADR0 => romeaddro3_s(1),
      ADR1 => romeaddro3_s(0),
      ADR2 => romeaddro3_s(3),
      ADR3 => romeaddro3_s(2),
      O => nx54672z219
    );
  ix54672z45319 : X_LUT4
    generic map(
      INIT => X"A578"
    )
    port map (
      ADR0 => romoaddro7_s(2),
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1173
    );
  ix54672z28521 : X_LUT4
    generic map(
      INIT => X"39E6"
    )
    port map (
      ADR0 => romoaddro7_s(2),
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1185
    );
  ix54672z23208 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => romoaddro7_s(2),
      ADR2 => romoaddro7_s(3),
      ADR3 => romoaddro7_s(0),
      O => nx54672z1178
    );
  ix54672z62512 : X_LUT4
    generic map(
      INIT => X"EA80"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => romoaddro7_s(2),
      ADR2 => romoaddro7_s(3),
      ADR3 => romoaddro7_s(0),
      O => nx54672z1182
    );
  ix54672z21769 : X_LUT4
    generic map(
      INIT => X"495A"
    )
    port map (
      ADR0 => romoaddro7_s(2),
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1187
    );
  ix54672z38869 : X_LUT4
    generic map(
      INIT => X"A424"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => romoaddro7_s(2),
      ADR2 => romoaddro7_s(3),
      ADR3 => romoaddro7_s(0),
      O => nx54672z1179
    );
  ix54672z37398 : X_LUT4
    generic map(
      INIT => X"943C"
    )
    port map (
      ADR0 => romoaddro7_s(2),
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1188
    );
  ix54672z28656 : X_LUT4
    generic map(
      INIT => X"22CC"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => romoaddro3_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro3_s(1),
      O => nx54672z847
    );
  ix54672z20064 : X_LUT4
    generic map(
      INIT => X"18A6"
    )
    port map (
      ADR0 => romoaddro7_s(2),
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1184
    );
  ix54672z23331 : X_LUT4
    generic map(
      INIT => X"3432"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(1),
      O => nx54672z844
    );
  ix54672z9426 : X_LUT4
    generic map(
      INIT => X"3942"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(2),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z572
    );
  ix54672z24941 : X_LUT4
    generic map(
      INIT => X"6158"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(2),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z569
    );
  ix54672z55105 : X_LUT4
    generic map(
      INIT => X"A5B4"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(2),
      O => nx54672z1070
    );
  ix54672z19239 : X_LUT4
    generic map(
      INIT => X"4D24"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(2),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z577
    );
  ix54672z34616 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(2),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z574
    );
  ix54672z28142 : X_LUT4
    generic map(
      INIT => X"5A96"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(2),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z578
    );
  ix54672z25989 : X_LUT4
    generic map(
      INIT => X"37C8"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(2),
      O => nx54672z1072
    );
  ix54672z17639 : X_LUT4
    generic map(
      INIT => X"39C6"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(2),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z575
    );
  ix54672z41384 : X_LUT4
    generic map(
      INIT => X"C36C"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(2),
      O => nx54672z1073
    );
  ix54672z10730 : X_LUT4
    generic map(
      INIT => X"56A8"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(2),
      O => nx54672z1069
    );
  ix54672z59447 : X_LUT4
    generic map(
      INIT => X"A6A6"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(1),
      ADR3 => VCC,
      O => nx54672z1078
    );
  ix54672z43182 : X_LUT4
    generic map(
      INIT => X"CF32"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(2),
      ADR3 => romoaddro6_s(1),
      O => nx54672z1075
    );
  ix54672z25925 : X_LUT4
    generic map(
      INIT => X"7130"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z563
    );
  ix54672z61902 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro8_s(1),
      ADR1 => romeaddro8_s(3),
      ADR2 => romeaddro8_s(0),
      ADR3 => romeaddro8_s(2),
      O => nx54672z556
    );
  ix54672z14574 : X_LUT4
    generic map(
      INIT => X"7510"
    )
    port map (
      ADR0 => romeaddro8_s(1),
      ADR1 => romeaddro8_s(3),
      ADR2 => romeaddro8_s(0),
      ADR3 => romeaddro8_s(2),
      O => nx54672z560
    );
  ix54672z19159 : X_LUT4
    generic map(
      INIT => X"2942"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z565
    );
  ix54672z4327 : X_LUT4
    generic map(
      INIT => X"30B2"
    )
    port map (
      ADR0 => romeaddro8_s(1),
      ADR1 => romeaddro8_s(3),
      ADR2 => romeaddro8_s(0),
      ADR3 => romeaddro8_s(2),
      O => nx54672z557
    );
  ix54672z5330 : X_LUT4
    generic map(
      INIT => X"5D04"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z566
    );
  ix54672z12685 : X_LUT4
    generic map(
      INIT => X"2492"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(2),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z571
    );
  ix54672z34600 : X_LUT4
    generic map(
      INIT => X"7EE8"
    )
    port map (
      ADR0 => romeaddro8_s(2),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z562
    );
  ix54672z61918 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro8_s(0),
      ADR1 => romeaddro8_s(2),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(1),
      O => nx54672z568
    );
  ix54672z24883 : X_LUT4
    generic map(
      INIT => X"05FA"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro7_s(3),
      ADR3 => romoaddro7_s(0),
      O => nx54672z1209
    );
  ix54672z26161 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romoaddro7_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro7_s(2),
      ADR3 => VCC,
      O => nx54672z1213
    );
  ix54672z7108 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romoaddro7_s(2),
      ADR3 => romoaddro7_s(3),
      O => U1_ROMO7_modgen_rom_ix0_nx_rm64_16_u
    );
  ix54672z29246 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romoaddro7_s(0),
      ADR1 => romoaddro7_s(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z1214
    );
  ix54672z16289 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro7_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro7_s(3),
      O => U1_ROMO7_modgen_rom_ix0_nx_rm64_16_l
    );
  ix54672z26049 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romoaddro6_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro6_s(2),
      ADR3 => VCC,
      O => nx54672z1134
    );
  ix54672z29134 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romoaddro6_s(0),
      ADR1 => romoaddro6_s(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z1135
    );
  ix54672z6996 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romoaddro6_s(2),
      ADR3 => romoaddro6_s(3),
      O => U1_ROMO6_modgen_rom_ix0_nx_rm64_16_u
    );
  ix54672z25766 : X_LUT4
    generic map(
      INIT => X"5A6A"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(1),
      ADR2 => romoaddro4_s(0),
      ADR3 => romoaddro4_s(3),
      O => nx54672z914
    );
  ix54672z16177 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro6_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro6_s(3),
      O => U1_ROMO6_modgen_rom_ix0_nx_rm64_16_l
    );
  ix54672z15138 : X_LUT4
    generic map(
      INIT => X"1818"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(1),
      ADR3 => VCC,
      O => nx54672z1079
    );
  ix54672z4441 : X_LUT4
    generic map(
      INIT => X"5566"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(2),
      ADR2 => VCC,
      ADR3 => romoaddro6_s(0),
      O => nx54672z1132
    );
  ix54672z24675 : X_LUT4
    generic map(
      INIT => X"3232"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => romoaddro6_s(0),
      ADR2 => romoaddro6_s(2),
      ADR3 => VCC,
      O => nx54672z1076
    );
  ix54672z10622 : X_LUT4
    generic map(
      INIT => X"333C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro6_s(2),
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(0),
      O => nx54672z1133
    );
  ix54672z56785 : X_LUT4
    generic map(
      INIT => X"A5F0"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(2),
      O => nx54672z1129
    );
  ix54672z24770 : X_LUT4
    generic map(
      INIT => X"05FA"
    )
    port map (
      ADR0 => romoaddro6_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro6_s(1),
      ADR3 => romoaddro6_s(0),
      O => nx54672z1130
    );
  ix54672z12592 : X_LUT4
    generic map(
      INIT => X"4924"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(2),
      ADR3 => romeaddro7_s(0),
      O => nx54672z506
    );
  ix54672z61825 : X_LUT4
    generic map(
      INIT => X"E996"
    )
    port map (
      ADR0 => romeaddro7_s(1),
      ADR1 => romeaddro7_s(3),
      ADR2 => romeaddro7_s(2),
      ADR3 => romeaddro7_s(0),
      O => nx54672z503
    );
  ready_OUTPUT_OFF_O1INV_7641 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlcn339,
      O => ready_OUTPUT_OFF_O1INV
    );
  ready_OUTPUT_OFF_OCEINV_7642 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_istate_reg(0),
      O => ready_OUTPUT_OFF_OCEINV
    );
  ready_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ready_repl0,
      O => ready_O
    );
  ready_OUTPUT_OTCLK1INV_7643 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => ready_OUTPUT_OTCLK1INV
    );
  U_DCT1D_reg_ready_reg_repl0 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ready_OUTPUT_OFF_O1INV,
      CE => ready_OUTPUT_OFF_OCEINV,
      CLK => ready_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => ready_OUTPUT_OFF_OFF1_RST,
      O => ready_repl0
    );
  ready_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => ready_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => ready_OUTPUT_OFF_OFF1_RST
    );
  ready_OUTPUT_OFF_OFF1_RSTAND_7644 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ready_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto_10_OUTPUT_OTCLK1INV_7645 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto_10_OUTPUT_OTCLK1INV
    );
  dcto_10_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_dup0(10),
      O => dcto_10_O
    );
  dcto_10_OUTPUT_OFF_OCEINV_7646 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => dcto_10_OUTPUT_OFF_OCEINV
    );
  dcto_10_OUTPUT_OFF_O1INV_7647 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491(22),
      O => dcto_10_OUTPUT_OFF_O1INV
    );
  U_DCT2D_reg_dcto_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto_10_OUTPUT_OFF_O1INV,
      CE => dcto_10_OUTPUT_OFF_OCEINV,
      CLK => dcto_10_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto_10_OUTPUT_OFF_OFF1_RST,
      O => dcto_dup0(10)
    );
  dcto_10_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto_10_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto_10_OUTPUT_OFF_OFF1_RST
    );
  dcto_10_OUTPUT_OFF_OFF1_RSTAND_7648 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto_10_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto_11_OUTPUT_OFF_O1INV_7649 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491(23),
      O => dcto_11_OUTPUT_OFF_O1INV
    );
  dcto_11_OUTPUT_OFF_OCEINV_7650 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => dcto_11_OUTPUT_OFF_OCEINV
    );
  dcto_11_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_dup0(11),
      O => dcto_11_O
    );
  dcto_11_OUTPUT_OTCLK1INV_7651 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto_11_OUTPUT_OTCLK1INV
    );
  U_DCT2D_reg_dcto_11_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto_11_OUTPUT_OFF_O1INV,
      CE => dcto_11_OUTPUT_OFF_OCEINV,
      CLK => dcto_11_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto_11_OUTPUT_OFF_OFF1_RST,
      O => dcto_dup0(11)
    );
  dcto_11_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto_11_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto_11_OUTPUT_OFF_OFF1_RST
    );
  dcto_11_OUTPUT_OFF_OFF1_RSTAND_7652 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto_11_OUTPUT_OFF_OFF1_RSTAND
    );
  ix54672z38981 : X_LUT4
    generic map(
      INIT => X"A244"
    )
    port map (
      ADR0 => romoaddro8_s(1),
      ADR1 => romoaddro8_s(2),
      ADR2 => romoaddro8_s(0),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1258
    );
  ix54672z58782 : X_LUT4
    generic map(
      INIT => X"E836"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => romoaddro8_s(0),
      ADR2 => romoaddro8_s(2),
      ADR3 => romoaddro8_s(1),
      O => nx54672z1251
    );
  ix54672z45431 : X_LUT4
    generic map(
      INIT => X"96C6"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => romoaddro8_s(0),
      ADR2 => romoaddro8_s(2),
      ADR3 => romoaddro8_s(1),
      O => nx54672z1252
    );
  ix54672z53068 : X_LUT4
    generic map(
      INIT => X"9966"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => romoaddro8_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro8_s(2),
      O => nx54672z1255
    );
  ix54672z44471 : X_LUT4
    generic map(
      INIT => X"C1C0"
    )
    port map (
      ADR0 => romoaddro8_s(1),
      ADR1 => romoaddro8_s(2),
      ADR2 => romoaddro8_s(0),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1260
    );
  ix54672z62624 : X_LUT4
    generic map(
      INIT => X"E8A0"
    )
    port map (
      ADR0 => romoaddro8_s(1),
      ADR1 => romoaddro8_s(2),
      ADR2 => romoaddro8_s(0),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1261
    );
  ix54672z21881 : X_LUT4
    generic map(
      INIT => X"31C6"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => romoaddro8_s(0),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1266
    );
  ix54672z23320 : X_LUT4
    generic map(
      INIT => X"3B02"
    )
    port map (
      ADR0 => romoaddro8_s(1),
      ADR1 => romoaddro8_s(2),
      ADR2 => romoaddro8_s(0),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1257
    );
  ix54672z20176 : X_LUT4
    generic map(
      INIT => X"6518"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => romoaddro8_s(0),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1263
    );
  ix54672z26157 : X_LUT4
    generic map(
      INIT => X"37C8"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1191
    );
  ix54672z60276 : X_LUT4
    generic map(
      INIT => X"A800"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1142
    );
  ix54672z48690 : X_LUT4
    generic map(
      INIT => X"CF4C"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1146
    );
  ix54672z40835 : X_LUT4
    generic map(
      INIT => X"D25A"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1193
    );
  ix54672z55411 : X_LUT4
    generic map(
      INIT => X"F5F4"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1143
    );
  ix54672z11160 : X_LUT4
    generic map(
      INIT => X"56AA"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1194
    );
  ix54672z26207 : X_LUT4
    generic map(
      INIT => X"3CC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro7_s(2),
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1199
    );
  ix54672z29978 : X_LUT4
    generic map(
      INIT => X"3C96"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1190
    );
  ix54672z7036 : X_LUT4
    generic map(
      INIT => X"3388"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => romoaddro7_s(2),
      ADR2 => VCC,
      ADR3 => romoaddro7_s(3),
      O => nx54672z1196
    );
  ix54672z37510 : X_LUT4
    generic map(
      INIT => X"943C"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => romoaddro8_s(0),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1267
    );
  ix54672z28633 : X_LUT4
    generic map(
      INIT => X"6D5A"
    )
    port map (
      ADR0 => romoaddro8_s(3),
      ADR1 => romoaddro8_s(0),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1264
    );
  ix54672z55402 : X_LUT4
    generic map(
      INIT => X"DDDC"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1137
    );
  ix54672z40947 : X_LUT4
    generic map(
      INIT => X"B43C"
    )
    port map (
      ADR0 => romoaddro8_s(2),
      ADR1 => romoaddro8_s(3),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(0),
      O => nx54672z1272
    );
  ix54672z30090 : X_LUT4
    generic map(
      INIT => X"4BB4"
    )
    port map (
      ADR0 => romoaddro8_s(2),
      ADR1 => romoaddro8_s(3),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(0),
      O => nx54672z1269
    );
  ix54672z11272 : X_LUT4
    generic map(
      INIT => X"666C"
    )
    port map (
      ADR0 => romoaddro8_s(2),
      ADR1 => romoaddro8_s(3),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(0),
      O => nx54672z1273
    );
  ix54672z23519 : X_LUT4
    generic map(
      INIT => X"1F00"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1139
    );
  ix54672z26269 : X_LUT4
    generic map(
      INIT => X"56AA"
    )
    port map (
      ADR0 => romoaddro8_s(2),
      ADR1 => romoaddro8_s(3),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(0),
      O => nx54672z1270
    );
  ix54672z48682 : X_LUT4
    generic map(
      INIT => X"F370"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(1),
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1140
    );
  ix54672z23527 : X_LUT4
    generic map(
      INIT => X"3700"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(1),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1145
    );
  ix54672z2307 : X_LUT4
    generic map(
      INIT => X"0C0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(3),
      ADR3 => VCC,
      O => nx54672z580
    );
  ix54672z23630 : X_LUT4
    generic map(
      INIT => X"444C"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => romoaddro8_s(2),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1218
    );
  ix54672z48793 : X_LUT4
    generic map(
      INIT => X"8EAE"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => romoaddro8_s(2),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1219
    );
  ix54672z55514 : X_LUT4
    generic map(
      INIT => X"F0FE"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => romoaddro8_s(2),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1216
    );
  ix54672z26319 : X_LUT4
    generic map(
      INIT => X"5AA0"
    )
    port map (
      ADR0 => romoaddro8_s(2),
      ADR1 => VCC,
      ADR2 => romoaddro8_s(3),
      ADR3 => romoaddro8_s(0),
      O => nx54672z1278
    );
  ix54672z42184 : X_LUT4
    generic map(
      INIT => X"CC22"
    )
    port map (
      ADR0 => romoaddro8_s(2),
      ADR1 => romoaddro8_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro8_s(0),
      O => nx54672z1279
    );
  ix54672z7148 : X_LUT4
    generic map(
      INIT => X"5858"
    )
    port map (
      ADR0 => romoaddro8_s(2),
      ADR1 => romoaddro8_s(1),
      ADR2 => romoaddro8_s(3),
      ADR3 => VCC,
      O => nx54672z1275
    );
  ix54672z55375 : X_LUT4
    generic map(
      INIT => X"A5A0"
    )
    port map (
      ADR0 => romoaddro8_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro8_s(3),
      ADR3 => romoaddro8_s(0),
      O => nx54672z1276
    );
  ix54672z3377 : X_LUT4
    generic map(
      INIT => X"3322"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => romoaddro8_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro8_s(2),
      O => nx54672z1284
    );
  ix54672z42072 : X_LUT4
    generic map(
      INIT => X"AA44"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => romoaddro7_s(2),
      ADR2 => VCC,
      ADR3 => romoaddro7_s(0),
      O => nx54672z1200
    );
  ix54672z55263 : X_LUT4
    generic map(
      INIT => X"AA50"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro7_s(0),
      ADR3 => romoaddro7_s(3),
      O => nx54672z1197
    );
  ix54672z3265 : X_LUT4
    generic map(
      INIT => X"5454"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => romoaddro7_s(2),
      ADR3 => VCC,
      O => nx54672z1205
    );
  ix54672z2758 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romoaddro7_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro7_s(2),
      ADR3 => romoaddro7_s(1),
      O => nx54672z1206
    );
  ix54672z3060 : X_LUT4
    generic map(
      INIT => X"0050"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro7_s(2),
      ADR3 => romoaddro7_s(1),
      O => nx54672z1202
    );
  ix54672z2995 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro7_s(1),
      O => nx54672z1203
    );
  ix54672z4553 : X_LUT4
    generic map(
      INIT => X"5566"
    )
    port map (
      ADR0 => romoaddro7_s(3),
      ADR1 => romoaddro7_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro7_s(2),
      O => nx54672z1211
    );
  ix54672z10734 : X_LUT4
    generic map(
      INIT => X"11EE"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => romoaddro7_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro7_s(2),
      O => nx54672z1212
    );
  ix54672z55304 : X_LUT4
    generic map(
      INIT => X"A5AA"
    )
    port map (
      ADR0 => romoaddro7_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro7_s(3),
      ADR3 => romoaddro7_s(2),
      O => nx54672z1208
    );
  ix54672z10507 : X_LUT4
    generic map(
      INIT => X"56A8"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(1),
      ADR2 => romoaddro4_s(0),
      ADR3 => romoaddro4_s(3),
      O => nx54672z911
    );
  ix54672z41161 : X_LUT4
    generic map(
      INIT => X"96D2"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(1),
      ADR2 => romoaddro4_s(0),
      ADR3 => romoaddro4_s(3),
      O => nx54672z915
    );
  ix54672z41540 : X_LUT4
    generic map(
      INIT => X"9964"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(1),
      O => nx54672z859
    );
  ix54672z54882 : X_LUT4
    generic map(
      INIT => X"CC36"
    )
    port map (
      ADR0 => romoaddro4_s(2),
      ADR1 => romoaddro4_s(1),
      ADR2 => romoaddro4_s(0),
      ADR3 => romoaddro4_s(3),
      O => nx54672z912
    );
  ix54672z44870 : X_LUT4
    generic map(
      INIT => X"96C6"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(1),
      O => nx54672z857
    );
  ix54672z52507 : X_LUT4
    generic map(
      INIT => X"A55A"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => VCC,
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(1),
      O => nx54672z860
    );
  ix54672z25758 : X_LUT4
    generic map(
      INIT => X"3CC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro3_s(2),
      ADR2 => romoaddro3_s(0),
      ADR3 => romoaddro3_s(3),
      O => nx54672z883
    );
  ix54672z58221 : X_LUT4
    generic map(
      INIT => X"E836"
    )
    port map (
      ADR0 => romoaddro3_s(3),
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(1),
      O => nx54672z856
    );
  ix54672z6587 : X_LUT4
    generic map(
      INIT => X"3388"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(2),
      ADR2 => VCC,
      ADR3 => romoaddro3_s(3),
      O => nx54672z880
    );
  ix54672z41623 : X_LUT4
    generic map(
      INIT => X"9988"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro3_s(2),
      O => nx54672z884
    );
  ix54672z54814 : X_LUT4
    generic map(
      INIT => X"AA44"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro3_s(3),
      O => nx54672z881
    );
  ix54672z4104 : X_LUT4
    generic map(
      INIT => X"03FC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro3_s(0),
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(3),
      O => nx54672z895
    );
  ix54672z10285 : X_LUT4
    generic map(
      INIT => X"11EE"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro3_s(2),
      O => nx54672z896
    );
  ix54672z54855 : X_LUT4
    generic map(
      INIT => X"AA5A"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => VCC,
      ADR2 => romoaddro3_s(2),
      ADR3 => romoaddro3_s(3),
      O => nx54672z892
    );
  ix54672z24434 : X_LUT4
    generic map(
      INIT => X"3366"
    )
    port map (
      ADR0 => romoaddro3_s(1),
      ADR1 => romoaddro3_s(0),
      ADR2 => VCC,
      ADR3 => romoaddro3_s(3),
      O => nx54672z893
    );
  ix54672z29169 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro8_s(1),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(2),
      O => nx54672z582
    );
  ix54672z29166 : X_LUT4
    generic map(
      INIT => X"6996"
    )
    port map (
      ADR0 => romeaddro8_s(1),
      ADR1 => romeaddro8_s(0),
      ADR2 => romeaddro8_s(3),
      ADR3 => romeaddro8_s(2),
      O => U1_ROME8_modgen_rom_ix2_nx_rm64_16_u
    );
  ix54672z14476 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => romeaddro8_s(1),
      ADR1 => romeaddro8_s(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z583
    );
  dcto_4_OUTPUT_OFF_O1INV_7653 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491(16),
      O => dcto_4_OUTPUT_OFF_O1INV
    );
  dcto_4_OUTPUT_OFF_OCEINV_7654 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => dcto_4_OUTPUT_OFF_OCEINV
    );
  dcto_4_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_dup0(4),
      O => dcto_4_O
    );
  dcto_4_OUTPUT_OTCLK1INV_7655 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto_4_OUTPUT_OTCLK1INV
    );
  U_DCT2D_reg_dcto_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto_4_OUTPUT_OFF_O1INV,
      CE => dcto_4_OUTPUT_OFF_OCEINV,
      CLK => dcto_4_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto_4_OUTPUT_OFF_OFF1_RST,
      O => dcto_dup0(4)
    );
  dcto_4_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto_4_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto_4_OUTPUT_OFF_OFF1_RST
    );
  dcto_4_OUTPUT_OFF_OFF1_RSTAND_7656 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto_4_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto_5_OUTPUT_OFF_O1INV_7657 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491(17),
      O => dcto_5_OUTPUT_OFF_O1INV
    );
  dcto_5_OUTPUT_OFF_OCEINV_7658 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => dcto_5_OUTPUT_OFF_OCEINV
    );
  dcto_5_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_dup0(5),
      O => dcto_5_O
    );
  dcto_5_OUTPUT_OTCLK1INV_7659 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto_5_OUTPUT_OTCLK1INV
    );
  U_DCT2D_reg_dcto_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto_5_OUTPUT_OFF_O1INV,
      CE => dcto_5_OUTPUT_OFF_OCEINV,
      CLK => dcto_5_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto_5_OUTPUT_OFF_OFF1_RST,
      O => dcto_dup0(5)
    );
  dcto_5_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto_5_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto_5_OUTPUT_OFF_OFF1_RST
    );
  dcto_5_OUTPUT_OFF_OFF1_RSTAND_7660 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto_5_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto_6_OUTPUT_OFF_O1INV_7661 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491(18),
      O => dcto_6_OUTPUT_OFF_O1INV
    );
  dcto_6_OUTPUT_OFF_OCEINV_7662 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => dcto_6_OUTPUT_OFF_OCEINV
    );
  dcto_6_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_dup0(6),
      O => dcto_6_O
    );
  dcto_6_OUTPUT_OTCLK1INV_7663 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto_6_OUTPUT_OTCLK1INV
    );
  U_DCT2D_reg_dcto_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto_6_OUTPUT_OFF_O1INV,
      CE => dcto_6_OUTPUT_OFF_OCEINV,
      CLK => dcto_6_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto_6_OUTPUT_OFF_OFF1_RST,
      O => dcto_dup0(6)
    );
  dcto_6_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto_6_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto_6_OUTPUT_OFF_OFF1_RST
    );
  dcto_6_OUTPUT_OFF_OFF1_RSTAND_7664 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto_6_OUTPUT_OFF_OFF1_RSTAND
    );
  ix54672z3172 : X_LUT4
    generic map(
      INIT => X"0300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romoaddro8_s(3),
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1281
    );
  ix54672z2870 : X_LUT4
    generic map(
      INIT => X"FFFA"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro8_s(1),
      ADR3 => romoaddro8_s(2),
      O => nx54672z1285
    );
  ix54672z3107 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => romoaddro8_s(3),
      ADR2 => VCC,
      ADR3 => romoaddro8_s(1),
      O => nx54672z1282
    );
  ix54672z4666 : X_LUT4
    generic map(
      INIT => X"05FA"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro8_s(2),
      ADR3 => romoaddro8_s(3),
      O => nx54672z1290
    );
  ix54672z10847 : X_LUT4
    generic map(
      INIT => X"0F5A"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => VCC,
      ADR2 => romoaddro8_s(2),
      ADR3 => romoaddro8_s(1),
      O => nx54672z1291
    );
  ix54672z57237 : X_LUT4
    generic map(
      INIT => X"CC66"
    )
    port map (
      ADR0 => romoaddro8_s(2),
      ADR1 => romoaddro8_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro8_s(3),
      O => nx54672z1287
    );
  ix54672z24996 : X_LUT4
    generic map(
      INIT => X"5566"
    )
    port map (
      ADR0 => romoaddro8_s(0),
      ADR1 => romoaddro8_s(1),
      ADR2 => VCC,
      ADR3 => romoaddro8_s(3),
      O => nx54672z1288
    );
  dcto1_10_OUTPUT_OFF_O1INV_7665 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n2651,
      O => dcto1_10_OUTPUT_OFF_O1INV
    );
  dcto1_10_OUTPUT_OFF_OCEINV_7666 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => dcto1_10_OUTPUT_OFF_OCEINV
    );
  dcto1_10_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_9_repl1,
      O => dcto1_10_O
    );
  dcto1_10_OUTPUT_OTCLK1INV_7667 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto1_10_OUTPUT_OTCLK1INV
    );
  U_DCT1D_reg_ramdatai_s_9_repl1 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto1_10_OUTPUT_OFF_O1INV,
      CE => dcto1_10_OUTPUT_OFF_OCEINV,
      CLK => dcto1_10_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto1_10_OUTPUT_OFF_OFF1_RST,
      O => ramdatai_9_repl1
    );
  dcto1_10_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto1_10_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto1_10_OUTPUT_OFF_OFF1_RST
    );
  dcto1_10_OUTPUT_OFF_OFF1_RSTAND_7668 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto1_10_OUTPUT_OFF_OFF1_RSTAND
    );
  U_DCT1D_reg_istate_reg_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_istate_reg_1_DYMUX,
      CE => U_DCT1D_istate_reg_1_CEINV,
      CLK => U_DCT1D_istate_reg_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_istate_reg_1_FFY_RST,
      O => U_DCT1D_istate_reg(0)
    );
  U_DCT1D_istate_reg_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_istate_reg_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_istate_reg_1_FFY_RST
    );
  U_DCT1D_ix1822z1318 : X_LUT4
    generic map(
      INIT => X"5050"
    )
    port map (
      ADR0 => reqwrfail_s,
      ADR1 => VCC,
      ADR2 => U_DCT1D_istate_reg(0),
      ADR3 => VCC,
      O => U_DCT1D_rtlcn403
    );
  U_DCT1D_ix59993z1420 : X_LUT4
    generic map(
      INIT => X"7788"
    )
    port map (
      ADR0 => U_DCT1D_inpcnt_reg(1),
      ADR1 => U_DCT1D_inpcnt_reg(0),
      ADR2 => VCC,
      ADR3 => U_DCT1D_inpcnt_reg(2),
      O => U_DCT1D_nx59993z1
    );
  U_DCT1D_reg_istate_reg_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_istate_reg_1_DXMUX,
      CE => U_DCT1D_istate_reg_1_CEINV,
      CLK => U_DCT1D_istate_reg_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_istate_reg_1_FFX_RST,
      O => U_DCT1D_istate_reg(1)
    );
  U_DCT1D_istate_reg_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_istate_reg_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_istate_reg_1_FFX_RST
    );
  U_DCT1D_modgen_counter_inpcnt_reg_reg_q_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_inpcnt_reg_2_DYMUX,
      CE => U_DCT1D_inpcnt_reg_2_CEINV,
      CLK => U_DCT1D_inpcnt_reg_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_inpcnt_reg_2_FFY_RST,
      O => U_DCT1D_inpcnt_reg(2)
    );
  U_DCT1D_inpcnt_reg_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_inpcnt_reg_2_FFY_RSTAND,
      I1 => GSR,
      O => U_DCT1D_inpcnt_reg_2_FFY_RST
    );
  U_DCT1D_inpcnt_reg_2_FFY_RSTAND_7669 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_inpcnt_reg_2_FFY_RSTAND
    );
  ix57510z64083 : X_LUT4
    generic map(
      INIT => X"F351"
    )
    port map (
      ADR0 => U_DBUFCTL_mem1_full_reg,
      ADR1 => U_DBUFCTL_mem2_full_reg,
      ADR2 => U_DBUFCTL_mem2_lock_reg,
      ADR3 => U_DBUFCTL_mem1_lock_reg,
      O => U_DBUFCTL_rtlcn7
    );
  U_DBUFCTL_reg_reqrdfail : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => reqrdfail_s_DYMUX,
      CE => reqrdfail_s_CEINV,
      CLK => reqrdfail_s_CLKINV,
      SET => GND,
      RST => reqrdfail_s_FFY_RST,
      O => reqrdfail_s
    );
  reqrdfail_s_FFY_RSTOR : X_OR2
    port map (
      I0 => reqrdfail_s_FFY_RSTAND,
      I1 => GSR,
      O => reqrdfail_s_FFY_RST
    );
  reqrdfail_s_FFY_RSTAND_7670 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => reqrdfail_s_FFY_RSTAND
    );
  ix12221z65514 : X_LUT4
    generic map(
      INIT => X"FAC8"
    )
    port map (
      ADR0 => U_DBUFCTL_mem1_full_reg,
      ADR1 => U_DBUFCTL_mem2_full_reg,
      ADR2 => U_DBUFCTL_mem1_lock_reg,
      ADR3 => U_DBUFCTL_mem2_lock_reg,
      O => U_DBUFCTL_rtlc4n197
    );
  ix40249z1997 : X_LUT4
    generic map(
      INIT => X"5700"
    )
    port map (
      ADR0 => U_DBUFCTL_rtlcn1,
      ADR1 => U_DBUFCTL_mem2_full_reg,
      ADR2 => U_DBUFCTL_mem2_lock_reg,
      ADR3 => requestwr_s,
      O => reqrdfail_s_F
    );
  dcto_1_OUTPUT_OTCLK1INV_7671 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto_1_OUTPUT_OTCLK1INV
    );
  dcto_1_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_dup0(1),
      O => dcto_1_O
    );
  dcto_1_OUTPUT_OFF_OCEINV_7672 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => dcto_1_OUTPUT_OFF_OCEINV
    );
  dcto_1_OUTPUT_OFF_O1INV_7673 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491(13),
      O => dcto_1_OUTPUT_OFF_O1INV
    );
  U_DCT2D_reg_dcto_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto_1_OUTPUT_OFF_O1INV,
      CE => dcto_1_OUTPUT_OFF_OCEINV,
      CLK => dcto_1_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto_1_OUTPUT_OFF_OFF1_RST,
      O => dcto_dup0(1)
    );
  dcto_1_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto_1_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto_1_OUTPUT_OFF_OFF1_RST
    );
  dcto_1_OUTPUT_OFF_OFF1_RSTAND_7674 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto_1_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto_2_OUTPUT_OFF_O1INV_7675 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491(14),
      O => dcto_2_OUTPUT_OFF_O1INV
    );
  dcto_2_OUTPUT_OFF_OCEINV_7676 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => dcto_2_OUTPUT_OFF_OCEINV
    );
  dcto_2_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_dup0(2),
      O => dcto_2_O
    );
  dcto_2_OUTPUT_OTCLK1INV_7677 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto_2_OUTPUT_OTCLK1INV
    );
  U_DCT2D_reg_dcto_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto_2_OUTPUT_OFF_O1INV,
      CE => dcto_2_OUTPUT_OFF_OCEINV,
      CLK => dcto_2_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto_2_OUTPUT_OFF_OFF1_RST,
      O => dcto_dup0(2)
    );
  dcto_2_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto_2_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto_2_OUTPUT_OFF_OFF1_RST
    );
  dcto_2_OUTPUT_OFF_OFF1_RSTAND_7678 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto_2_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto_3_OUTPUT_OFF_O1INV_7679 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491(15),
      O => dcto_3_OUTPUT_OFF_O1INV
    );
  dcto_3_OUTPUT_OFF_OCEINV_7680 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => dcto_3_OUTPUT_OFF_OCEINV
    );
  dcto_3_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_dup0(3),
      O => dcto_3_O
    );
  dcto_3_OUTPUT_OTCLK1INV_7681 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto_3_OUTPUT_OTCLK1INV
    );
  U_DCT2D_reg_dcto_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto_3_OUTPUT_OFF_O1INV,
      CE => dcto_3_OUTPUT_OFF_OCEINV,
      CLK => dcto_3_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto_3_OUTPUT_OFF_OFF1_RST,
      O => dcto_dup0(3)
    );
  dcto_3_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto_3_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto_3_OUTPUT_OFF_OFF1_RST
    );
  dcto_3_OUTPUT_OFF_OFF1_RSTAND_7682 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto_3_OUTPUT_OFF_OFF1_RSTAND
    );
  dcti_6_IFF_IFFDMUX_7683 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti_6_INBUF,
      O => dcti_6_IFF_IFFDMUX
    );
  dcti_6_IFF_ICLK1INV_7684 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcti_6_IFF_ICLK1INV
    );
  dcti_6_IFF_ICEINV_7685 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => dcti_6_IFF_ICEINV
    );
  U_DCT1D_reg_latchbuf_reg_7_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcti_6_IFF_IFFDMUX,
      CE => dcti_6_IFF_ICEINV,
      CLK => dcti_6_IFF_ICLK1INV,
      SET => GND,
      RST => dcti_6_IFF_IFF1_RST,
      O => U_DCT1D_latchbuf_reg_7_Q(6)
    );
  dcti_6_IFF_IFF1_RSTOR : X_OR2
    port map (
      I0 => dcti_6_IFF_IFF1_RSTAND,
      I1 => GSR,
      O => dcti_6_IFF_IFF1_RST
    );
  dcti_6_IFF_IFF1_RSTAND_7686 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcti_6_IFF_IFF1_RSTAND
    );
  dcto_0_OUTPUT_OTCLK1INV_7687 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto_0_OUTPUT_OTCLK1INV
    );
  dcto_0_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_dup0(0),
      O => dcto_0_O
    );
  dcto_0_OUTPUT_OFF_OCEINV_7688 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => dcto_0_OUTPUT_OFF_OCEINV
    );
  dcto_0_OUTPUT_OFF_O1INV_7689 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491(12),
      O => dcto_0_OUTPUT_OFF_O1INV
    );
  U_DCT2D_reg_dcto_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto_0_OUTPUT_OFF_O1INV,
      CE => dcto_0_OUTPUT_OFF_OCEINV,
      CLK => dcto_0_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto_0_OUTPUT_OFF_OFF1_RST,
      O => dcto_dup0(0)
    );
  dcto_0_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto_0_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto_0_OUTPUT_OFF_OFF1_RST
    );
  dcto_0_OUTPUT_OFF_OFF1_RSTAND_7690 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto_0_OUTPUT_OFF_OFF1_RSTAND
    );
  U_DCT2D_reg_romeaddro1_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro1_s_1_DYMUX,
      CE => rome2addro1_s_1_CEINV,
      CLK => rome2addro1_s_1_CLKINV,
      SET => GND,
      RST => rome2addro1_s_1_FFY_RST,
      O => rome2addro1_s(0)
    );
  rome2addro1_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro1_s_1_SRINV,
      I1 => GSR,
      O => rome2addro1_s_1_FFY_RST
    );
  U_DCT2D_reg_romeaddro1_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro1_s_1_DXMUX,
      CE => rome2addro1_s_1_CEINV,
      CLK => rome2addro1_s_1_CLKINV,
      SET => GND,
      RST => rome2addro1_s_1_FFX_RST,
      O => rome2addro1_s(1)
    );
  rome2addro1_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro1_s_1_SRINV,
      I1 => GSR,
      O => rome2addro1_s_1_FFX_RST
    );
  U_DCT2D_reg_romeaddro1_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro1_s_3_DYMUX,
      CE => rome2addro1_s_3_CEINV,
      CLK => rome2addro1_s_3_CLKINV,
      SET => GND,
      RST => rome2addro1_s_3_FFY_RST,
      O => rome2addro1_s(2)
    );
  rome2addro1_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro1_s_3_SRINV,
      I1 => GSR,
      O => rome2addro1_s_3_FFY_RST
    );
  U_DCT2D_reg_romeaddro1_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro1_s_3_DXMUX,
      CE => rome2addro1_s_3_CEINV,
      CLK => rome2addro1_s_3_CLKINV,
      SET => GND,
      RST => rome2addro1_s_3_FFX_RST,
      O => rome2addro1_s(3)
    );
  rome2addro1_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro1_s_3_SRINV,
      I1 => GSR,
      O => rome2addro1_s_3_FFX_RST
    );
  U_DCT2D_reg_romeaddro2_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro2_s_1_DYMUX,
      CE => rome2addro2_s_1_CEINV,
      CLK => rome2addro2_s_1_CLKINV,
      SET => GND,
      RST => rome2addro2_s_1_FFY_RST,
      O => rome2addro2_s(0)
    );
  rome2addro2_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro2_s_1_SRINV,
      I1 => GSR,
      O => rome2addro2_s_1_FFY_RST
    );
  U_DCT2D_reg_romeaddro2_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro2_s_1_DXMUX,
      CE => rome2addro2_s_1_CEINV,
      CLK => rome2addro2_s_1_CLKINV,
      SET => GND,
      RST => rome2addro2_s_1_FFX_RST,
      O => rome2addro2_s(1)
    );
  rome2addro2_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro2_s_1_SRINV,
      I1 => GSR,
      O => rome2addro2_s_1_FFX_RST
    );
  dcto1_11_OUTPUT_OFF_O1INV_7691 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n2651,
      O => dcto1_11_OUTPUT_OFF_O1INV
    );
  dcto1_11_OUTPUT_OFF_OCEINV_7692 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => dcto1_11_OUTPUT_OFF_OCEINV
    );
  dcto1_11_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_9_repl2,
      O => dcto1_11_O
    );
  dcto1_11_OUTPUT_OTCLK1INV_7693 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto1_11_OUTPUT_OTCLK1INV
    );
  U_DCT1D_reg_ramdatai_s_9_repl2 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto1_11_OUTPUT_OFF_O1INV,
      CE => dcto1_11_OUTPUT_OFF_OCEINV,
      CLK => dcto1_11_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto1_11_OUTPUT_OFF_OFF1_RST,
      O => ramdatai_9_repl2
    );
  dcto1_11_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto1_11_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto1_11_OUTPUT_OFF_OFF1_RST
    );
  dcto1_11_OUTPUT_OFF_OFF1_RSTAND_7694 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto1_11_OUTPUT_OFF_OFF1_RSTAND
    );
  odv_OUTPUT_OTCLK1INV_7695 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => odv_OUTPUT_OTCLK1INV
    );
  odv_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => odv_dup0,
      O => odv_O
    );
  odv_OUTPUT_OFF_OCEINV_7696 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1854,
      O => odv_OUTPUT_OFF_OCEINV
    );
  odv_OUTPUT_OFF_O1INV_7697 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => odv_OUTPUT_OFF_O1INV
    );
  U_DCT2D_reg_odv : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => odv_OUTPUT_OFF_O1INV,
      CE => odv_OUTPUT_OFF_OCEINV,
      CLK => odv_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => odv_OUTPUT_OFF_OFF1_RST,
      O => odv_dup0
    );
  odv_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => odv_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => odv_OUTPUT_OFF_OFF1_RST
    );
  odv_OUTPUT_OFF_OFF1_RSTAND_7698 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => odv_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto1_0_OUTPUT_OFF_O1INV_7699 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n2660,
      O => dcto1_0_OUTPUT_OFF_O1INV
    );
  dcto1_0_OUTPUT_OFF_OCEINV_7700 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => dcto1_0_OUTPUT_OFF_OCEINV
    );
  dcto1_0_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_0_repl0,
      O => dcto1_0_O
    );
  dcto1_0_OUTPUT_OTCLK1INV_7701 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto1_0_OUTPUT_OTCLK1INV
    );
  U_DCT1D_reg_ramdatai_s_0_repl0 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto1_0_OUTPUT_OFF_O1INV,
      CE => dcto1_0_OUTPUT_OFF_OCEINV,
      CLK => dcto1_0_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto1_0_OUTPUT_OFF_OFF1_RST,
      O => ramdatai_0_repl0
    );
  dcto1_0_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto1_0_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto1_0_OUTPUT_OFF_OFF1_RST
    );
  dcto1_0_OUTPUT_OFF_OFF1_RSTAND_7702 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto1_0_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto1_1_OUTPUT_OFF_O1INV_7703 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n2659,
      O => dcto1_1_OUTPUT_OFF_O1INV
    );
  dcto1_1_OUTPUT_OFF_OCEINV_7704 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => dcto1_1_OUTPUT_OFF_OCEINV
    );
  dcto1_1_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_1_repl0,
      O => dcto1_1_O
    );
  dcto1_1_OUTPUT_OTCLK1INV_7705 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto1_1_OUTPUT_OTCLK1INV
    );
  U_DCT1D_reg_ramdatai_s_1_repl0 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto1_1_OUTPUT_OFF_O1INV,
      CE => dcto1_1_OUTPUT_OFF_OCEINV,
      CLK => dcto1_1_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto1_1_OUTPUT_OFF_OFF1_RST,
      O => ramdatai_1_repl0
    );
  dcto1_1_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto1_1_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto1_1_OUTPUT_OFF_OFF1_RST
    );
  dcto1_1_OUTPUT_OFF_OFF1_RSTAND_7706 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto1_1_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto1_2_OUTPUT_OFF_O1INV_7707 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n2658,
      O => dcto1_2_OUTPUT_OFF_O1INV
    );
  dcto1_2_OUTPUT_OFF_OCEINV_7708 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => dcto1_2_OUTPUT_OFF_OCEINV
    );
  dcto1_2_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_2_repl0,
      O => dcto1_2_O
    );
  dcto1_2_OUTPUT_OTCLK1INV_7709 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto1_2_OUTPUT_OTCLK1INV
    );
  U_DCT1D_reg_ramdatai_s_2_repl0 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto1_2_OUTPUT_OFF_O1INV,
      CE => dcto1_2_OUTPUT_OFF_OCEINV,
      CLK => dcto1_2_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto1_2_OUTPUT_OFF_OFF1_RST,
      O => ramdatai_2_repl0
    );
  dcto1_2_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto1_2_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto1_2_OUTPUT_OFF_OFF1_RST
    );
  dcto1_2_OUTPUT_OFF_OFF1_RSTAND_7710 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto1_2_OUTPUT_OFF_OFF1_RSTAND
    );
  dcti_2_IFF_IFFDMUX_7711 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti_2_INBUF,
      O => dcti_2_IFF_IFFDMUX
    );
  dcti_2_IFF_ICLK1INV_7712 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcti_2_IFF_ICLK1INV
    );
  dcti_2_IFF_ICEINV_7713 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => dcti_2_IFF_ICEINV
    );
  U_DCT1D_reg_latchbuf_reg_7_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcti_2_IFF_IFFDMUX,
      CE => dcti_2_IFF_ICEINV,
      CLK => dcti_2_IFF_ICLK1INV,
      SET => GND,
      RST => dcti_2_IFF_IFF1_RST,
      O => U_DCT1D_latchbuf_reg_7_Q(2)
    );
  dcti_2_IFF_IFF1_RSTOR : X_OR2
    port map (
      I0 => dcti_2_IFF_IFF1_RSTAND,
      I1 => GSR,
      O => dcti_2_IFF_IFF1_RST
    );
  dcti_2_IFF_IFF1_RSTAND_7714 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcti_2_IFF_IFF1_RSTAND
    );
  dcti_3_IFF_IFFDMUX_7715 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti_3_INBUF,
      O => dcti_3_IFF_IFFDMUX
    );
  dcti_3_IFF_ICLK1INV_7716 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcti_3_IFF_ICLK1INV
    );
  dcti_3_IFF_ICEINV_7717 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => dcti_3_IFF_ICEINV
    );
  U_DCT1D_reg_latchbuf_reg_7_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcti_3_IFF_IFFDMUX,
      CE => dcti_3_IFF_ICEINV,
      CLK => dcti_3_IFF_ICLK1INV,
      SET => GND,
      RST => dcti_3_IFF_IFF1_RST,
      O => U_DCT1D_latchbuf_reg_7_Q(3)
    );
  dcti_3_IFF_IFF1_RSTOR : X_OR2
    port map (
      I0 => dcti_3_IFF_IFF1_RSTAND,
      I1 => GSR,
      O => dcti_3_IFF_IFF1_RST
    );
  dcti_3_IFF_IFF1_RSTAND_7718 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcti_3_IFF_IFF1_RSTAND
    );
  dcti_5_IFF_IFF1_RSTOR : X_OR2
    port map (
      I0 => dcti_5_IFF_ISR_USED,
      I1 => GSR,
      O => dcti_5_IFF_IFF1_RST
    );
  U_DCT1D_reg_latchbuf_reg_7_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcti_5_IFF_IFFDMUX,
      CE => dcti_5_IFF_ICEINV,
      CLK => dcti_5_IFF_ICLK1INV,
      SET => GND,
      RST => dcti_5_IFF_IFF1_RST,
      O => U_DCT1D_latchbuf_reg_7_Q(5)
    );
  dcti_5_IFF_IFFDMUX_7719 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti_5_INBUF,
      O => dcti_5_IFF_IFFDMUX
    );
  dcti_5_IFF_ISR_USED_7720 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcti_5_IFF_ISR_USED
    );
  dcti_5_IFF_ICLK1INV_7721 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcti_5_IFF_ICLK1INV
    );
  dcti_5_IFF_ICEINV_7722 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => dcti_5_IFF_ICEINV
    );
  dcti_4_IFF_IFFDMUX_7723 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti_4_INBUF,
      O => dcti_4_IFF_IFFDMUX
    );
  dcti_4_IFF_ICLK1INV_7724 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcti_4_IFF_ICLK1INV
    );
  dcti_4_IFF_ICEINV_7725 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc2n465,
      O => dcti_4_IFF_ICEINV
    );
  U_DCT1D_reg_latchbuf_reg_7_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcti_4_IFF_IFFDMUX,
      CE => dcti_4_IFF_ICEINV,
      CLK => dcti_4_IFF_ICLK1INV,
      SET => GND,
      RST => dcti_4_IFF_IFF1_RST,
      O => U_DCT1D_latchbuf_reg_7_Q(4)
    );
  dcti_4_IFF_IFF1_RSTOR : X_OR2
    port map (
      I0 => dcti_4_IFF_IFF1_RSTAND,
      I1 => GSR,
      O => dcti_4_IFF_IFF1_RST
    );
  dcti_4_IFF_IFF1_RSTAND_7726 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcti_4_IFF_IFF1_RSTAND
    );
  dcto_7_OUTPUT_OFF_O1INV_7727 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491(19),
      O => dcto_7_OUTPUT_OFF_O1INV
    );
  dcto_7_OUTPUT_OFF_OCEINV_7728 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => dcto_7_OUTPUT_OFF_OCEINV
    );
  dcto_7_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_dup0(7),
      O => dcto_7_O
    );
  dcto_7_OUTPUT_OTCLK1INV_7729 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto_7_OUTPUT_OTCLK1INV
    );
  U_DCT2D_reg_dcto_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto_7_OUTPUT_OFF_O1INV,
      CE => dcto_7_OUTPUT_OFF_OCEINV,
      CLK => dcto_7_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto_7_OUTPUT_OFF_OFF1_RST,
      O => dcto_dup0(7)
    );
  dcto_7_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto_7_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto_7_OUTPUT_OFF_OFF1_RST
    );
  dcto_7_OUTPUT_OFF_OFF1_RSTAND_7730 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto_7_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto_8_OUTPUT_OFF_O1INV_7731 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491(20),
      O => dcto_8_OUTPUT_OFF_O1INV
    );
  dcto_8_OUTPUT_OFF_OCEINV_7732 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => dcto_8_OUTPUT_OFF_OCEINV
    );
  dcto_8_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_dup0(8),
      O => dcto_8_O
    );
  dcto_8_OUTPUT_OTCLK1INV_7733 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto_8_OUTPUT_OTCLK1INV
    );
  U_DCT2D_reg_dcto_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto_8_OUTPUT_OFF_O1INV,
      CE => dcto_8_OUTPUT_OFF_OCEINV,
      CLK => dcto_8_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto_8_OUTPUT_OFF_OFF1_RST,
      O => dcto_dup0(8)
    );
  dcto_8_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto_8_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto_8_OUTPUT_OFF_OFF1_RST
    );
  dcto_8_OUTPUT_OFF_OFF1_RSTAND_7734 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto_8_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto_9_OUTPUT_OFF_O1INV_7735 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_rtlc5n1491(21),
      O => dcto_9_OUTPUT_OFF_O1INV
    );
  dcto_9_OUTPUT_OFF_OCEINV_7736 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT2D_state_reg(1),
      O => dcto_9_OUTPUT_OFF_OCEINV
    );
  dcto_9_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcto_dup0(9),
      O => dcto_9_O
    );
  dcto_9_OUTPUT_OTCLK1INV_7737 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto_9_OUTPUT_OTCLK1INV
    );
  U_DCT2D_reg_dcto_9_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto_9_OUTPUT_OFF_O1INV,
      CE => dcto_9_OUTPUT_OFF_OCEINV,
      CLK => dcto_9_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto_9_OUTPUT_OFF_OFF1_RST,
      O => dcto_dup0(9)
    );
  dcto_9_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto_9_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto_9_OUTPUT_OFF_OFF1_RST
    );
  dcto_9_OUTPUT_OFF_OFF1_RSTAND_7738 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto_9_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto1_3_OUTPUT_OFF_O1INV_7739 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n2657,
      O => dcto1_3_OUTPUT_OFF_O1INV
    );
  dcto1_3_OUTPUT_OFF_OCEINV_7740 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => dcto1_3_OUTPUT_OFF_OCEINV
    );
  dcto1_3_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_3_repl0,
      O => dcto1_3_O
    );
  dcto1_3_OUTPUT_OTCLK1INV_7741 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto1_3_OUTPUT_OTCLK1INV
    );
  U_DCT1D_reg_ramdatai_s_3_repl0 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto1_3_OUTPUT_OFF_O1INV,
      CE => dcto1_3_OUTPUT_OFF_OCEINV,
      CLK => dcto1_3_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto1_3_OUTPUT_OFF_OFF1_RST,
      O => ramdatai_3_repl0
    );
  dcto1_3_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto1_3_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto1_3_OUTPUT_OFF_OFF1_RST
    );
  dcto1_3_OUTPUT_OFF_OFF1_RSTAND_7742 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto1_3_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto1_4_OUTPUT_OFF_O1INV_7743 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n2656,
      O => dcto1_4_OUTPUT_OFF_O1INV
    );
  dcto1_4_OUTPUT_OFF_OCEINV_7744 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => dcto1_4_OUTPUT_OFF_OCEINV
    );
  dcto1_4_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_4_repl0,
      O => dcto1_4_O
    );
  dcto1_4_OUTPUT_OTCLK1INV_7745 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto1_4_OUTPUT_OTCLK1INV
    );
  U_DCT1D_reg_ramdatai_s_4_repl0 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto1_4_OUTPUT_OFF_O1INV,
      CE => dcto1_4_OUTPUT_OFF_OCEINV,
      CLK => dcto1_4_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto1_4_OUTPUT_OFF_OFF1_RST,
      O => ramdatai_4_repl0
    );
  dcto1_4_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto1_4_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto1_4_OUTPUT_OFF_OFF1_RST
    );
  dcto1_4_OUTPUT_OFF_OFF1_RSTAND_7746 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto1_4_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto1_5_OUTPUT_OFF_O1INV_7747 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n2655,
      O => dcto1_5_OUTPUT_OFF_O1INV
    );
  dcto1_5_OUTPUT_OFF_OCEINV_7748 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => dcto1_5_OUTPUT_OFF_OCEINV
    );
  dcto1_5_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_5_repl0,
      O => dcto1_5_O
    );
  dcto1_5_OUTPUT_OTCLK1INV_7749 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto1_5_OUTPUT_OTCLK1INV
    );
  dcto1_9_OUTPUT_OFF_O1INV_7750 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n2651,
      O => dcto1_9_OUTPUT_OFF_O1INV
    );
  dcto1_9_OUTPUT_OFF_OCEINV_7751 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => dcto1_9_OUTPUT_OFF_OCEINV
    );
  dcto1_9_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_9_repl0,
      O => dcto1_9_O
    );
  dcto1_9_OUTPUT_OTCLK1INV_7752 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto1_9_OUTPUT_OTCLK1INV
    );
  U_DCT1D_reg_ramdatai_s_9_repl0 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto1_9_OUTPUT_OFF_O1INV,
      CE => dcto1_9_OUTPUT_OFF_OCEINV,
      CLK => dcto1_9_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto1_9_OUTPUT_OFF_OFF1_RST,
      O => ramdatai_9_repl0
    );
  dcto1_9_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto1_9_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto1_9_OUTPUT_OFF_OFF1_RST
    );
  dcto1_9_OUTPUT_OFF_OFF1_RSTAND_7753 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto1_9_OUTPUT_OFF_OFF1_RSTAND
    );
  U_DCT2D_ix1822z1331 : X_LUT4
    generic map(
      INIT => X"0302"
    )
    port map (
      ADR0 => requestrd_s,
      ADR1 => U_DCT2D_state_reg(1),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => U_DCT2D_istate_reg(1),
      O => U_DCT2D_nx1822z2
    );
  U_DCT1D_reg_ramdatai_s_5_repl0 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto1_5_OUTPUT_OFF_O1INV,
      CE => dcto1_5_OUTPUT_OFF_OCEINV,
      CLK => dcto1_5_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto1_5_OUTPUT_OFF_OFF1_RST,
      O => ramdatai_5_repl0
    );
  dcto1_5_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto1_5_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto1_5_OUTPUT_OFF_OFF1_RST
    );
  dcto1_5_OUTPUT_OFF_OFF1_RSTAND_7754 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto1_5_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto1_6_OUTPUT_OFF_O1INV_7755 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n2654,
      O => dcto1_6_OUTPUT_OFF_O1INV
    );
  dcto1_6_OUTPUT_OFF_OCEINV_7756 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => dcto1_6_OUTPUT_OFF_OCEINV
    );
  dcto1_6_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_6_repl0,
      O => dcto1_6_O
    );
  dcto1_6_OUTPUT_OTCLK1INV_7757 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto1_6_OUTPUT_OTCLK1INV
    );
  U_DCT1D_reg_ramdatai_s_6_repl0 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto1_6_OUTPUT_OFF_O1INV,
      CE => dcto1_6_OUTPUT_OFF_OCEINV,
      CLK => dcto1_6_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto1_6_OUTPUT_OFF_OFF1_RST,
      O => ramdatai_6_repl0
    );
  dcto1_6_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto1_6_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto1_6_OUTPUT_OFF_OFF1_RST
    );
  dcto1_6_OUTPUT_OFF_OFF1_RSTAND_7758 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto1_6_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto1_7_OUTPUT_OFF_O1INV_7759 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n2653,
      O => dcto1_7_OUTPUT_OFF_O1INV
    );
  dcto1_7_OUTPUT_OFF_OCEINV_7760 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => dcto1_7_OUTPUT_OFF_OCEINV
    );
  dcto1_7_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_7_repl0,
      O => dcto1_7_O
    );
  dcto1_7_OUTPUT_OTCLK1INV_7761 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto1_7_OUTPUT_OTCLK1INV
    );
  U_DCT1D_reg_ramdatai_s_7_repl0 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto1_7_OUTPUT_OFF_O1INV,
      CE => dcto1_7_OUTPUT_OFF_OCEINV,
      CLK => dcto1_7_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto1_7_OUTPUT_OFF_OFF1_RST,
      O => ramdatai_7_repl0
    );
  dcto1_7_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto1_7_OUTPUT_OFF_OFF1_RSTAND,
      I1 => GSR,
      O => dcto1_7_OUTPUT_OFF_OFF1_RST
    );
  dcto1_7_OUTPUT_OFF_OFF1_RSTAND_7762 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto1_7_OUTPUT_OFF_OFF1_RSTAND
    );
  dcto1_8_OUTPUT_OFF_OFF1_RSTOR : X_OR2
    port map (
      I0 => dcto1_8_OUTPUT_OFF_OSR_USED,
      I1 => GSR,
      O => dcto1_8_OUTPUT_OFF_OFF1_RST
    );
  U_DCT1D_reg_ramdatai_s_8_repl0 : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => dcto1_8_OUTPUT_OFF_O1INV,
      CE => dcto1_8_OUTPUT_OFF_OCEINV,
      CLK => dcto1_8_OUTPUT_OTCLK1INV,
      SET => GND,
      RST => dcto1_8_OUTPUT_OFF_OFF1_RST,
      O => ramdatai_8_repl0
    );
  dcto1_8_OUTPUT_OFF_O1INV_7763 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_rtlc5n2652,
      O => dcto1_8_OUTPUT_OFF_O1INV
    );
  dcto1_8_OUTPUT_OFF_OCEINV_7764 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => U_DCT1D_state_reg(1),
      O => dcto1_8_OUTPUT_OFF_OCEINV
    );
  dcto1_8_OUTPUT_OFF_OSR_USED_7765 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => dcto1_8_OUTPUT_OFF_OSR_USED
    );
  dcto1_8_OUTPUT_OFF_OMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => ramdatai_8_repl0,
      O => dcto1_8_O
    );
  dcto1_8_OUTPUT_OTCLK1INV_7766 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_int,
      O => dcto1_8_OUTPUT_OTCLK1INV
    );
  U_DCT2D_reg_istate_reg_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_istate_reg_1_DYMUX,
      CE => U_DCT2D_istate_reg_1_CEINV,
      CLK => U_DCT2D_istate_reg_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_istate_reg_1_FFY_RST,
      O => U_DCT2D_istate_reg(0)
    );
  U_DCT2D_istate_reg_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_istate_reg_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_istate_reg_1_FFY_RST
    );
  U_DCT2D_ix1822z14465 : X_LUT4
    generic map(
      INIT => X"335F"
    )
    port map (
      ADR0 => U_DCT2D_istate_reg(1),
      ADR1 => U_DCT2D_completed_reg,
      ADR2 => reqrdfail_s,
      ADR3 => U_DCT2D_istate_reg(0),
      O => U_DCT2D_rtlcn348
    );
  ix60496z1327 : X_LUT4
    generic map(
      INIT => X"F5F5"
    )
    port map (
      ADR0 => U_DBUFCTL_mem1_full_reg,
      ADR1 => VCC,
      ADR2 => U_DBUFCTL_mem1_lock_reg,
      ADR3 => VCC,
      O => memswitchrd_s_F
    );
  U_DCT2D_reg_istate_reg_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_istate_reg_1_DXMUX,
      CE => U_DCT2D_istate_reg_1_CEINV,
      CLK => U_DCT2D_istate_reg_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_istate_reg_1_FFX_RST,
      O => U_DCT2D_istate_reg(1)
    );
  U_DCT2D_istate_reg_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_istate_reg_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_istate_reg_1_FFX_RST
    );
  U_DBUFCTL_reg_memswitchrd_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => memswitchrd_s_DXMUX,
      CE => memswitchrd_s_CEINV,
      CLK => memswitchrd_s_CLKINV,
      SET => GND,
      RST => memswitchrd_s_FFX_RST,
      O => memswitchrd_s
    );
  memswitchrd_s_FFX_RSTOR : X_OR2
    port map (
      I0 => memswitchrd_s_FFX_RSTAND,
      I1 => GSR,
      O => memswitchrd_s_FFX_RST
    );
  memswitchrd_s_FFX_RSTAND_7767 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => memswitchrd_s_FFX_RSTAND
    );
  U_DCT2D_ix50410z1320 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => ramraddro_s(4),
      ADR2 => ramraddro_s(3),
      ADR3 => VCC,
      O => U_DCT2D_nx50410z1
    );
  U_DCT2D_modgen_counter_ramraddro_reg_q_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramraddro_s_5_DYMUX,
      CE => ramraddro_s_5_CEINV,
      CLK => ramraddro_s_5_CLKINV,
      SET => GND,
      RST => ramraddro_s_5_FFY_RST,
      O => ramraddro_s(4)
    );
  ramraddro_s_5_FFY_RSTOR : X_OR2
    port map (
      I0 => ramraddro_s_5_SRINV,
      I1 => GSR,
      O => ramraddro_s_5_FFY_RST
    );
  U_DCT2D_ix6411z13778 : X_LUT4
    generic map(
      INIT => X"20F0"
    )
    port map (
      ADR0 => U_DCT2D_completed_reg,
      ADR1 => U_DCT2D_rtlcn65,
      ADR2 => U_DCT2D_rtlc2n582,
      ADR3 => U_DCT2D_istate_reg(0),
      O => U_DCT2D_rtlc2n580_F
    );
  U_DCT2D_ix14976z1321 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_4_10_Q,
      ADR3 => U_DCT2D_latchbuf_reg_3_10_Q,
      O => U_DCT2D_nx14976z1_F
    );
  U_DCT2D_ix36450z1320 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT2D_col_reg(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_col_reg(1),
      O => U_DCT2D_nx36450z1
    );
  U_DCT2D_modgen_counter_col_reg_reg_q_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_col_reg_0_DYMUX,
      CE => U_DCT2D_col_reg_0_CEINV,
      CLK => U_DCT2D_col_reg_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_col_reg_0_FFY_RST,
      O => U_DCT2D_col_reg(1)
    );
  U_DCT2D_col_reg_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_col_reg_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_col_reg_0_FFY_RST
    );
  U_DCT2D_modgen_counter_col_reg_reg_q_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_col_reg_0_DXMUX,
      CE => U_DCT2D_col_reg_0_CEINV,
      CLK => U_DCT2D_col_reg_0_CLKINV,
      SET => GND,
      RST => U_DCT2D_col_reg_0_FFX_RST,
      O => U_DCT2D_col_reg(0)
    );
  U_DCT2D_col_reg_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_col_reg_0_SRINV,
      I1 => GSR,
      O => U_DCT2D_col_reg_0_FFX_RST
    );
  U_DCT1D_ix36450z1320 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_col_reg(1),
      ADR2 => U_DCT1D_col_reg(0),
      ADR3 => VCC,
      O => U_DCT1D_nx36450z1
    );
  U_DCT1D_modgen_counter_col_reg_reg_q_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_col_reg_0_DYMUX,
      CE => U_DCT1D_col_reg_0_CEINV,
      CLK => U_DCT1D_col_reg_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_col_reg_0_FFY_RST,
      O => U_DCT1D_col_reg(1)
    );
  U_DCT1D_col_reg_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_col_reg_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_col_reg_0_FFY_RST
    );
  U_DCT2D_ix22763z1321 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_2_10_Q,
      ADR2 => U_DCT2D_latchbuf_reg_5_10_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx8385z1_G
    );
  ix53675z3790 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => memswitchrd_s,
      ADR2 => ramdatao1_s(8),
      ADR3 => ramdatao2_s(8),
      O => ramdatao_s(8)
    );
  U_DCT2D_reg_latchbuf_reg_7_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_5_DYMUX,
      CE => U_DCT2D_latchbuf_reg_7_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_7_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_7_5_FFY_RST,
      O => U_DCT2D_latchbuf_reg_7_4_Q
    );
  U_DCT2D_latchbuf_reg_7_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_7_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_7_5_FFY_RST
    );
  ix53675z3792 : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => ramdatao1_s(6),
      ADR1 => VCC,
      ADR2 => memswitchrd_s,
      ADR3 => ramdatao2_s(6),
      O => ramdatao_s(6)
    );
  ix53675z3793 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => memswitchrd_s,
      ADR1 => ramdatao1_s(5),
      ADR2 => ramdatao2_s(5),
      ADR3 => VCC,
      O => ramdatao_s(5)
    );
  U_DCT2D_reg_latchbuf_reg_7_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_5_DXMUX,
      CE => U_DCT2D_latchbuf_reg_7_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_7_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_7_5_FFX_RST,
      O => U_DCT2D_latchbuf_reg_7_5_Q
    );
  U_DCT2D_latchbuf_reg_7_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_7_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_7_5_FFX_RST
    );
  U_DCT2D_ix65206z45474 : X_LUT4
    generic map(
      INIT => X"E14B"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => rome2datao10_s(13),
      ADR2 => U_DCT2D_rtlc5n1484(23),
      ADR3 => romo2datao10_s(13),
      O => U_DCT2D_nx65206z571_G
    );
  U_DCT2D_reg_latchbuf_reg_7_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_7_DYMUX,
      CE => U_DCT2D_latchbuf_reg_7_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_7_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_7_7_FFY_RST,
      O => U_DCT2D_latchbuf_reg_7_6_Q
    );
  U_DCT2D_latchbuf_reg_7_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_7_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_7_7_FFY_RST
    );
  ix53675z3791 : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => ramdatao2_s(7),
      ADR1 => VCC,
      ADR2 => memswitchrd_s,
      ADR3 => ramdatao1_s(7),
      O => ramdatao_s(7)
    );
  U_DCT2D_reg_latchbuf_reg_7_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_7_DXMUX,
      CE => U_DCT2D_latchbuf_reg_7_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_7_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_7_7_FFX_RST,
      O => U_DCT2D_latchbuf_reg_7_7_Q
    );
  U_DCT2D_latchbuf_reg_7_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_7_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_7_7_FFX_RST
    );
  U_DCT2D_ix65206z31069 : X_LUT4
    generic map(
      INIT => X"3CAA"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1498(22),
      ADR1 => U_DCT2D_rtlc5n1482(19),
      ADR2 => U_DCT2D_rtlc5n1483(21),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z252_G
    );
  ix31259z1396 : X_LUT4
    generic map(
      INIT => X"7733"
    )
    port map (
      ADR0 => memswitchwr_s,
      ADR1 => U_DBUFCTL_rtlcn38,
      ADR2 => VCC,
      ADR3 => releasewr_s,
      O => nx31259z2
    );
  U_DCT2D_ix2819z1318 : X_LUT4
    generic map(
      INIT => X"0202"
    )
    port map (
      ADR0 => U_DCT2D_istate_reg(1),
      ADR1 => U_DCT2D_istate_reg(0),
      ADR2 => reqrdfail_s,
      ADR3 => VCC,
      O => U_DCT2D_rtlc2_istate_reg_fsm_SS9_n171(0)
    );
  U_DCT2D_ix35453z1420 : X_LUT4
    generic map(
      INIT => X"66CC"
    )
    port map (
      ADR0 => U_DCT2D_col_reg(1),
      ADR1 => U_DCT2D_col_reg(2),
      ADR2 => VCC,
      ADR3 => U_DCT2D_col_reg(0),
      O => U_DCT2D_nx35453z1
    );
  U_DCT2D_modgen_counter_col_reg_reg_q_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_col_reg_2_DYMUX,
      CE => U_DCT2D_col_reg_2_CEINV,
      CLK => U_DCT2D_col_reg_2_CLKINV,
      SET => GND,
      RST => U_DCT2D_col_reg_2_FFY_RST,
      O => U_DCT2D_col_reg(2)
    );
  U_DCT2D_col_reg_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_col_reg_2_FFY_RSTAND,
      I1 => GSR,
      O => U_DCT2D_col_reg_2_FFY_RST
    );
  U_DCT2D_col_reg_2_FFY_RSTAND_7768 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_col_reg_2_FFY_RSTAND
    );
  U_DCT1D_ix35453z1420 : X_LUT4
    generic map(
      INIT => X"3FC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_col_reg(0),
      ADR2 => U_DCT1D_col_reg(1),
      ADR3 => U_DCT1D_col_reg(2),
      O => U_DCT1D_nx35453z1
    );
  U_DCT1D_modgen_counter_col_reg_reg_q_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_col_reg_2_DYMUX,
      CE => U_DCT1D_col_reg_2_CEINV,
      CLK => U_DCT1D_col_reg_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_col_reg_2_FFY_RST,
      O => U_DCT1D_col_reg(2)
    );
  U_DCT1D_col_reg_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_col_reg_2_FFY_RSTAND,
      I1 => GSR,
      O => U_DCT1D_col_reg_2_FFY_RST
    );
  U_DCT1D_col_reg_2_FFY_RSTAND_7769 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_col_reg_2_FFY_RSTAND
    );
  U_DCT1D_ix9237z10020 : X_LUT4
    generic map(
      INIT => X"4050"
    )
    port map (
      ADR0 => reqwrfail_s,
      ADR1 => U_DCT1D_NOT_rtlcs1,
      ADR2 => idv_int,
      ADR3 => U_DCT1D_ready,
      O => U_DCT1D_ready_G
    );
  U_DCT1D_reg_ready_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_ready_DYMUX,
      CE => U_DCT1D_ready_CEINV,
      CLK => U_DCT1D_ready_CLKINV,
      SET => GND,
      RST => U_DCT1D_ready_FFY_RST,
      O => U_DCT1D_ready
    );
  U_DCT1D_ready_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_ready_FFY_RSTAND,
      I1 => GSR,
      O => U_DCT1D_ready_FFY_RST
    );
  U_DCT1D_ready_FFY_RSTAND_7770 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_ready_FFY_RSTAND
    );
  U_DCT1D_ix13345z1442 : X_LUT4
    generic map(
      INIT => X"A000"
    )
    port map (
      ADR0 => U_DCT1D_istate_reg(0),
      ADR1 => VCC,
      ADR2 => idv_int,
      ADR3 => U_DCT1D_ready,
      O => U_DCT1D_ready_F
    );
  U_DCT1D_ix53037z1420 : X_LUT4
    generic map(
      INIT => X"7788"
    )
    port map (
      ADR0 => U_DCT1D_row_reg(0),
      ADR1 => U_DCT1D_row_reg(1),
      ADR2 => VCC,
      ADR3 => U_DCT1D_row_reg(2),
      O => U_DCT1D_nx53037z1
    );
  ix31259z53283 : X_LUT4
    generic map(
      INIT => X"F3BB"
    )
    port map (
      ADR0 => requestwr_s,
      ADR1 => U_DBUFCTL_rtlcn38,
      ADR2 => requestrd_s,
      ADR3 => U_DBUFCTL_mem1_full_reg,
      O => nx31259z1
    );
  ix40249z1328 : X_LUT4
    generic map(
      INIT => X"FFF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DBUFCTL_mem1_lock_reg,
      ADR3 => U_DBUFCTL_mem1_full_reg,
      O => memswitchwr_s_G
    );
  U_DCT2D_ix51407z1420 : X_LUT4
    generic map(
      INIT => X"3FC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => ramraddro_s(4),
      ADR2 => ramraddro_s(3),
      ADR3 => ramraddro_s(5),
      O => U_DCT2D_nx51407z1
    );
  U_DCT2D_modgen_counter_ramraddro_reg_q_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramraddro_s_5_DXMUX,
      CE => ramraddro_s_5_CEINV,
      CLK => ramraddro_s_5_CLKINV,
      SET => GND,
      RST => ramraddro_s_5_FFX_RST,
      O => ramraddro_s(5)
    );
  ramraddro_s_5_FFX_RSTOR : X_OR2
    port map (
      I0 => ramraddro_s_5_SRINV,
      I1 => GSR,
      O => ramraddro_s_5_FFX_RST
    );
  U_DBUFCTL_reg_memswitchwr_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => memswitchwr_s_DYMUX,
      CE => memswitchwr_s_CEINV,
      CLK => memswitchwr_s_CLKINV,
      SET => GND,
      RST => memswitchwr_s_FFY_RST,
      O => memswitchwr_s
    );
  memswitchwr_s_FFY_RSTOR : X_OR2
    port map (
      I0 => memswitchwr_s_FFY_RSTAND,
      I1 => GSR,
      O => memswitchwr_s_FFY_RST
    );
  memswitchwr_s_FFY_RSTAND_7771 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => memswitchwr_s_FFY_RSTAND
    );
  ix43562z803 : X_LUT4
    generic map(
      INIT => X"FDFF"
    )
    port map (
      ADR0 => requestwr_s,
      ADR1 => U_DBUFCTL_mem2_lock_reg,
      ADR2 => U_DBUFCTL_mem2_full_reg,
      ADR3 => U_DBUFCTL_rtlcn1,
      O => memswitchwr_s_F
    );
  ix24581z1505 : X_LUT4
    generic map(
      INIT => X"F3FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => releaserd_s,
      ADR2 => memswitchrd_s,
      ADR3 => U_DBUFCTL_mem1_lock_reg,
      O => U_DBUFCTL_mem1_full_reg_G
    );
  U_DBUFCTL_reg_mem1_full_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DBUFCTL_mem1_full_reg_DYMUX,
      CE => U_DBUFCTL_mem1_full_reg_CEINV,
      CLK => U_DBUFCTL_mem1_full_reg_CLKINV,
      SET => GND,
      RST => U_DBUFCTL_mem1_full_reg_FFY_RST,
      O => U_DBUFCTL_mem1_full_reg
    );
  U_DBUFCTL_mem1_full_reg_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DBUFCTL_mem1_full_reg_FFY_RSTAND,
      I1 => GSR,
      O => U_DBUFCTL_mem1_full_reg_FFY_RST
    );
  U_DBUFCTL_mem1_full_reg_FFY_RSTAND_7772 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DBUFCTL_mem1_full_reg_FFY_RSTAND
    );
  ix24581z17954 : X_LUT4
    generic map(
      INIT => X"2F0F"
    )
    port map (
      ADR0 => U_DBUFCTL_mem1_lock_reg,
      ADR1 => memswitchwr_s,
      ADR2 => U_DBUFCTL_rtlcn38,
      ADR3 => releasewr_s,
      O => U_DBUFCTL_mem1_full_reg_F
    );
  U_DCT1D_modgen_counter_row_reg_reg_q_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_row_reg_2_DYMUX,
      CE => U_DCT1D_row_reg_2_CEINV,
      CLK => U_DCT1D_row_reg_2_CLKINV,
      SET => GND,
      RST => U_DCT1D_row_reg_2_FFY_RST,
      O => U_DCT1D_row_reg(2)
    );
  U_DCT1D_row_reg_2_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_row_reg_2_FFY_RSTAND,
      I1 => GSR,
      O => U_DCT1D_row_reg_2_FFY_RST
    );
  U_DCT1D_row_reg_2_FFY_RSTAND_7773 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_row_reg_2_FFY_RSTAND
    );
  U_DCT2D_ix46656z1540 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(1),
      ADR1 => U_DCT2D_col_tmp_reg(1),
      ADR2 => VCC,
      ADR3 => U_DCT2D_col_reg(1),
      O => U_DCT2D_rtlc5_romeaddro0_SS3_n342(4)
    );
  U_DCT2D_reg_romeaddro10_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro0_s_5_DYMUX,
      CE => rome2addro0_s_5_CEINV,
      CLK => rome2addro0_s_5_CLKINV,
      SET => GND,
      RST => rome2addro0_s_5_FFY_RST,
      O => rome2addro0_s(4)
    );
  rome2addro0_s_5_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro0_s_5_SRINV,
      I1 => GSR,
      O => rome2addro0_s_5_FFY_RST
    );
  U_DCT2D_ix45659z1540 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(1),
      ADR1 => VCC,
      ADR2 => U_DCT2D_col_reg(2),
      ADR3 => U_DCT2D_col_tmp_reg(2),
      O => U_DCT2D_rtlc5_romeaddro0_SS3_n342(5)
    );
  U_DCT1D_ix54913z1540 : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => U_DCT1D_col_reg(1),
      ADR1 => U_DCT1D_col_tmp_reg(1),
      ADR2 => U_DCT1D_state_reg(1),
      ADR3 => VCC,
      O => U_DCT1D_rtlc5_romeaddro0_SS4_n350(4)
    );
  U_DCT2D_reg_romeaddro10_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro0_s_5_DXMUX,
      CE => rome2addro0_s_5_CEINV,
      CLK => rome2addro0_s_5_CLKINV,
      SET => GND,
      RST => rome2addro0_s_5_FFX_RST,
      O => rome2addro0_s(5)
    );
  rome2addro0_s_5_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro0_s_5_SRINV,
      I1 => GSR,
      O => rome2addro0_s_5_FFX_RST
    );
  U_DCT1D_reg_romeaddro8_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro0_s_5_DYMUX,
      CE => romeaddro0_s_5_CEINV,
      CLK => romeaddro0_s_5_CLKINV,
      SET => GND,
      RST => romeaddro0_s_5_FFY_RST,
      O => romeaddro0_s(4)
    );
  romeaddro0_s_5_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro0_s_5_SRINV,
      I1 => GSR,
      O => romeaddro0_s_5_FFY_RST
    );
  U_DCT1D_ix53916z1540 : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => U_DCT1D_col_reg(2),
      ADR1 => VCC,
      ADR2 => U_DCT1D_state_reg(1),
      ADR3 => U_DCT1D_col_tmp_reg(2),
      O => U_DCT1D_rtlc5_romeaddro0_SS4_n350(5)
    );
  U_DCT1D_reg_romeaddro8_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro0_s_5_DXMUX,
      CE => romeaddro0_s_5_CEINV,
      CLK => romeaddro0_s_5_CLKINV,
      SET => GND,
      RST => romeaddro0_s_5_FFX_RST,
      O => romeaddro0_s(5)
    );
  romeaddro0_s_5_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro0_s_5_SRINV,
      I1 => GSR,
      O => romeaddro0_s_5_FFX_RST
    );
  ix50240z1441 : X_LUT4
    generic map(
      INIT => X"77FF"
    )
    port map (
      ADR0 => U_DBUFCTL_mem2_lock_reg,
      ADR1 => memswitchrd_s,
      ADR2 => VCC,
      ADR3 => releaserd_s,
      O => U_DBUFCTL_mem2_full_reg_G
    );
  U_DBUFCTL_reg_mem1_lock_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DBUFCTL_mem1_lock_reg_DYMUX,
      CE => U_DBUFCTL_mem1_lock_reg_CEINV,
      CLK => U_DBUFCTL_mem1_lock_reg_CLKINV,
      SET => GND,
      RST => U_DBUFCTL_mem1_lock_reg_FFY_RST,
      O => U_DBUFCTL_mem1_lock_reg
    );
  U_DBUFCTL_mem1_lock_reg_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DBUFCTL_mem1_lock_reg_FFY_RSTAND,
      I1 => GSR,
      O => U_DBUFCTL_mem1_lock_reg_FFY_RST
    );
  U_DBUFCTL_mem1_lock_reg_FFY_RSTAND_7774 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DBUFCTL_mem1_lock_reg_FFY_RSTAND
    );
  ix1552z1322 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => ramwe_s,
      ADR2 => VCC,
      ADR3 => memswitchwr_s,
      O => U_DBUFCTL_mem1_lock_reg_F
    );
  U_DBUFCTL_reg_mem2_full_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DBUFCTL_mem2_full_reg_DYMUX,
      CE => U_DBUFCTL_mem2_full_reg_CEINV,
      CLK => U_DBUFCTL_mem2_full_reg_CLKINV,
      SET => GND,
      RST => U_DBUFCTL_mem2_full_reg_FFY_RST,
      O => U_DBUFCTL_mem2_full_reg
    );
  U_DBUFCTL_mem2_full_reg_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DBUFCTL_mem2_full_reg_FFY_RSTAND,
      I1 => GSR,
      O => U_DBUFCTL_mem2_full_reg_FFY_RST
    );
  U_DBUFCTL_mem2_full_reg_FFY_RSTAND_7775 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DBUFCTL_mem2_full_reg_FFY_RSTAND
    );
  ix43562z12236 : X_LUT4
    generic map(
      INIT => X"4CCC"
    )
    port map (
      ADR0 => releasewr_s,
      ADR1 => U_DBUFCTL_rtlcn42,
      ADR2 => memswitchwr_s,
      ADR3 => U_DBUFCTL_mem2_lock_reg,
      O => U_DBUFCTL_rtlcn76
    );
  ix43562z34340 : X_LUT4
    generic map(
      INIT => X"8F0F"
    )
    port map (
      ADR0 => U_DBUFCTL_mem2_lock_reg,
      ADR1 => memswitchwr_s,
      ADR2 => U_DBUFCTL_rtlcn42,
      ADR3 => releasewr_s,
      O => U_DBUFCTL_mem2_full_reg_F
    );
  U_DBUFCTL_reg_mem2_lock_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DBUFCTL_mem2_lock_reg_DYMUX,
      CE => U_DBUFCTL_mem2_lock_reg_CEINV,
      CLK => U_DBUFCTL_mem2_lock_reg_CLKINV,
      SET => GND,
      RST => U_DBUFCTL_mem2_lock_reg_FFY_RST,
      O => U_DBUFCTL_mem2_lock_reg
    );
  U_DBUFCTL_mem2_lock_reg_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DBUFCTL_mem2_lock_reg_FFY_RSTAND,
      I1 => GSR,
      O => U_DBUFCTL_mem2_lock_reg_FFY_RST
    );
  U_DBUFCTL_mem2_lock_reg_FFY_RSTAND_7776 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DBUFCTL_mem2_lock_reg_FFY_RSTAND
    );
  ix21201z1316 : X_LUT4
    generic map(
      INIT => X"4444"
    )
    port map (
      ADR0 => memswitchwr_s,
      ADR1 => ramwe_s,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DBUFCTL_mem2_lock_reg_F
    );
  U_DCT2D_ix39898z14165 : X_LUT4
    generic map(
      INIT => X"3233"
    )
    port map (
      ADR0 => ramraddro_s(2),
      ADR1 => ramraddro_s(1),
      ADR2 => ramraddro_s(0),
      ADR3 => U_DCT2D_colram_reg(3),
      O => U_DCT2D_nx39898z1
    );
  U_DCT2D_modgen_counter_colram_reg_reg_q_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramraddro_s_0_DYMUX,
      CE => ramraddro_s_0_CEINV,
      CLK => ramraddro_s_0_CLKINV,
      SET => GND,
      RST => ramraddro_s_0_FFY_RST,
      O => ramraddro_s(0)
    );
  ramraddro_s_0_FFY_RSTOR : X_OR2
    port map (
      I0 => ramraddro_s_0_FFY_RSTAND,
      I1 => GSR,
      O => ramraddro_s_0_FFY_RST
    );
  ramraddro_s_0_FFY_RSTAND_7777 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramraddro_s_0_FFY_RSTAND
    );
  U_DCT2D_ix13345z62978 : X_LUT4
    generic map(
      INIT => X"AAA8"
    )
    port map (
      ADR0 => U_DCT2D_NOT_rtlc2n488,
      ADR1 => ramraddro_s(2),
      ADR2 => U_DCT2D_nx49413z1,
      ADR3 => U_DCT2D_colram_reg(3),
      O => ramraddro_s_0_F
    );
  U_DCT2D_modgen_counter_colram_reg_reg_q_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramraddro_s_1_DYMUX,
      CE => ramraddro_s_1_CEINV,
      CLK => ramraddro_s_1_CLKINV,
      SET => GND,
      RST => ramraddro_s_1_FFY_RST,
      O => ramraddro_s(1)
    );
  ramraddro_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => ramraddro_s_1_FFY_RSTAND,
      I1 => GSR,
      O => ramraddro_s_1_FFY_RST
    );
  ramraddro_s_1_FFY_RSTAND_7778 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramraddro_s_1_FFY_RSTAND
    );
  U_DCT2D_ix40895z22903 : X_LUT4
    generic map(
      INIT => X"00FD"
    )
    port map (
      ADR0 => U_DCT2D_colram_reg(3),
      ADR1 => ramraddro_s(0),
      ADR2 => ramraddro_s(1),
      ADR3 => ramraddro_s(2),
      O => U_DCT2D_nx40895z1
    );
  U_DCT2D_ix39898z4643 : X_LUT4
    generic map(
      INIT => X"4404"
    )
    port map (
      ADR0 => U_DCT2D_istate_reg(0),
      ADR1 => U_DCT2D_istate_reg(1),
      ADR2 => U_DCT2D_NOT_rtlcs2,
      ADR3 => ramraddro_s(0),
      O => ramraddro_s_1_F
    );
  U_DCT2D_modgen_counter_colram_reg_reg_q_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramraddro_s_2_DYMUX,
      CE => ramraddro_s_2_CEINV,
      CLK => ramraddro_s_2_CLKINV,
      SET => GND,
      RST => ramraddro_s_2_FFY_RST,
      O => ramraddro_s(2)
    );
  ramraddro_s_2_FFY_RSTOR : X_OR2
    port map (
      I0 => ramraddro_s_2_FFY_RSTAND,
      I1 => GSR,
      O => ramraddro_s_2_FFY_RST
    );
  ramraddro_s_2_FFY_RSTAND_7779 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramraddro_s_2_FFY_RSTAND
    );
  U_DCT1D_ix2819z1321 : X_LUT4
    generic map(
      INIT => X"050F"
    )
    port map (
      ADR0 => U_DCT1D_istate_reg(1),
      ADR1 => VCC,
      ADR2 => U_DCT1D_istate_reg(0),
      ADR3 => U_DCT1D_completed_reg,
      O => U_DCT1D_rtlcn349
    );
  U_DCT1D_reg_latchbuf_reg_4_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_1_DYMUX,
      CE => U_DCT1D_latchbuf_reg_4_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_4_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_4_1_FFY_RST,
      O => U_DCT1D_latchbuf_reg_4_Q(0)
    );
  U_DCT1D_latchbuf_reg_4_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_4_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_4_1_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_4_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_1_DXMUX,
      CE => U_DCT1D_latchbuf_reg_4_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_4_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_4_1_FFX_RST,
      O => U_DCT1D_latchbuf_reg_4_Q(1)
    );
  U_DCT1D_latchbuf_reg_4_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_4_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_4_1_FFX_RST
    );
  U_DCT2D_reg_romoaddro3_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro3_s_1_DYMUX,
      CE => romo2addro3_s_1_CEINV,
      CLK => romo2addro3_s_1_CLKINV,
      SET => GND,
      RST => romo2addro3_s_1_FFY_RST,
      O => romo2addro3_s(0)
    );
  romo2addro3_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro3_s_1_SRINV,
      I1 => GSR,
      O => romo2addro3_s_1_FFY_RST
    );
  U_DCT2D_reg_romoaddro3_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro3_s_1_DXMUX,
      CE => romo2addro3_s_1_CEINV,
      CLK => romo2addro3_s_1_CLKINV,
      SET => GND,
      RST => romo2addro3_s_1_FFX_RST,
      O => romo2addro3_s(1)
    );
  romo2addro3_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro3_s_1_SRINV,
      I1 => GSR,
      O => romo2addro3_s_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_4_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_3_DYMUX,
      CE => U_DCT1D_latchbuf_reg_4_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_4_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_4_3_FFY_RST,
      O => U_DCT1D_latchbuf_reg_4_Q(2)
    );
  U_DCT1D_latchbuf_reg_4_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_4_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_4_3_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_4_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_3_DXMUX,
      CE => U_DCT1D_latchbuf_reg_4_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_4_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_4_3_FFX_RST,
      O => U_DCT1D_latchbuf_reg_4_Q(3)
    );
  U_DCT1D_latchbuf_reg_4_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_4_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_4_3_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_7_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_10_DYMUX,
      CE => U_DCT2D_latchbuf_reg_7_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_7_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_7_10_FFY_RST,
      O => U_DCT2D_latchbuf_reg_7_8_Q
    );
  U_DCT2D_latchbuf_reg_7_10_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_7_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_7_10_FFY_RST
    );
  ix53675z3789 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => memswitchrd_s,
      ADR1 => ramdatao1_s(9),
      ADR2 => ramdatao2_s(9),
      ADR3 => VCC,
      O => ramdatao_s(9)
    );
  U_DCT2D_reg_latchbuf_reg_7_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_10_DXMUX,
      CE => U_DCT2D_latchbuf_reg_7_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_7_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_7_10_FFX_RST,
      O => U_DCT2D_latchbuf_reg_7_10_Q
    );
  U_DCT2D_latchbuf_reg_7_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_7_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_7_10_FFX_RST
    );
  U_DCT1D_ix57999z3363 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => U_DCT1D_istate_reg(0),
      ADR1 => idv_int,
      ADR2 => U_DCT1D_istate_reg(1),
      ADR3 => U_DCT1D_ready,
      O => U_DCT1D_rtlc2n469_G
    );
  U_DCT1D_ix64092z1329 : X_LUT4
    generic map(
      INIT => X"0054"
    )
    port map (
      ADR0 => U_DCT1D_istate_reg(1),
      ADR1 => idv_int,
      ADR2 => requestwr_s,
      ADR3 => U_DCT1D_istate_reg(0),
      O => U_DCT1D_rtlc2n469_F
    );
  U_DCT2D_ix65206z58514 : X_LUT4
    generic map(
      INIT => X"F606"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1492(4),
      ADR1 => rome2datao2_s(2),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => U_DCT2D_rtlc5n1485(4),
      O => U_DCT2D_nx65206z251_G
    );
  U_DCT2D_ix65206z1895 : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1492(4),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => U_DCT2D_rtlc5n1485(4),
      O => U_DCT2D_nx65206z251_F
    );
  U_DCT2D_ix65206z49979 : X_LUT4
    generic map(
      INIT => X"A3AC"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1485(18),
      ADR1 => U_DCT2D_rtlc5n1493(17),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => U_DCT2D_rtlc5n1492(15),
      O => U_DCT2D_nx65206z218_G
    );
  U_DCT2D_ix65206z1830 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => VCC,
      ADR2 => U_DCT2D_rtlc5n1485(15),
      ADR3 => U_DCT2D_rtlc5n1492(15),
      O => U_DCT2D_nx65206z218_F
    );
  U_DCT2D_modgen_counter_ramraddro_reg_q_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramraddro_s_3_DYMUX,
      CE => ramraddro_s_3_CEINV,
      CLK => ramraddro_s_3_CLKINV,
      SET => GND,
      RST => ramraddro_s_3_FFY_RST,
      O => ramraddro_s(3)
    );
  ramraddro_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => ramraddro_s_3_FFY_RSTAND,
      I1 => GSR,
      O => ramraddro_s_3_FFY_RST
    );
  ramraddro_s_3_FFY_RSTAND_7780 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramraddro_s_3_FFY_RSTAND
    );
  U_DCT1D_reg_requestwr_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => requestwr_s_DYMUX,
      CE => requestwr_s_CEINV,
      CLK => requestwr_s_CLKINV,
      SET => GND,
      RST => requestwr_s_FFY_RST,
      O => requestwr_s
    );
  requestwr_s_FFY_RSTOR : X_OR2
    port map (
      I0 => requestwr_s_FFY_RSTAND,
      I1 => GSR,
      O => requestwr_s_FFY_RST
    );
  requestwr_s_FFY_RSTAND_7781 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => requestwr_s_FFY_RSTAND
    );
  ix43562z9510 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => U_DBUFCTL_mem2_full_reg,
      ADR1 => NOT_U_DBUFCTL_rtlc0n25,
      ADR2 => U_DBUFCTL_mem2_lock_reg,
      ADR3 => requestrd_s,
      O => U_DBUFCTL_rtlc4n378_G
    );
  ix60496z1323 : X_LUT4
    generic map(
      INIT => X"CC00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => nx53675z1582,
      ADR2 => VCC,
      ADR3 => requestrd_s,
      O => U_DBUFCTL_rtlc4n374_G
    );
  ix43562z1568 : X_LUT4
    generic map(
      INIT => X"FFBB"
    )
    port map (
      ADR0 => nx43562z1,
      ADR1 => U_DBUFCTL_rtlc4n202,
      ADR2 => VCC,
      ADR3 => nx43562z2,
      O => U_DBUFCTL_rtlc4n378_F
    );
  U_DCT2D_ix15104z1569 : X_LUT4
    generic map(
      INIT => X"FFEE"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(1),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => VCC,
      ADR3 => U_DCT2D_latch_done_reg,
      O => U_DCT2D_rtlc5n1702_G
    );
  U_DCT2D_ix60980z1318 : X_LUT4
    generic map(
      INIT => X"1100"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(1),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => VCC,
      ADR3 => U_DCT2D_latch_done_reg,
      O => U_DCT2D_rtlc5n1702_F
    );
  U_DCT2D_ix30550z1321 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_6_10_Q,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_1_10_Q,
      O => U_DCT2D_nx64938z1_G
    );
  U_DCT1D_ix16101z1442 : X_LUT4
    generic map(
      INIT => X"77FF"
    )
    port map (
      ADR0 => U_DCT1D_col_reg(1),
      ADR1 => U_DCT1D_col_reg(0),
      ADR2 => VCC,
      ADR3 => U_DCT1D_col_reg(2),
      O => U_DCT1D_state_reg_1_G
    );
  ix53675z6340 : X_LUT4
    generic map(
      INIT => X"7530"
    )
    port map (
      ADR0 => U_DBUFCTL_mem1_lock_reg,
      ADR1 => U_DBUFCTL_mem2_lock_reg,
      ADR2 => U_DBUFCTL_mem2_full_reg,
      ADR3 => U_DBUFCTL_mem1_full_reg,
      O => U_DCT2D_rtlc2n581_G
    );
  U_DBUFCTL_reg_reqwrfail : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => reqwrfail_s_DYMUX,
      CE => reqwrfail_s_CEINV,
      CLK => reqwrfail_s_CLKINV,
      SET => GND,
      RST => reqwrfail_s_FFY_RST,
      O => reqwrfail_s
    );
  reqwrfail_s_FFY_RSTOR : X_OR2
    port map (
      I0 => reqwrfail_s_FFY_RSTAND,
      I1 => GSR,
      O => reqwrfail_s_FFY_RST
    );
  reqwrfail_s_FFY_RSTAND_7782 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => reqwrfail_s_FFY_RSTAND
    );
  ix53675z3799 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => memswitchrd_s,
      ADR1 => ramdatao1_s(0),
      ADR2 => ramdatao2_s(0),
      ADR3 => VCC,
      O => ramdatao_s(0)
    );
  U_DCT2D_reg_latchbuf_reg_7_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_1_DYMUX,
      CE => U_DCT2D_latchbuf_reg_7_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_7_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_7_1_FFY_RST,
      O => U_DCT2D_latchbuf_reg_7_0_Q
    );
  U_DCT2D_latchbuf_reg_7_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_7_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_7_1_FFY_RST
    );
  ix53675z3794 : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => ramdatao2_s(4),
      ADR1 => ramdatao1_s(4),
      ADR2 => memswitchrd_s,
      ADR3 => VCC,
      O => ramdatao_s(4)
    );
  ix53675z3798 : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => ramdatao2_s(1),
      ADR1 => ramdatao1_s(1),
      ADR2 => memswitchrd_s,
      ADR3 => VCC,
      O => ramdatao_s(1)
    );
  ix53675z3797 : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => ramdatao1_s(2),
      ADR1 => VCC,
      ADR2 => memswitchrd_s,
      ADR3 => ramdatao2_s(2),
      O => ramdatao_s(2)
    );
  U_DCT2D_reg_latchbuf_reg_7_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_1_DXMUX,
      CE => U_DCT2D_latchbuf_reg_7_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_7_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_7_1_FFX_RST,
      O => U_DCT2D_latchbuf_reg_7_1_Q
    );
  U_DCT2D_latchbuf_reg_7_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_7_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_7_1_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_7_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_3_DYMUX,
      CE => U_DCT2D_latchbuf_reg_7_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_7_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_7_3_FFY_RST,
      O => U_DCT2D_latchbuf_reg_7_2_Q
    );
  U_DCT2D_latchbuf_reg_7_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_7_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_7_3_FFY_RST
    );
  ix53675z6053 : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => ramdatao2_s(3),
      ADR1 => VCC,
      ADR2 => memswitchrd_s,
      ADR3 => ramdatao1_s(3),
      O => ramdatao_s(3)
    );
  U_DCT2D_reg_latchbuf_reg_7_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_7_3_DXMUX,
      CE => U_DCT2D_latchbuf_reg_7_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_7_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_7_3_FFX_RST,
      O => U_DCT2D_latchbuf_reg_7_3_Q
    );
  U_DCT2D_latchbuf_reg_7_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_7_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_7_3_FFX_RST
    );
  U_DCT1D_modgen_counter_col_reg_reg_q_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_col_reg_0_DXMUX,
      CE => U_DCT1D_col_reg_0_CEINV,
      CLK => U_DCT1D_col_reg_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_col_reg_0_FFX_RST,
      O => U_DCT1D_col_reg(0)
    );
  U_DCT1D_col_reg_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_col_reg_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_col_reg_0_FFX_RST
    );
  U_DCT2D_ix8385z1324 : X_LUT4
    generic map(
      INIT => X"C3C3"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_2_10_Q,
      ADR2 => U_DCT2D_latchbuf_reg_5_10_Q,
      ADR3 => VCC,
      O => U_DCT2D_nx8385z1_F
    );
  U_DCT1D_reg_completed_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_completed_reg_DYMUX,
      CE => U_DCT1D_completed_reg_CEINV,
      CLK => U_DCT1D_completed_reg_CLKINV,
      SET => GND,
      RST => U_DCT1D_completed_reg_FFY_RST,
      O => U_DCT1D_completed_reg
    );
  U_DCT1D_completed_reg_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_completed_reg_FFY_RSTAND,
      I1 => GSR,
      O => U_DCT1D_completed_reg_FFY_RST
    );
  U_DCT1D_completed_reg_FFY_RSTAND_7783 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_completed_reg_FFY_RSTAND
    );
  U_DCT2D_ix7189z1324 : X_LUT4
    generic map(
      INIT => X"CC33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_7_10_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_0_10_Q,
      O => U_DCT2D_nx38337z1_G
    );
  U_DCT2D_ix38337z1321 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_latchbuf_reg_7_10_Q,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_0_10_Q,
      O => U_DCT2D_nx38337z1_F
    );
  U_DCT1D_ix2262z1321 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_5_Q(7),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_2_Q(7),
      ADR3 => VCC,
      O => U_DCT1D_nx47258z1_G
    );
  U_DCT1D_ix47258z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_5_Q(7),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_2_Q(7),
      ADR3 => VCC,
      O => U_DCT1D_nx47258z1_F
    );
  U_DCT1D_reg_state_reg_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_state_reg_1_DYMUX,
      CE => U_DCT1D_state_reg_1_CEINV,
      CLK => U_DCT1D_state_reg_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_state_reg_1_FFY_RST,
      O => U_DCT1D_state_reg(0)
    );
  U_DCT1D_state_reg_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_state_reg_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_state_reg_1_FFY_RST
    );
  U_DCT2D_ix43845z1329 : X_LUT4
    generic map(
      INIT => X"0302"
    )
    port map (
      ADR0 => requestrd_s,
      ADR1 => U_DCT2D_istate_reg(0),
      ADR2 => U_DCT2D_istate_reg(1),
      ADR3 => nx53675z1582,
      O => U_DCT2D_rtlc2n581_F
    );
  U_DCT1D_ix16101z1544 : X_LUT4
    generic map(
      INIT => X"FC3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_state_reg(1),
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_NOT_rtlcs7,
      O => U_DCT1D_rtlc5_state_reg_fsm_SS4_n374(1)
    );
  U_DCT1D_reg_state_reg_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_state_reg_1_DXMUX,
      CE => U_DCT1D_state_reg_1_CEINV,
      CLK => U_DCT1D_state_reg_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_state_reg_1_FFX_RST,
      O => U_DCT1D_state_reg(1)
    );
  U_DCT1D_state_reg_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_state_reg_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_state_reg_1_FFX_RST
    );
  U_DCT2D_ix64938z1324 : X_LUT4
    generic map(
      INIT => X"AA55"
    )
    port map (
      ADR0 => U_DCT2D_latchbuf_reg_6_10_Q,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_latchbuf_reg_1_10_Q,
      O => U_DCT2D_nx64938z1_F
    );
  U_DCT2D_ix6411z1331 : X_LUT4
    generic map(
      INIT => X"FFCC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => VCC,
      ADR3 => U_DCT2D_state_reg(1),
      O => U_DCT2D_rtlcs5_G
    );
  U_DCT2D_ix31471z1317 : X_LUT4
    generic map(
      INIT => X"3300"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => VCC,
      ADR3 => U_DCT2D_state_reg(1),
      O => U_DCT2D_rtlcs5_F
    );
  U_DCT2D_ix16172z1324 : X_LUT4
    generic map(
      INIT => X"F00F"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT2D_latchbuf_reg_4_10_Q,
      ADR3 => U_DCT2D_latchbuf_reg_3_10_Q,
      O => U_DCT2D_nx14976z1_G
    );
  U_DCT2D_ix6411z1483 : X_LUT4
    generic map(
      INIT => X"AAA0"
    )
    port map (
      ADR0 => U_DCT2D_istate_reg(1),
      ADR1 => VCC,
      ADR2 => U_DCT2D_istate_reg(0),
      ADR3 => U_DCT2D_nx6411z1,
      O => U_DCT2D_rtlc2n580_G
    );
  U_DCT1D_reg_latchbuf_reg_0_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_1_DYMUX,
      CE => U_DCT1D_latchbuf_reg_0_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_0_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_0_1_FFY_RST,
      O => U_DCT1D_latchbuf_reg_0_Q(0)
    );
  U_DCT1D_latchbuf_reg_0_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_0_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_0_1_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_0_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_1_DXMUX,
      CE => U_DCT1D_latchbuf_reg_0_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_0_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_0_1_FFX_RST,
      O => U_DCT1D_latchbuf_reg_0_Q(1)
    );
  U_DCT1D_latchbuf_reg_0_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_0_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_0_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_0_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_3_DYMUX,
      CE => U_DCT1D_latchbuf_reg_0_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_0_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_0_3_FFY_RST,
      O => U_DCT1D_latchbuf_reg_0_Q(2)
    );
  U_DCT1D_latchbuf_reg_0_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_0_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_0_3_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_0_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_3_DXMUX,
      CE => U_DCT1D_latchbuf_reg_0_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_0_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_0_3_FFX_RST,
      O => U_DCT1D_latchbuf_reg_0_Q(3)
    );
  U_DCT1D_latchbuf_reg_0_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_0_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_0_3_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_0_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_5_DYMUX,
      CE => U_DCT1D_latchbuf_reg_0_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_0_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_0_5_FFY_RST,
      O => U_DCT1D_latchbuf_reg_0_Q(4)
    );
  U_DCT1D_latchbuf_reg_0_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_0_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_0_5_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_0_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_5_DXMUX,
      CE => U_DCT1D_latchbuf_reg_0_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_0_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_0_5_FFX_RST,
      O => U_DCT1D_latchbuf_reg_0_Q(5)
    );
  U_DCT1D_latchbuf_reg_0_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_0_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_0_5_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_0_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_7_DYMUX,
      CE => U_DCT1D_latchbuf_reg_0_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_0_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_0_7_FFY_RST,
      O => U_DCT1D_latchbuf_reg_0_Q(6)
    );
  U_DCT1D_latchbuf_reg_0_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_0_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_0_7_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_0_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_0_7_DXMUX,
      CE => U_DCT1D_latchbuf_reg_0_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_0_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_0_7_FFX_RST,
      O => U_DCT1D_latchbuf_reg_0_Q(7)
    );
  U_DCT1D_latchbuf_reg_0_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_0_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_0_7_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_1_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_1_DYMUX,
      CE => U_DCT1D_latchbuf_reg_1_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_1_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_1_1_FFY_RST,
      O => U_DCT1D_latchbuf_reg_1_Q(0)
    );
  U_DCT1D_latchbuf_reg_1_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_1_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_1_1_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_1_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_1_DXMUX,
      CE => U_DCT1D_latchbuf_reg_1_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_1_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_1_1_FFX_RST,
      O => U_DCT1D_latchbuf_reg_1_Q(1)
    );
  U_DCT1D_latchbuf_reg_1_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_1_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_1_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_1_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_3_DYMUX,
      CE => U_DCT1D_latchbuf_reg_1_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_1_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_1_3_FFY_RST,
      O => U_DCT1D_latchbuf_reg_1_Q(2)
    );
  U_DCT1D_latchbuf_reg_1_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_1_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_1_3_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_1_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_3_DXMUX,
      CE => U_DCT1D_latchbuf_reg_1_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_1_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_1_3_FFX_RST,
      O => U_DCT1D_latchbuf_reg_1_Q(3)
    );
  U_DCT1D_latchbuf_reg_1_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_1_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_1_3_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_1_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_1_5_DYMUX,
      CE => U_DCT1D_latchbuf_reg_1_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_1_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_1_5_FFY_RST,
      O => U_DCT1D_latchbuf_reg_1_Q(4)
    );
  U_DCT1D_latchbuf_reg_1_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_1_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_1_5_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_2_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_7_DXMUX,
      CE => U_DCT1D_latchbuf_reg_2_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_2_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_2_7_FFX_RST,
      O => U_DCT1D_latchbuf_reg_2_Q(7)
    );
  U_DCT1D_latchbuf_reg_2_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_2_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_2_7_FFX_RST
    );
  U_DCT2D_reg_romoaddro0_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro0_s_3_DYMUX,
      CE => romo2addro0_s_3_CEINV,
      CLK => romo2addro0_s_3_CLKINV,
      SET => GND,
      RST => romo2addro0_s_3_FFY_RST,
      O => romo2addro0_s(2)
    );
  romo2addro0_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro0_s_3_SRINV,
      I1 => GSR,
      O => romo2addro0_s_3_FFY_RST
    );
  U_DCT2D_reg_romoaddro0_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro0_s_3_DXMUX,
      CE => romo2addro0_s_3_CEINV,
      CLK => romo2addro0_s_3_CLKINV,
      SET => GND,
      RST => romo2addro0_s_3_FFX_RST,
      O => romo2addro0_s(3)
    );
  romo2addro0_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro0_s_3_SRINV,
      I1 => GSR,
      O => romo2addro0_s_3_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_3_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_1_DYMUX,
      CE => U_DCT1D_latchbuf_reg_3_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_3_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_3_1_FFY_RST,
      O => U_DCT1D_latchbuf_reg_3_Q(0)
    );
  U_DCT1D_latchbuf_reg_3_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_3_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_3_1_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_3_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_1_DXMUX,
      CE => U_DCT1D_latchbuf_reg_3_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_3_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_3_1_FFX_RST,
      O => U_DCT1D_latchbuf_reg_3_Q(1)
    );
  U_DCT1D_latchbuf_reg_3_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_3_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_3_1_FFX_RST
    );
  U_DCT2D_reg_romoaddro1_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro1_s_1_DYMUX,
      CE => romo2addro1_s_1_CEINV,
      CLK => romo2addro1_s_1_CLKINV,
      SET => GND,
      RST => romo2addro1_s_1_FFY_RST,
      O => romo2addro1_s(0)
    );
  romo2addro1_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro1_s_1_SRINV,
      I1 => GSR,
      O => romo2addro1_s_1_FFY_RST
    );
  U_DCT2D_reg_romoaddro1_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro1_s_1_DXMUX,
      CE => romo2addro1_s_1_CEINV,
      CLK => romo2addro1_s_1_CLKINV,
      SET => GND,
      RST => romo2addro1_s_1_FFX_RST,
      O => romo2addro1_s(1)
    );
  romo2addro1_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro1_s_1_SRINV,
      I1 => GSR,
      O => romo2addro1_s_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_3_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_3_DYMUX,
      CE => U_DCT1D_latchbuf_reg_3_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_3_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_3_3_FFY_RST,
      O => U_DCT1D_latchbuf_reg_3_Q(2)
    );
  U_DCT1D_latchbuf_reg_3_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_3_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_3_3_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_3_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_3_DXMUX,
      CE => U_DCT1D_latchbuf_reg_3_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_3_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_3_3_FFX_RST,
      O => U_DCT1D_latchbuf_reg_3_Q(3)
    );
  U_DCT1D_latchbuf_reg_3_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_3_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_3_3_FFX_RST
    );
  U_DCT2D_reg_romoaddro1_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro1_s_3_DYMUX,
      CE => romo2addro1_s_3_CEINV,
      CLK => romo2addro1_s_3_CLKINV,
      SET => GND,
      RST => romo2addro1_s_3_FFY_RST,
      O => romo2addro1_s(2)
    );
  romo2addro1_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro1_s_3_SRINV,
      I1 => GSR,
      O => romo2addro1_s_3_FFY_RST
    );
  U_DCT2D_reg_romoaddro1_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro1_s_3_DXMUX,
      CE => romo2addro1_s_3_CEINV,
      CLK => romo2addro1_s_3_CLKINV,
      SET => GND,
      RST => romo2addro1_s_3_FFX_RST,
      O => romo2addro1_s(3)
    );
  romo2addro1_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro1_s_3_SRINV,
      I1 => GSR,
      O => romo2addro1_s_3_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_3_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_5_DYMUX,
      CE => U_DCT1D_latchbuf_reg_3_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_3_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_3_5_FFY_RST,
      O => U_DCT1D_latchbuf_reg_3_Q(4)
    );
  U_DCT1D_latchbuf_reg_3_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_3_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_3_5_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_3_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_5_DXMUX,
      CE => U_DCT1D_latchbuf_reg_3_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_3_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_3_5_FFX_RST,
      O => U_DCT1D_latchbuf_reg_3_Q(5)
    );
  U_DCT1D_latchbuf_reg_3_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_3_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_3_5_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_2_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_3_DXMUX,
      CE => U_DCT1D_latchbuf_reg_2_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_2_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_2_3_FFX_RST,
      O => U_DCT1D_latchbuf_reg_2_Q(3)
    );
  U_DCT1D_latchbuf_reg_2_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_2_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_2_3_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_2_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_5_DYMUX,
      CE => U_DCT1D_latchbuf_reg_2_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_2_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_2_5_FFY_RST,
      O => U_DCT1D_latchbuf_reg_2_Q(4)
    );
  U_DCT1D_latchbuf_reg_2_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_2_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_2_5_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_2_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_5_DXMUX,
      CE => U_DCT1D_latchbuf_reg_2_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_2_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_2_5_FFX_RST,
      O => U_DCT1D_latchbuf_reg_2_Q(5)
    );
  U_DCT1D_latchbuf_reg_2_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_2_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_2_5_FFX_RST
    );
  U_DCT2D_reg_romoaddro0_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro0_s_1_DYMUX,
      CE => romo2addro0_s_1_CEINV,
      CLK => romo2addro0_s_1_CLKINV,
      SET => GND,
      RST => romo2addro0_s_1_FFY_RST,
      O => romo2addro0_s(0)
    );
  romo2addro0_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro0_s_1_SRINV,
      I1 => GSR,
      O => romo2addro0_s_1_FFY_RST
    );
  U_DCT2D_reg_romoaddro0_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro0_s_1_DXMUX,
      CE => romo2addro0_s_1_CEINV,
      CLK => romo2addro0_s_1_CLKINV,
      SET => GND,
      RST => romo2addro0_s_1_FFX_RST,
      O => romo2addro0_s(1)
    );
  romo2addro0_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro0_s_1_SRINV,
      I1 => GSR,
      O => romo2addro0_s_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_2_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_2_7_DYMUX,
      CE => U_DCT1D_latchbuf_reg_2_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_2_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_2_7_FFY_RST,
      O => U_DCT1D_latchbuf_reg_2_Q(6)
    );
  U_DCT1D_latchbuf_reg_2_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_2_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_2_7_FFY_RST
    );
  U_DCT2D_reg_romoaddro8_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro8_s_1_DXMUX,
      CE => romo2addro8_s_1_CEINV,
      CLK => romo2addro8_s_1_CLKINV,
      SET => GND,
      RST => romo2addro8_s_1_FFX_RST,
      O => romo2addro8_s(1)
    );
  romo2addro8_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro8_s_1_SRINV,
      I1 => GSR,
      O => romo2addro8_s_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_6_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_7_DYMUX,
      CE => U_DCT1D_latchbuf_reg_6_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_6_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_6_7_FFY_RST,
      O => U_DCT1D_latchbuf_reg_6_Q(6)
    );
  U_DCT1D_latchbuf_reg_6_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_6_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_6_7_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_6_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_7_DXMUX,
      CE => U_DCT1D_latchbuf_reg_6_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_6_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_6_7_FFX_RST,
      O => U_DCT1D_latchbuf_reg_6_Q(7)
    );
  U_DCT1D_latchbuf_reg_6_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_6_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_6_7_FFX_RST
    );
  U_DCT2D_reg_romoaddro8_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro8_s_3_DYMUX,
      CE => romo2addro8_s_3_CEINV,
      CLK => romo2addro8_s_3_CLKINV,
      SET => GND,
      RST => romo2addro8_s_3_FFY_RST,
      O => romo2addro8_s(2)
    );
  romo2addro8_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro8_s_3_SRINV,
      I1 => GSR,
      O => romo2addro8_s_3_FFY_RST
    );
  U_DCT2D_reg_romoaddro8_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro8_s_3_DXMUX,
      CE => romo2addro8_s_3_CEINV,
      CLK => romo2addro8_s_3_CLKINV,
      SET => GND,
      RST => romo2addro8_s_3_FFX_RST,
      O => romo2addro8_s(3)
    );
  romo2addro8_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro8_s_3_SRINV,
      I1 => GSR,
      O => romo2addro8_s_3_FFX_RST
    );
  U_DCT2D_reg_romoaddro9_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro9_s_1_DYMUX,
      CE => romo2addro9_s_1_CEINV,
      CLK => romo2addro9_s_1_CLKINV,
      SET => GND,
      RST => romo2addro9_s_1_FFY_RST,
      O => romo2addro9_s(0)
    );
  romo2addro9_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro9_s_1_SRINV,
      I1 => GSR,
      O => romo2addro9_s_1_FFY_RST
    );
  U_DCT2D_reg_romoaddro2_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro2_s_1_DYMUX,
      CE => romo2addro2_s_1_CEINV,
      CLK => romo2addro2_s_1_CLKINV,
      SET => GND,
      RST => romo2addro2_s_1_FFY_RST,
      O => romo2addro2_s(0)
    );
  romo2addro2_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro2_s_1_SRINV,
      I1 => GSR,
      O => romo2addro2_s_1_FFY_RST
    );
  U_DCT2D_reg_romoaddro2_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro2_s_1_DXMUX,
      CE => romo2addro2_s_1_CEINV,
      CLK => romo2addro2_s_1_CLKINV,
      SET => GND,
      RST => romo2addro2_s_1_FFX_RST,
      O => romo2addro2_s(1)
    );
  romo2addro2_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro2_s_1_SRINV,
      I1 => GSR,
      O => romo2addro2_s_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_3_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_7_DYMUX,
      CE => U_DCT1D_latchbuf_reg_3_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_3_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_3_7_FFY_RST,
      O => U_DCT1D_latchbuf_reg_3_Q(6)
    );
  U_DCT1D_latchbuf_reg_3_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_3_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_3_7_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_3_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_3_7_DXMUX,
      CE => U_DCT1D_latchbuf_reg_3_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_3_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_3_7_FFX_RST,
      O => U_DCT1D_latchbuf_reg_3_Q(7)
    );
  U_DCT1D_latchbuf_reg_3_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_3_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_3_7_FFX_RST
    );
  U_DCT2D_reg_romoaddro2_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro2_s_3_DYMUX,
      CE => romo2addro2_s_3_CEINV,
      CLK => romo2addro2_s_3_CLKINV,
      SET => GND,
      RST => romo2addro2_s_3_FFY_RST,
      O => romo2addro2_s(2)
    );
  romo2addro2_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro2_s_3_SRINV,
      I1 => GSR,
      O => romo2addro2_s_3_FFY_RST
    );
  U_DCT2D_reg_romoaddro2_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro2_s_3_DXMUX,
      CE => romo2addro2_s_3_CEINV,
      CLK => romo2addro2_s_3_CLKINV,
      SET => GND,
      RST => romo2addro2_s_3_FFX_RST,
      O => romo2addro2_s(3)
    );
  romo2addro2_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro2_s_3_SRINV,
      I1 => GSR,
      O => romo2addro2_s_3_FFX_RST
    );
  U_DCT2D_reg_romoaddro3_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro3_s_3_DYMUX,
      CE => romo2addro3_s_3_CEINV,
      CLK => romo2addro3_s_3_CLKINV,
      SET => GND,
      RST => romo2addro3_s_3_FFY_RST,
      O => romo2addro3_s(2)
    );
  romo2addro3_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro3_s_3_SRINV,
      I1 => GSR,
      O => romo2addro3_s_3_FFY_RST
    );
  U_DCT2D_reg_romoaddro3_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro3_s_3_DXMUX,
      CE => romo2addro3_s_3_CEINV,
      CLK => romo2addro3_s_3_CLKINV,
      SET => GND,
      RST => romo2addro3_s_3_FFX_RST,
      O => romo2addro3_s(3)
    );
  romo2addro3_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro3_s_3_SRINV,
      I1 => GSR,
      O => romo2addro3_s_3_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_4_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_5_DYMUX,
      CE => U_DCT1D_latchbuf_reg_4_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_4_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_4_5_FFY_RST,
      O => U_DCT1D_latchbuf_reg_4_Q(4)
    );
  U_DCT1D_latchbuf_reg_4_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_4_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_4_5_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_4_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_5_DXMUX,
      CE => U_DCT1D_latchbuf_reg_4_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_4_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_4_5_FFX_RST,
      O => U_DCT1D_latchbuf_reg_4_Q(5)
    );
  U_DCT1D_latchbuf_reg_4_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_4_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_4_5_FFX_RST
    );
  U_DCT2D_reg_romoaddro4_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro4_s_1_DYMUX,
      CE => romo2addro4_s_1_CEINV,
      CLK => romo2addro4_s_1_CLKINV,
      SET => GND,
      RST => romo2addro4_s_1_FFY_RST,
      O => romo2addro4_s(0)
    );
  romo2addro4_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro4_s_1_SRINV,
      I1 => GSR,
      O => romo2addro4_s_1_FFY_RST
    );
  U_DCT2D_reg_romoaddro4_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro4_s_1_DXMUX,
      CE => romo2addro4_s_1_CEINV,
      CLK => romo2addro4_s_1_CLKINV,
      SET => GND,
      RST => romo2addro4_s_1_FFX_RST,
      O => romo2addro4_s(1)
    );
  romo2addro4_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro4_s_1_SRINV,
      I1 => GSR,
      O => romo2addro4_s_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_5_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_5_DXMUX,
      CE => U_DCT1D_latchbuf_reg_5_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_5_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_5_5_FFX_RST,
      O => U_DCT1D_latchbuf_reg_5_Q(5)
    );
  U_DCT1D_latchbuf_reg_5_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_5_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_5_5_FFX_RST
    );
  U_DCT2D_reg_romoaddro6_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro6_s_1_DYMUX,
      CE => romo2addro6_s_1_CEINV,
      CLK => romo2addro6_s_1_CLKINV,
      SET => GND,
      RST => romo2addro6_s_1_FFY_RST,
      O => romo2addro6_s(0)
    );
  romo2addro6_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro6_s_1_SRINV,
      I1 => GSR,
      O => romo2addro6_s_1_FFY_RST
    );
  U_DCT2D_reg_romoaddro6_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro6_s_1_DXMUX,
      CE => romo2addro6_s_1_CEINV,
      CLK => romo2addro6_s_1_CLKINV,
      SET => GND,
      RST => romo2addro6_s_1_FFX_RST,
      O => romo2addro6_s(1)
    );
  romo2addro6_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro6_s_1_SRINV,
      I1 => GSR,
      O => romo2addro6_s_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_5_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_7_DYMUX,
      CE => U_DCT1D_latchbuf_reg_5_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_5_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_5_7_FFY_RST,
      O => U_DCT1D_latchbuf_reg_5_Q(6)
    );
  U_DCT1D_latchbuf_reg_5_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_5_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_5_7_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_5_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_7_DXMUX,
      CE => U_DCT1D_latchbuf_reg_5_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_5_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_5_7_FFX_RST,
      O => U_DCT1D_latchbuf_reg_5_Q(7)
    );
  U_DCT1D_latchbuf_reg_5_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_5_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_5_7_FFX_RST
    );
  U_DCT2D_reg_romoaddro6_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro6_s_3_DYMUX,
      CE => romo2addro6_s_3_CEINV,
      CLK => romo2addro6_s_3_CLKINV,
      SET => GND,
      RST => romo2addro6_s_3_FFY_RST,
      O => romo2addro6_s(2)
    );
  romo2addro6_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro6_s_3_SRINV,
      I1 => GSR,
      O => romo2addro6_s_3_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_4_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_7_DYMUX,
      CE => U_DCT1D_latchbuf_reg_4_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_4_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_4_7_FFY_RST,
      O => U_DCT1D_latchbuf_reg_4_Q(6)
    );
  U_DCT1D_latchbuf_reg_4_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_4_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_4_7_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_4_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_4_7_DXMUX,
      CE => U_DCT1D_latchbuf_reg_4_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_4_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_4_7_FFX_RST,
      O => U_DCT1D_latchbuf_reg_4_Q(7)
    );
  U_DCT1D_latchbuf_reg_4_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_4_7_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_4_7_FFX_RST
    );
  U_DCT2D_reg_romoaddro4_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro4_s_3_DYMUX,
      CE => romo2addro4_s_3_CEINV,
      CLK => romo2addro4_s_3_CLKINV,
      SET => GND,
      RST => romo2addro4_s_3_FFY_RST,
      O => romo2addro4_s(2)
    );
  romo2addro4_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro4_s_3_SRINV,
      I1 => GSR,
      O => romo2addro4_s_3_FFY_RST
    );
  U_DCT2D_reg_romoaddro4_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro4_s_3_DXMUX,
      CE => romo2addro4_s_3_CEINV,
      CLK => romo2addro4_s_3_CLKINV,
      SET => GND,
      RST => romo2addro4_s_3_FFX_RST,
      O => romo2addro4_s(3)
    );
  romo2addro4_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro4_s_3_SRINV,
      I1 => GSR,
      O => romo2addro4_s_3_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_5_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_1_DYMUX,
      CE => U_DCT1D_latchbuf_reg_5_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_5_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_5_1_FFY_RST,
      O => U_DCT1D_latchbuf_reg_5_Q(0)
    );
  U_DCT1D_latchbuf_reg_5_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_5_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_5_1_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_5_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_5_1_DXMUX,
      CE => U_DCT1D_latchbuf_reg_5_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_5_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_5_1_FFX_RST,
      O => U_DCT1D_latchbuf_reg_5_Q(1)
    );
  U_DCT1D_latchbuf_reg_5_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_5_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_5_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_6_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_3_DXMUX,
      CE => U_DCT1D_latchbuf_reg_6_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_6_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_6_3_FFX_RST,
      O => U_DCT1D_latchbuf_reg_6_Q(3)
    );
  U_DCT1D_latchbuf_reg_6_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_6_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_6_3_FFX_RST
    );
  U_DCT2D_reg_romoaddro7_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro7_s_3_DYMUX,
      CE => romo2addro7_s_3_CEINV,
      CLK => romo2addro7_s_3_CLKINV,
      SET => GND,
      RST => romo2addro7_s_3_FFY_RST,
      O => romo2addro7_s(2)
    );
  romo2addro7_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro7_s_3_SRINV,
      I1 => GSR,
      O => romo2addro7_s_3_FFY_RST
    );
  U_DCT2D_reg_romoaddro7_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro7_s_3_DXMUX,
      CE => romo2addro7_s_3_CEINV,
      CLK => romo2addro7_s_3_CLKINV,
      SET => GND,
      RST => romo2addro7_s_3_FFX_RST,
      O => romo2addro7_s(3)
    );
  romo2addro7_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro7_s_3_SRINV,
      I1 => GSR,
      O => romo2addro7_s_3_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_6_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_5_DYMUX,
      CE => U_DCT1D_latchbuf_reg_6_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_6_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_6_5_FFY_RST,
      O => U_DCT1D_latchbuf_reg_6_Q(4)
    );
  U_DCT1D_latchbuf_reg_6_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_6_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_6_5_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_6_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_5_DXMUX,
      CE => U_DCT1D_latchbuf_reg_6_5_CEINV,
      CLK => U_DCT1D_latchbuf_reg_6_5_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_6_5_FFX_RST,
      O => U_DCT1D_latchbuf_reg_6_Q(5)
    );
  U_DCT1D_latchbuf_reg_6_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_6_5_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_6_5_FFX_RST
    );
  U_DCT2D_reg_romoaddro8_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro8_s_1_DYMUX,
      CE => romo2addro8_s_1_CEINV,
      CLK => romo2addro8_s_1_CLKINV,
      SET => GND,
      RST => romo2addro8_s_1_FFY_RST,
      O => romo2addro8_s(0)
    );
  romo2addro8_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro8_s_1_SRINV,
      I1 => GSR,
      O => romo2addro8_s_1_FFY_RST
    );
  U_DCT2D_reg_romoaddro9_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro9_s_1_DXMUX,
      CE => romo2addro9_s_1_CEINV,
      CLK => romo2addro9_s_1_CLKINV,
      SET => GND,
      RST => romo2addro9_s_1_FFX_RST,
      O => romo2addro9_s(1)
    );
  romo2addro9_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro9_s_1_SRINV,
      I1 => GSR,
      O => romo2addro9_s_1_FFX_RST
    );
  U_DCT2D_reg_romoaddro9_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro9_s_3_DYMUX,
      CE => romo2addro9_s_3_CEINV,
      CLK => romo2addro9_s_3_CLKINV,
      SET => GND,
      RST => romo2addro9_s_3_FFY_RST,
      O => romo2addro9_s(2)
    );
  romo2addro9_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro9_s_3_SRINV,
      I1 => GSR,
      O => romo2addro9_s_3_FFY_RST
    );
  U_DCT2D_reg_romoaddro9_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro9_s_3_DXMUX,
      CE => romo2addro9_s_3_CEINV,
      CLK => romo2addro9_s_3_CLKINV,
      SET => GND,
      RST => romo2addro9_s_3_FFX_RST,
      O => romo2addro9_s(3)
    );
  romo2addro9_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro9_s_3_SRINV,
      I1 => GSR,
      O => romo2addro9_s_3_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_7_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_7_7_DYMUX,
      CE => U_DCT1D_latchbuf_reg_7_7_CEINV,
      CLK => U_DCT1D_latchbuf_reg_7_7_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_7_7_FFY_RST,
      O => U_DCT1D_latchbuf_reg_7_Q(7)
    );
  U_DCT1D_latchbuf_reg_7_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_7_7_FFY_RSTAND,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_7_7_FFY_RST
    );
  U_DCT1D_latchbuf_reg_7_7_FFY_RSTAND_7784 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latchbuf_reg_7_7_FFY_RSTAND
    );
  U_DCT2D_ix7599z3405 : X_LUT4
    generic map(
      INIT => X"1D00"
    )
    port map (
      ADR0 => U_DCT2D_NOT_rtlcs2,
      ADR1 => U_DCT2D_istate_reg(0),
      ADR2 => U_DCT2D_rtlcn65,
      ADR3 => U_DCT2D_istate_reg(1),
      O => U_DCT2D_rtlc2n579_G
    );
  U_DCT2D_reg_latch_done_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latch_done_reg_DYMUX,
      CE => U_DCT2D_latch_done_reg_CEINV,
      CLK => U_DCT2D_latch_done_reg_CLKINV,
      SET => GND,
      RST => U_DCT2D_latch_done_reg_FFY_RST,
      O => U_DCT2D_latch_done_reg
    );
  U_DCT2D_latch_done_reg_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latch_done_reg_FFY_RSTAND,
      I1 => GSR,
      O => U_DCT2D_latch_done_reg_FFY_RST
    );
  U_DCT2D_latch_done_reg_FFY_RSTAND_7785 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_latch_done_reg_FFY_RSTAND
    );
  U_DCT2D_ix41892z1059 : X_LUT4
    generic map(
      INIT => X"FEFF"
    )
    port map (
      ADR0 => ramraddro_s(2),
      ADR1 => ramraddro_s(1),
      ADR2 => ramraddro_s(0),
      ADR3 => U_DCT2D_colram_reg(3),
      O => U_DCT2D_nx6411z1_G
    );
  U_DCT2D_ix41892z1324 : X_LUT4
    generic map(
      INIT => X"55FF"
    )
    port map (
      ADR0 => ramraddro_s(0),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => ramraddro_s(1),
      O => U_DCT2D_nx41892z2_G
    );
  U_DCT2D_ix6411z1444 : X_LUT4
    generic map(
      INIT => X"0800"
    )
    port map (
      ADR0 => ramraddro_s(5),
      ADR1 => ramraddro_s(3),
      ADR2 => U_DCT2D_NOT_rtlcs2,
      ADR3 => ramraddro_s(4),
      O => U_DCT2D_nx6411z1_F
    );
  U_DCT1D_reg_romeaddro6_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro6_s_3_DXMUX,
      CE => romeaddro6_s_3_CEINV,
      CLK => romeaddro6_s_3_CLKINV,
      SET => GND,
      RST => romeaddro6_s_3_FFX_RST,
      O => romeaddro6_s(3)
    );
  romeaddro6_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro6_s_3_SRINV,
      I1 => GSR,
      O => romeaddro6_s_3_FFX_RST
    );
  U_DCT2D_reg_romoaddro10_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro0_s_5_DYMUX,
      CE => romo2addro0_s_5_CEINV,
      CLK => romo2addro0_s_5_CLKINV,
      SET => GND,
      RST => romo2addro0_s_5_FFY_RST,
      O => romo2addro0_s(4)
    );
  romo2addro0_s_5_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro0_s_5_SRINV,
      I1 => GSR,
      O => romo2addro0_s_5_FFY_RST
    );
  U_DCT2D_reg_romoaddro10_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro0_s_5_DXMUX,
      CE => romo2addro0_s_5_CEINV,
      CLK => romo2addro0_s_5_CLKINV,
      SET => GND,
      RST => romo2addro0_s_5_FFX_RST,
      O => romo2addro0_s(5)
    );
  romo2addro0_s_5_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro0_s_5_SRINV,
      I1 => GSR,
      O => romo2addro0_s_5_FFX_RST
    );
  U_DCT1D_reg_romeaddro7_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro7_s_1_DYMUX,
      CE => romeaddro7_s_1_CEINV,
      CLK => romeaddro7_s_1_CLKINV,
      SET => GND,
      RST => romeaddro7_s_1_FFY_RST,
      O => romeaddro7_s(0)
    );
  romeaddro7_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro7_s_1_SRINV,
      I1 => GSR,
      O => romeaddro7_s_1_FFY_RST
    );
  U_DCT1D_reg_romeaddro7_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro7_s_1_DXMUX,
      CE => romeaddro7_s_1_CEINV,
      CLK => romeaddro7_s_1_CLKINV,
      SET => GND,
      RST => romeaddro7_s_1_FFX_RST,
      O => romeaddro7_s(1)
    );
  romeaddro7_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro7_s_1_SRINV,
      I1 => GSR,
      O => romeaddro7_s_1_FFX_RST
    );
  U_DCT1D_reg_romeaddro7_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro7_s_3_DYMUX,
      CE => romeaddro7_s_3_CEINV,
      CLK => romeaddro7_s_3_CLKINV,
      SET => GND,
      RST => romeaddro7_s_3_FFY_RST,
      O => romeaddro7_s(2)
    );
  romeaddro7_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro7_s_3_SRINV,
      I1 => GSR,
      O => romeaddro7_s_3_FFY_RST
    );
  U_DCT1D_reg_romeaddro7_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro7_s_3_DXMUX,
      CE => romeaddro7_s_3_CEINV,
      CLK => romeaddro7_s_3_CLKINV,
      SET => GND,
      RST => romeaddro7_s_3_FFX_RST,
      O => romeaddro7_s(3)
    );
  romeaddro7_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro7_s_3_SRINV,
      I1 => GSR,
      O => romeaddro7_s_3_FFX_RST
    );
  U_DCT1D_reg_romoaddro1_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro1_s_3_DXMUX,
      CE => romoaddro1_s_3_CEINV,
      CLK => romoaddro1_s_3_CLKINV,
      SET => GND,
      RST => romoaddro1_s_3_FFX_RST,
      O => romoaddro1_s(3)
    );
  romoaddro1_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro1_s_3_SRINV,
      I1 => GSR,
      O => romoaddro1_s_3_FFX_RST
    );
  U_DCT1D_reg_romoaddro2_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro2_s_1_DYMUX,
      CE => romoaddro2_s_1_CEINV,
      CLK => romoaddro2_s_1_CLKINV,
      SET => GND,
      RST => romoaddro2_s_1_FFY_RST,
      O => romoaddro2_s(0)
    );
  romoaddro2_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro2_s_1_SRINV,
      I1 => GSR,
      O => romoaddro2_s_1_FFY_RST
    );
  U_DCT1D_reg_romoaddro2_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro2_s_1_DXMUX,
      CE => romoaddro2_s_1_CEINV,
      CLK => romoaddro2_s_1_CLKINV,
      SET => GND,
      RST => romoaddro2_s_1_FFX_RST,
      O => romoaddro2_s(1)
    );
  romoaddro2_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro2_s_1_SRINV,
      I1 => GSR,
      O => romoaddro2_s_1_FFX_RST
    );
  U_DCT1D_reg_romoaddro2_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro2_s_3_DYMUX,
      CE => romoaddro2_s_3_CEINV,
      CLK => romoaddro2_s_3_CLKINV,
      SET => GND,
      RST => romoaddro2_s_3_FFY_RST,
      O => romoaddro2_s(2)
    );
  romoaddro2_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro2_s_3_SRINV,
      I1 => GSR,
      O => romoaddro2_s_3_FFY_RST
    );
  U_DCT1D_reg_romoaddro2_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro2_s_3_DXMUX,
      CE => romoaddro2_s_3_CEINV,
      CLK => romoaddro2_s_3_CLKINV,
      SET => GND,
      RST => romoaddro2_s_3_FFX_RST,
      O => romoaddro2_s(3)
    );
  romoaddro2_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro2_s_3_SRINV,
      I1 => GSR,
      O => romoaddro2_s_3_FFX_RST
    );
  U_DCT1D_reg_romoaddro3_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro3_s_1_DYMUX,
      CE => romoaddro3_s_1_CEINV,
      CLK => romoaddro3_s_1_CLKINV,
      SET => GND,
      RST => romoaddro3_s_1_FFY_RST,
      O => romoaddro3_s(0)
    );
  romoaddro3_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro3_s_1_SRINV,
      I1 => GSR,
      O => romoaddro3_s_1_FFY_RST
    );
  U_DCT1D_reg_romoaddro3_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro3_s_1_DXMUX,
      CE => romoaddro3_s_1_CEINV,
      CLK => romoaddro3_s_1_CLKINV,
      SET => GND,
      RST => romoaddro3_s_1_FFX_RST,
      O => romoaddro3_s(1)
    );
  romoaddro3_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro3_s_1_SRINV,
      I1 => GSR,
      O => romoaddro3_s_1_FFX_RST
    );
  U_DCT2D_reg_romoaddro6_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro6_s_3_DXMUX,
      CE => romo2addro6_s_3_CEINV,
      CLK => romo2addro6_s_3_CLKINV,
      SET => GND,
      RST => romo2addro6_s_3_FFX_RST,
      O => romo2addro6_s(3)
    );
  romo2addro6_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro6_s_3_SRINV,
      I1 => GSR,
      O => romo2addro6_s_3_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_6_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_1_DYMUX,
      CE => U_DCT1D_latchbuf_reg_6_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_6_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_6_1_FFY_RST,
      O => U_DCT1D_latchbuf_reg_6_Q(0)
    );
  U_DCT1D_latchbuf_reg_6_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_6_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_6_1_FFY_RST
    );
  U_DCT1D_reg_latchbuf_reg_6_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_1_DXMUX,
      CE => U_DCT1D_latchbuf_reg_6_1_CEINV,
      CLK => U_DCT1D_latchbuf_reg_6_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_6_1_FFX_RST,
      O => U_DCT1D_latchbuf_reg_6_Q(1)
    );
  U_DCT1D_latchbuf_reg_6_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_6_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_6_1_FFX_RST
    );
  U_DCT2D_reg_romoaddro7_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro7_s_1_DYMUX,
      CE => romo2addro7_s_1_CEINV,
      CLK => romo2addro7_s_1_CLKINV,
      SET => GND,
      RST => romo2addro7_s_1_FFY_RST,
      O => romo2addro7_s(0)
    );
  romo2addro7_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro7_s_1_SRINV,
      I1 => GSR,
      O => romo2addro7_s_1_FFY_RST
    );
  U_DCT2D_reg_romoaddro7_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro7_s_1_DXMUX,
      CE => romo2addro7_s_1_CEINV,
      CLK => romo2addro7_s_1_CLKINV,
      SET => GND,
      RST => romo2addro7_s_1_FFX_RST,
      O => romo2addro7_s(1)
    );
  romo2addro7_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro7_s_1_SRINV,
      I1 => GSR,
      O => romo2addro7_s_1_FFX_RST
    );
  U_DCT1D_reg_latchbuf_reg_6_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latchbuf_reg_6_3_DYMUX,
      CE => U_DCT1D_latchbuf_reg_6_3_CEINV,
      CLK => U_DCT1D_latchbuf_reg_6_3_CLKINV,
      SET => GND,
      RST => U_DCT1D_latchbuf_reg_6_3_FFY_RST,
      O => U_DCT1D_latchbuf_reg_6_Q(2)
    );
  U_DCT1D_latchbuf_reg_6_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latchbuf_reg_6_3_SRINV,
      I1 => GSR,
      O => U_DCT1D_latchbuf_reg_6_3_FFY_RST
    );
  U_DCT1D_reg_romeaddro3_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro3_s_1_DXMUX,
      CE => romeaddro3_s_1_CEINV,
      CLK => romeaddro3_s_1_CLKINV,
      SET => GND,
      RST => romeaddro3_s_1_FFX_RST,
      O => romeaddro3_s(1)
    );
  romeaddro3_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro3_s_1_SRINV,
      I1 => GSR,
      O => romeaddro3_s_1_FFX_RST
    );
  U_DCT1D_reg_romeaddro3_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro3_s_3_DYMUX,
      CE => romeaddro3_s_3_CEINV,
      CLK => romeaddro3_s_3_CLKINV,
      SET => GND,
      RST => romeaddro3_s_3_FFY_RST,
      O => romeaddro3_s(2)
    );
  romeaddro3_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro3_s_3_SRINV,
      I1 => GSR,
      O => romeaddro3_s_3_FFY_RST
    );
  U_DCT1D_reg_romeaddro3_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro3_s_3_DXMUX,
      CE => romeaddro3_s_3_CEINV,
      CLK => romeaddro3_s_3_CLKINV,
      SET => GND,
      RST => romeaddro3_s_3_FFX_RST,
      O => romeaddro3_s(3)
    );
  romeaddro3_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro3_s_3_SRINV,
      I1 => GSR,
      O => romeaddro3_s_3_FFX_RST
    );
  U_DCT1D_reg_romeaddro4_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro4_s_1_DYMUX,
      CE => romeaddro4_s_1_CEINV,
      CLK => romeaddro4_s_1_CLKINV,
      SET => GND,
      RST => romeaddro4_s_1_FFY_RST,
      O => romeaddro4_s(0)
    );
  romeaddro4_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro4_s_1_SRINV,
      I1 => GSR,
      O => romeaddro4_s_1_FFY_RST
    );
  U_DCT1D_reg_romeaddro4_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro4_s_1_DXMUX,
      CE => romeaddro4_s_1_CEINV,
      CLK => romeaddro4_s_1_CLKINV,
      SET => GND,
      RST => romeaddro4_s_1_FFX_RST,
      O => romeaddro4_s(1)
    );
  romeaddro4_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro4_s_1_SRINV,
      I1 => GSR,
      O => romeaddro4_s_1_FFX_RST
    );
  U_DCT1D_reg_romeaddro4_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro4_s_3_DYMUX,
      CE => romeaddro4_s_3_CEINV,
      CLK => romeaddro4_s_3_CLKINV,
      SET => GND,
      RST => romeaddro4_s_3_FFY_RST,
      O => romeaddro4_s(2)
    );
  romeaddro4_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro4_s_3_SRINV,
      I1 => GSR,
      O => romeaddro4_s_3_FFY_RST
    );
  U_DCT2D_ix41892z13779 : X_LUT4
    generic map(
      INIT => X"0A8A"
    )
    port map (
      ADR0 => U_DCT2D_NOT_rtlc2n488,
      ADR1 => ramraddro_s(2),
      ADR2 => U_DCT2D_NOT_rtlcs2,
      ADR3 => U_DCT2D_nx41892z3,
      O => U_DCT2D_nx41892z2_F
    );
  U_DCT1D_ix52040z1320 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_row_reg(0),
      ADR1 => U_DCT1D_row_reg(1),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx52040z1
    );
  U_DCT1D_modgen_counter_row_reg_reg_q_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_row_reg_0_DYMUX,
      CE => U_DCT1D_row_reg_0_CEINV,
      CLK => U_DCT1D_row_reg_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_row_reg_0_FFY_RST,
      O => U_DCT1D_row_reg(1)
    );
  U_DCT1D_row_reg_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_row_reg_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_row_reg_0_FFY_RST
    );
  U_DCT1D_modgen_counter_row_reg_reg_q_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_row_reg_0_DXMUX,
      CE => U_DCT1D_row_reg_0_CEINV,
      CLK => U_DCT1D_row_reg_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_row_reg_0_FFX_RST,
      O => U_DCT1D_row_reg(0)
    );
  U_DCT1D_row_reg_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_row_reg_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_row_reg_0_FFX_RST
    );
  U_DCT2D_ix16101z1442 : X_LUT4
    generic map(
      INIT => X"5FFF"
    )
    port map (
      ADR0 => U_DCT2D_col_reg(2),
      ADR1 => VCC,
      ADR2 => U_DCT2D_col_reg(0),
      ADR3 => U_DCT2D_col_reg(1),
      O => U_DCT2D_state_reg_1_G
    );
  U_DCT2D_reg_state_reg_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_state_reg_1_DYMUX,
      CE => U_DCT2D_state_reg_1_CEINV,
      CLK => U_DCT2D_state_reg_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_state_reg_1_FFY_RST,
      O => U_DCT2D_state_reg(0)
    );
  U_DCT2D_state_reg_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_state_reg_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_state_reg_1_FFY_RST
    );
  U_DCT2D_ix16101z1544 : X_LUT4
    generic map(
      INIT => X"EE66"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_state_reg(1),
      ADR2 => VCC,
      ADR3 => U_DCT2D_NOT_rtlcs7,
      O => U_DCT2D_rtlc5_state_reg_fsm_SS3_n367(1)
    );
  U_DCT2D_reg_romeaddro4_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro4_s_1_DYMUX,
      CE => rome2addro4_s_1_CEINV,
      CLK => rome2addro4_s_1_CLKINV,
      SET => GND,
      RST => rome2addro4_s_1_FFY_RST,
      O => rome2addro4_s(0)
    );
  rome2addro4_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro4_s_1_SRINV,
      I1 => GSR,
      O => rome2addro4_s_1_FFY_RST
    );
  U_DCT2D_reg_romeaddro4_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro4_s_1_DXMUX,
      CE => rome2addro4_s_1_CEINV,
      CLK => rome2addro4_s_1_CLKINV,
      SET => GND,
      RST => rome2addro4_s_1_FFX_RST,
      O => rome2addro4_s(1)
    );
  rome2addro4_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro4_s_1_SRINV,
      I1 => GSR,
      O => rome2addro4_s_1_FFX_RST
    );
  U_DCT2D_reg_romeaddro4_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro4_s_3_DYMUX,
      CE => rome2addro4_s_3_CEINV,
      CLK => rome2addro4_s_3_CLKINV,
      SET => GND,
      RST => rome2addro4_s_3_FFY_RST,
      O => rome2addro4_s(2)
    );
  rome2addro4_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro4_s_3_SRINV,
      I1 => GSR,
      O => rome2addro4_s_3_FFY_RST
    );
  U_DCT2D_reg_romeaddro4_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro4_s_3_DXMUX,
      CE => rome2addro4_s_3_CEINV,
      CLK => rome2addro4_s_3_CLKINV,
      SET => GND,
      RST => rome2addro4_s_3_FFX_RST,
      O => rome2addro4_s(3)
    );
  rome2addro4_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro4_s_3_SRINV,
      I1 => GSR,
      O => rome2addro4_s_3_FFX_RST
    );
  U_DCT2D_reg_romeaddro5_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro5_s_1_DYMUX,
      CE => rome2addro5_s_1_CEINV,
      CLK => rome2addro5_s_1_CLKINV,
      SET => GND,
      RST => rome2addro5_s_1_FFY_RST,
      O => rome2addro5_s(0)
    );
  rome2addro5_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro5_s_1_SRINV,
      I1 => GSR,
      O => rome2addro5_s_1_FFY_RST
    );
  U_DCT2D_reg_romeaddro5_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro5_s_1_DXMUX,
      CE => rome2addro5_s_1_CEINV,
      CLK => rome2addro5_s_1_CLKINV,
      SET => GND,
      RST => rome2addro5_s_1_FFX_RST,
      O => rome2addro5_s(1)
    );
  rome2addro5_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro5_s_1_SRINV,
      I1 => GSR,
      O => rome2addro5_s_1_FFX_RST
    );
  U_DCT1D_reg_romeaddro8_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro8_s_1_DYMUX,
      CE => romeaddro8_s_1_CEINV,
      CLK => romeaddro8_s_1_CLKINV,
      SET => GND,
      RST => romeaddro8_s_1_FFY_RST,
      O => romeaddro8_s(0)
    );
  romeaddro8_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro8_s_1_SRINV,
      I1 => GSR,
      O => romeaddro8_s_1_FFY_RST
    );
  U_DCT1D_reg_romeaddro8_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro8_s_1_DXMUX,
      CE => romeaddro8_s_1_CEINV,
      CLK => romeaddro8_s_1_CLKINV,
      SET => GND,
      RST => romeaddro8_s_1_FFX_RST,
      O => romeaddro8_s(1)
    );
  romeaddro8_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro8_s_1_SRINV,
      I1 => GSR,
      O => romeaddro8_s_1_FFX_RST
    );
  U_DCT1D_reg_romeaddro8_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro8_s_3_DYMUX,
      CE => romeaddro8_s_3_CEINV,
      CLK => romeaddro8_s_3_CLKINV,
      SET => GND,
      RST => romeaddro8_s_3_FFY_RST,
      O => romeaddro8_s(2)
    );
  romeaddro8_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro8_s_3_SRINV,
      I1 => GSR,
      O => romeaddro8_s_3_FFY_RST
    );
  U_DCT2D_ix45659z1511 : X_LUT4
    generic map(
      INIT => X"A0AA"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => VCC,
      ADR2 => U_DCT2D_NOT_rtlcs7,
      ADR3 => U_DCT2D_state_reg(1),
      O => U_DCT2D_rtlc5n1854_G
    );
  U_DCT1D_reg_romeaddro8_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro8_s_3_DXMUX,
      CE => romeaddro8_s_3_CEINV,
      CLK => romeaddro8_s_3_CLKINV,
      SET => GND,
      RST => romeaddro8_s_3_FFX_RST,
      O => romeaddro8_s(3)
    );
  romeaddro8_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro8_s_3_SRINV,
      I1 => GSR,
      O => romeaddro8_s_3_FFX_RST
    );
  U_DCT2D_ix62982z1321 : X_LUT4
    generic map(
      INIT => X"33FF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => VCC,
      ADR3 => U_DCT2D_state_reg(1),
      O => U_DCT2D_rtlc5n1854_F
    );
  U_DCT2D_ix65206z2037 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao7_s(13),
      ADR2 => romo2datao6_s(13),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z253_G
    );
  U_DCT2D_ix65206z1321 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT2D_rtlc5n1499(23),
      ADR3 => U_DCT2D_rtlc5n1501(23),
      O => U_DCT2D_nx65206z1_G
    );
  U_DCT2D_ix65206z1327 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao2_s(13),
      ADR2 => VCC,
      ADR3 => rome2datao3_s(13),
      O => U_DCT2D_nx65206z5_G
    );
  U_DCT1D_reg_romeaddro4_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro4_s_3_DXMUX,
      CE => romeaddro4_s_3_CEINV,
      CLK => romeaddro4_s_3_CLKINV,
      SET => GND,
      RST => romeaddro4_s_3_FFX_RST,
      O => romeaddro4_s(3)
    );
  romeaddro4_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro4_s_3_SRINV,
      I1 => GSR,
      O => romeaddro4_s_3_FFX_RST
    );
  U_DCT1D_reg_romeaddro5_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro5_s_1_DYMUX,
      CE => romeaddro5_s_1_CEINV,
      CLK => romeaddro5_s_1_CLKINV,
      SET => GND,
      RST => romeaddro5_s_1_FFY_RST,
      O => romeaddro5_s(0)
    );
  romeaddro5_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro5_s_1_SRINV,
      I1 => GSR,
      O => romeaddro5_s_1_FFY_RST
    );
  U_DCT1D_reg_romeaddro5_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro5_s_1_DXMUX,
      CE => romeaddro5_s_1_CEINV,
      CLK => romeaddro5_s_1_CLKINV,
      SET => GND,
      RST => romeaddro5_s_1_FFX_RST,
      O => romeaddro5_s(1)
    );
  romeaddro5_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro5_s_1_SRINV,
      I1 => GSR,
      O => romeaddro5_s_1_FFX_RST
    );
  U_DCT1D_reg_romeaddro5_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro5_s_3_DYMUX,
      CE => romeaddro5_s_3_CEINV,
      CLK => romeaddro5_s_3_CLKINV,
      SET => GND,
      RST => romeaddro5_s_3_FFY_RST,
      O => romeaddro5_s(2)
    );
  romeaddro5_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro5_s_3_SRINV,
      I1 => GSR,
      O => romeaddro5_s_3_FFY_RST
    );
  U_DCT1D_reg_romeaddro5_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro5_s_3_DXMUX,
      CE => romeaddro5_s_3_CEINV,
      CLK => romeaddro5_s_3_CLKINV,
      SET => GND,
      RST => romeaddro5_s_3_FFX_RST,
      O => romeaddro5_s(3)
    );
  romeaddro5_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro5_s_3_SRINV,
      I1 => GSR,
      O => romeaddro5_s_3_FFX_RST
    );
  U_DCT2D_reg_romoaddro10_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro10_s_1_DYMUX,
      CE => romo2addro10_s_1_CEINV,
      CLK => romo2addro10_s_1_CLKINV,
      SET => GND,
      RST => romo2addro10_s_1_FFY_RST,
      O => romo2addro10_s(0)
    );
  romo2addro10_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro10_s_1_SRINV,
      I1 => GSR,
      O => romo2addro10_s_1_FFY_RST
    );
  U_DCT2D_reg_state_reg_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_state_reg_1_DXMUX,
      CE => U_DCT2D_state_reg_1_CEINV,
      CLK => U_DCT2D_state_reg_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_state_reg_1_FFX_RST,
      O => U_DCT2D_state_reg(1)
    );
  U_DCT2D_state_reg_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_state_reg_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_state_reg_1_FFX_RST
    );
  U_DCT2D_reg_romeaddro10_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro10_s_1_DYMUX,
      CE => rome2addro10_s_1_CEINV,
      CLK => rome2addro10_s_1_CLKINV,
      SET => GND,
      RST => rome2addro10_s_1_FFY_RST,
      O => rome2addro10_s(0)
    );
  rome2addro10_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro10_s_1_SRINV,
      I1 => GSR,
      O => rome2addro10_s_1_FFY_RST
    );
  U_DCT2D_reg_romeaddro10_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro10_s_1_DXMUX,
      CE => rome2addro10_s_1_CEINV,
      CLK => rome2addro10_s_1_CLKINV,
      SET => GND,
      RST => rome2addro10_s_1_FFX_RST,
      O => rome2addro10_s(1)
    );
  rome2addro10_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro10_s_1_SRINV,
      I1 => GSR,
      O => rome2addro10_s_1_FFX_RST
    );
  U_DCT2D_reg_romeaddro10_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro10_s_3_DYMUX,
      CE => rome2addro10_s_3_CEINV,
      CLK => rome2addro10_s_3_CLKINV,
      SET => GND,
      RST => rome2addro10_s_3_FFY_RST,
      O => rome2addro10_s(2)
    );
  rome2addro10_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro10_s_3_SRINV,
      I1 => GSR,
      O => rome2addro10_s_3_FFY_RST
    );
  U_DCT1D_ix6411z1186 : X_LUT4
    generic map(
      INIT => X"FF7F"
    )
    port map (
      ADR0 => U_DCT1D_row_reg(2),
      ADR1 => U_DCT1D_row_reg(0),
      ADR2 => U_DCT1D_row_reg(1),
      ADR3 => U_DCT1D_NOT_rtlcs7,
      O => U_DCT1D_rtlc5n1684_G
    );
  U_DCT2D_reg_romeaddro10_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro10_s_3_DXMUX,
      CE => rome2addro10_s_3_CEINV,
      CLK => rome2addro10_s_3_CLKINV,
      SET => GND,
      RST => rome2addro10_s_3_FFX_RST,
      O => rome2addro10_s(3)
    );
  rome2addro10_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro10_s_3_SRINV,
      I1 => GSR,
      O => rome2addro10_s_3_FFX_RST
    );
  U_DCT1D_ix932z1339 : X_LUT4
    generic map(
      INIT => X"0C33"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_state_reg(1),
      ADR2 => U_DCT1D_rtlc5n1311,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_rtlc5n1684_F
    );
  U_DCT2D_ix65206z1468 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romo2datao3_s(13),
      ADR1 => romo2datao2_s(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z121_G
    );
  U_DCT2D_ix65206z1825 : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1485(16),
      ADR1 => VCC,
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => U_DCT2D_rtlc5n1492(15),
      O => U_DCT2D_nx65206z215_F
    );
  U_DCT2D_ix65206z1732 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => rome2datao5_s(13),
      ADR1 => rome2datao4_s(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z297_G
    );
  U_DCT2D_ix65206z2372 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => rome2datao8_s(7),
      ADR3 => romo2datao8_s(7),
      O => U_DCT2D_nx65206z595_F
    );
  U_DCT2D_ix65206z2381 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => rome2datao8_s(4),
      ADR2 => romo2datao8_s(4),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z604_F
    );
  U_DCT2D_ix65206z2357 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => romo2datao8_s(12),
      ADR2 => VCC,
      ADR3 => rome2datao8_s(12),
      O => U_DCT2D_nx65206z580_F
    );
  U_DCT2D_ix65206z2366 : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => rome2datao8_s(9),
      ADR1 => VCC,
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => romo2datao8_s(9),
      O => U_DCT2D_nx65206z589_F
    );
  U_DCT2D_ix65206z2375 : X_LUT4
    generic map(
      INIT => X"ACAC"
    )
    port map (
      ADR0 => romo2datao8_s(6),
      ADR1 => rome2datao8_s(6),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z598_F
    );
  U_DCT2D_ix65206z2384 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao8_s(3),
      ADR2 => romo2datao8_s(3),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z607_F
    );
  U_DCT2D_ix65206z2473 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => romo2datao5_s(13),
      ADR3 => romo2datao4_s(13),
      O => U_DCT2D_nx65206z413_G
    );
  U_DCT1D_reg_romeaddro1_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro1_s_3_DXMUX,
      CE => romeaddro1_s_3_CEINV,
      CLK => romeaddro1_s_3_CLKINV,
      SET => GND,
      RST => romeaddro1_s_3_FFX_RST,
      O => romeaddro1_s(3)
    );
  romeaddro1_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro1_s_3_SRINV,
      I1 => GSR,
      O => romeaddro1_s_3_FFX_RST
    );
  U_DCT1D_reg_romeaddro2_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro2_s_1_DYMUX,
      CE => romeaddro2_s_1_CEINV,
      CLK => romeaddro2_s_1_CLKINV,
      SET => GND,
      RST => romeaddro2_s_1_FFY_RST,
      O => romeaddro2_s(0)
    );
  romeaddro2_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro2_s_1_SRINV,
      I1 => GSR,
      O => romeaddro2_s_1_FFY_RST
    );
  U_DCT1D_reg_romeaddro2_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro2_s_1_DXMUX,
      CE => romeaddro2_s_1_CEINV,
      CLK => romeaddro2_s_1_CLKINV,
      SET => GND,
      RST => romeaddro2_s_1_FFX_RST,
      O => romeaddro2_s(1)
    );
  romeaddro2_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro2_s_1_SRINV,
      I1 => GSR,
      O => romeaddro2_s_1_FFX_RST
    );
  U_DCT1D_reg_romeaddro2_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro2_s_3_DYMUX,
      CE => romeaddro2_s_3_CEINV,
      CLK => romeaddro2_s_3_CLKINV,
      SET => GND,
      RST => romeaddro2_s_3_FFY_RST,
      O => romeaddro2_s(2)
    );
  romeaddro2_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro2_s_3_SRINV,
      I1 => GSR,
      O => romeaddro2_s_3_FFY_RST
    );
  U_DCT1D_reg_romeaddro2_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro2_s_3_DXMUX,
      CE => romeaddro2_s_3_CEINV,
      CLK => romeaddro2_s_3_CLKINV,
      SET => GND,
      RST => romeaddro2_s_3_FFX_RST,
      O => romeaddro2_s(3)
    );
  romeaddro2_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro2_s_3_SRINV,
      I1 => GSR,
      O => romeaddro2_s_3_FFX_RST
    );
  U_DCT1D_reg_romeaddro3_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro3_s_1_DYMUX,
      CE => romeaddro3_s_1_CEINV,
      CLK => romeaddro3_s_1_CLKINV,
      SET => GND,
      RST => romeaddro3_s_1_FFY_RST,
      O => romeaddro3_s(0)
    );
  romeaddro3_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro3_s_1_SRINV,
      I1 => GSR,
      O => romeaddro3_s_1_FFY_RST
    );
  U_DCT1D_reg_romeaddro0_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro0_s_1_DYMUX,
      CE => romeaddro0_s_1_CEINV,
      CLK => romeaddro0_s_1_CLKINV,
      SET => GND,
      RST => romeaddro0_s_1_FFY_RST,
      O => romeaddro0_s(0)
    );
  romeaddro0_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro0_s_1_SRINV,
      I1 => GSR,
      O => romeaddro0_s_1_FFY_RST
    );
  U_DCT1D_reg_romeaddro0_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro0_s_1_DXMUX,
      CE => romeaddro0_s_1_CEINV,
      CLK => romeaddro0_s_1_CLKINV,
      SET => GND,
      RST => romeaddro0_s_1_FFX_RST,
      O => romeaddro0_s(1)
    );
  romeaddro0_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro0_s_1_SRINV,
      I1 => GSR,
      O => romeaddro0_s_1_FFX_RST
    );
  U_DCT1D_reg_romeaddro0_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro0_s_3_DYMUX,
      CE => romeaddro0_s_3_CEINV,
      CLK => romeaddro0_s_3_CLKINV,
      SET => GND,
      RST => romeaddro0_s_3_FFY_RST,
      O => romeaddro0_s(2)
    );
  romeaddro0_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro0_s_3_SRINV,
      I1 => GSR,
      O => romeaddro0_s_3_FFY_RST
    );
  U_DCT1D_reg_romeaddro0_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro0_s_3_DXMUX,
      CE => romeaddro0_s_3_CEINV,
      CLK => romeaddro0_s_3_CLKINV,
      SET => GND,
      RST => romeaddro0_s_3_FFX_RST,
      O => romeaddro0_s(3)
    );
  romeaddro0_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro0_s_3_SRINV,
      I1 => GSR,
      O => romeaddro0_s_3_FFX_RST
    );
  U_DCT1D_reg_romeaddro1_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro1_s_1_DYMUX,
      CE => romeaddro1_s_1_CEINV,
      CLK => romeaddro1_s_1_CLKINV,
      SET => GND,
      RST => romeaddro1_s_1_FFY_RST,
      O => romeaddro1_s(0)
    );
  romeaddro1_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro1_s_1_SRINV,
      I1 => GSR,
      O => romeaddro1_s_1_FFY_RST
    );
  U_DCT1D_reg_romeaddro1_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro1_s_1_DXMUX,
      CE => romeaddro1_s_1_CEINV,
      CLK => romeaddro1_s_1_CLKINV,
      SET => GND,
      RST => romeaddro1_s_1_FFX_RST,
      O => romeaddro1_s(1)
    );
  romeaddro1_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro1_s_1_SRINV,
      I1 => GSR,
      O => romeaddro1_s_1_FFX_RST
    );
  U_DCT1D_reg_romeaddro1_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro1_s_3_DYMUX,
      CE => romeaddro1_s_3_CEINV,
      CLK => romeaddro1_s_3_CLKINV,
      SET => GND,
      RST => romeaddro1_s_3_FFY_RST,
      O => romeaddro1_s(2)
    );
  romeaddro1_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro1_s_3_SRINV,
      I1 => GSR,
      O => romeaddro1_s_3_FFY_RST
    );
  U_DCT2D_reg_romoaddro10_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro10_s_1_DXMUX,
      CE => romo2addro10_s_1_CEINV,
      CLK => romo2addro10_s_1_CLKINV,
      SET => GND,
      RST => romo2addro10_s_1_FFX_RST,
      O => romo2addro10_s(1)
    );
  romo2addro10_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro10_s_1_SRINV,
      I1 => GSR,
      O => romo2addro10_s_1_FFX_RST
    );
  U_DCT1D_reg_romeaddro6_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro6_s_1_DYMUX,
      CE => romeaddro6_s_1_CEINV,
      CLK => romeaddro6_s_1_CLKINV,
      SET => GND,
      RST => romeaddro6_s_1_FFY_RST,
      O => romeaddro6_s(0)
    );
  romeaddro6_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro6_s_1_SRINV,
      I1 => GSR,
      O => romeaddro6_s_1_FFY_RST
    );
  U_DCT1D_reg_romeaddro6_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro6_s_1_DXMUX,
      CE => romeaddro6_s_1_CEINV,
      CLK => romeaddro6_s_1_CLKINV,
      SET => GND,
      RST => romeaddro6_s_1_FFX_RST,
      O => romeaddro6_s(1)
    );
  romeaddro6_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romeaddro6_s_1_SRINV,
      I1 => GSR,
      O => romeaddro6_s_1_FFX_RST
    );
  U_DCT2D_reg_romoaddro10_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro10_s_3_DYMUX,
      CE => romo2addro10_s_3_CEINV,
      CLK => romo2addro10_s_3_CLKINV,
      SET => GND,
      RST => romo2addro10_s_3_FFY_RST,
      O => romo2addro10_s(2)
    );
  romo2addro10_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romo2addro10_s_3_SRINV,
      I1 => GSR,
      O => romo2addro10_s_3_FFY_RST
    );
  U_DCT2D_reg_romoaddro10_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romo2addro10_s_3_DXMUX,
      CE => romo2addro10_s_3_CEINV,
      CLK => romo2addro10_s_3_CLKINV,
      SET => GND,
      RST => romo2addro10_s_3_FFX_RST,
      O => romo2addro10_s(3)
    );
  romo2addro10_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romo2addro10_s_3_SRINV,
      I1 => GSR,
      O => romo2addro10_s_3_FFX_RST
    );
  U_DCT1D_reg_romeaddro6_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romeaddro6_s_3_DYMUX,
      CE => romeaddro6_s_3_CEINV,
      CLK => romeaddro6_s_3_CLKINV,
      SET => GND,
      RST => romeaddro6_s_3_FFY_RST,
      O => romeaddro6_s(2)
    );
  romeaddro6_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romeaddro6_s_3_SRINV,
      I1 => GSR,
      O => romeaddro6_s_3_FFY_RST
    );
  U_DCT2D_ix65206z1416 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1480(15),
      ADR1 => VCC,
      ADR2 => U_DCT2D_rtlc5n1481(17),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z78_G
    );
  U_DCT2D_ix65206z1418 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romo2datao1_s(13),
      ADR2 => VCC,
      ADR3 => romo2datao0_s(13),
      O => U_DCT2D_nx65206z79_G
    );
  U_DCT2D_ix65206z1371 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao0_s(13),
      ADR2 => rome2datao1_s(13),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z42_G
    );
  U_DCT2D_ix65206z2350 : X_LUT4
    generic map(
      INIT => X"D8D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => romo2datao8_s(13),
      ADR2 => rome2datao8_s(13),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z572_G
    );
  U_DCT2D_ix65206z24305 : X_LUT4
    generic map(
      INIT => X"27D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => romo2datao9_s(13),
      ADR2 => rome2datao9_s(13),
      ADR3 => U_DCT2D_nx65206z573,
      O => U_DCT2D_nx65206z572_F
    );
  U_DCT2D_ix65206z1730 : X_LUT4
    generic map(
      INIT => X"55AA"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1494(19),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT2D_rtlc5n1495(21),
      O => U_DCT2D_nx65206z296_G
    );
  U_DCT2D_ix65206z2360 : X_LUT4
    generic map(
      INIT => X"D8D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => romo2datao8_s(11),
      ADR2 => rome2datao8_s(11),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z583_F
    );
  U_DCT2D_ix65206z2363 : X_LUT4
    generic map(
      INIT => X"EE22"
    )
    port map (
      ADR0 => rome2datao8_s(10),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => VCC,
      ADR3 => romo2datao8_s(10),
      O => U_DCT2D_nx65206z586_F
    );
  U_DCT2D_ix65206z1820 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1485(17),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => U_DCT2D_rtlc5n1492(15),
      O => U_DCT2D_nx65206z215_G
    );
  U_DCT1D_modgen_counter_inpcnt_reg_reg_q_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_inpcnt_reg_0_DXMUX,
      CE => U_DCT1D_inpcnt_reg_0_CEINV,
      CLK => U_DCT1D_inpcnt_reg_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_inpcnt_reg_0_FFX_RST,
      O => U_DCT1D_inpcnt_reg(0)
    );
  U_DCT1D_inpcnt_reg_0_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_inpcnt_reg_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_inpcnt_reg_0_FFX_RST
    );
  U_DCT1D_reg_ramwe_s : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramwe_s_DYMUX,
      CE => ramwe_s_CEINV,
      CLK => ramwe_s_CLKINV,
      SET => GND,
      RST => ramwe_s_FFY_RST,
      O => ramwe_s
    );
  ramwe_s_FFY_RSTOR : X_OR2
    port map (
      I0 => ramwe_s_FFY_RSTAND,
      I1 => GSR,
      O => ramwe_s_FFY_RST
    );
  ramwe_s_FFY_RSTAND_7786 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => ramwe_s_FFY_RSTAND
    );
  U_DCT2D_reg_romeaddro0_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro0_s_1_DYMUX,
      CE => rome2addro0_s_1_CEINV,
      CLK => rome2addro0_s_1_CLKINV,
      SET => GND,
      RST => rome2addro0_s_1_FFY_RST,
      O => rome2addro0_s(0)
    );
  rome2addro0_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro0_s_1_SRINV,
      I1 => GSR,
      O => rome2addro0_s_1_FFY_RST
    );
  U_DCT2D_reg_romeaddro0_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro0_s_1_DXMUX,
      CE => rome2addro0_s_1_CEINV,
      CLK => rome2addro0_s_1_CLKINV,
      SET => GND,
      RST => rome2addro0_s_1_FFX_RST,
      O => rome2addro0_s(1)
    );
  rome2addro0_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro0_s_1_SRINV,
      I1 => GSR,
      O => rome2addro0_s_1_FFX_RST
    );
  U_DCT2D_reg_romeaddro0_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro0_s_3_DYMUX,
      CE => rome2addro0_s_3_CEINV,
      CLK => rome2addro0_s_3_CLKINV,
      SET => GND,
      RST => rome2addro0_s_3_FFY_RST,
      O => rome2addro0_s(2)
    );
  rome2addro0_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro0_s_3_SRINV,
      I1 => GSR,
      O => rome2addro0_s_3_FFY_RST
    );
  U_DCT2D_reg_romeaddro0_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro0_s_3_DXMUX,
      CE => rome2addro0_s_3_CEINV,
      CLK => rome2addro0_s_3_CLKINV,
      SET => GND,
      RST => rome2addro0_s_3_FFX_RST,
      O => rome2addro0_s(3)
    );
  rome2addro0_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro0_s_3_SRINV,
      I1 => GSR,
      O => rome2addro0_s_3_FFX_RST
    );
  U_DCT2D_ix65206z1866 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => VCC,
      ADR2 => U_DCT2D_rtlc5n1492(9),
      ADR3 => U_DCT2D_rtlc5n1485(9),
      O => U_DCT2D_nx65206z236_G
    );
  U_DCT2D_ix65206z1884 : X_LUT4
    generic map(
      INIT => X"E2E2"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1492(6),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => U_DCT2D_rtlc5n1485(6),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z245_G
    );
  U_DCT2D_ix65206z1878 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1485(7),
      ADR2 => U_DCT2D_rtlc5n1492(7),
      ADR3 => U_DCT2D_state_reg(0),
      O => U_DCT2D_nx65206z242_G
    );
  U_DCT2D_reg_requestrd_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => requestrd_s_DYMUX,
      CE => requestrd_s_CEINV,
      CLK => requestrd_s_CLKINV,
      SET => GND,
      RST => requestrd_s_FFY_RST,
      O => requestrd_s
    );
  requestrd_s_FFY_RSTOR : X_OR2
    port map (
      I0 => requestrd_s_FFY_RSTAND,
      I1 => GSR,
      O => requestrd_s_FFY_RST
    );
  requestrd_s_FFY_RSTAND_7787 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => requestrd_s_FFY_RSTAND
    );
  U_DCT2D_ix49413z1331 : X_LUT4
    generic map(
      INIT => X"FFAA"
    )
    port map (
      ADR0 => ramraddro_s(1),
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => ramraddro_s(0),
      O => U_DCT2D_rtlc2n446_G
    );
  U_DCT2D_ix49413z1827 : X_LUT4
    generic map(
      INIT => X"0200"
    )
    port map (
      ADR0 => U_DCT2D_colram_reg(3),
      ADR1 => U_DCT2D_nx49413z1,
      ADR2 => ramraddro_s(2),
      ADR3 => U_DCT2D_NOT_rtlc2n488,
      O => U_DCT2D_rtlc2n446_F
    );
  U_DCT1D_ix7397z1321 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_6_Q(7),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_1_Q(7),
      ADR3 => VCC,
      O => U_DCT1D_nx52393z1_G
    );
  U_DCT2D_ix49413z1318 : X_LUT4
    generic map(
      INIT => X"00F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT2D_istate_reg(1),
      ADR3 => U_DCT2D_istate_reg(0),
      O => U_DCT2D_nx40895z2_G
    );
  U_DCT2D_ix40895z37923 : X_LUT4
    generic map(
      INIT => X"B030"
    )
    port map (
      ADR0 => ramraddro_s(0),
      ADR1 => U_DCT2D_NOT_rtlcs2,
      ADR2 => U_DCT2D_NOT_rtlc2n488,
      ADR3 => ramraddro_s(1),
      O => U_DCT2D_nx40895z2_F
    );
  U_DCT1D_reg_ramwaddro_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramwaddro_s_1_DXMUX,
      CE => ramwaddro_s_1_CEINV,
      CLK => ramwaddro_s_1_CLKINV,
      SET => GND,
      RST => ramwaddro_s_1_FFX_RST,
      O => ramwaddro_s(1)
    );
  ramwaddro_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => ramwaddro_s_1_SRINV,
      I1 => GSR,
      O => ramwaddro_s_1_FFX_RST
    );
  U_DCT1D_reg_ramwaddro_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramwaddro_s_3_DYMUX,
      CE => ramwaddro_s_3_CEINV,
      CLK => ramwaddro_s_3_CLKINV,
      SET => GND,
      RST => ramwaddro_s_3_FFY_RST,
      O => ramwaddro_s(2)
    );
  ramwaddro_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => ramwaddro_s_3_SRINV,
      I1 => GSR,
      O => ramwaddro_s_3_FFY_RST
    );
  U_DCT1D_reg_ramwaddro_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramwaddro_s_3_DXMUX,
      CE => ramwaddro_s_3_CEINV,
      CLK => ramwaddro_s_3_CLKINV,
      SET => GND,
      RST => ramwaddro_s_3_FFX_RST,
      O => ramwaddro_s(3)
    );
  ramwaddro_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => ramwaddro_s_3_SRINV,
      I1 => GSR,
      O => ramwaddro_s_3_FFX_RST
    );
  U_DCT1D_reg_ramwaddro_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramwaddro_s_5_DYMUX,
      CE => ramwaddro_s_5_CEINV,
      CLK => ramwaddro_s_5_CLKINV,
      SET => GND,
      RST => ramwaddro_s_5_FFY_RST,
      O => ramwaddro_s(4)
    );
  ramwaddro_s_5_FFY_RSTOR : X_OR2
    port map (
      I0 => ramwaddro_s_5_SRINV,
      I1 => GSR,
      O => ramwaddro_s_5_FFY_RST
    );
  U_DCT1D_reg_ramwaddro_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramwaddro_s_5_DXMUX,
      CE => ramwaddro_s_5_CEINV,
      CLK => ramwaddro_s_5_CLKINV,
      SET => GND,
      RST => ramwaddro_s_5_FFX_RST,
      O => ramwaddro_s(5)
    );
  ramwaddro_s_5_FFX_RSTOR : X_OR2
    port map (
      I0 => ramwaddro_s_5_SRINV,
      I1 => GSR,
      O => ramwaddro_s_5_FFX_RST
    );
  U_DCT1D_ix58996z1320 : X_LUT4
    generic map(
      INIT => X"0FF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT1D_inpcnt_reg(0),
      ADR3 => U_DCT1D_inpcnt_reg(1),
      O => U_DCT1D_nx58996z1
    );
  U_DCT1D_modgen_counter_inpcnt_reg_reg_q_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_inpcnt_reg_0_DYMUX,
      CE => U_DCT1D_inpcnt_reg_0_CEINV,
      CLK => U_DCT1D_inpcnt_reg_0_CLKINV,
      SET => GND,
      RST => U_DCT1D_inpcnt_reg_0_FFY_RST,
      O => U_DCT1D_inpcnt_reg(1)
    );
  U_DCT1D_inpcnt_reg_0_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_inpcnt_reg_0_SRINV,
      I1 => GSR,
      O => U_DCT1D_inpcnt_reg_0_FFY_RST
    );
  U_DCT2D_reg_completed_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_completed_reg_DYMUX,
      CE => U_DCT2D_completed_reg_CEINV,
      CLK => U_DCT2D_completed_reg_CLKINV,
      SET => GND,
      RST => U_DCT2D_completed_reg_FFY_RST,
      O => U_DCT2D_completed_reg
    );
  U_DCT2D_completed_reg_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_completed_reg_FFY_RSTAND,
      I1 => GSR,
      O => U_DCT2D_completed_reg_FFY_RST
    );
  U_DCT2D_completed_reg_FFY_RSTAND_7788 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_completed_reg_FFY_RSTAND
    );
  U_DCT2D_ix31471z1320 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT2D_col_reg(1),
      ADR1 => U_DCT2D_col_reg(2),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_rtlc5n942(2)
    );
  U_DCT2D_reg_col_tmp_reg_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_col_tmp_reg_1_DYMUX,
      CE => U_DCT2D_col_tmp_reg_1_CEINV,
      CLK => U_DCT2D_col_tmp_reg_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_col_tmp_reg_1_FFY_RST,
      O => U_DCT2D_col_tmp_reg(2)
    );
  U_DCT2D_col_tmp_reg_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_col_tmp_reg_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_col_tmp_reg_1_FFY_RST
    );
  U_DCT1D_ix53004z1321 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_7_Q(7),
      ADR1 => U_DCT1D_latchbuf_reg_0_Q(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx57528z1_G
    );
  U_DCT2D_reg_col_tmp_reg_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_col_tmp_reg_1_DXMUX,
      CE => U_DCT2D_col_tmp_reg_1_CEINV,
      CLK => U_DCT2D_col_tmp_reg_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_col_tmp_reg_1_FFX_RST,
      O => U_DCT2D_col_tmp_reg(1)
    );
  U_DCT2D_col_tmp_reg_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_col_tmp_reg_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_col_tmp_reg_1_FFX_RST
    );
  U_DCT1D_ix57528z1324 : X_LUT4
    generic map(
      INIT => X"9999"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_7_Q(7),
      ADR1 => U_DCT1D_latchbuf_reg_0_Q(7),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx57528z1_F
    );
  U_DCT1D_reg_ramwaddro_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => ramwaddro_s_1_DYMUX,
      CE => ramwaddro_s_1_CEINV,
      CLK => ramwaddro_s_1_CLKINV,
      SET => GND,
      RST => ramwaddro_s_1_FFY_RST,
      O => ramwaddro_s(0)
    );
  ramwaddro_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => ramwaddro_s_1_SRINV,
      I1 => GSR,
      O => ramwaddro_s_1_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_5_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_1_DYMUX,
      CE => U_DCT2D_latchbuf_reg_5_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_5_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_5_1_FFY_RST,
      O => U_DCT2D_latchbuf_reg_5_0_Q
    );
  U_DCT2D_latchbuf_reg_5_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_5_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_5_1_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_5_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_1_DXMUX,
      CE => U_DCT2D_latchbuf_reg_5_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_5_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_5_1_FFX_RST,
      O => U_DCT2D_latchbuf_reg_5_1_Q
    );
  U_DCT2D_latchbuf_reg_5_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_5_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_5_1_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_5_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_3_DYMUX,
      CE => U_DCT2D_latchbuf_reg_5_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_5_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_5_3_FFY_RST,
      O => U_DCT2D_latchbuf_reg_5_2_Q
    );
  U_DCT2D_latchbuf_reg_5_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_5_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_5_3_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_5_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_3_DXMUX,
      CE => U_DCT2D_latchbuf_reg_5_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_5_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_5_3_FFX_RST,
      O => U_DCT2D_latchbuf_reg_5_3_Q
    );
  U_DCT2D_latchbuf_reg_5_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_5_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_5_3_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_5_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_5_DYMUX,
      CE => U_DCT2D_latchbuf_reg_5_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_5_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_5_5_FFY_RST,
      O => U_DCT2D_latchbuf_reg_5_4_Q
    );
  U_DCT2D_latchbuf_reg_5_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_5_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_5_5_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_5_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_5_DXMUX,
      CE => U_DCT2D_latchbuf_reg_5_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_5_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_5_5_FFX_RST,
      O => U_DCT2D_latchbuf_reg_5_5_Q
    );
  U_DCT2D_latchbuf_reg_5_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_5_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_5_5_FFX_RST
    );
  U_DCT1D_reg_releasewr_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => releasewr_s_DYMUX,
      CE => releasewr_s_CEINV,
      CLK => releasewr_s_CLKINV,
      SET => GND,
      RST => releasewr_s_FFY_RST,
      O => releasewr_s
    );
  releasewr_s_FFY_RSTOR : X_OR2
    port map (
      I0 => releasewr_s_FFY_RSTAND,
      I1 => GSR,
      O => releasewr_s_FFY_RST
    );
  releasewr_s_FFY_RSTAND_7789 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => releasewr_s_FFY_RSTAND
    );
  U_DCT1D_reg_latch_done_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_latch_done_reg_DYMUX,
      CE => U_DCT1D_latch_done_reg_CEINV,
      CLK => U_DCT1D_latch_done_reg_CLKINV,
      SET => GND,
      RST => U_DCT1D_latch_done_reg_FFY_RST,
      O => U_DCT1D_latch_done_reg
    );
  U_DCT1D_latch_done_reg_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_latch_done_reg_FFY_RSTAND,
      I1 => GSR,
      O => U_DCT1D_latch_done_reg_FFY_RST
    );
  U_DCT1D_latch_done_reg_FFY_RSTAND_7790 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT1D_latch_done_reg_FFY_RSTAND
    );
  U_DCT1D_ix31471z1317 : X_LUT4
    generic map(
      INIT => X"0F00"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_state_reg(1),
      O => U_DCT1D_NOT_rtlcs2_G
    );
  U_DCT1D_ix55759z1321 : X_LUT4
    generic map(
      INIT => X"0FFF"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_state_reg(1),
      O => U_DCT1D_NOT_rtlcs2_F
    );
  U_DCT1D_ix42123z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_3_Q(7),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_4_Q(7),
      ADR3 => VCC,
      O => U_DCT1D_nx62663z1_G
    );
  U_DCT1D_ix62663z1321 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_3_Q(7),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_4_Q(7),
      ADR3 => VCC,
      O => U_DCT1D_nx62663z1_F
    );
  U_DCT1D_ix51043z1379 : X_LUT4
    generic map(
      INIT => X"2020"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(1),
      ADR1 => U_DCT1D_NOT_rtlcs7,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => VCC,
      O => U_DCT1D_rtlc5n1612_G
    );
  U_DCT1D_ix53916z1511 : X_LUT4
    generic map(
      INIT => X"D0D0"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(1),
      ADR1 => U_DCT1D_NOT_rtlcs7,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => VCC,
      O => U_DCT1D_rtlc5n1612_F
    );
  U_DCT2D_reg_latchbuf_reg_3_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_7_DXMUX,
      CE => U_DCT2D_latchbuf_reg_3_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_3_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_3_7_FFX_RST,
      O => U_DCT2D_latchbuf_reg_3_7_Q
    );
  U_DCT2D_latchbuf_reg_3_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_3_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_3_7_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_3_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_10_DYMUX,
      CE => U_DCT2D_latchbuf_reg_3_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_3_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_3_10_FFY_RST,
      O => U_DCT2D_latchbuf_reg_3_8_Q
    );
  U_DCT2D_latchbuf_reg_3_10_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_3_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_3_10_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_3_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_10_DXMUX,
      CE => U_DCT2D_latchbuf_reg_3_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_3_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_3_10_FFX_RST,
      O => U_DCT2D_latchbuf_reg_3_10_Q
    );
  U_DCT2D_latchbuf_reg_3_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_3_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_3_10_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_4_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_1_DYMUX,
      CE => U_DCT2D_latchbuf_reg_4_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_4_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_4_1_FFY_RST,
      O => U_DCT2D_latchbuf_reg_4_0_Q
    );
  U_DCT2D_latchbuf_reg_4_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_4_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_4_1_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_4_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_1_DXMUX,
      CE => U_DCT2D_latchbuf_reg_4_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_4_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_4_1_FFX_RST,
      O => U_DCT2D_latchbuf_reg_4_1_Q
    );
  U_DCT2D_latchbuf_reg_4_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_4_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_4_1_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_4_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_4_3_DYMUX,
      CE => U_DCT2D_latchbuf_reg_4_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_4_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_4_3_FFY_RST,
      O => U_DCT2D_latchbuf_reg_4_2_Q
    );
  U_DCT2D_latchbuf_reg_4_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_4_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_4_3_FFY_RST
    );
  U_DCT2D_ix65206z2369 : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => rome2datao8_s(8),
      ADR1 => romo2datao8_s(8),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z592_F
    );
  U_DCT2D_ix65206z1842 : X_LUT4
    generic map(
      INIT => X"D8D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1485(13),
      ADR2 => U_DCT2D_rtlc5n1492(13),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z224_G
    );
  U_DCT2D_ix65206z2378 : X_LUT4
    generic map(
      INIT => X"BB88"
    )
    port map (
      ADR0 => romo2datao8_s(5),
      ADR1 => U_DCT2D_state_reg(0),
      ADR2 => VCC,
      ADR3 => rome2datao8_s(5),
      O => U_DCT2D_nx65206z601_F
    );
  U_DCT2D_ix65206z1860 : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1492(10),
      ADR1 => U_DCT2D_rtlc5n1485(10),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z233_G
    );
  U_DCT2D_ix65206z1836 : X_LUT4
    generic map(
      INIT => X"CACA"
    )
    port map (
      ADR0 => U_DCT2D_rtlc5n1492(14),
      ADR1 => U_DCT2D_rtlc5n1485(14),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z221_G
    );
  U_DCT2D_ix65206z1854 : X_LUT4
    generic map(
      INIT => X"D8D8"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1485(11),
      ADR2 => U_DCT2D_rtlc5n1492(11),
      ADR3 => VCC,
      O => U_DCT2D_nx65206z230_G
    );
  U_DCT2D_ix65206z1872 : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT2D_rtlc5n1492(8),
      ADR2 => U_DCT2D_state_reg(0),
      ADR3 => U_DCT2D_rtlc5n1485(8),
      O => U_DCT2D_nx65206z239_G
    );
  U_DCT2D_ix65206z1848 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1492(12),
      ADR2 => VCC,
      ADR3 => U_DCT2D_rtlc5n1485(12),
      O => U_DCT2D_nx65206z227_G
    );
  U_DCT2D_ix65206z1776 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => rome2datao6_s(13),
      ADR2 => VCC,
      ADR3 => rome2datao7_s(13),
      O => U_DCT2D_nx65206z334_G
    );
  U_DCT2D_ix65206z1890 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => U_DCT2D_state_reg(0),
      ADR1 => U_DCT2D_rtlc5n1492(5),
      ADR2 => VCC,
      ADR3 => U_DCT2D_rtlc5n1485(5),
      O => U_DCT2D_nx65206z248_G
    );
  U_DCT1D_ix9237z1442 : X_LUT4
    generic map(
      INIT => X"77FF"
    )
    port map (
      ADR0 => U_DCT1D_inpcnt_reg(1),
      ADR1 => U_DCT1D_inpcnt_reg(0),
      ADR2 => VCC,
      ADR3 => U_DCT1D_inpcnt_reg(2),
      O => U_DCT1D_rtlc2n293_G
    );
  U_DCT1D_ix52393z1324 : X_LUT4
    generic map(
      INIT => X"A5A5"
    )
    port map (
      ADR0 => U_DCT1D_latchbuf_reg_6_Q(7),
      ADR1 => VCC,
      ADR2 => U_DCT1D_latchbuf_reg_1_Q(7),
      ADR3 => VCC,
      O => U_DCT1D_nx52393z1_F
    );
  U_DCT1D_ix7599z1563 : X_LUT4
    generic map(
      INIT => X"FF5F"
    )
    port map (
      ADR0 => U_DCT1D_ready,
      ADR1 => VCC,
      ADR2 => idv_int,
      ADR3 => U_DCT1D_NOT_rtlcs1,
      O => U_DCT1D_rtlc2n293_F
    );
  U_DCT1D_ix7599z1404 : X_LUT4
    generic map(
      INIT => X"3737"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => U_DCT1D_istate_reg(1),
      ADR2 => U_DCT1D_state_reg(1),
      ADR3 => VCC,
      O => U_DCT1D_rtlc2n468_G
    );
  U_DCT1D_ix7599z13091 : X_LUT4
    generic map(
      INIT => X"50C0"
    )
    port map (
      ADR0 => U_DCT1D_rtlc2n293,
      ADR1 => U_DCT1D_istate_reg(1),
      ADR2 => U_DCT1D_nx7599z1,
      ADR3 => U_DCT1D_istate_reg(0),
      O => U_DCT1D_rtlc2n468_F
    );
  U_DCT2D_modgen_counter_colram_reg_reg_q_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_colram_reg_3_DYMUX,
      CE => U_DCT2D_colram_reg_3_CEINV,
      CLK => U_DCT2D_colram_reg_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_colram_reg_3_FFY_RST,
      O => U_DCT2D_colram_reg(3)
    );
  U_DCT2D_colram_reg_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_colram_reg_3_FFY_RSTAND,
      I1 => GSR,
      O => U_DCT2D_colram_reg_3_FFY_RST
    );
  U_DCT2D_colram_reg_3_FFY_RSTAND_7791 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => U_DCT2D_colram_reg_3_FFY_RSTAND
    );
  U_DCT1D_ix15104z1569 : X_LUT4
    generic map(
      INIT => X"FFFC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latch_done_reg,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_state_reg(1),
      O => U_DCT1D_rtlc5n1558_G
    );
  U_DCT1D_ix60980z1320 : X_LUT4
    generic map(
      INIT => X"000C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_latch_done_reg,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_state_reg(1),
      O => U_DCT1D_rtlc5n1558_F
    );
  U_DCT2D_reg_romeaddro5_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro5_s_3_DYMUX,
      CE => rome2addro5_s_3_CEINV,
      CLK => rome2addro5_s_3_CLKINV,
      SET => GND,
      RST => rome2addro5_s_3_FFY_RST,
      O => rome2addro5_s(2)
    );
  rome2addro5_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro5_s_3_SRINV,
      I1 => GSR,
      O => rome2addro5_s_3_FFY_RST
    );
  U_DCT2D_reg_romeaddro5_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro5_s_3_DXMUX,
      CE => rome2addro5_s_3_CEINV,
      CLK => rome2addro5_s_3_CLKINV,
      SET => GND,
      RST => rome2addro5_s_3_FFX_RST,
      O => rome2addro5_s(3)
    );
  rome2addro5_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro5_s_3_SRINV,
      I1 => GSR,
      O => rome2addro5_s_3_FFX_RST
    );
  U_DCT2D_reg_romeaddro6_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro6_s_1_DYMUX,
      CE => rome2addro6_s_1_CEINV,
      CLK => rome2addro6_s_1_CLKINV,
      SET => GND,
      RST => rome2addro6_s_1_FFY_RST,
      O => rome2addro6_s(0)
    );
  rome2addro6_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro6_s_1_SRINV,
      I1 => GSR,
      O => rome2addro6_s_1_FFY_RST
    );
  U_DCT2D_reg_romeaddro6_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro6_s_1_DXMUX,
      CE => rome2addro6_s_1_CEINV,
      CLK => rome2addro6_s_1_CLKINV,
      SET => GND,
      RST => rome2addro6_s_1_FFX_RST,
      O => rome2addro6_s(1)
    );
  rome2addro6_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro6_s_1_SRINV,
      I1 => GSR,
      O => rome2addro6_s_1_FFX_RST
    );
  U_DCT2D_reg_romeaddro6_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro6_s_3_DYMUX,
      CE => rome2addro6_s_3_CEINV,
      CLK => rome2addro6_s_3_CLKINV,
      SET => GND,
      RST => rome2addro6_s_3_FFY_RST,
      O => rome2addro6_s(2)
    );
  rome2addro6_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro6_s_3_SRINV,
      I1 => GSR,
      O => rome2addro6_s_3_FFY_RST
    );
  U_DCT2D_reg_romeaddro6_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro6_s_3_DXMUX,
      CE => rome2addro6_s_3_CEINV,
      CLK => rome2addro6_s_3_CLKINV,
      SET => GND,
      RST => rome2addro6_s_3_FFX_RST,
      O => rome2addro6_s(3)
    );
  rome2addro6_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro6_s_3_SRINV,
      I1 => GSR,
      O => rome2addro6_s_3_FFX_RST
    );
  U_DCT2D_reg_romeaddro7_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro7_s_1_DYMUX,
      CE => rome2addro7_s_1_CEINV,
      CLK => rome2addro7_s_1_CLKINV,
      SET => GND,
      RST => rome2addro7_s_1_FFY_RST,
      O => rome2addro7_s(0)
    );
  rome2addro7_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro7_s_1_SRINV,
      I1 => GSR,
      O => rome2addro7_s_1_FFY_RST
    );
  U_DCT2D_reg_romeaddro2_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro2_s_3_DYMUX,
      CE => rome2addro2_s_3_CEINV,
      CLK => rome2addro2_s_3_CLKINV,
      SET => GND,
      RST => rome2addro2_s_3_FFY_RST,
      O => rome2addro2_s(2)
    );
  rome2addro2_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro2_s_3_SRINV,
      I1 => GSR,
      O => rome2addro2_s_3_FFY_RST
    );
  U_DCT2D_reg_romeaddro2_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro2_s_3_DXMUX,
      CE => rome2addro2_s_3_CEINV,
      CLK => rome2addro2_s_3_CLKINV,
      SET => GND,
      RST => rome2addro2_s_3_FFX_RST,
      O => rome2addro2_s(3)
    );
  rome2addro2_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro2_s_3_SRINV,
      I1 => GSR,
      O => rome2addro2_s_3_FFX_RST
    );
  U_DCT2D_reg_romeaddro3_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro3_s_1_DYMUX,
      CE => rome2addro3_s_1_CEINV,
      CLK => rome2addro3_s_1_CLKINV,
      SET => GND,
      RST => rome2addro3_s_1_FFY_RST,
      O => rome2addro3_s(0)
    );
  rome2addro3_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro3_s_1_SRINV,
      I1 => GSR,
      O => rome2addro3_s_1_FFY_RST
    );
  U_DCT2D_reg_romeaddro3_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro3_s_1_DXMUX,
      CE => rome2addro3_s_1_CEINV,
      CLK => rome2addro3_s_1_CLKINV,
      SET => GND,
      RST => rome2addro3_s_1_FFX_RST,
      O => rome2addro3_s(1)
    );
  rome2addro3_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro3_s_1_SRINV,
      I1 => GSR,
      O => rome2addro3_s_1_FFX_RST
    );
  U_DCT2D_reg_romeaddro3_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro3_s_3_DYMUX,
      CE => rome2addro3_s_3_CEINV,
      CLK => rome2addro3_s_3_CLKINV,
      SET => GND,
      RST => rome2addro3_s_3_FFY_RST,
      O => rome2addro3_s(2)
    );
  rome2addro3_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro3_s_3_SRINV,
      I1 => GSR,
      O => rome2addro3_s_3_FFY_RST
    );
  U_DCT2D_reg_romeaddro3_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro3_s_3_DXMUX,
      CE => rome2addro3_s_3_CEINV,
      CLK => rome2addro3_s_3_CLKINV,
      SET => GND,
      RST => rome2addro3_s_3_FFX_RST,
      O => rome2addro3_s(3)
    );
  rome2addro3_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro3_s_3_SRINV,
      I1 => GSR,
      O => rome2addro3_s_3_FFX_RST
    );
  U_DCT2D_reg_romeaddro7_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro7_s_1_DXMUX,
      CE => rome2addro7_s_1_CEINV,
      CLK => rome2addro7_s_1_CLKINV,
      SET => GND,
      RST => rome2addro7_s_1_FFX_RST,
      O => rome2addro7_s(1)
    );
  rome2addro7_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro7_s_1_SRINV,
      I1 => GSR,
      O => rome2addro7_s_1_FFX_RST
    );
  U_DCT2D_reg_romeaddro7_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro7_s_3_DYMUX,
      CE => rome2addro7_s_3_CEINV,
      CLK => rome2addro7_s_3_CLKINV,
      SET => GND,
      RST => rome2addro7_s_3_FFY_RST,
      O => rome2addro7_s(2)
    );
  rome2addro7_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro7_s_3_SRINV,
      I1 => GSR,
      O => rome2addro7_s_3_FFY_RST
    );
  U_DCT2D_reg_romeaddro7_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro7_s_3_DXMUX,
      CE => rome2addro7_s_3_CEINV,
      CLK => rome2addro7_s_3_CLKINV,
      SET => GND,
      RST => rome2addro7_s_3_FFX_RST,
      O => rome2addro7_s(3)
    );
  rome2addro7_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro7_s_3_SRINV,
      I1 => GSR,
      O => rome2addro7_s_3_FFX_RST
    );
  U_DCT2D_reg_romeaddro8_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro8_s_1_DYMUX,
      CE => rome2addro8_s_1_CEINV,
      CLK => rome2addro8_s_1_CLKINV,
      SET => GND,
      RST => rome2addro8_s_1_FFY_RST,
      O => rome2addro8_s(0)
    );
  rome2addro8_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro8_s_1_SRINV,
      I1 => GSR,
      O => rome2addro8_s_1_FFY_RST
    );
  U_DCT2D_reg_romeaddro8_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro8_s_1_DXMUX,
      CE => rome2addro8_s_1_CEINV,
      CLK => rome2addro8_s_1_CLKINV,
      SET => GND,
      RST => rome2addro8_s_1_FFX_RST,
      O => rome2addro8_s(1)
    );
  rome2addro8_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro8_s_1_SRINV,
      I1 => GSR,
      O => rome2addro8_s_1_FFX_RST
    );
  U_DCT2D_reg_romeaddro8_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro8_s_3_DYMUX,
      CE => rome2addro8_s_3_CEINV,
      CLK => rome2addro8_s_3_CLKINV,
      SET => GND,
      RST => rome2addro8_s_3_FFY_RST,
      O => rome2addro8_s(2)
    );
  rome2addro8_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro8_s_3_SRINV,
      I1 => GSR,
      O => rome2addro8_s_3_FFY_RST
    );
  U_DCT2D_reg_romeaddro8_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro8_s_3_DXMUX,
      CE => rome2addro8_s_3_CEINV,
      CLK => rome2addro8_s_3_CLKINV,
      SET => GND,
      RST => rome2addro8_s_3_FFX_RST,
      O => rome2addro8_s(3)
    );
  rome2addro8_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro8_s_3_SRINV,
      I1 => GSR,
      O => rome2addro8_s_3_FFX_RST
    );
  U_DCT2D_reg_romeaddro9_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro9_s_1_DYMUX,
      CE => rome2addro9_s_1_CEINV,
      CLK => rome2addro9_s_1_CLKINV,
      SET => GND,
      RST => rome2addro9_s_1_FFY_RST,
      O => rome2addro9_s(0)
    );
  rome2addro9_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro9_s_1_SRINV,
      I1 => GSR,
      O => rome2addro9_s_1_FFY_RST
    );
  U_DCT2D_reg_romeaddro9_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro9_s_1_DXMUX,
      CE => rome2addro9_s_1_CEINV,
      CLK => rome2addro9_s_1_CLKINV,
      SET => GND,
      RST => rome2addro9_s_1_FFX_RST,
      O => rome2addro9_s(1)
    );
  rome2addro9_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro9_s_1_SRINV,
      I1 => GSR,
      O => rome2addro9_s_1_FFX_RST
    );
  U_DCT2D_reg_romeaddro9_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro9_s_3_DYMUX,
      CE => rome2addro9_s_3_CEINV,
      CLK => rome2addro9_s_3_CLKINV,
      SET => GND,
      RST => rome2addro9_s_3_FFY_RST,
      O => rome2addro9_s(2)
    );
  rome2addro9_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => rome2addro9_s_3_SRINV,
      I1 => GSR,
      O => rome2addro9_s_3_FFY_RST
    );
  U_DCT1D_ix2819z17955 : X_LUT4
    generic map(
      INIT => X"08FF"
    )
    port map (
      ADR0 => U_DCT1D_rtlc2n293,
      ADR1 => U_DCT1D_istate_reg(0),
      ADR2 => reqwrfail_s,
      ADR3 => U_DCT1D_nx7599z1,
      O => U_DCT1D_rtlc2n471_G
    );
  U_DCT2D_reg_romeaddro9_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => rome2addro9_s_3_DXMUX,
      CE => rome2addro9_s_3_CEINV,
      CLK => rome2addro9_s_3_CLKINV,
      SET => GND,
      RST => rome2addro9_s_3_FFX_RST,
      O => rome2addro9_s(3)
    );
  rome2addro9_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => rome2addro9_s_3_SRINV,
      I1 => GSR,
      O => rome2addro9_s_3_FFX_RST
    );
  U_DCT1D_ix2819z1569 : X_LUT4
    generic map(
      INIT => X"00FE"
    )
    port map (
      ADR0 => U_DCT1D_istate_reg(0),
      ADR1 => U_DCT1D_istate_reg(1),
      ADR2 => requestwr_s,
      ADR3 => U_DCT1D_nx2819z1,
      O => U_DCT1D_rtlc2n471_F
    );
  U_DCT2D_reg_latchbuf_reg_1_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_3_DYMUX,
      CE => U_DCT2D_latchbuf_reg_1_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_1_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_1_3_FFY_RST,
      O => U_DCT2D_latchbuf_reg_1_2_Q
    );
  U_DCT2D_latchbuf_reg_1_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_1_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_1_3_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_1_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_3_DXMUX,
      CE => U_DCT2D_latchbuf_reg_1_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_1_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_1_3_FFX_RST,
      O => U_DCT2D_latchbuf_reg_1_3_Q
    );
  U_DCT2D_latchbuf_reg_1_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_1_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_1_3_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_1_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_5_DYMUX,
      CE => U_DCT2D_latchbuf_reg_1_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_1_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_1_5_FFY_RST,
      O => U_DCT2D_latchbuf_reg_1_4_Q
    );
  U_DCT2D_latchbuf_reg_1_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_1_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_1_5_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_1_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_5_DXMUX,
      CE => U_DCT2D_latchbuf_reg_1_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_1_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_1_5_FFX_RST,
      O => U_DCT2D_latchbuf_reg_1_5_Q
    );
  U_DCT2D_latchbuf_reg_1_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_1_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_1_5_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_1_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_7_DYMUX,
      CE => U_DCT2D_latchbuf_reg_1_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_1_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_1_7_FFY_RST,
      O => U_DCT2D_latchbuf_reg_1_6_Q
    );
  U_DCT2D_latchbuf_reg_1_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_1_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_1_7_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_1_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_7_DXMUX,
      CE => U_DCT2D_latchbuf_reg_1_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_1_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_1_7_FFX_RST,
      O => U_DCT2D_latchbuf_reg_1_7_Q
    );
  U_DCT2D_latchbuf_reg_1_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_1_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_1_7_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_1_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_10_DYMUX,
      CE => U_DCT2D_latchbuf_reg_1_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_1_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_1_10_FFY_RST,
      O => U_DCT2D_latchbuf_reg_1_8_Q
    );
  U_DCT2D_latchbuf_reg_1_10_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_1_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_1_10_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_0_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_1_DYMUX,
      CE => U_DCT2D_latchbuf_reg_0_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_0_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_0_1_FFY_RST,
      O => U_DCT2D_latchbuf_reg_0_0_Q
    );
  U_DCT2D_latchbuf_reg_0_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_0_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_0_1_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_0_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_1_DXMUX,
      CE => U_DCT2D_latchbuf_reg_0_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_0_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_0_1_FFX_RST,
      O => U_DCT2D_latchbuf_reg_0_1_Q
    );
  U_DCT2D_latchbuf_reg_0_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_0_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_0_1_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_0_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_3_DYMUX,
      CE => U_DCT2D_latchbuf_reg_0_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_0_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_0_3_FFY_RST,
      O => U_DCT2D_latchbuf_reg_0_2_Q
    );
  U_DCT2D_latchbuf_reg_0_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_0_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_0_3_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_0_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_3_DXMUX,
      CE => U_DCT2D_latchbuf_reg_0_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_0_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_0_3_FFX_RST,
      O => U_DCT2D_latchbuf_reg_0_3_Q
    );
  U_DCT2D_latchbuf_reg_0_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_0_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_0_3_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_0_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_5_DYMUX,
      CE => U_DCT2D_latchbuf_reg_0_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_0_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_0_5_FFY_RST,
      O => U_DCT2D_latchbuf_reg_0_4_Q
    );
  U_DCT2D_latchbuf_reg_0_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_0_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_0_5_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_0_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_5_DXMUX,
      CE => U_DCT2D_latchbuf_reg_0_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_0_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_0_5_FFX_RST,
      O => U_DCT2D_latchbuf_reg_0_5_Q
    );
  U_DCT2D_latchbuf_reg_0_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_0_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_0_5_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_0_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_7_DYMUX,
      CE => U_DCT2D_latchbuf_reg_0_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_0_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_0_7_FFY_RST,
      O => U_DCT2D_latchbuf_reg_0_6_Q
    );
  U_DCT2D_latchbuf_reg_0_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_0_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_0_7_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_0_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_7_DXMUX,
      CE => U_DCT2D_latchbuf_reg_0_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_0_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_0_7_FFX_RST,
      O => U_DCT2D_latchbuf_reg_0_7_Q
    );
  U_DCT2D_latchbuf_reg_0_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_0_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_0_7_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_0_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_10_DYMUX,
      CE => U_DCT2D_latchbuf_reg_0_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_0_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_0_10_FFY_RST,
      O => U_DCT2D_latchbuf_reg_0_8_Q
    );
  U_DCT2D_latchbuf_reg_0_10_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_0_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_0_10_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_0_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_0_10_DXMUX,
      CE => U_DCT2D_latchbuf_reg_0_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_0_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_0_10_FFX_RST,
      O => U_DCT2D_latchbuf_reg_0_10_Q
    );
  U_DCT2D_latchbuf_reg_0_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_0_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_0_10_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_1_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_1_DYMUX,
      CE => U_DCT2D_latchbuf_reg_1_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_1_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_1_1_FFY_RST,
      O => U_DCT2D_latchbuf_reg_1_0_Q
    );
  U_DCT2D_latchbuf_reg_1_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_1_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_1_1_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_1_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_1_DXMUX,
      CE => U_DCT2D_latchbuf_reg_1_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_1_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_1_1_FFX_RST,
      O => U_DCT2D_latchbuf_reg_1_1_Q
    );
  U_DCT2D_latchbuf_reg_1_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_1_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_1_1_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_2_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_5_DXMUX,
      CE => U_DCT2D_latchbuf_reg_2_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_2_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_2_5_FFX_RST,
      O => U_DCT2D_latchbuf_reg_2_5_Q
    );
  U_DCT2D_latchbuf_reg_2_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_2_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_2_5_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_2_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_7_DYMUX,
      CE => U_DCT2D_latchbuf_reg_2_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_2_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_2_7_FFY_RST,
      O => U_DCT2D_latchbuf_reg_2_6_Q
    );
  U_DCT2D_latchbuf_reg_2_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_2_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_2_7_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_2_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_7_DXMUX,
      CE => U_DCT2D_latchbuf_reg_2_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_2_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_2_7_FFX_RST,
      O => U_DCT2D_latchbuf_reg_2_7_Q
    );
  U_DCT2D_latchbuf_reg_2_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_2_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_2_7_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_2_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_10_DYMUX,
      CE => U_DCT2D_latchbuf_reg_2_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_2_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_2_10_FFY_RST,
      O => U_DCT2D_latchbuf_reg_2_8_Q
    );
  U_DCT2D_latchbuf_reg_2_10_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_2_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_2_10_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_2_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_10_DXMUX,
      CE => U_DCT2D_latchbuf_reg_2_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_2_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_2_10_FFX_RST,
      O => U_DCT2D_latchbuf_reg_2_10_Q
    );
  U_DCT2D_latchbuf_reg_2_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_2_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_2_10_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_3_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_1_DYMUX,
      CE => U_DCT2D_latchbuf_reg_3_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_3_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_3_1_FFY_RST,
      O => U_DCT2D_latchbuf_reg_3_0_Q
    );
  U_DCT2D_latchbuf_reg_3_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_3_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_3_1_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_1_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_1_10_DXMUX,
      CE => U_DCT2D_latchbuf_reg_1_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_1_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_1_10_FFX_RST,
      O => U_DCT2D_latchbuf_reg_1_10_Q
    );
  U_DCT2D_latchbuf_reg_1_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_1_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_1_10_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_2_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_1_DYMUX,
      CE => U_DCT2D_latchbuf_reg_2_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_2_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_2_1_FFY_RST,
      O => U_DCT2D_latchbuf_reg_2_0_Q
    );
  U_DCT2D_latchbuf_reg_2_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_2_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_2_1_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_2_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_1_DXMUX,
      CE => U_DCT2D_latchbuf_reg_2_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_2_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_2_1_FFX_RST,
      O => U_DCT2D_latchbuf_reg_2_1_Q
    );
  U_DCT2D_latchbuf_reg_2_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_2_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_2_1_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_2_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_3_DYMUX,
      CE => U_DCT2D_latchbuf_reg_2_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_2_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_2_3_FFY_RST,
      O => U_DCT2D_latchbuf_reg_2_2_Q
    );
  U_DCT2D_latchbuf_reg_2_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_2_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_2_3_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_2_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_3_DXMUX,
      CE => U_DCT2D_latchbuf_reg_2_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_2_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_2_3_FFX_RST,
      O => U_DCT2D_latchbuf_reg_2_3_Q
    );
  U_DCT2D_latchbuf_reg_2_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_2_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_2_3_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_2_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_2_5_DYMUX,
      CE => U_DCT2D_latchbuf_reg_2_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_2_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_2_5_FFY_RST,
      O => U_DCT2D_latchbuf_reg_2_4_Q
    );
  U_DCT2D_latchbuf_reg_2_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_2_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_2_5_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_5_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_7_DYMUX,
      CE => U_DCT2D_latchbuf_reg_5_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_5_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_5_7_FFY_RST,
      O => U_DCT2D_latchbuf_reg_5_6_Q
    );
  U_DCT2D_latchbuf_reg_5_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_5_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_5_7_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_5_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_7_DXMUX,
      CE => U_DCT2D_latchbuf_reg_5_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_5_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_5_7_FFX_RST,
      O => U_DCT2D_latchbuf_reg_5_7_Q
    );
  U_DCT2D_latchbuf_reg_5_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_5_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_5_7_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_5_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_10_DYMUX,
      CE => U_DCT2D_latchbuf_reg_5_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_5_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_5_10_FFY_RST,
      O => U_DCT2D_latchbuf_reg_5_8_Q
    );
  U_DCT2D_latchbuf_reg_5_10_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_5_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_5_10_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_5_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_5_10_DXMUX,
      CE => U_DCT2D_latchbuf_reg_5_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_5_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_5_10_FFX_RST,
      O => U_DCT2D_latchbuf_reg_5_10_Q
    );
  U_DCT2D_latchbuf_reg_5_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_5_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_5_10_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_6_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_1_DYMUX,
      CE => U_DCT2D_latchbuf_reg_6_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_6_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_6_1_FFY_RST,
      O => U_DCT2D_latchbuf_reg_6_0_Q
    );
  U_DCT2D_latchbuf_reg_6_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_6_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_6_1_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_6_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_1_DXMUX,
      CE => U_DCT2D_latchbuf_reg_6_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_6_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_6_1_FFX_RST,
      O => U_DCT2D_latchbuf_reg_6_1_Q
    );
  U_DCT2D_latchbuf_reg_6_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_6_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_6_1_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_3_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_1_DXMUX,
      CE => U_DCT2D_latchbuf_reg_3_1_CEINV,
      CLK => U_DCT2D_latchbuf_reg_3_1_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_3_1_FFX_RST,
      O => U_DCT2D_latchbuf_reg_3_1_Q
    );
  U_DCT2D_latchbuf_reg_3_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_3_1_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_3_1_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_3_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_3_DYMUX,
      CE => U_DCT2D_latchbuf_reg_3_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_3_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_3_3_FFY_RST,
      O => U_DCT2D_latchbuf_reg_3_2_Q
    );
  U_DCT2D_latchbuf_reg_3_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_3_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_3_3_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_3_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_3_DXMUX,
      CE => U_DCT2D_latchbuf_reg_3_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_3_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_3_3_FFX_RST,
      O => U_DCT2D_latchbuf_reg_3_3_Q
    );
  U_DCT2D_latchbuf_reg_3_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_3_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_3_3_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_3_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_5_DYMUX,
      CE => U_DCT2D_latchbuf_reg_3_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_3_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_3_5_FFY_RST,
      O => U_DCT2D_latchbuf_reg_3_4_Q
    );
  U_DCT2D_latchbuf_reg_3_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_3_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_3_5_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_3_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_5_DXMUX,
      CE => U_DCT2D_latchbuf_reg_3_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_3_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_3_5_FFX_RST,
      O => U_DCT2D_latchbuf_reg_3_5_Q
    );
  U_DCT2D_latchbuf_reg_3_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_3_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_3_5_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_3_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_3_7_DYMUX,
      CE => U_DCT2D_latchbuf_reg_3_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_3_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_3_7_FFY_RST,
      O => U_DCT2D_latchbuf_reg_3_6_Q
    );
  U_DCT2D_latchbuf_reg_3_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_3_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_3_7_FFY_RST
    );
  U_DCT1D_ix59700z1986 : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => romedatao4_s(3),
      ADR1 => U_DCT1D_rtlc5n1346(7),
      ADR2 => VCC,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z333_F
    );
  U_DCT1D_ix59700z1895 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => U_DCT1D_rtlc5n1354(4),
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1348(4),
      O => U_DCT1D_nx59700z251_F
    );
  U_DCT1D_ix59700z49979 : X_LUT4
    generic map(
      INIT => X"BE14"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => U_DCT1D_rtlc5n1355(17),
      ADR2 => U_DCT1D_rtlc5n1354(15),
      ADR3 => U_DCT1D_rtlc5n1348(18),
      O => U_DCT1D_nx59700z218_G
    );
  U_DCT1D_ix59700z1830 : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1348(15),
      ADR1 => VCC,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_rtlc5n1354(15),
      O => U_DCT1D_nx59700z218_F
    );
  U_DCT1D_ix59700z2021 : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => romedatao6_s(7),
      ADR1 => romodatao6_s(7),
      ADR2 => VCC,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z357_F
    );
  U_DCT1D_ix59700z2012 : X_LUT4
    generic map(
      INIT => X"CFC0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao6_s(10),
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => romedatao6_s(10),
      O => U_DCT1D_nx59700z348_F
    );
  U_DCT1D_ix59700z2030 : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => romodatao6_s(4),
      ADR1 => VCC,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => romedatao6_s(4),
      O => U_DCT1D_nx59700z366_F
    );
  U_DCT1D_ix59700z2006 : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => romedatao6_s(12),
      ADR1 => romodatao6_s(12),
      ADR2 => VCC,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z342_F
    );
  U_DCT1D_ix59700z2015 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => romedatao6_s(9),
      ADR2 => VCC,
      ADR3 => romodatao6_s(9),
      O => U_DCT1D_nx59700z351_F
    );
  U_DCT1D_ix59700z2024 : X_LUT4
    generic map(
      INIT => X"AAF0"
    )
    port map (
      ADR0 => romodatao6_s(6),
      ADR1 => VCC,
      ADR2 => romedatao6_s(6),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z360_F
    );
  U_DCT1D_ix59700z1966 : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => romedatao4_s(8),
      ADR1 => U_DCT1D_rtlc5n1346(12),
      ADR2 => VCC,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z318_G
    );
  U_DCT1D_ix59700z1958 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => VCC,
      ADR2 => romedatao4_s(10),
      ADR3 => U_DCT1D_rtlc5n1346(14),
      O => U_DCT1D_nx59700z312_G
    );
  U_DCT1D_ix59700z1978 : X_LUT4
    generic map(
      INIT => X"CCF0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_rtlc5n1346(9),
      ADR2 => romedatao4_s(5),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z327_G
    );
  U_DCT1D_ix59700z1999 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => VCC,
      ADR2 => romedatao6_s(13),
      ADR3 => romodatao6_s(13),
      O => U_DCT1D_nx59700z334_G
    );
  U_DCT1D_ix59700z23954 : X_LUT4
    generic map(
      INIT => X"3C5A"
    )
    port map (
      ADR0 => romedatao7_s(13),
      ADR1 => romodatao7_s(13),
      ADR2 => U_DCT1D_nx59700z335,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z334_F
    );
  U_DCT2D_reg_releaserd_reg : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => releaserd_s_DYMUX,
      CE => releaserd_s_CEINV,
      CLK => releaserd_s_CLKINV,
      SET => GND,
      RST => releaserd_s_FFY_RST,
      O => releaserd_s
    );
  releaserd_s_FFY_RSTOR : X_OR2
    port map (
      I0 => releaserd_s_FFY_RSTAND,
      I1 => GSR,
      O => releaserd_s_FFY_RST
    );
  releaserd_s_FFY_RSTAND_7792 : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_int,
      O => releaserd_s_FFY_RSTAND
    );
  U_DCT1D_reg_romoaddro0_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro0_s_1_DYMUX,
      CE => romoaddro0_s_1_CEINV,
      CLK => romoaddro0_s_1_CLKINV,
      SET => GND,
      RST => romoaddro0_s_1_FFY_RST,
      O => romoaddro0_s(0)
    );
  romoaddro0_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro0_s_1_SRINV,
      I1 => GSR,
      O => romoaddro0_s_1_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_6_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_3_DYMUX,
      CE => U_DCT2D_latchbuf_reg_6_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_6_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_6_3_FFY_RST,
      O => U_DCT2D_latchbuf_reg_6_2_Q
    );
  U_DCT2D_latchbuf_reg_6_3_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_6_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_6_3_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_6_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_3_DXMUX,
      CE => U_DCT2D_latchbuf_reg_6_3_CEINV,
      CLK => U_DCT2D_latchbuf_reg_6_3_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_6_3_FFX_RST,
      O => U_DCT2D_latchbuf_reg_6_3_Q
    );
  U_DCT2D_latchbuf_reg_6_3_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_6_3_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_6_3_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_6_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_5_DYMUX,
      CE => U_DCT2D_latchbuf_reg_6_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_6_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_6_5_FFY_RST,
      O => U_DCT2D_latchbuf_reg_6_4_Q
    );
  U_DCT2D_latchbuf_reg_6_5_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_6_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_6_5_FFY_RST
    );
  U_DCT1D_ix6411z18530 : X_LUT4
    generic map(
      INIT => X"0C22"
    )
    port map (
      ADR0 => U_DCT1D_latch_done_reg,
      ADR1 => U_DCT1D_state_reg(1),
      ADR2 => U_DCT1D_rtlc5n1311,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_rtlc5n1685_G
    );
  U_DCT2D_reg_latchbuf_reg_6_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_5_DXMUX,
      CE => U_DCT2D_latchbuf_reg_6_5_CEINV,
      CLK => U_DCT2D_latchbuf_reg_6_5_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_6_5_FFX_RST,
      O => U_DCT2D_latchbuf_reg_6_5_Q
    );
  U_DCT2D_latchbuf_reg_6_5_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_6_5_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_6_5_FFX_RST
    );
  U_DCT2D_reg_latchbuf_reg_6_6_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_7_DYMUX,
      CE => U_DCT2D_latchbuf_reg_6_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_6_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_6_7_FFY_RST,
      O => U_DCT2D_latchbuf_reg_6_6_Q
    );
  U_DCT2D_latchbuf_reg_6_7_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_6_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_6_7_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_6_7_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_7_DXMUX,
      CE => U_DCT2D_latchbuf_reg_6_7_CEINV,
      CLK => U_DCT2D_latchbuf_reg_6_7_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_6_7_FFX_RST,
      O => U_DCT2D_latchbuf_reg_6_7_Q
    );
  U_DCT2D_latchbuf_reg_6_7_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_6_7_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_6_7_FFX_RST
    );
  U_DCT1D_ix59700z2033 : X_LUT4
    generic map(
      INIT => X"F0CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao6_s(3),
      ADR2 => romodatao6_s(3),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z369_F
    );
  U_DCT1D_ix59700z2009 : X_LUT4
    generic map(
      INIT => X"CCAA"
    )
    port map (
      ADR0 => romedatao6_s(11),
      ADR1 => romodatao6_s(11),
      ADR2 => VCC,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z345_F
    );
  U_DCT1D_ix59700z2018 : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => romodatao6_s(8),
      ADR1 => VCC,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => romedatao6_s(8),
      O => U_DCT1D_nx59700z354_F
    );
  U_DCT1D_ix59700z2027 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => romodatao6_s(5),
      ADR2 => VCC,
      ADR3 => romedatao6_s(5),
      O => U_DCT1D_nx59700z363_F
    );
  U_DCT1D_ix59700z1327 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romedatao3_s(13),
      ADR2 => romedatao2_s(13),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z5_G
    );
  U_DCT1D_ix59700z1416 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1344(15),
      ADR1 => VCC,
      ADR2 => U_DCT1D_rtlc5n1345(17),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z78_G
    );
  U_DCT1D_ix59700z1418 : X_LUT4
    generic map(
      INIT => X"5A5A"
    )
    port map (
      ADR0 => romodatao1_s(13),
      ADR1 => VCC,
      ADR2 => romodatao0_s(13),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z79_G
    );
  U_DCT1D_ix59700z1371 : X_LUT4
    generic map(
      INIT => X"6666"
    )
    port map (
      ADR0 => romedatao1_s(13),
      ADR1 => romedatao0_s(13),
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z42_G
    );
  U_DCT1D_ix59700z1820 : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1348(17),
      ADR1 => U_DCT1D_rtlc5n1354(15),
      ADR2 => VCC,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z215_G
    );
  U_DCT1D_ix59700z1468 : X_LUT4
    generic map(
      INIT => X"3C3C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao3_s(13),
      ADR2 => romodatao2_s(13),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z121_G
    );
  U_DCT1D_ix59700z1890 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => VCC,
      ADR2 => U_DCT1D_rtlc5n1354(5),
      ADR3 => U_DCT1D_rtlc5n1348(5),
      O => U_DCT1D_nx59700z248_G
    );
  U_DCT1D_ix59700z1866 : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1348(9),
      ADR1 => U_DCT1D_rtlc5n1354(9),
      ADR2 => VCC,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z236_G
    );
  U_DCT1D_ix59700z1970 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => VCC,
      ADR2 => romedatao4_s(7),
      ADR3 => U_DCT1D_rtlc5n1346(11),
      O => U_DCT1D_nx59700z321_G
    );
  U_DCT1D_ix59700z1962 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => U_DCT1D_rtlc5n1346(13),
      ADR2 => VCC,
      ADR3 => romedatao4_s(9),
      O => U_DCT1D_nx59700z315_G
    );
  U_DCT1D_ix59700z1954 : X_LUT4
    generic map(
      INIT => X"FA50"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => VCC,
      ADR2 => romedatao4_s(11),
      ADR3 => U_DCT1D_rtlc5n1346(15),
      O => U_DCT1D_nx59700z309_G
    );
  U_DCT1D_ix59700z1884 : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1354(6),
      ADR1 => VCC,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_rtlc5n1348(6),
      O => U_DCT1D_nx59700z245_G
    );
  U_DCT1D_ix59700z1878 : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1354(7),
      ADR1 => VCC,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_rtlc5n1348(7),
      O => U_DCT1D_nx59700z242_G
    );
  U_DCT1D_ix59700z1982 : X_LUT4
    generic map(
      INIT => X"E4E4"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => romedatao4_s(4),
      ADR2 => U_DCT1D_rtlc5n1346(8),
      ADR3 => VCC,
      O => U_DCT1D_nx59700z330_G
    );
  U_DCT1D_ix59700z1974 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => VCC,
      ADR2 => U_DCT1D_rtlc5n1346(10),
      ADR3 => romedatao4_s(6),
      O => U_DCT1D_nx59700z324_G
    );
  U_DCT1D_ix59700z55401 : X_LUT4
    generic map(
      INIT => X"B1E4"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => romedatao5_s(13),
      ADR2 => U_DCT1D_rtlc5n1346(19),
      ADR3 => romedatao4_s(13),
      O => U_DCT1D_nx59700z303_G
    );
  U_DCT2D_reg_latchbuf_reg_6_8_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_10_DYMUX,
      CE => U_DCT2D_latchbuf_reg_6_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_6_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_6_10_FFY_RST,
      O => U_DCT2D_latchbuf_reg_6_8_Q
    );
  U_DCT2D_latchbuf_reg_6_10_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_6_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_6_10_FFY_RST
    );
  U_DCT2D_reg_latchbuf_reg_6_10_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT2D_latchbuf_reg_6_10_DXMUX,
      CE => U_DCT2D_latchbuf_reg_6_10_CEINV,
      CLK => U_DCT2D_latchbuf_reg_6_10_CLKINV,
      SET => GND,
      RST => U_DCT2D_latchbuf_reg_6_10_FFX_RST,
      O => U_DCT2D_latchbuf_reg_6_10_Q
    );
  U_DCT2D_latchbuf_reg_6_10_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT2D_latchbuf_reg_6_10_SRINV,
      I1 => GSR,
      O => U_DCT2D_latchbuf_reg_6_10_FFX_RST
    );
  U_DCT1D_ix59700z1946 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => VCC,
      ADR2 => U_DCT1D_rtlc5n1346(17),
      ADR3 => romedatao4_s(13),
      O => U_DCT1D_nx59700z303_F
    );
  U_DCT1D_ix59700z44668 : X_LUT4
    generic map(
      INIT => X"C693"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => U_DCT1D_rtlc5n1350(21),
      ADR2 => romodatao8_s(13),
      ADR3 => romedatao8_s(13),
      O => U_DCT1D_nx59700z1_G
    );
  U_DCT1D_ix59700z58514 : X_LUT4
    generic map(
      INIT => X"B1E4"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => romedatao2_s(2),
      ADR2 => U_DCT1D_rtlc5n1348(4),
      ADR3 => U_DCT1D_rtlc5n1354(4),
      O => U_DCT1D_nx59700z251_G
    );
  U_DCT1D_ix31471z1320 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_col_reg(2),
      ADR2 => VCC,
      ADR3 => U_DCT1D_col_reg(1),
      O => U_DCT1D_rtlc5n875(2)
    );
  U_DCT1D_reg_col_tmp_reg_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_col_tmp_reg_1_DYMUX,
      CE => U_DCT1D_col_tmp_reg_1_CEINV,
      CLK => U_DCT1D_col_tmp_reg_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_col_tmp_reg_1_FFY_RST,
      O => U_DCT1D_col_tmp_reg(2)
    );
  U_DCT1D_col_tmp_reg_1_FFY_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_col_tmp_reg_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_col_tmp_reg_1_FFY_RST
    );
  U_DCT1D_ix59700z55498 : X_LUT4
    generic map(
      INIT => X"CC5A"
    )
    port map (
      ADR0 => romedatao4_s(3),
      ADR1 => U_DCT1D_rtlc5n1346(7),
      ADR2 => romedatao5_s(2),
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z333_G
    );
  U_DCT1D_reg_col_tmp_reg_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => U_DCT1D_col_tmp_reg_1_DXMUX,
      CE => U_DCT1D_col_tmp_reg_1_CEINV,
      CLK => U_DCT1D_col_tmp_reg_1_CLKINV,
      SET => GND,
      RST => U_DCT1D_col_tmp_reg_1_FFX_RST,
      O => U_DCT1D_col_tmp_reg(1)
    );
  U_DCT1D_col_tmp_reg_1_FFX_RSTOR : X_OR2
    port map (
      I0 => U_DCT1D_col_tmp_reg_1_SRINV,
      I1 => GSR,
      O => U_DCT1D_col_tmp_reg_1_FFX_RST
    );
  U_DCT1D_ix59700z1825 : X_LUT4
    generic map(
      INIT => X"FA0A"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1354(15),
      ADR1 => VCC,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_rtlc5n1348(16),
      O => U_DCT1D_nx59700z215_F
    );
  U_DCT1D_ix59700z1842 : X_LUT4
    generic map(
      INIT => X"AACC"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1348(13),
      ADR1 => U_DCT1D_rtlc5n1354(13),
      ADR2 => VCC,
      ADR3 => U_DCT1D_state_reg(0),
      O => U_DCT1D_nx59700z224_G
    );
  U_DCT1D_ix59700z1860 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => U_DCT1D_rtlc5n1348(10),
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1354(10),
      O => U_DCT1D_nx59700z233_G
    );
  U_DCT1D_ix59700z1836 : X_LUT4
    generic map(
      INIT => X"DD88"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => U_DCT1D_rtlc5n1348(14),
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1354(14),
      O => U_DCT1D_nx59700z221_G
    );
  U_DCT1D_ix59700z1854 : X_LUT4
    generic map(
      INIT => X"AFA0"
    )
    port map (
      ADR0 => U_DCT1D_rtlc5n1348(11),
      ADR1 => VCC,
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_rtlc5n1354(11),
      O => U_DCT1D_nx59700z230_G
    );
  U_DCT1D_ix59700z1950 : X_LUT4
    generic map(
      INIT => X"EE44"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => romedatao4_s(12),
      ADR2 => VCC,
      ADR3 => U_DCT1D_rtlc5n1346(16),
      O => U_DCT1D_nx59700z306_G
    );
  U_DCT1D_ix59700z1942 : X_LUT4
    generic map(
      INIT => X"F5A0"
    )
    port map (
      ADR0 => U_DCT1D_state_reg(0),
      ADR1 => VCC,
      ADR2 => U_DCT1D_rtlc5n1346(18),
      ADR3 => romedatao4_s(13),
      O => U_DCT1D_nx59700z300_G
    );
  U_DCT1D_ix59700z1679 : X_LUT4
    generic map(
      INIT => X"33CC"
    )
    port map (
      ADR0 => VCC,
      ADR1 => romodatao5_s(13),
      ADR2 => VCC,
      ADR3 => romodatao4_s(13),
      O => U_DCT1D_nx59700z255_G
    );
  U_DCT1D_ix59700z1872 : X_LUT4
    generic map(
      INIT => X"FC0C"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_rtlc5n1354(8),
      ADR2 => U_DCT1D_state_reg(0),
      ADR3 => U_DCT1D_rtlc5n1348(8),
      O => U_DCT1D_nx59700z239_G
    );
  U_DCT1D_ix59700z1848 : X_LUT4
    generic map(
      INIT => X"FC30"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_state_reg(0),
      ADR2 => U_DCT1D_rtlc5n1354(12),
      ADR3 => U_DCT1D_rtlc5n1348(12),
      O => U_DCT1D_nx59700z227_G
    );
  U_DCT1D_reg_romoaddro0_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro0_s_1_DXMUX,
      CE => romoaddro0_s_1_CEINV,
      CLK => romoaddro0_s_1_CLKINV,
      SET => GND,
      RST => romoaddro0_s_1_FFX_RST,
      O => romoaddro0_s(1)
    );
  romoaddro0_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro0_s_1_SRINV,
      I1 => GSR,
      O => romoaddro0_s_1_FFX_RST
    );
  U_DCT1D_reg_romoaddro0_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro0_s_3_DYMUX,
      CE => romoaddro0_s_3_CEINV,
      CLK => romoaddro0_s_3_CLKINV,
      SET => GND,
      RST => romoaddro0_s_3_FFY_RST,
      O => romoaddro0_s(2)
    );
  romoaddro0_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro0_s_3_SRINV,
      I1 => GSR,
      O => romoaddro0_s_3_FFY_RST
    );
  U_DCT1D_reg_romoaddro0_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro0_s_3_DXMUX,
      CE => romoaddro0_s_3_CEINV,
      CLK => romoaddro0_s_3_CLKINV,
      SET => GND,
      RST => romoaddro0_s_3_FFX_RST,
      O => romoaddro0_s(3)
    );
  romoaddro0_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro0_s_3_SRINV,
      I1 => GSR,
      O => romoaddro0_s_3_FFX_RST
    );
  U_DCT1D_reg_romoaddro1_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro1_s_1_DYMUX,
      CE => romoaddro1_s_1_CEINV,
      CLK => romoaddro1_s_1_CLKINV,
      SET => GND,
      RST => romoaddro1_s_1_FFY_RST,
      O => romoaddro1_s(0)
    );
  romoaddro1_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro1_s_1_SRINV,
      I1 => GSR,
      O => romoaddro1_s_1_FFY_RST
    );
  U_DCT1D_reg_romoaddro1_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro1_s_1_DXMUX,
      CE => romoaddro1_s_1_CEINV,
      CLK => romoaddro1_s_1_CLKINV,
      SET => GND,
      RST => romoaddro1_s_1_FFX_RST,
      O => romoaddro1_s(1)
    );
  romoaddro1_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro1_s_1_SRINV,
      I1 => GSR,
      O => romoaddro1_s_1_FFX_RST
    );
  U_DCT1D_reg_romoaddro1_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro1_s_3_DYMUX,
      CE => romoaddro1_s_3_CEINV,
      CLK => romoaddro1_s_3_CLKINV,
      SET => GND,
      RST => romoaddro1_s_3_FFY_RST,
      O => romoaddro1_s(2)
    );
  romoaddro1_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro1_s_3_SRINV,
      I1 => GSR,
      O => romoaddro1_s_3_FFY_RST
    );
  U_DCT1D_reg_romoaddro6_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro6_s_3_DYMUX,
      CE => romoaddro6_s_3_CEINV,
      CLK => romoaddro6_s_3_CLKINV,
      SET => GND,
      RST => romoaddro6_s_3_FFY_RST,
      O => romoaddro6_s(2)
    );
  romoaddro6_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro6_s_3_SRINV,
      I1 => GSR,
      O => romoaddro6_s_3_FFY_RST
    );
  U_DCT1D_reg_romoaddro6_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro6_s_3_DXMUX,
      CE => romoaddro6_s_3_CEINV,
      CLK => romoaddro6_s_3_CLKINV,
      SET => GND,
      RST => romoaddro6_s_3_FFX_RST,
      O => romoaddro6_s(3)
    );
  romoaddro6_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro6_s_3_SRINV,
      I1 => GSR,
      O => romoaddro6_s_3_FFX_RST
    );
  U_DCT1D_reg_romoaddro7_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro7_s_1_DYMUX,
      CE => romoaddro7_s_1_CEINV,
      CLK => romoaddro7_s_1_CLKINV,
      SET => GND,
      RST => romoaddro7_s_1_FFY_RST,
      O => romoaddro7_s(0)
    );
  romoaddro7_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro7_s_1_SRINV,
      I1 => GSR,
      O => romoaddro7_s_1_FFY_RST
    );
  U_DCT1D_reg_romoaddro7_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro7_s_1_DXMUX,
      CE => romoaddro7_s_1_CEINV,
      CLK => romoaddro7_s_1_CLKINV,
      SET => GND,
      RST => romoaddro7_s_1_FFX_RST,
      O => romoaddro7_s(1)
    );
  romoaddro7_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro7_s_1_SRINV,
      I1 => GSR,
      O => romoaddro7_s_1_FFX_RST
    );
  U_DCT1D_reg_romoaddro7_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro7_s_3_DYMUX,
      CE => romoaddro7_s_3_CEINV,
      CLK => romoaddro7_s_3_CLKINV,
      SET => GND,
      RST => romoaddro7_s_3_FFY_RST,
      O => romoaddro7_s(2)
    );
  romoaddro7_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro7_s_3_SRINV,
      I1 => GSR,
      O => romoaddro7_s_3_FFY_RST
    );
  U_DCT1D_reg_romoaddro7_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro7_s_3_DXMUX,
      CE => romoaddro7_s_3_CEINV,
      CLK => romoaddro7_s_3_CLKINV,
      SET => GND,
      RST => romoaddro7_s_3_FFX_RST,
      O => romoaddro7_s(3)
    );
  romoaddro7_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro7_s_3_SRINV,
      I1 => GSR,
      O => romoaddro7_s_3_FFX_RST
    );
  U_DCT1D_reg_romoaddro8_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro8_s_1_DYMUX,
      CE => romoaddro8_s_1_CEINV,
      CLK => romoaddro8_s_1_CLKINV,
      SET => GND,
      RST => romoaddro8_s_1_FFY_RST,
      O => romoaddro8_s(0)
    );
  romoaddro8_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro8_s_1_SRINV,
      I1 => GSR,
      O => romoaddro8_s_1_FFY_RST
    );
  U_DCT1D_reg_romoaddro8_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro8_s_1_DXMUX,
      CE => romoaddro8_s_1_CEINV,
      CLK => romoaddro8_s_1_CLKINV,
      SET => GND,
      RST => romoaddro8_s_1_FFX_RST,
      O => romoaddro8_s(1)
    );
  romoaddro8_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro8_s_1_SRINV,
      I1 => GSR,
      O => romoaddro8_s_1_FFX_RST
    );
  U_DCT1D_reg_romoaddro8_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro8_s_3_DYMUX,
      CE => romoaddro8_s_3_CEINV,
      CLK => romoaddro8_s_3_CLKINV,
      SET => GND,
      RST => romoaddro8_s_3_FFY_RST,
      O => romoaddro8_s(2)
    );
  romoaddro8_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro8_s_3_SRINV,
      I1 => GSR,
      O => romoaddro8_s_3_FFY_RST
    );
  U_DCT1D_reg_romoaddro8_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro8_s_3_DXMUX,
      CE => romoaddro8_s_3_CEINV,
      CLK => romoaddro8_s_3_CLKINV,
      SET => GND,
      RST => romoaddro8_s_3_FFX_RST,
      O => romoaddro8_s(3)
    );
  romoaddro8_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro8_s_3_SRINV,
      I1 => GSR,
      O => romoaddro8_s_3_FFX_RST
    );
  U_DCT1D_reg_romoaddro8_4_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro0_s_5_DYMUX,
      CE => romoaddro0_s_5_CEINV,
      CLK => romoaddro0_s_5_CLKINV,
      SET => GND,
      RST => romoaddro0_s_5_FFY_RST,
      O => romoaddro0_s(4)
    );
  romoaddro0_s_5_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro0_s_5_SRINV,
      I1 => GSR,
      O => romoaddro0_s_5_FFY_RST
    );
  U_DCT1D_reg_romoaddro8_5_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro0_s_5_DXMUX,
      CE => romoaddro0_s_5_CEINV,
      CLK => romoaddro0_s_5_CLKINV,
      SET => GND,
      RST => romoaddro0_s_5_FFX_RST,
      O => romoaddro0_s(5)
    );
  romoaddro0_s_5_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro0_s_5_SRINV,
      I1 => GSR,
      O => romoaddro0_s_5_FFX_RST
    );
  U_DCT1D_reg_romoaddro5_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro5_s_1_DYMUX,
      CE => romoaddro5_s_1_CEINV,
      CLK => romoaddro5_s_1_CLKINV,
      SET => GND,
      RST => romoaddro5_s_1_FFY_RST,
      O => romoaddro5_s(0)
    );
  romoaddro5_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro5_s_1_SRINV,
      I1 => GSR,
      O => romoaddro5_s_1_FFY_RST
    );
  U_DCT1D_reg_romoaddro5_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro5_s_1_DXMUX,
      CE => romoaddro5_s_1_CEINV,
      CLK => romoaddro5_s_1_CLKINV,
      SET => GND,
      RST => romoaddro5_s_1_FFX_RST,
      O => romoaddro5_s(1)
    );
  romoaddro5_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro5_s_1_SRINV,
      I1 => GSR,
      O => romoaddro5_s_1_FFX_RST
    );
  U_DCT1D_reg_romoaddro5_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro5_s_3_DYMUX,
      CE => romoaddro5_s_3_CEINV,
      CLK => romoaddro5_s_3_CLKINV,
      SET => GND,
      RST => romoaddro5_s_3_FFY_RST,
      O => romoaddro5_s(2)
    );
  romoaddro5_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro5_s_3_SRINV,
      I1 => GSR,
      O => romoaddro5_s_3_FFY_RST
    );
  U_DCT1D_reg_romoaddro5_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro5_s_3_DXMUX,
      CE => romoaddro5_s_3_CEINV,
      CLK => romoaddro5_s_3_CLKINV,
      SET => GND,
      RST => romoaddro5_s_3_FFX_RST,
      O => romoaddro5_s(3)
    );
  romoaddro5_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro5_s_3_SRINV,
      I1 => GSR,
      O => romoaddro5_s_3_FFX_RST
    );
  U_DCT1D_reg_romoaddro6_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro6_s_1_DYMUX,
      CE => romoaddro6_s_1_CEINV,
      CLK => romoaddro6_s_1_CLKINV,
      SET => GND,
      RST => romoaddro6_s_1_FFY_RST,
      O => romoaddro6_s(0)
    );
  romoaddro6_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro6_s_1_SRINV,
      I1 => GSR,
      O => romoaddro6_s_1_FFY_RST
    );
  U_DCT1D_reg_romoaddro6_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro6_s_1_DXMUX,
      CE => romoaddro6_s_1_CEINV,
      CLK => romoaddro6_s_1_CLKINV,
      SET => GND,
      RST => romoaddro6_s_1_FFX_RST,
      O => romoaddro6_s(1)
    );
  romoaddro6_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro6_s_1_SRINV,
      I1 => GSR,
      O => romoaddro6_s_1_FFX_RST
    );
  U_DCT1D_reg_romoaddro3_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro3_s_3_DYMUX,
      CE => romoaddro3_s_3_CEINV,
      CLK => romoaddro3_s_3_CLKINV,
      SET => GND,
      RST => romoaddro3_s_3_FFY_RST,
      O => romoaddro3_s(2)
    );
  romoaddro3_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro3_s_3_SRINV,
      I1 => GSR,
      O => romoaddro3_s_3_FFY_RST
    );
  U_DCT1D_reg_romoaddro3_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro3_s_3_DXMUX,
      CE => romoaddro3_s_3_CEINV,
      CLK => romoaddro3_s_3_CLKINV,
      SET => GND,
      RST => romoaddro3_s_3_FFX_RST,
      O => romoaddro3_s(3)
    );
  romoaddro3_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro3_s_3_SRINV,
      I1 => GSR,
      O => romoaddro3_s_3_FFX_RST
    );
  U_DCT1D_reg_romoaddro4_0_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro4_s_1_DYMUX,
      CE => romoaddro4_s_1_CEINV,
      CLK => romoaddro4_s_1_CLKINV,
      SET => GND,
      RST => romoaddro4_s_1_FFY_RST,
      O => romoaddro4_s(0)
    );
  romoaddro4_s_1_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro4_s_1_SRINV,
      I1 => GSR,
      O => romoaddro4_s_1_FFY_RST
    );
  U_DCT1D_reg_romoaddro4_1_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro4_s_1_DXMUX,
      CE => romoaddro4_s_1_CEINV,
      CLK => romoaddro4_s_1_CLKINV,
      SET => GND,
      RST => romoaddro4_s_1_FFX_RST,
      O => romoaddro4_s(1)
    );
  romoaddro4_s_1_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro4_s_1_SRINV,
      I1 => GSR,
      O => romoaddro4_s_1_FFX_RST
    );
  U_DCT1D_reg_romoaddro4_2_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro4_s_3_DYMUX,
      CE => romoaddro4_s_3_CEINV,
      CLK => romoaddro4_s_3_CLKINV,
      SET => GND,
      RST => romoaddro4_s_3_FFY_RST,
      O => romoaddro4_s(2)
    );
  romoaddro4_s_3_FFY_RSTOR : X_OR2
    port map (
      I0 => romoaddro4_s_3_SRINV,
      I1 => GSR,
      O => romoaddro4_s_3_FFY_RST
    );
  U_DCT1D_reg_romoaddro4_3_Q : X_FF
    generic map(
      INIT => '0'
    )
    port map (
      I => romoaddro4_s_3_DXMUX,
      CE => romoaddro4_s_3_CEINV,
      CLK => romoaddro4_s_3_CLKINV,
      SET => GND,
      RST => romoaddro4_s_3_FFX_RST,
      O => romoaddro4_s(3)
    );
  romoaddro4_s_3_FFX_RSTOR : X_OR2
    port map (
      I0 => romoaddro4_s_3_SRINV,
      I1 => GSR,
      O => romoaddro4_s_3_FFX_RST
    );
  PWR_VCC_0_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1
    );
  PWR_VCC_1_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_0
    );
  PWR_VCC_2_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_1
    );
  PWR_VCC_3_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_2
    );
  PWR_VCC_4_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_3
    );
  PWR_VCC_5_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_4
    );
  PWR_VCC_6_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_5
    );
  PWR_VCC_7_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_6
    );
  PWR_VCC_8_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_7
    );
  PWR_VCC_9_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_8
    );
  PWR_VCC_10_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_9
    );
  PWR_VCC_11_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_10
    );
  PWR_VCC_12_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_11
    );
  PWR_VCC_13_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_12
    );
  PWR_VCC_14_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_13
    );
  PWR_VCC_15_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_14
    );
  PWR_VCC_16_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_15
    );
  PWR_VCC_17_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_16
    );
  PWR_VCC_18_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_17
    );
  PWR_VCC_19_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_18
    );
  PWR_VCC_20_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_19
    );
  PWR_VCC_21_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_20
    );
  PWR_VCC_22_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_21
    );
  PWR_VCC_23_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_22
    );
  PWR_VCC_24_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_23
    );
  PWR_VCC_25_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_24
    );
  PWR_VCC_26_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_25
    );
  PWR_VCC_27_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_26
    );
  PWR_VCC_28_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_27
    );
  PWR_VCC_29_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_28
    );
  PWR_VCC_30_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_29
    );
  PWR_VCC_31_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_30
    );
  PWR_VCC_32_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_31
    );
  PWR_VCC_33_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_32
    );
  PWR_VCC_34_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_33
    );
  PWR_VCC_35_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_34
    );
  PWR_VCC_36_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_35
    );
  PWR_VCC_37_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_36
    );
  PWR_VCC_38_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_37
    );
  PWR_VCC_39_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_38
    );
  PWR_VCC_40_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_39
    );
  PWR_VCC_41_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_40
    );
  PWR_VCC_42_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_41
    );
  PWR_VCC_43_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_42
    );
  PWR_VCC_44_LOGICAL_ONE : X_ONE
    port map (
      O => GLOBAL_LOGIC1_43
    );
  PWR_GND_0_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => PWR_GND_0_G,
      O => GLOBAL_LOGIC0
    );
  PWR_GND_0_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_0_G
    );
  PWR_GND_1_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => PWR_GND_1_G,
      O => GLOBAL_LOGIC0_0
    );
  PWR_GND_1_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_1_G
    );
  PWR_GND_2_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => PWR_GND_2_G,
      O => GLOBAL_LOGIC0_1
    );
  PWR_GND_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_2_G
    );
  PWR_GND_3_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => PWR_GND_3_G,
      O => GLOBAL_LOGIC0_2
    );
  PWR_GND_3_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_3_G
    );
  PWR_GND_4_YUSED : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => PWR_GND_4_G,
      O => GLOBAL_LOGIC0_3
    );
  PWR_GND_4_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => PWR_GND_4_G
    );
  nx54672z899_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z899_G
    );
  nx54672z820_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z820_G
    );
  nx54672z390_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z390_G
    );
  U_DCT1D_nx59700z428_F_X_LUT4 : X_LUT4
    generic map(
      INIT => X"F0F0"
    )
    port map (
      ADR0 => VCC,
      ADR1 => U_DCT1D_nx59700z333,
      ADR2 => U_DCT1D_nx59700z332,
      ADR3 => VCC,
      O => U_DCT1D_nx59700z428_F
    );
  U_DCT2D_nx65206z570_F_X_LUT4 : X_LUT4
    generic map(
      INIT => X"CCCC"
    )
    port map (
      ADR0 => U_DCT2D_nx65206z251,
      ADR1 => U_DCT2D_nx65206z250,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U_DCT2D_nx65206z570_F
    );
  U_DCT1D_nx59700z493_F_X_LUT4 : X_LUT4
    generic map(
      INIT => X"FF00"
    )
    port map (
      ADR0 => U_DCT1D_nx59700z251,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => U_DCT1D_nx59700z250,
      O => U_DCT1D_nx59700z493_F
    );
  rome2datao5_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rome2datao5_s_2_G
    );
  U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROME5_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx53675z1345_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1345_G
    );
  rome2datao7_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rome2datao7_s_2_G
    );
  U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROME7_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx53675z585_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z585_G
    );
  rome2datao8_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rome2datao8_s_2_G
    );
  U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROME8_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx53675z792_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z792_G
    );
  nx53675z130_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z130_G
    );
  nx53675z1424_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1424_G
    );
  nx53675z650_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z650_G
    );
  nx53675z65_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z65_G
    );
  rome2datao1_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rome2datao1_s_2_G
    );
  U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROME1_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx53675z1_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1_G
    );
  nx53675z871_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z871_G
    );
  rome2datao3_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rome2datao3_s_2_G
    );
  U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROME3_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx53675z195_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z195_G
    );
  rome2datao10_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rome2datao10_s_2_G
    );
  U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROME10_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx53675z325_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z325_G
    );
  rome2datao2_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rome2datao2_s_2_G
    );
  U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROME2_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx53675z390_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z390_G
    );
  rome2datao4_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rome2datao4_s_2_G
    );
  U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROME4_modgen_rom_ix2_nx_ro64_32_u_G
    );
  rome2datao9_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rome2datao9_s_2_G
    );
  U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROME9_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx53675z1503_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1503_G
    );
  nx53675z950_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z950_G
    );
  rome2datao6_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => rome2datao6_s_2_G
    );
  U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U2_ROME6_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx53675z715_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z715_G
    );
  nx53675z1029_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1029_G
    );
  nx53675z455_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z455_G
    );
  nx53675z1108_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1108_G
    );
  nx53675z260_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z260_G
    );
  nx53675z520_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z520_G
    );
  nx53675z1187_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1187_G
    );
  nx53675z1266_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx53675z1266_G
    );
  nx54672z585_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z585_G
    );
  romedatao8_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => romedatao8_s_2_G
    );
  U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U1_ROME8_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx54672z662_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z662_G
    );
  nx54672z130_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z130_G
    );
  nx54672z741_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z741_G
    );
  nx54672z65_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z65_G
    );
  romedatao1_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => romedatao1_s_2_G
    );
  U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U1_ROME1_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx54672z1_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z1_G
    );
  romedatao3_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => romedatao3_s_2_G
    );
  U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U1_ROME3_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx54672z195_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z195_G
    );
  nx54672z325_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z325_G
    );
  romedatao2_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => romedatao2_s_2_G
    );
  U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U1_ROME2_modgen_rom_ix2_nx_ro64_32_u_G
    );
  romedatao4_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => romedatao4_s_2_G
    );
  U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U1_ROME4_modgen_rom_ix2_nx_ro64_32_u_G
    );
  romedatao6_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => romedatao6_s_2_G
    );
  U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U1_ROME6_modgen_rom_ix2_nx_ro64_32_u_G
    );
  romedatao5_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => romedatao5_s_2_G
    );
  U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U1_ROME5_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx54672z978_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z978_G
    );
  romedatao7_s_2_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => romedatao7_s_2_G
    );
  U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => U1_ROME7_modgen_rom_ix2_nx_ro64_32_u_G
    );
  nx54672z455_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z455_G
    );
  nx54672z260_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z260_G
    );
  nx54672z520_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z520_G
    );
  nx54672z1057_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z1057_G
    );
  nx54672z1136_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z1136_G
    );
  nx54672z1215_G_X_LUT4 : X_LUT4
    generic map(
      INIT => X"0000"
    )
    port map (
      ADR0 => VCC,
      ADR1 => VCC,
      ADR2 => VCC,
      ADR3 => VCC,
      O => nx54672z1215_G
    );
  clk_IFF_IMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => clk_INBUF,
      O => clk_ibuf_IBUFG
    );
  idv_IFF_IMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => idv_INBUF,
      O => idv_int
    );
  rst_IFF_IMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => rst_INBUF,
      O => rst_int
    );
  dcti_7_IFF_IMUX : X_BUF_PP
    generic map(
      PATHPULSE => 757 ps
    )
    port map (
      I => dcti_7_INBUF,
      O => dcti_int(7)
    );
  NlwBlock_MDCT_GND : X_ZERO
    port map (
      O => GND
    );
  NlwBlock_MDCT_VCC : X_ONE
    port map (
      O => VCC
    );
  NlwBlockROC : X_ROC
    generic map (ROC_WIDTH => 100 ns)
    port map (O => GSR);
  NlwBlockTOC : X_TOC
    port map (O => GTS);

end STRUCTURE;

