
library IEEE;
use     IEEE.STD_LOGIC_1164.ALL;
use     IEEE.STD_LOGIC_UNSIGNED.all;

use work.AGCPACK.all;

entity agc_erasable is
  port (
    clka  : in  std_logic;
	 wea   : in  std_logic_vector(  0 downto 0 );
	 addra : in  std_logic_vector( 10 downto 0 );
	 dina  : in  std_logic_vector( 15 downto 0 );
	 clkb  : in  std_logic;
	 addrb : in  std_logic_vector( 10 downto 0 );
	 doutb : out std_logic_vector( 15 downto 0 )
  );
end agc_erasable;

architecture Rtl of agc_erasable is

  type t_CORES is array( 0 to 2047 ) of AGCBITARRAY( 15 downto 0 );
  
  signal CORES : t_CORES := (
    "0000000000000001", -- 000000 (00000)  0    0 000000
    "0000000000000001", -- 000000 (00000)  0    1 000001
    "0000000000000001", -- 000000 (00000)  0    2 000002
    "0000000000000001", -- 000000 (00000)  0    3 000003
    "0000000000000001", -- 000000 (00000)  0    4 000004
    "0000000000000001", -- 000000 (00000)  0    5 000005
    "0000000000000001", -- 000000 (00000)  0    6 000006
    "0000000000000001", -- 000000 (00000)  0    7 000007
    "0000000000000001", -- 000000 (00000)  0    8 000010
    "0000000000000001", -- 000000 (00000)  0    9 000011
    "0000000000000001", -- 000000 (00000)  0   10 000012
    "0000000000000001", -- 000000 (00000)  0   11 000013
    "0000000000000001", -- 000000 (00000)  0   12 000014
    "0000000000000001", -- 000000 (00000)  0   13 000015
    "0000000000000001", -- 000000 (00000)  0   14 000016
    "0000000000000001", -- 000000 (00000)  0   15 000017
    "0000000000000001", -- 000000 (00000)  0   16 000020
    "0000000000000001", -- 000000 (00000)  0   17 000021
    "0000000000000001", -- 000000 (00000)  0   18 000022
    "0000000000000001", -- 000000 (00000)  0   19 000023
    "0000000000000001", -- 000000 (00000)  0   20 000024
    "0000000000000001", -- 000000 (00000)  0   21 000025
    "0000000000000001", -- 000000 (00000)  0   22 000026
    "0000000000000001", -- 000000 (00000)  0   23 000027
    "0000000000000001", -- 000000 (00000)  0   24 000030
    "0000000000000001", -- 000000 (00000)  0   25 000031
    "0000000000000001", -- 000000 (00000)  0   26 000032
    "0000000000000001", -- 000000 (00000)  0   27 000033
    "0000000000000001", -- 000000 (00000)  0   28 000034
    "0000000000000001", -- 000000 (00000)  0   29 000035
    "0000000000000001", -- 000000 (00000)  0   30 000036
    "0000000000000001", -- 000000 (00000)  0   31 000037
    "0000000000000001", -- 000000 (00000)  0   32 000040
    "0000000000000001", -- 000000 (00000)  0   33 000041
    "0000000000000001", -- 000000 (00000)  0   34 000042
    "0000000000000001", -- 000000 (00000)  0   35 000043
    "0000000000000001", -- 000000 (00000)  0   36 000044
    "0000000000000001", -- 000000 (00000)  0   37 000045
    "0000000000000001", -- 000000 (00000)  0   38 000046
    "0000000000000001", -- 000000 (00000)  0   39 000047
    "0000000000000001", -- 000000 (00000)  0   40 000050
    "0000000000000001", -- 000000 (00000)  0   41 000051
    "0000000000000001", -- 000000 (00000)  0   42 000052
    "0000000000000001", -- 000000 (00000)  0   43 000053
    "0000000000000001", -- 000000 (00000)  0   44 000054
    "0000000000000001", -- 000000 (00000)  0   45 000055
    "0000000000000001", -- 000000 (00000)  0   46 000056
    "0000000000000001", -- 000000 (00000)  0   47 000057
    "0000000000000001", -- 000000 (00000)  0   48 000060
    "0000000000000001", -- 000000 (00000)  0   49 000061
    "0000000000000001", -- 000000 (00000)  0   50 000062
    "0000000000000001", -- 000000 (00000)  0   51 000063
    "0000000000000001", -- 000000 (00000)  0   52 000064
    "0000000000000001", -- 000000 (00000)  0   53 000065
    "0000000000000001", -- 000000 (00000)  0   54 000066
    "0000000000000001", -- 000000 (00000)  0   55 000067
    "0000000000000001", -- 000000 (00000)  0   56 000070
    "0000000000000001", -- 000000 (00000)  0   57 000071
    "0000000000000001", -- 000000 (00000)  0   58 000072
    "0000000000000001", -- 000000 (00000)  0   59 000073
    "0000000000000001", -- 000000 (00000)  0   60 000074
    "0000000000000001", -- 000000 (00000)  0   61 000075
    "0000000000000001", -- 000000 (00000)  0   62 000076
    "0000000000000001", -- 000000 (00000)  0   63 000077
    "0000000000000001", -- 000000 (00000)  0   64 000100
    "0000000000000001", -- 000000 (00000)  0   65 000101
    "0000000000000001", -- 000000 (00000)  0   66 000102
    "0000000000000001", -- 000000 (00000)  0   67 000103
    "0000000000000001", -- 000000 (00000)  0   68 000104
    "0000000000000001", -- 000000 (00000)  0   69 000105
    "0000000000000001", -- 000000 (00000)  0   70 000106
    "0000000000000001", -- 000000 (00000)  0   71 000107
    "0000000000000001", -- 000000 (00000)  0   72 000110
    "0000000000000001", -- 000000 (00000)  0   73 000111
    "0000000000000001", -- 000000 (00000)  0   74 000112
    "0000000000000001", -- 000000 (00000)  0   75 000113
    "0000000000000001", -- 000000 (00000)  0   76 000114
    "0000000000000001", -- 000000 (00000)  0   77 000115
    "0000000000000001", -- 000000 (00000)  0   78 000116
    "0000000000000001", -- 000000 (00000)  0   79 000117
    "0000000000000001", -- 000000 (00000)  0   80 000120
    "0000000000000001", -- 000000 (00000)  0   81 000121
    "0000000000000001", -- 000000 (00000)  0   82 000122
    "0000000000000001", -- 000000 (00000)  0   83 000123
    "0000000000000001", -- 000000 (00000)  0   84 000124
    "0000000000000001", -- 000000 (00000)  0   85 000125
    "0000000000000001", -- 000000 (00000)  0   86 000126
    "0000000000000001", -- 000000 (00000)  0   87 000127
    "0000000000000001", -- 000000 (00000)  0   88 000130
    "0000000000000001", -- 000000 (00000)  0   89 000131
    "0000000000000001", -- 000000 (00000)  0   90 000132
    "0000000000000001", -- 000000 (00000)  0   91 000133
    "0000000000000001", -- 000000 (00000)  0   92 000134
    "0000000000000001", -- 000000 (00000)  0   93 000135
    "0000000000000001", -- 000000 (00000)  0   94 000136
    "0000000000000001", -- 000000 (00000)  0   95 000137
    "0000000000000001", -- 000000 (00000)  0   96 000140
    "0000000000000001", -- 000000 (00000)  0   97 000141
    "0000000000000001", -- 000000 (00000)  0   98 000142
    "0000000000000001", -- 000000 (00000)  0   99 000143
    "0000000000000001", -- 000000 (00000)  0  100 000144
    "0000000000000001", -- 000000 (00000)  0  101 000145
    "0000000000000001", -- 000000 (00000)  0  102 000146
    "0000000000000001", -- 000000 (00000)  0  103 000147
    "0000000000000001", -- 000000 (00000)  0  104 000150
    "0000000000000001", -- 000000 (00000)  0  105 000151
    "0000000000000001", -- 000000 (00000)  0  106 000152
    "0000000000000001", -- 000000 (00000)  0  107 000153
    "0000000000000001", -- 000000 (00000)  0  108 000154
    "0000000000000001", -- 000000 (00000)  0  109 000155
    "0000000000000001", -- 000000 (00000)  0  110 000156
    "0000000000000001", -- 000000 (00000)  0  111 000157
    "0000000000000001", -- 000000 (00000)  0  112 000160
    "0000000000000001", -- 000000 (00000)  0  113 000161
    "0000000000000001", -- 000000 (00000)  0  114 000162
    "0000000000000001", -- 000000 (00000)  0  115 000163
    "0000000000000001", -- 000000 (00000)  0  116 000164
    "0000000000000001", -- 000000 (00000)  0  117 000165
    "0000000000000001", -- 000000 (00000)  0  118 000166
    "0000000000000001", -- 000000 (00000)  0  119 000167
    "0000000000000001", -- 000000 (00000)  0  120 000170
    "0000000000000001", -- 000000 (00000)  0  121 000171
    "0000000000000001", -- 000000 (00000)  0  122 000172
    "0000000000000001", -- 000000 (00000)  0  123 000173
    "0000000000000001", -- 000000 (00000)  0  124 000174
    "0000000000000001", -- 000000 (00000)  0  125 000175
    "0000000000000001", -- 000000 (00000)  0  126 000176
    "0000000000000001", -- 000000 (00000)  0  127 000177
    "0000000000000001", -- 000000 (00000)  0  128 000200
    "0000000000000001", -- 000000 (00000)  0  129 000201
    "0000000000000001", -- 000000 (00000)  0  130 000202
    "0000000000000001", -- 000000 (00000)  0  131 000203
    "0000000000000001", -- 000000 (00000)  0  132 000204
    "0000000000000001", -- 000000 (00000)  0  133 000205
    "0000000000000001", -- 000000 (00000)  0  134 000206
    "0000000000000001", -- 000000 (00000)  0  135 000207
    "0000000000000001", -- 000000 (00000)  0  136 000210
    "0000000000000001", -- 000000 (00000)  0  137 000211
    "0000000000000001", -- 000000 (00000)  0  138 000212
    "0000000000000001", -- 000000 (00000)  0  139 000213
    "0000000000000001", -- 000000 (00000)  0  140 000214
    "0000000000000001", -- 000000 (00000)  0  141 000215
    "0000000000000001", -- 000000 (00000)  0  142 000216
    "0000000000000001", -- 000000 (00000)  0  143 000217
    "0000000000000001", -- 000000 (00000)  0  144 000220
    "0000000000000001", -- 000000 (00000)  0  145 000221
    "0000000000000001", -- 000000 (00000)  0  146 000222
    "0000000000000001", -- 000000 (00000)  0  147 000223
    "0000000000000001", -- 000000 (00000)  0  148 000224
    "0000000000000001", -- 000000 (00000)  0  149 000225
    "0000000000000001", -- 000000 (00000)  0  150 000226
    "0000000000000001", -- 000000 (00000)  0  151 000227
    "0000000000000001", -- 000000 (00000)  0  152 000230
    "0000000000000001", -- 000000 (00000)  0  153 000231
    "0000000000000001", -- 000000 (00000)  0  154 000232
    "0000000000000001", -- 000000 (00000)  0  155 000233
    "0000000000000001", -- 000000 (00000)  0  156 000234
    "0000000000000001", -- 000000 (00000)  0  157 000235
    "0000000000000001", -- 000000 (00000)  0  158 000236
    "0000000000000001", -- 000000 (00000)  0  159 000237
    "0000000000000001", -- 000000 (00000)  0  160 000240
    "0000000000000001", -- 000000 (00000)  0  161 000241
    "0000000000000001", -- 000000 (00000)  0  162 000242
    "0000000000000001", -- 000000 (00000)  0  163 000243
    "0000000000000001", -- 000000 (00000)  0  164 000244
    "0000000000000001", -- 000000 (00000)  0  165 000245
    "0000000000000001", -- 000000 (00000)  0  166 000246
    "0000000000000001", -- 000000 (00000)  0  167 000247
    "0000000000000001", -- 000000 (00000)  0  168 000250
    "0000000000000001", -- 000000 (00000)  0  169 000251
    "0000000000000001", -- 000000 (00000)  0  170 000252
    "0000000000000001", -- 000000 (00000)  0  171 000253
    "0000000000000001", -- 000000 (00000)  0  172 000254
    "0000000000000001", -- 000000 (00000)  0  173 000255
    "0000000000000001", -- 000000 (00000)  0  174 000256
    "0000000000000001", -- 000000 (00000)  0  175 000257
    "0000000000000001", -- 000000 (00000)  0  176 000260
    "0000000000000001", -- 000000 (00000)  0  177 000261
    "0000000000000001", -- 000000 (00000)  0  178 000262
    "0000000000000001", -- 000000 (00000)  0  179 000263
    "0000000000000001", -- 000000 (00000)  0  180 000264
    "0000000000000001", -- 000000 (00000)  0  181 000265
    "0000000000000001", -- 000000 (00000)  0  182 000266
    "0000000000000001", -- 000000 (00000)  0  183 000267
    "0000000000000001", -- 000000 (00000)  0  184 000270
    "0000000000000001", -- 000000 (00000)  0  185 000271
    "0000000000000001", -- 000000 (00000)  0  186 000272
    "0000000000000001", -- 000000 (00000)  0  187 000273
    "0000000000000001", -- 000000 (00000)  0  188 000274
    "0000000000000001", -- 000000 (00000)  0  189 000275
    "0000000000000001", -- 000000 (00000)  0  190 000276
    "0000000000000001", -- 000000 (00000)  0  191 000277
    "0000000000000001", -- 000000 (00000)  0  192 000300
    "0000000000000001", -- 000000 (00000)  0  193 000301
    "0000000000000001", -- 000000 (00000)  0  194 000302
    "0000000000000001", -- 000000 (00000)  0  195 000303
    "0000000000000001", -- 000000 (00000)  0  196 000304
    "0000000000000001", -- 000000 (00000)  0  197 000305
    "0000000000000001", -- 000000 (00000)  0  198 000306
    "0000000000000001", -- 000000 (00000)  0  199 000307
    "0000000000000001", -- 000000 (00000)  0  200 000310
    "0000000000000001", -- 000000 (00000)  0  201 000311
    "0000000000000001", -- 000000 (00000)  0  202 000312
    "0000000000000001", -- 000000 (00000)  0  203 000313
    "0000000000000001", -- 000000 (00000)  0  204 000314
    "0000000000000001", -- 000000 (00000)  0  205 000315
    "0000000000000001", -- 000000 (00000)  0  206 000316
    "0000000000000001", -- 000000 (00000)  0  207 000317
    "0000000000000001", -- 000000 (00000)  0  208 000320
    "0000000000000001", -- 000000 (00000)  0  209 000321
    "0000000000000001", -- 000000 (00000)  0  210 000322
    "0000000000000001", -- 000000 (00000)  0  211 000323
    "0000000000000001", -- 000000 (00000)  0  212 000324
    "0000000000000001", -- 000000 (00000)  0  213 000325
    "0000000000000001", -- 000000 (00000)  0  214 000326
    "0000000000000001", -- 000000 (00000)  0  215 000327
    "0000000000000001", -- 000000 (00000)  0  216 000330
    "0000000000000001", -- 000000 (00000)  0  217 000331
    "0000000000000001", -- 000000 (00000)  0  218 000332
    "0000000000000001", -- 000000 (00000)  0  219 000333
    "0000000000000001", -- 000000 (00000)  0  220 000334
    "0000000000000001", -- 000000 (00000)  0  221 000335
    "0000000000000001", -- 000000 (00000)  0  222 000336
    "0000000000000001", -- 000000 (00000)  0  223 000337
    "0000000000000001", -- 000000 (00000)  0  224 000340
    "0000000000000001", -- 000000 (00000)  0  225 000341
    "0000000000000001", -- 000000 (00000)  0  226 000342
    "0000000000000001", -- 000000 (00000)  0  227 000343
    "0000000000000001", -- 000000 (00000)  0  228 000344
    "0000000000000001", -- 000000 (00000)  0  229 000345
    "0000000000000001", -- 000000 (00000)  0  230 000346
    "0000000000000001", -- 000000 (00000)  0  231 000347
    "0000000000000001", -- 000000 (00000)  0  232 000350
    "0000000000000001", -- 000000 (00000)  0  233 000351
    "0000000000000001", -- 000000 (00000)  0  234 000352
    "0000000000000001", -- 000000 (00000)  0  235 000353
    "0000000000000001", -- 000000 (00000)  0  236 000354
    "0000000000000001", -- 000000 (00000)  0  237 000355
    "0000000000000001", -- 000000 (00000)  0  238 000356
    "0000000000000001", -- 000000 (00000)  0  239 000357
    "0000000000000001", -- 000000 (00000)  0  240 000360
    "0000000000000001", -- 000000 (00000)  0  241 000361
    "0000000000000001", -- 000000 (00000)  0  242 000362
    "0000000000000001", -- 000000 (00000)  0  243 000363
    "0000000000000001", -- 000000 (00000)  0  244 000364
    "0000000000000001", -- 000000 (00000)  0  245 000365
    "0000000000000001", -- 000000 (00000)  0  246 000366
    "0000000000000001", -- 000000 (00000)  0  247 000367
    "0000000000000001", -- 000000 (00000)  0  248 000370
    "0000000000000001", -- 000000 (00000)  0  249 000371
    "0000000000000001", -- 000000 (00000)  0  250 000372
    "0000000000000001", -- 000000 (00000)  0  251 000373
    "0000000000000001", -- 000000 (00000)  0  252 000374
    "0000000000000001", -- 000000 (00000)  0  253 000375
    "0000000000000001", -- 000000 (00000)  0  254 000376
    "0000000000000001", -- 000000 (00000)  0  255 000377
    "0000000000000001", -- 000000 (00000)  1    0 000400
    "0000000000000001", -- 000000 (00000)  1    1 000401
    "0000000000000001", -- 000000 (00000)  1    2 000402
    "0000000000000001", -- 000000 (00000)  1    3 000403
    "0000000000000001", -- 000000 (00000)  1    4 000404
    "0000000000000001", -- 000000 (00000)  1    5 000405
    "0000000000000001", -- 000000 (00000)  1    6 000406
    "0000000000000001", -- 000000 (00000)  1    7 000407
    "0000000000000001", -- 000000 (00000)  1    8 000410
    "0000000000000001", -- 000000 (00000)  1    9 000411
    "0000000000000001", -- 000000 (00000)  1   10 000412
    "0000000000000001", -- 000000 (00000)  1   11 000413
    "0000000000000001", -- 000000 (00000)  1   12 000414
    "0000000000000001", -- 000000 (00000)  1   13 000415
    "0000000000000001", -- 000000 (00000)  1   14 000416
    "0000000000000001", -- 000000 (00000)  1   15 000417
    "0000000000000001", -- 000000 (00000)  1   16 000420
    "0000000000000001", -- 000000 (00000)  1   17 000421
    "0000000000000001", -- 000000 (00000)  1   18 000422
    "0000000000000001", -- 000000 (00000)  1   19 000423
    "0000000000000001", -- 000000 (00000)  1   20 000424
    "0000000000000001", -- 000000 (00000)  1   21 000425
    "0000000000000001", -- 000000 (00000)  1   22 000426
    "0000000000000001", -- 000000 (00000)  1   23 000427
    "0000000000000001", -- 000000 (00000)  1   24 000430
    "0000000000000001", -- 000000 (00000)  1   25 000431
    "0000000000000001", -- 000000 (00000)  1   26 000432
    "0000000000000001", -- 000000 (00000)  1   27 000433
    "0000000000000001", -- 000000 (00000)  1   28 000434
    "0000000000000001", -- 000000 (00000)  1   29 000435
    "0000000000000001", -- 000000 (00000)  1   30 000436
    "0000000000000001", -- 000000 (00000)  1   31 000437
    "0000000000000001", -- 000000 (00000)  1   32 000440
    "0000000000000001", -- 000000 (00000)  1   33 000441
    "0000000000000001", -- 000000 (00000)  1   34 000442
    "0000000000000001", -- 000000 (00000)  1   35 000443
    "0000000000000001", -- 000000 (00000)  1   36 000444
    "0000000000000001", -- 000000 (00000)  1   37 000445
    "0000000000000001", -- 000000 (00000)  1   38 000446
    "0000000000000001", -- 000000 (00000)  1   39 000447
    "0000000000000001", -- 000000 (00000)  1   40 000450
    "0000000000000001", -- 000000 (00000)  1   41 000451
    "0000000000000001", -- 000000 (00000)  1   42 000452
    "0000000000000001", -- 000000 (00000)  1   43 000453
    "0000000000000001", -- 000000 (00000)  1   44 000454
    "0000000000000001", -- 000000 (00000)  1   45 000455
    "0000000000000001", -- 000000 (00000)  1   46 000456
    "0000000000000001", -- 000000 (00000)  1   47 000457
    "0000000000000001", -- 000000 (00000)  1   48 000460
    "0000000000000001", -- 000000 (00000)  1   49 000461
    "0000000000000001", -- 000000 (00000)  1   50 000462
    "0000000000000001", -- 000000 (00000)  1   51 000463
    "0000000000000001", -- 000000 (00000)  1   52 000464
    "0000000000000001", -- 000000 (00000)  1   53 000465
    "0000000000000001", -- 000000 (00000)  1   54 000466
    "0000000000000001", -- 000000 (00000)  1   55 000467
    "0000000000000001", -- 000000 (00000)  1   56 000470
    "0000000000000001", -- 000000 (00000)  1   57 000471
    "0000000000000001", -- 000000 (00000)  1   58 000472
    "0000000000000001", -- 000000 (00000)  1   59 000473
    "0000000000000001", -- 000000 (00000)  1   60 000474
    "0000000000000001", -- 000000 (00000)  1   61 000475
    "0000000000000001", -- 000000 (00000)  1   62 000476
    "0000000000000001", -- 000000 (00000)  1   63 000477
    "0000000000000001", -- 000000 (00000)  1   64 000500
    "0000000000000001", -- 000000 (00000)  1   65 000501
    "0000000000000001", -- 000000 (00000)  1   66 000502
    "0000000000000001", -- 000000 (00000)  1   67 000503
    "0000000000000001", -- 000000 (00000)  1   68 000504
    "0000000000000001", -- 000000 (00000)  1   69 000505
    "0000000000000001", -- 000000 (00000)  1   70 000506
    "0000000000000001", -- 000000 (00000)  1   71 000507
    "0000000000000001", -- 000000 (00000)  1   72 000510
    "0000000000000001", -- 000000 (00000)  1   73 000511
    "0000000000000001", -- 000000 (00000)  1   74 000512
    "0000000000000001", -- 000000 (00000)  1   75 000513
    "0000000000000001", -- 000000 (00000)  1   76 000514
    "0000000000000001", -- 000000 (00000)  1   77 000515
    "0000000000000001", -- 000000 (00000)  1   78 000516
    "0000000000000001", -- 000000 (00000)  1   79 000517
    "0000000000000001", -- 000000 (00000)  1   80 000520
    "0000000000000001", -- 000000 (00000)  1   81 000521
    "0000000000000001", -- 000000 (00000)  1   82 000522
    "0000000000000001", -- 000000 (00000)  1   83 000523
    "0000000000000001", -- 000000 (00000)  1   84 000524
    "0000000000000001", -- 000000 (00000)  1   85 000525
    "0000000000000001", -- 000000 (00000)  1   86 000526
    "0000000000000001", -- 000000 (00000)  1   87 000527
    "0000000000000001", -- 000000 (00000)  1   88 000530
    "0000000000000001", -- 000000 (00000)  1   89 000531
    "0000000000000001", -- 000000 (00000)  1   90 000532
    "0000000000000001", -- 000000 (00000)  1   91 000533
    "0000000000000001", -- 000000 (00000)  1   92 000534
    "0000000000000001", -- 000000 (00000)  1   93 000535
    "0000000000000001", -- 000000 (00000)  1   94 000536
    "0000000000000001", -- 000000 (00000)  1   95 000537
    "0000000000000001", -- 000000 (00000)  1   96 000540
    "0000000000000001", -- 000000 (00000)  1   97 000541
    "0000000000000001", -- 000000 (00000)  1   98 000542
    "0000000000000001", -- 000000 (00000)  1   99 000543
    "0000000000000001", -- 000000 (00000)  1  100 000544
    "0000000000000001", -- 000000 (00000)  1  101 000545
    "0000000000000001", -- 000000 (00000)  1  102 000546
    "0000000000000001", -- 000000 (00000)  1  103 000547
    "0000000000000001", -- 000000 (00000)  1  104 000550
    "0000000000000001", -- 000000 (00000)  1  105 000551
    "0000000000000001", -- 000000 (00000)  1  106 000552
    "0000000000000001", -- 000000 (00000)  1  107 000553
    "0000000000000001", -- 000000 (00000)  1  108 000554
    "0000000000000001", -- 000000 (00000)  1  109 000555
    "0000000000000001", -- 000000 (00000)  1  110 000556
    "0000000000000001", -- 000000 (00000)  1  111 000557
    "0000000000000001", -- 000000 (00000)  1  112 000560
    "0000000000000001", -- 000000 (00000)  1  113 000561
    "0000000000000001", -- 000000 (00000)  1  114 000562
    "0000000000000001", -- 000000 (00000)  1  115 000563
    "0000000000000001", -- 000000 (00000)  1  116 000564
    "0000000000000001", -- 000000 (00000)  1  117 000565
    "0000000000000001", -- 000000 (00000)  1  118 000566
    "0000000000000001", -- 000000 (00000)  1  119 000567
    "0000000000000001", -- 000000 (00000)  1  120 000570
    "0000000000000001", -- 000000 (00000)  1  121 000571
    "0000000000000001", -- 000000 (00000)  1  122 000572
    "0000000000000001", -- 000000 (00000)  1  123 000573
    "0000000000000001", -- 000000 (00000)  1  124 000574
    "0000000000000001", -- 000000 (00000)  1  125 000575
    "0000000000000001", -- 000000 (00000)  1  126 000576
    "0000000000000001", -- 000000 (00000)  1  127 000577
    "0000000000000001", -- 000000 (00000)  1  128 000600
    "0000000000000001", -- 000000 (00000)  1  129 000601
    "0000000000000001", -- 000000 (00000)  1  130 000602
    "0000000000000001", -- 000000 (00000)  1  131 000603
    "0000000000000001", -- 000000 (00000)  1  132 000604
    "0000000000000001", -- 000000 (00000)  1  133 000605
    "0000000000000001", -- 000000 (00000)  1  134 000606
    "0000000000000001", -- 000000 (00000)  1  135 000607
    "0000000000000001", -- 000000 (00000)  1  136 000610
    "0000000000000001", -- 000000 (00000)  1  137 000611
    "0000000000000001", -- 000000 (00000)  1  138 000612
    "0000000000000001", -- 000000 (00000)  1  139 000613
    "0000000000000001", -- 000000 (00000)  1  140 000614
    "0000000000000001", -- 000000 (00000)  1  141 000615
    "0000000000000001", -- 000000 (00000)  1  142 000616
    "0000000000000001", -- 000000 (00000)  1  143 000617
    "0000000000000001", -- 000000 (00000)  1  144 000620
    "0000000000000001", -- 000000 (00000)  1  145 000621
    "0000000000000001", -- 000000 (00000)  1  146 000622
    "0000000000000001", -- 000000 (00000)  1  147 000623
    "0000000000000001", -- 000000 (00000)  1  148 000624
    "0000000000000001", -- 000000 (00000)  1  149 000625
    "0000000000000001", -- 000000 (00000)  1  150 000626
    "0000000000000001", -- 000000 (00000)  1  151 000627
    "0000000000000001", -- 000000 (00000)  1  152 000630
    "0000000000000001", -- 000000 (00000)  1  153 000631
    "0000000000000001", -- 000000 (00000)  1  154 000632
    "0000000000000001", -- 000000 (00000)  1  155 000633
    "0000000000000001", -- 000000 (00000)  1  156 000634
    "0000000000000001", -- 000000 (00000)  1  157 000635
    "0000000000000001", -- 000000 (00000)  1  158 000636
    "0000000000000001", -- 000000 (00000)  1  159 000637
    "0000000000000001", -- 000000 (00000)  1  160 000640
    "0000000000000001", -- 000000 (00000)  1  161 000641
    "0000000000000001", -- 000000 (00000)  1  162 000642
    "0000000000000001", -- 000000 (00000)  1  163 000643
    "0000000000000001", -- 000000 (00000)  1  164 000644
    "0000000000000001", -- 000000 (00000)  1  165 000645
    "0000000000000001", -- 000000 (00000)  1  166 000646
    "0000000000000001", -- 000000 (00000)  1  167 000647
    "0000000000000001", -- 000000 (00000)  1  168 000650
    "0000000000000001", -- 000000 (00000)  1  169 000651
    "0000000000000001", -- 000000 (00000)  1  170 000652
    "0000000000000001", -- 000000 (00000)  1  171 000653
    "0000000000000001", -- 000000 (00000)  1  172 000654
    "0000000000000001", -- 000000 (00000)  1  173 000655
    "0000000000000001", -- 000000 (00000)  1  174 000656
    "0000000000000001", -- 000000 (00000)  1  175 000657
    "0000000000000001", -- 000000 (00000)  1  176 000660
    "0000000000000001", -- 000000 (00000)  1  177 000661
    "0000000000000001", -- 000000 (00000)  1  178 000662
    "0000000000000001", -- 000000 (00000)  1  179 000663
    "0000000000000001", -- 000000 (00000)  1  180 000664
    "0000000000000001", -- 000000 (00000)  1  181 000665
    "0000000000000001", -- 000000 (00000)  1  182 000666
    "0000000000000001", -- 000000 (00000)  1  183 000667
    "0000000000000001", -- 000000 (00000)  1  184 000670
    "0000000000000001", -- 000000 (00000)  1  185 000671
    "0000000000000001", -- 000000 (00000)  1  186 000672
    "0000000000000001", -- 000000 (00000)  1  187 000673
    "0000000000000001", -- 000000 (00000)  1  188 000674
    "0000000000000001", -- 000000 (00000)  1  189 000675
    "0000000000000001", -- 000000 (00000)  1  190 000676
    "0000000000000001", -- 000000 (00000)  1  191 000677
    "0000000000000001", -- 000000 (00000)  1  192 000700
    "0000000000000001", -- 000000 (00000)  1  193 000701
    "0000000000000001", -- 000000 (00000)  1  194 000702
    "0000000000000001", -- 000000 (00000)  1  195 000703
    "0000000000000001", -- 000000 (00000)  1  196 000704
    "0000000000000001", -- 000000 (00000)  1  197 000705
    "0000000000000001", -- 000000 (00000)  1  198 000706
    "0000000000000001", -- 000000 (00000)  1  199 000707
    "0000000000000001", -- 000000 (00000)  1  200 000710
    "0000000000000001", -- 000000 (00000)  1  201 000711
    "0000000000000001", -- 000000 (00000)  1  202 000712
    "0000000000000001", -- 000000 (00000)  1  203 000713
    "0000000000000001", -- 000000 (00000)  1  204 000714
    "0000000000000001", -- 000000 (00000)  1  205 000715
    "0000000000000001", -- 000000 (00000)  1  206 000716
    "0000000000000001", -- 000000 (00000)  1  207 000717
    "0000000000000001", -- 000000 (00000)  1  208 000720
    "0000000000000001", -- 000000 (00000)  1  209 000721
    "0000000000000001", -- 000000 (00000)  1  210 000722
    "0000000000000001", -- 000000 (00000)  1  211 000723
    "0000000000000001", -- 000000 (00000)  1  212 000724
    "0000000000000001", -- 000000 (00000)  1  213 000725
    "0000000000000001", -- 000000 (00000)  1  214 000726
    "0000000000000001", -- 000000 (00000)  1  215 000727
    "0000000000000001", -- 000000 (00000)  1  216 000730
    "0000000000000001", -- 000000 (00000)  1  217 000731
    "0000000000000001", -- 000000 (00000)  1  218 000732
    "0000000000000001", -- 000000 (00000)  1  219 000733
    "0000000000000001", -- 000000 (00000)  1  220 000734
    "0000000000000001", -- 000000 (00000)  1  221 000735
    "0000000000000001", -- 000000 (00000)  1  222 000736
    "0000000000000001", -- 000000 (00000)  1  223 000737
    "0000000000000001", -- 000000 (00000)  1  224 000740
    "0000000000000001", -- 000000 (00000)  1  225 000741
    "0000000000000001", -- 000000 (00000)  1  226 000742
    "0000000000000001", -- 000000 (00000)  1  227 000743
    "0000000000000001", -- 000000 (00000)  1  228 000744
    "0000000000000001", -- 000000 (00000)  1  229 000745
    "0000000000000001", -- 000000 (00000)  1  230 000746
    "0000000000000001", -- 000000 (00000)  1  231 000747
    "0000000000000001", -- 000000 (00000)  1  232 000750
    "0000000000000001", -- 000000 (00000)  1  233 000751
    "0000000000000001", -- 000000 (00000)  1  234 000752
    "0000000000000001", -- 000000 (00000)  1  235 000753
    "0000000000000001", -- 000000 (00000)  1  236 000754
    "0000000000000001", -- 000000 (00000)  1  237 000755
    "0000000000000001", -- 000000 (00000)  1  238 000756
    "0000000000000001", -- 000000 (00000)  1  239 000757
    "0000000000000001", -- 000000 (00000)  1  240 000760
    "0000000000000001", -- 000000 (00000)  1  241 000761
    "0000000000000001", -- 000000 (00000)  1  242 000762
    "0000000000000001", -- 000000 (00000)  1  243 000763
    "0000000000000001", -- 000000 (00000)  1  244 000764
    "0000000000000001", -- 000000 (00000)  1  245 000765
    "0000000000000001", -- 000000 (00000)  1  246 000766
    "0000000000000001", -- 000000 (00000)  1  247 000767
    "0000000000000001", -- 000000 (00000)  1  248 000770
    "0000000000000001", -- 000000 (00000)  1  249 000771
    "0000000000000001", -- 000000 (00000)  1  250 000772
    "0000000000000001", -- 000000 (00000)  1  251 000773
    "0000000000000001", -- 000000 (00000)  1  252 000774
    "0000000000000001", -- 000000 (00000)  1  253 000775
    "0000000000000001", -- 000000 (00000)  1  254 000776
    "0000000000000001", -- 000000 (00000)  1  255 000777
    "0000000000000001", -- 000000 (00000)  2    0 001000
    "0000000000000001", -- 000000 (00000)  2    1 001001
    "0000000000000001", -- 000000 (00000)  2    2 001002
    "0000000000000001", -- 000000 (00000)  2    3 001003
    "0000000000000001", -- 000000 (00000)  2    4 001004
    "0000000000000001", -- 000000 (00000)  2    5 001005
    "0000000000000001", -- 000000 (00000)  2    6 001006
    "0000000000000001", -- 000000 (00000)  2    7 001007
    "0000000000000001", -- 000000 (00000)  2    8 001010
    "0000000000000001", -- 000000 (00000)  2    9 001011
    "0000000000000001", -- 000000 (00000)  2   10 001012
    "0000000000000001", -- 000000 (00000)  2   11 001013
    "0000000000000001", -- 000000 (00000)  2   12 001014
    "0000000000000001", -- 000000 (00000)  2   13 001015
    "0000000000000001", -- 000000 (00000)  2   14 001016
    "0000000000000001", -- 000000 (00000)  2   15 001017
    "0000000000000001", -- 000000 (00000)  2   16 001020
    "0000000000000001", -- 000000 (00000)  2   17 001021
    "0000000000000001", -- 000000 (00000)  2   18 001022
    "0000000000000001", -- 000000 (00000)  2   19 001023
    "0000000000000001", -- 000000 (00000)  2   20 001024
    "0000000000000001", -- 000000 (00000)  2   21 001025
    "0000000000000001", -- 000000 (00000)  2   22 001026
    "0000000000000001", -- 000000 (00000)  2   23 001027
    "0000000000000001", -- 000000 (00000)  2   24 001030
    "0000000000000001", -- 000000 (00000)  2   25 001031
    "0000000000000001", -- 000000 (00000)  2   26 001032
    "0000000000000001", -- 000000 (00000)  2   27 001033
    "0000000000000001", -- 000000 (00000)  2   28 001034
    "0000000000000001", -- 000000 (00000)  2   29 001035
    "0000000000000001", -- 000000 (00000)  2   30 001036
    "0000000000000001", -- 000000 (00000)  2   31 001037
    "0000000000000001", -- 000000 (00000)  2   32 001040
    "0000000000000001", -- 000000 (00000)  2   33 001041
    "0000000000000001", -- 000000 (00000)  2   34 001042
    "0000000000000001", -- 000000 (00000)  2   35 001043
    "0000000000000001", -- 000000 (00000)  2   36 001044
    "0000000000000001", -- 000000 (00000)  2   37 001045
    "0000000000000001", -- 000000 (00000)  2   38 001046
    "0000000000000001", -- 000000 (00000)  2   39 001047
    "0000000000000001", -- 000000 (00000)  2   40 001050
    "0000000000000001", -- 000000 (00000)  2   41 001051
    "0000000000000001", -- 000000 (00000)  2   42 001052
    "0000000000000001", -- 000000 (00000)  2   43 001053
    "0000000000000001", -- 000000 (00000)  2   44 001054
    "0000000000000001", -- 000000 (00000)  2   45 001055
    "0000000000000001", -- 000000 (00000)  2   46 001056
    "0000000000000001", -- 000000 (00000)  2   47 001057
    "0000000000000001", -- 000000 (00000)  2   48 001060
    "0000000000000001", -- 000000 (00000)  2   49 001061
    "0000000000000001", -- 000000 (00000)  2   50 001062
    "0000000000000001", -- 000000 (00000)  2   51 001063
    "0000000000000001", -- 000000 (00000)  2   52 001064
    "0000000000000001", -- 000000 (00000)  2   53 001065
    "0000000000000001", -- 000000 (00000)  2   54 001066
    "0000000000000001", -- 000000 (00000)  2   55 001067
    "0000000000000001", -- 000000 (00000)  2   56 001070
    "0000000000000001", -- 000000 (00000)  2   57 001071
    "0000000000000001", -- 000000 (00000)  2   58 001072
    "0000000000000001", -- 000000 (00000)  2   59 001073
    "0000000000000001", -- 000000 (00000)  2   60 001074
    "0000000000000001", -- 000000 (00000)  2   61 001075
    "0000000000000001", -- 000000 (00000)  2   62 001076
    "0000000000000001", -- 000000 (00000)  2   63 001077
    "0000000000000001", -- 000000 (00000)  2   64 001100
    "0000000000000001", -- 000000 (00000)  2   65 001101
    "0000000000000001", -- 000000 (00000)  2   66 001102
    "0000000000000001", -- 000000 (00000)  2   67 001103
    "0000000000000001", -- 000000 (00000)  2   68 001104
    "0000000000000001", -- 000000 (00000)  2   69 001105
    "0000000000000001", -- 000000 (00000)  2   70 001106
    "0000000000000001", -- 000000 (00000)  2   71 001107
    "0000000000000001", -- 000000 (00000)  2   72 001110
    "0000000000000001", -- 000000 (00000)  2   73 001111
    "0000000000000001", -- 000000 (00000)  2   74 001112
    "0000000000000001", -- 000000 (00000)  2   75 001113
    "0000000000000001", -- 000000 (00000)  2   76 001114
    "0000000000000001", -- 000000 (00000)  2   77 001115
    "0000000000000001", -- 000000 (00000)  2   78 001116
    "0000000000000001", -- 000000 (00000)  2   79 001117
    "0000000000000001", -- 000000 (00000)  2   80 001120
    "0000000000000001", -- 000000 (00000)  2   81 001121
    "0000000000000001", -- 000000 (00000)  2   82 001122
    "0000000000000001", -- 000000 (00000)  2   83 001123
    "0000000000000001", -- 000000 (00000)  2   84 001124
    "0000000000000001", -- 000000 (00000)  2   85 001125
    "0000000000000001", -- 000000 (00000)  2   86 001126
    "0000000000000001", -- 000000 (00000)  2   87 001127
    "0000000000000001", -- 000000 (00000)  2   88 001130
    "0000000000000001", -- 000000 (00000)  2   89 001131
    "0000000000000001", -- 000000 (00000)  2   90 001132
    "0000000000000001", -- 000000 (00000)  2   91 001133
    "0000000000000001", -- 000000 (00000)  2   92 001134
    "0000000000000001", -- 000000 (00000)  2   93 001135
    "0000000000000001", -- 000000 (00000)  2   94 001136
    "0000000000000001", -- 000000 (00000)  2   95 001137
    "0000000000000001", -- 000000 (00000)  2   96 001140
    "0000000000000001", -- 000000 (00000)  2   97 001141
    "0000000000000001", -- 000000 (00000)  2   98 001142
    "0000000000000001", -- 000000 (00000)  2   99 001143
    "0000000000000001", -- 000000 (00000)  2  100 001144
    "0000000000000001", -- 000000 (00000)  2  101 001145
    "0000000000000001", -- 000000 (00000)  2  102 001146
    "0000000000000001", -- 000000 (00000)  2  103 001147
    "0000000000000001", -- 000000 (00000)  2  104 001150
    "0000000000000001", -- 000000 (00000)  2  105 001151
    "0000000000000001", -- 000000 (00000)  2  106 001152
    "0000000000000001", -- 000000 (00000)  2  107 001153
    "0000000000000001", -- 000000 (00000)  2  108 001154
    "0000000000000001", -- 000000 (00000)  2  109 001155
    "0000000000000001", -- 000000 (00000)  2  110 001156
    "0000000000000001", -- 000000 (00000)  2  111 001157
    "0000000000000001", -- 000000 (00000)  2  112 001160
    "0000000000000001", -- 000000 (00000)  2  113 001161
    "0000000000000001", -- 000000 (00000)  2  114 001162
    "0000000000000001", -- 000000 (00000)  2  115 001163
    "0000000000000001", -- 000000 (00000)  2  116 001164
    "0000000000000001", -- 000000 (00000)  2  117 001165
    "0000000000000001", -- 000000 (00000)  2  118 001166
    "0000000000000001", -- 000000 (00000)  2  119 001167
    "0000000000000001", -- 000000 (00000)  2  120 001170
    "0000000000000001", -- 000000 (00000)  2  121 001171
    "0000000000000001", -- 000000 (00000)  2  122 001172
    "0000000000000001", -- 000000 (00000)  2  123 001173
    "0000000000000001", -- 000000 (00000)  2  124 001174
    "0000000000000001", -- 000000 (00000)  2  125 001175
    "0000000000000001", -- 000000 (00000)  2  126 001176
    "0000000000000001", -- 000000 (00000)  2  127 001177
    "0000000000000001", -- 000000 (00000)  2  128 001200
    "0000000000000001", -- 000000 (00000)  2  129 001201
    "0000000000000001", -- 000000 (00000)  2  130 001202
    "0000000000000001", -- 000000 (00000)  2  131 001203
    "0000000000000001", -- 000000 (00000)  2  132 001204
    "0000000000000001", -- 000000 (00000)  2  133 001205
    "0000000000000001", -- 000000 (00000)  2  134 001206
    "0000000000000001", -- 000000 (00000)  2  135 001207
    "0000000000000001", -- 000000 (00000)  2  136 001210
    "0000000000000001", -- 000000 (00000)  2  137 001211
    "0000000000000001", -- 000000 (00000)  2  138 001212
    "0000000000000001", -- 000000 (00000)  2  139 001213
    "0000000000000001", -- 000000 (00000)  2  140 001214
    "0000000000000001", -- 000000 (00000)  2  141 001215
    "0000000000000001", -- 000000 (00000)  2  142 001216
    "0000000000000001", -- 000000 (00000)  2  143 001217
    "0000000000000001", -- 000000 (00000)  2  144 001220
    "0000000000000001", -- 000000 (00000)  2  145 001221
    "0000000000000001", -- 000000 (00000)  2  146 001222
    "0000000000000001", -- 000000 (00000)  2  147 001223
    "0000000000000001", -- 000000 (00000)  2  148 001224
    "0000000000000001", -- 000000 (00000)  2  149 001225
    "0000000000000001", -- 000000 (00000)  2  150 001226
    "0000000000000001", -- 000000 (00000)  2  151 001227
    "0000000000000001", -- 000000 (00000)  2  152 001230
    "0000000000000001", -- 000000 (00000)  2  153 001231
    "0000000000000001", -- 000000 (00000)  2  154 001232
    "0000000000000001", -- 000000 (00000)  2  155 001233
    "0000000000000001", -- 000000 (00000)  2  156 001234
    "0000000000000001", -- 000000 (00000)  2  157 001235
    "0000000000000001", -- 000000 (00000)  2  158 001236
    "0000000000000001", -- 000000 (00000)  2  159 001237
    "0000000000000001", -- 000000 (00000)  2  160 001240
    "0000000000000001", -- 000000 (00000)  2  161 001241
    "0000000000000001", -- 000000 (00000)  2  162 001242
    "0000000000000001", -- 000000 (00000)  2  163 001243
    "0000000000000001", -- 000000 (00000)  2  164 001244
    "0000000000000001", -- 000000 (00000)  2  165 001245
    "0000000000000001", -- 000000 (00000)  2  166 001246
    "0000000000000001", -- 000000 (00000)  2  167 001247
    "0000000000000001", -- 000000 (00000)  2  168 001250
    "0000000000000001", -- 000000 (00000)  2  169 001251
    "0000000000000001", -- 000000 (00000)  2  170 001252
    "0000000000000001", -- 000000 (00000)  2  171 001253
    "0000000000000001", -- 000000 (00000)  2  172 001254
    "0000000000000001", -- 000000 (00000)  2  173 001255
    "0000000000000001", -- 000000 (00000)  2  174 001256
    "0000000000000001", -- 000000 (00000)  2  175 001257
    "0000000000000001", -- 000000 (00000)  2  176 001260
    "0000000000000001", -- 000000 (00000)  2  177 001261
    "0000000000000001", -- 000000 (00000)  2  178 001262
    "0000000000000001", -- 000000 (00000)  2  179 001263
    "0000000000000001", -- 000000 (00000)  2  180 001264
    "0000000000000001", -- 000000 (00000)  2  181 001265
    "0000000000000001", -- 000000 (00000)  2  182 001266
    "0000000000000001", -- 000000 (00000)  2  183 001267
    "0000000000000001", -- 000000 (00000)  2  184 001270
    "0000000000000001", -- 000000 (00000)  2  185 001271
    "0000000000000001", -- 000000 (00000)  2  186 001272
    "0000000000000001", -- 000000 (00000)  2  187 001273
    "0000000000000001", -- 000000 (00000)  2  188 001274
    "0000000000000001", -- 000000 (00000)  2  189 001275
    "0000000000000001", -- 000000 (00000)  2  190 001276
    "0000000000000001", -- 000000 (00000)  2  191 001277
    "0000000000000001", -- 000000 (00000)  2  192 001300
    "0000000000000001", -- 000000 (00000)  2  193 001301
    "0000000000000001", -- 000000 (00000)  2  194 001302
    "0000000000000001", -- 000000 (00000)  2  195 001303
    "0000000000000001", -- 000000 (00000)  2  196 001304
    "0000000000000001", -- 000000 (00000)  2  197 001305
    "0000000000000001", -- 000000 (00000)  2  198 001306
    "0000000000000001", -- 000000 (00000)  2  199 001307
    "0000000000000001", -- 000000 (00000)  2  200 001310
    "0000000000000001", -- 000000 (00000)  2  201 001311
    "0000000000000001", -- 000000 (00000)  2  202 001312
    "0000000000000001", -- 000000 (00000)  2  203 001313
    "0000000000000001", -- 000000 (00000)  2  204 001314
    "0000000000000001", -- 000000 (00000)  2  205 001315
    "0000000000000001", -- 000000 (00000)  2  206 001316
    "0000000000000001", -- 000000 (00000)  2  207 001317
    "0000000000000001", -- 000000 (00000)  2  208 001320
    "0000000000000001", -- 000000 (00000)  2  209 001321
    "0000000000000001", -- 000000 (00000)  2  210 001322
    "0000000000000001", -- 000000 (00000)  2  211 001323
    "0000000000000001", -- 000000 (00000)  2  212 001324
    "0000000000000001", -- 000000 (00000)  2  213 001325
    "0000000000000001", -- 000000 (00000)  2  214 001326
    "0000000000000001", -- 000000 (00000)  2  215 001327
    "0000000000000001", -- 000000 (00000)  2  216 001330
    "0000000000000001", -- 000000 (00000)  2  217 001331
    "0000000000000001", -- 000000 (00000)  2  218 001332
    "0000000000000001", -- 000000 (00000)  2  219 001333
    "0000000000000001", -- 000000 (00000)  2  220 001334
    "0000000000000001", -- 000000 (00000)  2  221 001335
    "0000000000000001", -- 000000 (00000)  2  222 001336
    "0000000000000001", -- 000000 (00000)  2  223 001337
    "0000000000000001", -- 000000 (00000)  2  224 001340
    "0000000000000001", -- 000000 (00000)  2  225 001341
    "0000000000000001", -- 000000 (00000)  2  226 001342
    "0000000000000001", -- 000000 (00000)  2  227 001343
    "0000000000000001", -- 000000 (00000)  2  228 001344
    "0000000000000001", -- 000000 (00000)  2  229 001345
    "0000000000000001", -- 000000 (00000)  2  230 001346
    "0000000000000001", -- 000000 (00000)  2  231 001347
    "0000000000000001", -- 000000 (00000)  2  232 001350
    "0000000000000001", -- 000000 (00000)  2  233 001351
    "0000000000000001", -- 000000 (00000)  2  234 001352
    "0000000000000001", -- 000000 (00000)  2  235 001353
    "0000000000000001", -- 000000 (00000)  2  236 001354
    "0000000000000001", -- 000000 (00000)  2  237 001355
    "0000000000000001", -- 000000 (00000)  2  238 001356
    "0000000000000001", -- 000000 (00000)  2  239 001357
    "0000000000000001", -- 000000 (00000)  2  240 001360
    "0000000000000001", -- 000000 (00000)  2  241 001361
    "0000000000000001", -- 000000 (00000)  2  242 001362
    "0000000000000001", -- 000000 (00000)  2  243 001363
    "0000000000000001", -- 000000 (00000)  2  244 001364
    "0000000000000001", -- 000000 (00000)  2  245 001365
    "0000000000000001", -- 000000 (00000)  2  246 001366
    "0000000000000001", -- 000000 (00000)  2  247 001367
    "0000000000000001", -- 000000 (00000)  2  248 001370
    "0000000000000001", -- 000000 (00000)  2  249 001371
    "0000000000000001", -- 000000 (00000)  2  250 001372
    "0000000000000001", -- 000000 (00000)  2  251 001373
    "0000000000000001", -- 000000 (00000)  2  252 001374
    "0000000000000001", -- 000000 (00000)  2  253 001375
    "0000000000000001", -- 000000 (00000)  2  254 001376
    "0000000000000001", -- 000000 (00000)  2  255 001377
    "0000000000000001", -- 000000 (00000)  3    0 001400
    "0000000000000001", -- 000000 (00000)  3    1 001401
    "0000000000000001", -- 000000 (00000)  3    2 001402
    "0000000000000001", -- 000000 (00000)  3    3 001403
    "0000000000000001", -- 000000 (00000)  3    4 001404
    "0000000000000001", -- 000000 (00000)  3    5 001405
    "0000000000000001", -- 000000 (00000)  3    6 001406
    "0000000000000001", -- 000000 (00000)  3    7 001407
    "0000000000000001", -- 000000 (00000)  3    8 001410
    "0000000000000001", -- 000000 (00000)  3    9 001411
    "0000000000000001", -- 000000 (00000)  3   10 001412
    "0000000000000001", -- 000000 (00000)  3   11 001413
    "0000000000000001", -- 000000 (00000)  3   12 001414
    "0000000000000001", -- 000000 (00000)  3   13 001415
    "0000000000000001", -- 000000 (00000)  3   14 001416
    "0000000000000001", -- 000000 (00000)  3   15 001417
    "0000000000000001", -- 000000 (00000)  3   16 001420
    "0000000000000001", -- 000000 (00000)  3   17 001421
    "0000000000000001", -- 000000 (00000)  3   18 001422
    "0000000000000001", -- 000000 (00000)  3   19 001423
    "0000000000000001", -- 000000 (00000)  3   20 001424
    "0000000000000001", -- 000000 (00000)  3   21 001425
    "0000000000000001", -- 000000 (00000)  3   22 001426
    "0000000000000001", -- 000000 (00000)  3   23 001427
    "0000000000000001", -- 000000 (00000)  3   24 001430
    "0000000000000001", -- 000000 (00000)  3   25 001431
    "0000000000000001", -- 000000 (00000)  3   26 001432
    "0000000000000001", -- 000000 (00000)  3   27 001433
    "0000000000000001", -- 000000 (00000)  3   28 001434
    "0000000000000001", -- 000000 (00000)  3   29 001435
    "0000000000000001", -- 000000 (00000)  3   30 001436
    "0000000000000001", -- 000000 (00000)  3   31 001437
    "0000000000000001", -- 000000 (00000)  3   32 001440
    "0000000000000001", -- 000000 (00000)  3   33 001441
    "0000000000000001", -- 000000 (00000)  3   34 001442
    "0000000000000001", -- 000000 (00000)  3   35 001443
    "0000000000000001", -- 000000 (00000)  3   36 001444
    "0000000000000001", -- 000000 (00000)  3   37 001445
    "0000000000000001", -- 000000 (00000)  3   38 001446
    "0000000000000001", -- 000000 (00000)  3   39 001447
    "0000000000000001", -- 000000 (00000)  3   40 001450
    "0000000000000001", -- 000000 (00000)  3   41 001451
    "0000000000000001", -- 000000 (00000)  3   42 001452
    "0000000000000001", -- 000000 (00000)  3   43 001453
    "0000000000000001", -- 000000 (00000)  3   44 001454
    "0000000000000001", -- 000000 (00000)  3   45 001455
    "0000000000000001", -- 000000 (00000)  3   46 001456
    "0000000000000001", -- 000000 (00000)  3   47 001457
    "0000000000000001", -- 000000 (00000)  3   48 001460
    "0000000000000001", -- 000000 (00000)  3   49 001461
    "0000000000000001", -- 000000 (00000)  3   50 001462
    "0000000000000001", -- 000000 (00000)  3   51 001463
    "0000000000000001", -- 000000 (00000)  3   52 001464
    "0000000000000001", -- 000000 (00000)  3   53 001465
    "0000000000000001", -- 000000 (00000)  3   54 001466
    "0000000000000001", -- 000000 (00000)  3   55 001467
    "0000000000000001", -- 000000 (00000)  3   56 001470
    "0000000000000001", -- 000000 (00000)  3   57 001471
    "0000000000000001", -- 000000 (00000)  3   58 001472
    "0000000000000001", -- 000000 (00000)  3   59 001473
    "0000000000000001", -- 000000 (00000)  3   60 001474
    "0000000000000001", -- 000000 (00000)  3   61 001475
    "0000000000000001", -- 000000 (00000)  3   62 001476
    "0000000000000001", -- 000000 (00000)  3   63 001477
    "0000000000000001", -- 000000 (00000)  3   64 001500
    "0000000000000001", -- 000000 (00000)  3   65 001501
    "0000000000000001", -- 000000 (00000)  3   66 001502
    "0000000000000001", -- 000000 (00000)  3   67 001503
    "0000000000000001", -- 000000 (00000)  3   68 001504
    "0000000000000001", -- 000000 (00000)  3   69 001505
    "0000000000000001", -- 000000 (00000)  3   70 001506
    "0000000000000001", -- 000000 (00000)  3   71 001507
    "0000000000000001", -- 000000 (00000)  3   72 001510
    "0000000000000001", -- 000000 (00000)  3   73 001511
    "0000000000000001", -- 000000 (00000)  3   74 001512
    "0000000000000001", -- 000000 (00000)  3   75 001513
    "0000000000000001", -- 000000 (00000)  3   76 001514
    "0000000000000001", -- 000000 (00000)  3   77 001515
    "0000000000000001", -- 000000 (00000)  3   78 001516
    "0000000000000001", -- 000000 (00000)  3   79 001517
    "0000000000000001", -- 000000 (00000)  3   80 001520
    "0000000000000001", -- 000000 (00000)  3   81 001521
    "0000000000000001", -- 000000 (00000)  3   82 001522
    "0000000000000001", -- 000000 (00000)  3   83 001523
    "0000000000000001", -- 000000 (00000)  3   84 001524
    "0000000000000001", -- 000000 (00000)  3   85 001525
    "0000000000000001", -- 000000 (00000)  3   86 001526
    "0000000000000001", -- 000000 (00000)  3   87 001527
    "0000000000000001", -- 000000 (00000)  3   88 001530
    "0000000000000001", -- 000000 (00000)  3   89 001531
    "0000000000000001", -- 000000 (00000)  3   90 001532
    "0000000000000001", -- 000000 (00000)  3   91 001533
    "0000000000000001", -- 000000 (00000)  3   92 001534
    "0000000000000001", -- 000000 (00000)  3   93 001535
    "0000000000000001", -- 000000 (00000)  3   94 001536
    "0000000000000001", -- 000000 (00000)  3   95 001537
    "0000000000000001", -- 000000 (00000)  3   96 001540
    "0000000000000001", -- 000000 (00000)  3   97 001541
    "0000000000000001", -- 000000 (00000)  3   98 001542
    "0000000000000001", -- 000000 (00000)  3   99 001543
    "0000000000000001", -- 000000 (00000)  3  100 001544
    "0000000000000001", -- 000000 (00000)  3  101 001545
    "0000000000000001", -- 000000 (00000)  3  102 001546
    "0000000000000001", -- 000000 (00000)  3  103 001547
    "0000000000000001", -- 000000 (00000)  3  104 001550
    "0000000000000001", -- 000000 (00000)  3  105 001551
    "0000000000000001", -- 000000 (00000)  3  106 001552
    "0000000000000001", -- 000000 (00000)  3  107 001553
    "0000000000000001", -- 000000 (00000)  3  108 001554
    "0000000000000001", -- 000000 (00000)  3  109 001555
    "0000000000000001", -- 000000 (00000)  3  110 001556
    "0000000000000001", -- 000000 (00000)  3  111 001557
    "0000000000000001", -- 000000 (00000)  3  112 001560
    "0000000000000001", -- 000000 (00000)  3  113 001561
    "0000000000000001", -- 000000 (00000)  3  114 001562
    "0000000000000001", -- 000000 (00000)  3  115 001563
    "0000000000000001", -- 000000 (00000)  3  116 001564
    "0000000000000001", -- 000000 (00000)  3  117 001565
    "0000000000000001", -- 000000 (00000)  3  118 001566
    "0000000000000001", -- 000000 (00000)  3  119 001567
    "0000000000000001", -- 000000 (00000)  3  120 001570
    "0000000000000001", -- 000000 (00000)  3  121 001571
    "0000000000000001", -- 000000 (00000)  3  122 001572
    "0000000000000001", -- 000000 (00000)  3  123 001573
    "0000000000000001", -- 000000 (00000)  3  124 001574
    "0000000000000001", -- 000000 (00000)  3  125 001575
    "0000000000000001", -- 000000 (00000)  3  126 001576
    "0000000000000001", -- 000000 (00000)  3  127 001577
    "0000000000000001", -- 000000 (00000)  3  128 001600
    "0000000000000001", -- 000000 (00000)  3  129 001601
    "0000000000000001", -- 000000 (00000)  3  130 001602
    "0000000000000001", -- 000000 (00000)  3  131 001603
    "0000000000000001", -- 000000 (00000)  3  132 001604
    "0000000000000001", -- 000000 (00000)  3  133 001605
    "0000000000000001", -- 000000 (00000)  3  134 001606
    "0000000000000001", -- 000000 (00000)  3  135 001607
    "0000000000000001", -- 000000 (00000)  3  136 001610
    "0000000000000001", -- 000000 (00000)  3  137 001611
    "0000000000000001", -- 000000 (00000)  3  138 001612
    "0000000000000001", -- 000000 (00000)  3  139 001613
    "0000000000000001", -- 000000 (00000)  3  140 001614
    "0000000000000001", -- 000000 (00000)  3  141 001615
    "0000000000000001", -- 000000 (00000)  3  142 001616
    "0000000000000001", -- 000000 (00000)  3  143 001617
    "0000000000000001", -- 000000 (00000)  3  144 001620
    "0000000000000001", -- 000000 (00000)  3  145 001621
    "0000000000000001", -- 000000 (00000)  3  146 001622
    "0000000000000001", -- 000000 (00000)  3  147 001623
    "0000000000000001", -- 000000 (00000)  3  148 001624
    "0000000000000001", -- 000000 (00000)  3  149 001625
    "0000000000000001", -- 000000 (00000)  3  150 001626
    "0000000000000001", -- 000000 (00000)  3  151 001627
    "0000000000000001", -- 000000 (00000)  3  152 001630
    "0000000000000001", -- 000000 (00000)  3  153 001631
    "0000000000000001", -- 000000 (00000)  3  154 001632
    "0000000000000001", -- 000000 (00000)  3  155 001633
    "0000000000000001", -- 000000 (00000)  3  156 001634
    "0000000000000001", -- 000000 (00000)  3  157 001635
    "0000000000000001", -- 000000 (00000)  3  158 001636
    "0000000000000001", -- 000000 (00000)  3  159 001637
    "0000000000000001", -- 000000 (00000)  3  160 001640
    "0000000000000001", -- 000000 (00000)  3  161 001641
    "0000000000000001", -- 000000 (00000)  3  162 001642
    "0000000000000001", -- 000000 (00000)  3  163 001643
    "0000000000000001", -- 000000 (00000)  3  164 001644
    "0000000000000001", -- 000000 (00000)  3  165 001645
    "0000000000000001", -- 000000 (00000)  3  166 001646
    "0000000000000001", -- 000000 (00000)  3  167 001647
    "0000000000000001", -- 000000 (00000)  3  168 001650
    "0000000000000001", -- 000000 (00000)  3  169 001651
    "0000000000000001", -- 000000 (00000)  3  170 001652
    "0000000000000001", -- 000000 (00000)  3  171 001653
    "0000000000000001", -- 000000 (00000)  3  172 001654
    "0000000000000001", -- 000000 (00000)  3  173 001655
    "0000000000000001", -- 000000 (00000)  3  174 001656
    "0000000000000001", -- 000000 (00000)  3  175 001657
    "0000000000000001", -- 000000 (00000)  3  176 001660
    "0000000000000001", -- 000000 (00000)  3  177 001661
    "0000000000000001", -- 000000 (00000)  3  178 001662
    "0000000000000001", -- 000000 (00000)  3  179 001663
    "0000000000000001", -- 000000 (00000)  3  180 001664
    "0000000000000001", -- 000000 (00000)  3  181 001665
    "0000000000000001", -- 000000 (00000)  3  182 001666
    "0000000000000001", -- 000000 (00000)  3  183 001667
    "0000000000000001", -- 000000 (00000)  3  184 001670
    "0000000000000001", -- 000000 (00000)  3  185 001671
    "0000000000000001", -- 000000 (00000)  3  186 001672
    "0000000000000001", -- 000000 (00000)  3  187 001673
    "0000000000000001", -- 000000 (00000)  3  188 001674
    "0000000000000001", -- 000000 (00000)  3  189 001675
    "0000000000000001", -- 000000 (00000)  3  190 001676
    "0000000000000001", -- 000000 (00000)  3  191 001677
    "0000000000000001", -- 000000 (00000)  3  192 001700
    "0000000000000001", -- 000000 (00000)  3  193 001701
    "0000000000000001", -- 000000 (00000)  3  194 001702
    "0000000000000001", -- 000000 (00000)  3  195 001703
    "0000000000000001", -- 000000 (00000)  3  196 001704
    "0000000000000001", -- 000000 (00000)  3  197 001705
    "0000000000000001", -- 000000 (00000)  3  198 001706
    "0000000000000001", -- 000000 (00000)  3  199 001707
    "0000000000000001", -- 000000 (00000)  3  200 001710
    "0000000000000001", -- 000000 (00000)  3  201 001711
    "0000000000000001", -- 000000 (00000)  3  202 001712
    "0000000000000001", -- 000000 (00000)  3  203 001713
    "0000000000000001", -- 000000 (00000)  3  204 001714
    "0000000000000001", -- 000000 (00000)  3  205 001715
    "0000000000000001", -- 000000 (00000)  3  206 001716
    "0000000000000001", -- 000000 (00000)  3  207 001717
    "0000000000000001", -- 000000 (00000)  3  208 001720
    "0000000000000001", -- 000000 (00000)  3  209 001721
    "0000000000000001", -- 000000 (00000)  3  210 001722
    "0000000000000001", -- 000000 (00000)  3  211 001723
    "0000000000000001", -- 000000 (00000)  3  212 001724
    "0000000000000001", -- 000000 (00000)  3  213 001725
    "0000000000000001", -- 000000 (00000)  3  214 001726
    "0000000000000001", -- 000000 (00000)  3  215 001727
    "0000000000000001", -- 000000 (00000)  3  216 001730
    "0000000000000001", -- 000000 (00000)  3  217 001731
    "0000000000000001", -- 000000 (00000)  3  218 001732
    "0000000000000001", -- 000000 (00000)  3  219 001733
    "0000000000000001", -- 000000 (00000)  3  220 001734
    "0000000000000001", -- 000000 (00000)  3  221 001735
    "0000000000000001", -- 000000 (00000)  3  222 001736
    "0000000000000001", -- 000000 (00000)  3  223 001737
    "0000000000000001", -- 000000 (00000)  3  224 001740
    "0000000000000001", -- 000000 (00000)  3  225 001741
    "0000000000000001", -- 000000 (00000)  3  226 001742
    "0000000000000001", -- 000000 (00000)  3  227 001743
    "0000000000000001", -- 000000 (00000)  3  228 001744
    "0000000000000001", -- 000000 (00000)  3  229 001745
    "0000000000000001", -- 000000 (00000)  3  230 001746
    "0000000000000001", -- 000000 (00000)  3  231 001747
    "0000000000000001", -- 000000 (00000)  3  232 001750
    "0000000000000001", -- 000000 (00000)  3  233 001751
    "0000000000000001", -- 000000 (00000)  3  234 001752
    "0000000000000001", -- 000000 (00000)  3  235 001753
    "0000000000000001", -- 000000 (00000)  3  236 001754
    "0000000000000001", -- 000000 (00000)  3  237 001755
    "0000000000000001", -- 000000 (00000)  3  238 001756
    "0000000000000001", -- 000000 (00000)  3  239 001757
    "0000000000000001", -- 000000 (00000)  3  240 001760
    "0000000000000001", -- 000000 (00000)  3  241 001761
    "0000000000000001", -- 000000 (00000)  3  242 001762
    "0000000000000001", -- 000000 (00000)  3  243 001763
    "0000000000000001", -- 000000 (00000)  3  244 001764
    "0000000000000001", -- 000000 (00000)  3  245 001765
    "0000000000000001", -- 000000 (00000)  3  246 001766
    "0000000000000001", -- 000000 (00000)  3  247 001767
    "0000000000000001", -- 000000 (00000)  3  248 001770
    "0000000000000001", -- 000000 (00000)  3  249 001771
    "0000000000000001", -- 000000 (00000)  3  250 001772
    "0000000000000001", -- 000000 (00000)  3  251 001773
    "0000000000000001", -- 000000 (00000)  3  252 001774
    "0000000000000001", -- 000000 (00000)  3  253 001775
    "0000000000000001", -- 000000 (00000)  3  254 001776
    "0000000000000001", -- 000000 (00000)  3  255 001777
    "0000000000000001", -- 000000 (00000)  4    0 002000
    "0000000000000001", -- 000000 (00000)  4    1 002001
    "0000000000000001", -- 000000 (00000)  4    2 002002
    "0000000000000001", -- 000000 (00000)  4    3 002003
    "0000000000000001", -- 000000 (00000)  4    4 002004
    "0000000000000001", -- 000000 (00000)  4    5 002005
    "0000000000000001", -- 000000 (00000)  4    6 002006
    "0000000000000001", -- 000000 (00000)  4    7 002007
    "0000000000000001", -- 000000 (00000)  4    8 002010
    "0000000000000001", -- 000000 (00000)  4    9 002011
    "0000000000000001", -- 000000 (00000)  4   10 002012
    "0000000000000001", -- 000000 (00000)  4   11 002013
    "0000000000000001", -- 000000 (00000)  4   12 002014
    "0000000000000001", -- 000000 (00000)  4   13 002015
    "0000000000000001", -- 000000 (00000)  4   14 002016
    "0000000000000001", -- 000000 (00000)  4   15 002017
    "0000000000000001", -- 000000 (00000)  4   16 002020
    "0000000000000001", -- 000000 (00000)  4   17 002021
    "0000000000000001", -- 000000 (00000)  4   18 002022
    "0000000000000001", -- 000000 (00000)  4   19 002023
    "0000000000000001", -- 000000 (00000)  4   20 002024
    "0000000000000001", -- 000000 (00000)  4   21 002025
    "0000000000000001", -- 000000 (00000)  4   22 002026
    "0000000000000001", -- 000000 (00000)  4   23 002027
    "0000000000000001", -- 000000 (00000)  4   24 002030
    "0000000000000001", -- 000000 (00000)  4   25 002031
    "0000000000000001", -- 000000 (00000)  4   26 002032
    "0000000000000001", -- 000000 (00000)  4   27 002033
    "0000000000000001", -- 000000 (00000)  4   28 002034
    "0000000000000001", -- 000000 (00000)  4   29 002035
    "0000000000000001", -- 000000 (00000)  4   30 002036
    "0000000000000001", -- 000000 (00000)  4   31 002037
    "0000000000000001", -- 000000 (00000)  4   32 002040
    "0000000000000001", -- 000000 (00000)  4   33 002041
    "0000000000000001", -- 000000 (00000)  4   34 002042
    "0000000000000001", -- 000000 (00000)  4   35 002043
    "0000000000000001", -- 000000 (00000)  4   36 002044
    "0000000000000001", -- 000000 (00000)  4   37 002045
    "0000000000000001", -- 000000 (00000)  4   38 002046
    "0000000000000001", -- 000000 (00000)  4   39 002047
    "0000000000000001", -- 000000 (00000)  4   40 002050
    "0000000000000001", -- 000000 (00000)  4   41 002051
    "0000000000000001", -- 000000 (00000)  4   42 002052
    "0000000000000001", -- 000000 (00000)  4   43 002053
    "0000000000000001", -- 000000 (00000)  4   44 002054
    "0000000000000001", -- 000000 (00000)  4   45 002055
    "0000000000000001", -- 000000 (00000)  4   46 002056
    "0000000000000001", -- 000000 (00000)  4   47 002057
    "0000000000000001", -- 000000 (00000)  4   48 002060
    "0000000000000001", -- 000000 (00000)  4   49 002061
    "0000000000000001", -- 000000 (00000)  4   50 002062
    "0000000000000001", -- 000000 (00000)  4   51 002063
    "0000000000000001", -- 000000 (00000)  4   52 002064
    "0000000000000001", -- 000000 (00000)  4   53 002065
    "0000000000000001", -- 000000 (00000)  4   54 002066
    "0000000000000001", -- 000000 (00000)  4   55 002067
    "0000000000000001", -- 000000 (00000)  4   56 002070
    "0000000000000001", -- 000000 (00000)  4   57 002071
    "0000000000000001", -- 000000 (00000)  4   58 002072
    "0000000000000001", -- 000000 (00000)  4   59 002073
    "0000000000000001", -- 000000 (00000)  4   60 002074
    "0000000000000001", -- 000000 (00000)  4   61 002075
    "0000000000000001", -- 000000 (00000)  4   62 002076
    "0000000000000001", -- 000000 (00000)  4   63 002077
    "0000000000000001", -- 000000 (00000)  4   64 002100
    "0000000000000001", -- 000000 (00000)  4   65 002101
    "0000000000000001", -- 000000 (00000)  4   66 002102
    "0000000000000001", -- 000000 (00000)  4   67 002103
    "0000000000000001", -- 000000 (00000)  4   68 002104
    "0000000000000001", -- 000000 (00000)  4   69 002105
    "0000000000000001", -- 000000 (00000)  4   70 002106
    "0000000000000001", -- 000000 (00000)  4   71 002107
    "0000000000000001", -- 000000 (00000)  4   72 002110
    "0000000000000001", -- 000000 (00000)  4   73 002111
    "0000000000000001", -- 000000 (00000)  4   74 002112
    "0000000000000001", -- 000000 (00000)  4   75 002113
    "0000000000000001", -- 000000 (00000)  4   76 002114
    "0000000000000001", -- 000000 (00000)  4   77 002115
    "0000000000000001", -- 000000 (00000)  4   78 002116
    "0000000000000001", -- 000000 (00000)  4   79 002117
    "0000000000000001", -- 000000 (00000)  4   80 002120
    "0000000000000001", -- 000000 (00000)  4   81 002121
    "0000000000000001", -- 000000 (00000)  4   82 002122
    "0000000000000001", -- 000000 (00000)  4   83 002123
    "0000000000000001", -- 000000 (00000)  4   84 002124
    "0000000000000001", -- 000000 (00000)  4   85 002125
    "0000000000000001", -- 000000 (00000)  4   86 002126
    "0000000000000001", -- 000000 (00000)  4   87 002127
    "0000000000000001", -- 000000 (00000)  4   88 002130
    "0000000000000001", -- 000000 (00000)  4   89 002131
    "0000000000000001", -- 000000 (00000)  4   90 002132
    "0000000000000001", -- 000000 (00000)  4   91 002133
    "0000000000000001", -- 000000 (00000)  4   92 002134
    "0000000000000001", -- 000000 (00000)  4   93 002135
    "0000000000000001", -- 000000 (00000)  4   94 002136
    "0000000000000001", -- 000000 (00000)  4   95 002137
    "0000000000000001", -- 000000 (00000)  4   96 002140
    "0000000000000001", -- 000000 (00000)  4   97 002141
    "0000000000000001", -- 000000 (00000)  4   98 002142
    "0000000000000001", -- 000000 (00000)  4   99 002143
    "0000000000000001", -- 000000 (00000)  4  100 002144
    "0000000000000001", -- 000000 (00000)  4  101 002145
    "0000000000000001", -- 000000 (00000)  4  102 002146
    "0000000000000001", -- 000000 (00000)  4  103 002147
    "0000000000000001", -- 000000 (00000)  4  104 002150
    "0000000000000001", -- 000000 (00000)  4  105 002151
    "0000000000000001", -- 000000 (00000)  4  106 002152
    "0000000000000001", -- 000000 (00000)  4  107 002153
    "0000000000000001", -- 000000 (00000)  4  108 002154
    "0000000000000001", -- 000000 (00000)  4  109 002155
    "0000000000000001", -- 000000 (00000)  4  110 002156
    "0000000000000001", -- 000000 (00000)  4  111 002157
    "0000000000000001", -- 000000 (00000)  4  112 002160
    "0000000000000001", -- 000000 (00000)  4  113 002161
    "0000000000000001", -- 000000 (00000)  4  114 002162
    "0000000000000001", -- 000000 (00000)  4  115 002163
    "0000000000000001", -- 000000 (00000)  4  116 002164
    "0000000000000001", -- 000000 (00000)  4  117 002165
    "0000000000000001", -- 000000 (00000)  4  118 002166
    "0000000000000001", -- 000000 (00000)  4  119 002167
    "0000000000000001", -- 000000 (00000)  4  120 002170
    "0000000000000001", -- 000000 (00000)  4  121 002171
    "0000000000000001", -- 000000 (00000)  4  122 002172
    "0000000000000001", -- 000000 (00000)  4  123 002173
    "0000000000000001", -- 000000 (00000)  4  124 002174
    "0000000000000001", -- 000000 (00000)  4  125 002175
    "0000000000000001", -- 000000 (00000)  4  126 002176
    "0000000000000001", -- 000000 (00000)  4  127 002177
    "0000000000000001", -- 000000 (00000)  4  128 002200
    "0000000000000001", -- 000000 (00000)  4  129 002201
    "0000000000000001", -- 000000 (00000)  4  130 002202
    "0000000000000001", -- 000000 (00000)  4  131 002203
    "0000000000000001", -- 000000 (00000)  4  132 002204
    "0000000000000001", -- 000000 (00000)  4  133 002205
    "0000000000000001", -- 000000 (00000)  4  134 002206
    "0000000000000001", -- 000000 (00000)  4  135 002207
    "0000000000000001", -- 000000 (00000)  4  136 002210
    "0000000000000001", -- 000000 (00000)  4  137 002211
    "0000000000000001", -- 000000 (00000)  4  138 002212
    "0000000000000001", -- 000000 (00000)  4  139 002213
    "0000000000000001", -- 000000 (00000)  4  140 002214
    "0000000000000001", -- 000000 (00000)  4  141 002215
    "0000000000000001", -- 000000 (00000)  4  142 002216
    "0000000000000001", -- 000000 (00000)  4  143 002217
    "0000000000000001", -- 000000 (00000)  4  144 002220
    "0000000000000001", -- 000000 (00000)  4  145 002221
    "0000000000000001", -- 000000 (00000)  4  146 002222
    "0000000000000001", -- 000000 (00000)  4  147 002223
    "0000000000000001", -- 000000 (00000)  4  148 002224
    "0000000000000001", -- 000000 (00000)  4  149 002225
    "0000000000000001", -- 000000 (00000)  4  150 002226
    "0000000000000001", -- 000000 (00000)  4  151 002227
    "0000000000000001", -- 000000 (00000)  4  152 002230
    "0000000000000001", -- 000000 (00000)  4  153 002231
    "0000000000000001", -- 000000 (00000)  4  154 002232
    "0000000000000001", -- 000000 (00000)  4  155 002233
    "0000000000000001", -- 000000 (00000)  4  156 002234
    "0000000000000001", -- 000000 (00000)  4  157 002235
    "0000000000000001", -- 000000 (00000)  4  158 002236
    "0000000000000001", -- 000000 (00000)  4  159 002237
    "0000000000000001", -- 000000 (00000)  4  160 002240
    "0000000000000001", -- 000000 (00000)  4  161 002241
    "0000000000000001", -- 000000 (00000)  4  162 002242
    "0000000000000001", -- 000000 (00000)  4  163 002243
    "0000000000000001", -- 000000 (00000)  4  164 002244
    "0000000000000001", -- 000000 (00000)  4  165 002245
    "0000000000000001", -- 000000 (00000)  4  166 002246
    "0000000000000001", -- 000000 (00000)  4  167 002247
    "0000000000000001", -- 000000 (00000)  4  168 002250
    "0000000000000001", -- 000000 (00000)  4  169 002251
    "0000000000000001", -- 000000 (00000)  4  170 002252
    "0000000000000001", -- 000000 (00000)  4  171 002253
    "0000000000000001", -- 000000 (00000)  4  172 002254
    "0000000000000001", -- 000000 (00000)  4  173 002255
    "0000000000000001", -- 000000 (00000)  4  174 002256
    "0000000000000001", -- 000000 (00000)  4  175 002257
    "0000000000000001", -- 000000 (00000)  4  176 002260
    "0000000000000001", -- 000000 (00000)  4  177 002261
    "0000000000000001", -- 000000 (00000)  4  178 002262
    "0000000000000001", -- 000000 (00000)  4  179 002263
    "0000000000000001", -- 000000 (00000)  4  180 002264
    "0000000000000001", -- 000000 (00000)  4  181 002265
    "0000000000000001", -- 000000 (00000)  4  182 002266
    "0000000000000001", -- 000000 (00000)  4  183 002267
    "0000000000000001", -- 000000 (00000)  4  184 002270
    "0000000000000001", -- 000000 (00000)  4  185 002271
    "0000000000000001", -- 000000 (00000)  4  186 002272
    "0000000000000001", -- 000000 (00000)  4  187 002273
    "0000000000000001", -- 000000 (00000)  4  188 002274
    "0000000000000001", -- 000000 (00000)  4  189 002275
    "0000000000000001", -- 000000 (00000)  4  190 002276
    "0000000000000001", -- 000000 (00000)  4  191 002277
    "0000000000000001", -- 000000 (00000)  4  192 002300
    "0000000000000001", -- 000000 (00000)  4  193 002301
    "0000000000000001", -- 000000 (00000)  4  194 002302
    "0000000000000001", -- 000000 (00000)  4  195 002303
    "0000000000000001", -- 000000 (00000)  4  196 002304
    "0000000000000001", -- 000000 (00000)  4  197 002305
    "0000000000000001", -- 000000 (00000)  4  198 002306
    "0000000000000001", -- 000000 (00000)  4  199 002307
    "0000000000000001", -- 000000 (00000)  4  200 002310
    "0000000000000001", -- 000000 (00000)  4  201 002311
    "0000000000000001", -- 000000 (00000)  4  202 002312
    "0000000000000001", -- 000000 (00000)  4  203 002313
    "0000000000000001", -- 000000 (00000)  4  204 002314
    "0000000000000001", -- 000000 (00000)  4  205 002315
    "0000000000000001", -- 000000 (00000)  4  206 002316
    "0000000000000001", -- 000000 (00000)  4  207 002317
    "0000000000000001", -- 000000 (00000)  4  208 002320
    "0000000000000001", -- 000000 (00000)  4  209 002321
    "0000000000000001", -- 000000 (00000)  4  210 002322
    "0000000000000001", -- 000000 (00000)  4  211 002323
    "0000000000000001", -- 000000 (00000)  4  212 002324
    "0000000000000001", -- 000000 (00000)  4  213 002325
    "0000000000000001", -- 000000 (00000)  4  214 002326
    "0000000000000001", -- 000000 (00000)  4  215 002327
    "0000000000000001", -- 000000 (00000)  4  216 002330
    "0000000000000001", -- 000000 (00000)  4  217 002331
    "0000000000000001", -- 000000 (00000)  4  218 002332
    "0000000000000001", -- 000000 (00000)  4  219 002333
    "0000000000000001", -- 000000 (00000)  4  220 002334
    "0000000000000001", -- 000000 (00000)  4  221 002335
    "0000000000000001", -- 000000 (00000)  4  222 002336
    "0000000000000001", -- 000000 (00000)  4  223 002337
    "0000000000000001", -- 000000 (00000)  4  224 002340
    "0000000000000001", -- 000000 (00000)  4  225 002341
    "0000000000000001", -- 000000 (00000)  4  226 002342
    "0000000000000001", -- 000000 (00000)  4  227 002343
    "0000000000000001", -- 000000 (00000)  4  228 002344
    "0000000000000001", -- 000000 (00000)  4  229 002345
    "0000000000000001", -- 000000 (00000)  4  230 002346
    "0000000000000001", -- 000000 (00000)  4  231 002347
    "0000000000000001", -- 000000 (00000)  4  232 002350
    "0000000000000001", -- 000000 (00000)  4  233 002351
    "0000000000000001", -- 000000 (00000)  4  234 002352
    "0000000000000001", -- 000000 (00000)  4  235 002353
    "0000000000000001", -- 000000 (00000)  4  236 002354
    "0000000000000001", -- 000000 (00000)  4  237 002355
    "0000000000000001", -- 000000 (00000)  4  238 002356
    "0000000000000001", -- 000000 (00000)  4  239 002357
    "0000000000000001", -- 000000 (00000)  4  240 002360
    "0000000000000001", -- 000000 (00000)  4  241 002361
    "0000000000000001", -- 000000 (00000)  4  242 002362
    "0000000000000001", -- 000000 (00000)  4  243 002363
    "0000000000000001", -- 000000 (00000)  4  244 002364
    "0000000000000001", -- 000000 (00000)  4  245 002365
    "0000000000000001", -- 000000 (00000)  4  246 002366
    "0000000000000001", -- 000000 (00000)  4  247 002367
    "0000000000000001", -- 000000 (00000)  4  248 002370
    "0000000000000001", -- 000000 (00000)  4  249 002371
    "0000000000000001", -- 000000 (00000)  4  250 002372
    "0000000000000001", -- 000000 (00000)  4  251 002373
    "0000000000000001", -- 000000 (00000)  4  252 002374
    "0000000000000001", -- 000000 (00000)  4  253 002375
    "0000000000000001", -- 000000 (00000)  4  254 002376
    "0000000000000001", -- 000000 (00000)  4  255 002377
    "0000000000000001", -- 000000 (00000)  5    0 002400
    "0000000000000001", -- 000000 (00000)  5    1 002401
    "0000000000000001", -- 000000 (00000)  5    2 002402
    "0000000000000001", -- 000000 (00000)  5    3 002403
    "0000000000000001", -- 000000 (00000)  5    4 002404
    "0000000000000001", -- 000000 (00000)  5    5 002405
    "0000000000000001", -- 000000 (00000)  5    6 002406
    "0000000000000001", -- 000000 (00000)  5    7 002407
    "0000000000000001", -- 000000 (00000)  5    8 002410
    "0000000000000001", -- 000000 (00000)  5    9 002411
    "0000000000000001", -- 000000 (00000)  5   10 002412
    "0000000000000001", -- 000000 (00000)  5   11 002413
    "0000000000000001", -- 000000 (00000)  5   12 002414
    "0000000000000001", -- 000000 (00000)  5   13 002415
    "0000000000000001", -- 000000 (00000)  5   14 002416
    "0000000000000001", -- 000000 (00000)  5   15 002417
    "0000000000000001", -- 000000 (00000)  5   16 002420
    "0000000000000001", -- 000000 (00000)  5   17 002421
    "0000000000000001", -- 000000 (00000)  5   18 002422
    "0000000000000001", -- 000000 (00000)  5   19 002423
    "0000000000000001", -- 000000 (00000)  5   20 002424
    "0000000000000001", -- 000000 (00000)  5   21 002425
    "0000000000000001", -- 000000 (00000)  5   22 002426
    "0000000000000001", -- 000000 (00000)  5   23 002427
    "0000000000000001", -- 000000 (00000)  5   24 002430
    "0000000000000001", -- 000000 (00000)  5   25 002431
    "0000000000000001", -- 000000 (00000)  5   26 002432
    "0000000000000001", -- 000000 (00000)  5   27 002433
    "0000000000000001", -- 000000 (00000)  5   28 002434
    "0000000000000001", -- 000000 (00000)  5   29 002435
    "0000000000000001", -- 000000 (00000)  5   30 002436
    "0000000000000001", -- 000000 (00000)  5   31 002437
    "0000000000000001", -- 000000 (00000)  5   32 002440
    "0000000000000001", -- 000000 (00000)  5   33 002441
    "0000000000000001", -- 000000 (00000)  5   34 002442
    "0000000000000001", -- 000000 (00000)  5   35 002443
    "0000000000000001", -- 000000 (00000)  5   36 002444
    "0000000000000001", -- 000000 (00000)  5   37 002445
    "0000000000000001", -- 000000 (00000)  5   38 002446
    "0000000000000001", -- 000000 (00000)  5   39 002447
    "0000000000000001", -- 000000 (00000)  5   40 002450
    "0000000000000001", -- 000000 (00000)  5   41 002451
    "0000000000000001", -- 000000 (00000)  5   42 002452
    "0000000000000001", -- 000000 (00000)  5   43 002453
    "0000000000000001", -- 000000 (00000)  5   44 002454
    "0000000000000001", -- 000000 (00000)  5   45 002455
    "0000000000000001", -- 000000 (00000)  5   46 002456
    "0000000000000001", -- 000000 (00000)  5   47 002457
    "0000000000000001", -- 000000 (00000)  5   48 002460
    "0000000000000001", -- 000000 (00000)  5   49 002461
    "0000000000000001", -- 000000 (00000)  5   50 002462
    "0000000000000001", -- 000000 (00000)  5   51 002463
    "0000000000000001", -- 000000 (00000)  5   52 002464
    "0000000000000001", -- 000000 (00000)  5   53 002465
    "0000000000000001", -- 000000 (00000)  5   54 002466
    "0000000000000001", -- 000000 (00000)  5   55 002467
    "0000000000000001", -- 000000 (00000)  5   56 002470
    "0000000000000001", -- 000000 (00000)  5   57 002471
    "0000000000000001", -- 000000 (00000)  5   58 002472
    "0000000000000001", -- 000000 (00000)  5   59 002473
    "0000000000000001", -- 000000 (00000)  5   60 002474
    "0000000000000001", -- 000000 (00000)  5   61 002475
    "0000000000000001", -- 000000 (00000)  5   62 002476
    "0000000000000001", -- 000000 (00000)  5   63 002477
    "0000000000000001", -- 000000 (00000)  5   64 002500
    "0000000000000001", -- 000000 (00000)  5   65 002501
    "0000000000000001", -- 000000 (00000)  5   66 002502
    "0000000000000001", -- 000000 (00000)  5   67 002503
    "0000000000000001", -- 000000 (00000)  5   68 002504
    "0000000000000001", -- 000000 (00000)  5   69 002505
    "0000000000000001", -- 000000 (00000)  5   70 002506
    "0000000000000001", -- 000000 (00000)  5   71 002507
    "0000000000000001", -- 000000 (00000)  5   72 002510
    "0000000000000001", -- 000000 (00000)  5   73 002511
    "0000000000000001", -- 000000 (00000)  5   74 002512
    "0000000000000001", -- 000000 (00000)  5   75 002513
    "0000000000000001", -- 000000 (00000)  5   76 002514
    "0000000000000001", -- 000000 (00000)  5   77 002515
    "0000000000000001", -- 000000 (00000)  5   78 002516
    "0000000000000001", -- 000000 (00000)  5   79 002517
    "0000000000000001", -- 000000 (00000)  5   80 002520
    "0000000000000001", -- 000000 (00000)  5   81 002521
    "0000000000000001", -- 000000 (00000)  5   82 002522
    "0000000000000001", -- 000000 (00000)  5   83 002523
    "0000000000000001", -- 000000 (00000)  5   84 002524
    "0000000000000001", -- 000000 (00000)  5   85 002525
    "0000000000000001", -- 000000 (00000)  5   86 002526
    "0000000000000001", -- 000000 (00000)  5   87 002527
    "0000000000000001", -- 000000 (00000)  5   88 002530
    "0000000000000001", -- 000000 (00000)  5   89 002531
    "0000000000000001", -- 000000 (00000)  5   90 002532
    "0000000000000001", -- 000000 (00000)  5   91 002533
    "0000000000000001", -- 000000 (00000)  5   92 002534
    "0000000000000001", -- 000000 (00000)  5   93 002535
    "0000000000000001", -- 000000 (00000)  5   94 002536
    "0000000000000001", -- 000000 (00000)  5   95 002537
    "0000000000000001", -- 000000 (00000)  5   96 002540
    "0000000000000001", -- 000000 (00000)  5   97 002541
    "0000000000000001", -- 000000 (00000)  5   98 002542
    "0000000000000001", -- 000000 (00000)  5   99 002543
    "0000000000000001", -- 000000 (00000)  5  100 002544
    "0000000000000001", -- 000000 (00000)  5  101 002545
    "0000000000000001", -- 000000 (00000)  5  102 002546
    "0000000000000001", -- 000000 (00000)  5  103 002547
    "0000000000000001", -- 000000 (00000)  5  104 002550
    "0000000000000001", -- 000000 (00000)  5  105 002551
    "0000000000000001", -- 000000 (00000)  5  106 002552
    "0000000000000001", -- 000000 (00000)  5  107 002553
    "0000000000000001", -- 000000 (00000)  5  108 002554
    "0000000000000001", -- 000000 (00000)  5  109 002555
    "0000000000000001", -- 000000 (00000)  5  110 002556
    "0000000000000001", -- 000000 (00000)  5  111 002557
    "0000000000000001", -- 000000 (00000)  5  112 002560
    "0000000000000001", -- 000000 (00000)  5  113 002561
    "0000000000000001", -- 000000 (00000)  5  114 002562
    "0000000000000001", -- 000000 (00000)  5  115 002563
    "0000000000000001", -- 000000 (00000)  5  116 002564
    "0000000000000001", -- 000000 (00000)  5  117 002565
    "0000000000000001", -- 000000 (00000)  5  118 002566
    "0000000000000001", -- 000000 (00000)  5  119 002567
    "0000000000000001", -- 000000 (00000)  5  120 002570
    "0000000000000001", -- 000000 (00000)  5  121 002571
    "0000000000000001", -- 000000 (00000)  5  122 002572
    "0000000000000001", -- 000000 (00000)  5  123 002573
    "0000000000000001", -- 000000 (00000)  5  124 002574
    "0000000000000001", -- 000000 (00000)  5  125 002575
    "0000000000000001", -- 000000 (00000)  5  126 002576
    "0000000000000001", -- 000000 (00000)  5  127 002577
    "0000000000000001", -- 000000 (00000)  5  128 002600
    "0000000000000001", -- 000000 (00000)  5  129 002601
    "0000000000000001", -- 000000 (00000)  5  130 002602
    "0000000000000001", -- 000000 (00000)  5  131 002603
    "0000000000000001", -- 000000 (00000)  5  132 002604
    "0000000000000001", -- 000000 (00000)  5  133 002605
    "0000000000000001", -- 000000 (00000)  5  134 002606
    "0000000000000001", -- 000000 (00000)  5  135 002607
    "0000000000000001", -- 000000 (00000)  5  136 002610
    "0000000000000001", -- 000000 (00000)  5  137 002611
    "0000000000000001", -- 000000 (00000)  5  138 002612
    "0000000000000001", -- 000000 (00000)  5  139 002613
    "0000000000000001", -- 000000 (00000)  5  140 002614
    "0000000000000001", -- 000000 (00000)  5  141 002615
    "0000000000000001", -- 000000 (00000)  5  142 002616
    "0000000000000001", -- 000000 (00000)  5  143 002617
    "0000000000000001", -- 000000 (00000)  5  144 002620
    "0000000000000001", -- 000000 (00000)  5  145 002621
    "0000000000000001", -- 000000 (00000)  5  146 002622
    "0000000000000001", -- 000000 (00000)  5  147 002623
    "0000000000000001", -- 000000 (00000)  5  148 002624
    "0000000000000001", -- 000000 (00000)  5  149 002625
    "0000000000000001", -- 000000 (00000)  5  150 002626
    "0000000000000001", -- 000000 (00000)  5  151 002627
    "0000000000000001", -- 000000 (00000)  5  152 002630
    "0000000000000001", -- 000000 (00000)  5  153 002631
    "0000000000000001", -- 000000 (00000)  5  154 002632
    "0000000000000001", -- 000000 (00000)  5  155 002633
    "0000000000000001", -- 000000 (00000)  5  156 002634
    "0000000000000001", -- 000000 (00000)  5  157 002635
    "0000000000000001", -- 000000 (00000)  5  158 002636
    "0000000000000001", -- 000000 (00000)  5  159 002637
    "0000000000000001", -- 000000 (00000)  5  160 002640
    "0000000000000001", -- 000000 (00000)  5  161 002641
    "0000000000000001", -- 000000 (00000)  5  162 002642
    "0000000000000001", -- 000000 (00000)  5  163 002643
    "0000000000000001", -- 000000 (00000)  5  164 002644
    "0000000000000001", -- 000000 (00000)  5  165 002645
    "0000000000000001", -- 000000 (00000)  5  166 002646
    "0000000000000001", -- 000000 (00000)  5  167 002647
    "0000000000000001", -- 000000 (00000)  5  168 002650
    "0000000000000001", -- 000000 (00000)  5  169 002651
    "0000000000000001", -- 000000 (00000)  5  170 002652
    "0000000000000001", -- 000000 (00000)  5  171 002653
    "0000000000000001", -- 000000 (00000)  5  172 002654
    "0000000000000001", -- 000000 (00000)  5  173 002655
    "0000000000000001", -- 000000 (00000)  5  174 002656
    "0000000000000001", -- 000000 (00000)  5  175 002657
    "0000000000000001", -- 000000 (00000)  5  176 002660
    "0000000000000001", -- 000000 (00000)  5  177 002661
    "0000000000000001", -- 000000 (00000)  5  178 002662
    "0000000000000001", -- 000000 (00000)  5  179 002663
    "0000000000000001", -- 000000 (00000)  5  180 002664
    "0000000000000001", -- 000000 (00000)  5  181 002665
    "0000000000000001", -- 000000 (00000)  5  182 002666
    "0000000000000001", -- 000000 (00000)  5  183 002667
    "0000000000000001", -- 000000 (00000)  5  184 002670
    "0000000000000001", -- 000000 (00000)  5  185 002671
    "0000000000000001", -- 000000 (00000)  5  186 002672
    "0000000000000001", -- 000000 (00000)  5  187 002673
    "0000000000000001", -- 000000 (00000)  5  188 002674
    "0000000000000001", -- 000000 (00000)  5  189 002675
    "0000000000000001", -- 000000 (00000)  5  190 002676
    "0000000000000001", -- 000000 (00000)  5  191 002677
    "0000000000000001", -- 000000 (00000)  5  192 002700
    "0000000000000001", -- 000000 (00000)  5  193 002701
    "0000000000000001", -- 000000 (00000)  5  194 002702
    "0000000000000001", -- 000000 (00000)  5  195 002703
    "0000000000000001", -- 000000 (00000)  5  196 002704
    "0000000000000001", -- 000000 (00000)  5  197 002705
    "0000000000000001", -- 000000 (00000)  5  198 002706
    "0000000000000001", -- 000000 (00000)  5  199 002707
    "0000000000000001", -- 000000 (00000)  5  200 002710
    "0000000000000001", -- 000000 (00000)  5  201 002711
    "0000000000000001", -- 000000 (00000)  5  202 002712
    "0000000000000001", -- 000000 (00000)  5  203 002713
    "0000000000000001", -- 000000 (00000)  5  204 002714
    "0000000000000001", -- 000000 (00000)  5  205 002715
    "0000000000000001", -- 000000 (00000)  5  206 002716
    "0000000000000001", -- 000000 (00000)  5  207 002717
    "0000000000000001", -- 000000 (00000)  5  208 002720
    "0000000000000001", -- 000000 (00000)  5  209 002721
    "0000000000000001", -- 000000 (00000)  5  210 002722
    "0000000000000001", -- 000000 (00000)  5  211 002723
    "0000000000000001", -- 000000 (00000)  5  212 002724
    "0000000000000001", -- 000000 (00000)  5  213 002725
    "0000000000000001", -- 000000 (00000)  5  214 002726
    "0000000000000001", -- 000000 (00000)  5  215 002727
    "0000000000000001", -- 000000 (00000)  5  216 002730
    "0000000000000001", -- 000000 (00000)  5  217 002731
    "0000000000000001", -- 000000 (00000)  5  218 002732
    "0000000000000001", -- 000000 (00000)  5  219 002733
    "0000000000000001", -- 000000 (00000)  5  220 002734
    "0000000000000001", -- 000000 (00000)  5  221 002735
    "0000000000000001", -- 000000 (00000)  5  222 002736
    "0000000000000001", -- 000000 (00000)  5  223 002737
    "0000000000000001", -- 000000 (00000)  5  224 002740
    "0000000000000001", -- 000000 (00000)  5  225 002741
    "0000000000000001", -- 000000 (00000)  5  226 002742
    "0000000000000001", -- 000000 (00000)  5  227 002743
    "0000000000000001", -- 000000 (00000)  5  228 002744
    "0000000000000001", -- 000000 (00000)  5  229 002745
    "0000000000000001", -- 000000 (00000)  5  230 002746
    "0000000000000001", -- 000000 (00000)  5  231 002747
    "0000000000000001", -- 000000 (00000)  5  232 002750
    "0000000000000001", -- 000000 (00000)  5  233 002751
    "0000000000000001", -- 000000 (00000)  5  234 002752
    "0000000000000001", -- 000000 (00000)  5  235 002753
    "0000000000000001", -- 000000 (00000)  5  236 002754
    "0000000000000001", -- 000000 (00000)  5  237 002755
    "0000000000000001", -- 000000 (00000)  5  238 002756
    "0000000000000001", -- 000000 (00000)  5  239 002757
    "0000000000000001", -- 000000 (00000)  5  240 002760
    "0000000000000001", -- 000000 (00000)  5  241 002761
    "0000000000000001", -- 000000 (00000)  5  242 002762
    "0000000000000001", -- 000000 (00000)  5  243 002763
    "0000000000000001", -- 000000 (00000)  5  244 002764
    "0000000000000001", -- 000000 (00000)  5  245 002765
    "0000000000000001", -- 000000 (00000)  5  246 002766
    "0000000000000001", -- 000000 (00000)  5  247 002767
    "0000000000000001", -- 000000 (00000)  5  248 002770
    "0000000000000001", -- 000000 (00000)  5  249 002771
    "0000000000000001", -- 000000 (00000)  5  250 002772
    "0000000000000001", -- 000000 (00000)  5  251 002773
    "0000000000000001", -- 000000 (00000)  5  252 002774
    "0000000000000001", -- 000000 (00000)  5  253 002775
    "0000000000000001", -- 000000 (00000)  5  254 002776
    "0000000000000001", -- 000000 (00000)  5  255 002777
    "0000000000000001", -- 000000 (00000)  6    0 003000
    "0000000000000001", -- 000000 (00000)  6    1 003001
    "0000000000000001", -- 000000 (00000)  6    2 003002
    "0000000000000001", -- 000000 (00000)  6    3 003003
    "0000000000000001", -- 000000 (00000)  6    4 003004
    "0000000000000001", -- 000000 (00000)  6    5 003005
    "0000000000000001", -- 000000 (00000)  6    6 003006
    "0000000000000001", -- 000000 (00000)  6    7 003007
    "0000000000000001", -- 000000 (00000)  6    8 003010
    "0000000000000001", -- 000000 (00000)  6    9 003011
    "0000000000000001", -- 000000 (00000)  6   10 003012
    "0000000000000001", -- 000000 (00000)  6   11 003013
    "0000000000000001", -- 000000 (00000)  6   12 003014
    "0000000000000001", -- 000000 (00000)  6   13 003015
    "0000000000000001", -- 000000 (00000)  6   14 003016
    "0000000000000001", -- 000000 (00000)  6   15 003017
    "0000000000000001", -- 000000 (00000)  6   16 003020
    "0000000000000001", -- 000000 (00000)  6   17 003021
    "0000000000000001", -- 000000 (00000)  6   18 003022
    "0000000000000001", -- 000000 (00000)  6   19 003023
    "0000000000000001", -- 000000 (00000)  6   20 003024
    "0000000000000001", -- 000000 (00000)  6   21 003025
    "0000000000000001", -- 000000 (00000)  6   22 003026
    "0000000000000001", -- 000000 (00000)  6   23 003027
    "0000000000000001", -- 000000 (00000)  6   24 003030
    "0000000000000001", -- 000000 (00000)  6   25 003031
    "0000000000000001", -- 000000 (00000)  6   26 003032
    "0000000000000001", -- 000000 (00000)  6   27 003033
    "0000000000000001", -- 000000 (00000)  6   28 003034
    "0000000000000001", -- 000000 (00000)  6   29 003035
    "0000000000000001", -- 000000 (00000)  6   30 003036
    "0000000000000001", -- 000000 (00000)  6   31 003037
    "0000000000000001", -- 000000 (00000)  6   32 003040
    "0000000000000001", -- 000000 (00000)  6   33 003041
    "0000000000000001", -- 000000 (00000)  6   34 003042
    "0000000000000001", -- 000000 (00000)  6   35 003043
    "0000000000000001", -- 000000 (00000)  6   36 003044
    "0000000000000001", -- 000000 (00000)  6   37 003045
    "0000000000000001", -- 000000 (00000)  6   38 003046
    "0000000000000001", -- 000000 (00000)  6   39 003047
    "0000000000000001", -- 000000 (00000)  6   40 003050
    "0000000000000001", -- 000000 (00000)  6   41 003051
    "0000000000000001", -- 000000 (00000)  6   42 003052
    "0000000000000001", -- 000000 (00000)  6   43 003053
    "0000000000000001", -- 000000 (00000)  6   44 003054
    "0000000000000001", -- 000000 (00000)  6   45 003055
    "0000000000000001", -- 000000 (00000)  6   46 003056
    "0000000000000001", -- 000000 (00000)  6   47 003057
    "0000000000000001", -- 000000 (00000)  6   48 003060
    "0000000000000001", -- 000000 (00000)  6   49 003061
    "0000000000000001", -- 000000 (00000)  6   50 003062
    "0000000000000001", -- 000000 (00000)  6   51 003063
    "0000000000000001", -- 000000 (00000)  6   52 003064
    "0000000000000001", -- 000000 (00000)  6   53 003065
    "0000000000000001", -- 000000 (00000)  6   54 003066
    "0000000000000001", -- 000000 (00000)  6   55 003067
    "0000000000000001", -- 000000 (00000)  6   56 003070
    "0000000000000001", -- 000000 (00000)  6   57 003071
    "0000000000000001", -- 000000 (00000)  6   58 003072
    "0000000000000001", -- 000000 (00000)  6   59 003073
    "0000000000000001", -- 000000 (00000)  6   60 003074
    "0000000000000001", -- 000000 (00000)  6   61 003075
    "0000000000000001", -- 000000 (00000)  6   62 003076
    "0000000000000001", -- 000000 (00000)  6   63 003077
    "0000000000000001", -- 000000 (00000)  6   64 003100
    "0000000000000001", -- 000000 (00000)  6   65 003101
    "0000000000000001", -- 000000 (00000)  6   66 003102
    "0000000000000001", -- 000000 (00000)  6   67 003103
    "0000000000000001", -- 000000 (00000)  6   68 003104
    "0000000000000001", -- 000000 (00000)  6   69 003105
    "0000000000000001", -- 000000 (00000)  6   70 003106
    "0000000000000001", -- 000000 (00000)  6   71 003107
    "0000000000000001", -- 000000 (00000)  6   72 003110
    "0000000000000001", -- 000000 (00000)  6   73 003111
    "0000000000000001", -- 000000 (00000)  6   74 003112
    "0000000000000001", -- 000000 (00000)  6   75 003113
    "0000000000000001", -- 000000 (00000)  6   76 003114
    "0000000000000001", -- 000000 (00000)  6   77 003115
    "0000000000000001", -- 000000 (00000)  6   78 003116
    "0000000000000001", -- 000000 (00000)  6   79 003117
    "0000000000000001", -- 000000 (00000)  6   80 003120
    "0000000000000001", -- 000000 (00000)  6   81 003121
    "0000000000000001", -- 000000 (00000)  6   82 003122
    "0000000000000001", -- 000000 (00000)  6   83 003123
    "0000000000000001", -- 000000 (00000)  6   84 003124
    "0000000000000001", -- 000000 (00000)  6   85 003125
    "0000000000000001", -- 000000 (00000)  6   86 003126
    "0000000000000001", -- 000000 (00000)  6   87 003127
    "0000000000000001", -- 000000 (00000)  6   88 003130
    "0000000000000001", -- 000000 (00000)  6   89 003131
    "0000000000000001", -- 000000 (00000)  6   90 003132
    "0000000000000001", -- 000000 (00000)  6   91 003133
    "0000000000000001", -- 000000 (00000)  6   92 003134
    "0000000000000001", -- 000000 (00000)  6   93 003135
    "0000000000000001", -- 000000 (00000)  6   94 003136
    "0000000000000001", -- 000000 (00000)  6   95 003137
    "0000000000000001", -- 000000 (00000)  6   96 003140
    "0000000000000001", -- 000000 (00000)  6   97 003141
    "0000000000000001", -- 000000 (00000)  6   98 003142
    "0000000000000001", -- 000000 (00000)  6   99 003143
    "0000000000000001", -- 000000 (00000)  6  100 003144
    "0000000000000001", -- 000000 (00000)  6  101 003145
    "0000000000000001", -- 000000 (00000)  6  102 003146
    "0000000000000001", -- 000000 (00000)  6  103 003147
    "0000000000000001", -- 000000 (00000)  6  104 003150
    "0000000000000001", -- 000000 (00000)  6  105 003151
    "0000000000000001", -- 000000 (00000)  6  106 003152
    "0000000000000001", -- 000000 (00000)  6  107 003153
    "0000000000000001", -- 000000 (00000)  6  108 003154
    "0000000000000001", -- 000000 (00000)  6  109 003155
    "0000000000000001", -- 000000 (00000)  6  110 003156
    "0000000000000001", -- 000000 (00000)  6  111 003157
    "0000000000000001", -- 000000 (00000)  6  112 003160
    "0000000000000001", -- 000000 (00000)  6  113 003161
    "0000000000000001", -- 000000 (00000)  6  114 003162
    "0000000000000001", -- 000000 (00000)  6  115 003163
    "0000000000000001", -- 000000 (00000)  6  116 003164
    "0000000000000001", -- 000000 (00000)  6  117 003165
    "0000000000000001", -- 000000 (00000)  6  118 003166
    "0000000000000001", -- 000000 (00000)  6  119 003167
    "0000000000000001", -- 000000 (00000)  6  120 003170
    "0000000000000001", -- 000000 (00000)  6  121 003171
    "0000000000000001", -- 000000 (00000)  6  122 003172
    "0000000000000001", -- 000000 (00000)  6  123 003173
    "0000000000000001", -- 000000 (00000)  6  124 003174
    "0000000000000001", -- 000000 (00000)  6  125 003175
    "0000000000000001", -- 000000 (00000)  6  126 003176
    "0000000000000001", -- 000000 (00000)  6  127 003177
    "0000000000000001", -- 000000 (00000)  6  128 003200
    "0000000000000001", -- 000000 (00000)  6  129 003201
    "0000000000000001", -- 000000 (00000)  6  130 003202
    "0000000000000001", -- 000000 (00000)  6  131 003203
    "0000000000000001", -- 000000 (00000)  6  132 003204
    "0000000000000001", -- 000000 (00000)  6  133 003205
    "0000000000000001", -- 000000 (00000)  6  134 003206
    "0000000000000001", -- 000000 (00000)  6  135 003207
    "0000000000000001", -- 000000 (00000)  6  136 003210
    "0000000000000001", -- 000000 (00000)  6  137 003211
    "0000000000000001", -- 000000 (00000)  6  138 003212
    "0000000000000001", -- 000000 (00000)  6  139 003213
    "0000000000000001", -- 000000 (00000)  6  140 003214
    "0000000000000001", -- 000000 (00000)  6  141 003215
    "0000000000000001", -- 000000 (00000)  6  142 003216
    "0000000000000001", -- 000000 (00000)  6  143 003217
    "0000000000000001", -- 000000 (00000)  6  144 003220
    "0000000000000001", -- 000000 (00000)  6  145 003221
    "0000000000000001", -- 000000 (00000)  6  146 003222
    "0000000000000001", -- 000000 (00000)  6  147 003223
    "0000000000000001", -- 000000 (00000)  6  148 003224
    "0000000000000001", -- 000000 (00000)  6  149 003225
    "0000000000000001", -- 000000 (00000)  6  150 003226
    "0000000000000001", -- 000000 (00000)  6  151 003227
    "0000000000000001", -- 000000 (00000)  6  152 003230
    "0000000000000001", -- 000000 (00000)  6  153 003231
    "0000000000000001", -- 000000 (00000)  6  154 003232
    "0000000000000001", -- 000000 (00000)  6  155 003233
    "0000000000000001", -- 000000 (00000)  6  156 003234
    "0000000000000001", -- 000000 (00000)  6  157 003235
    "0000000000000001", -- 000000 (00000)  6  158 003236
    "0000000000000001", -- 000000 (00000)  6  159 003237
    "0000000000000001", -- 000000 (00000)  6  160 003240
    "0000000000000001", -- 000000 (00000)  6  161 003241
    "0000000000000001", -- 000000 (00000)  6  162 003242
    "0000000000000001", -- 000000 (00000)  6  163 003243
    "0000000000000001", -- 000000 (00000)  6  164 003244
    "0000000000000001", -- 000000 (00000)  6  165 003245
    "0000000000000001", -- 000000 (00000)  6  166 003246
    "0000000000000001", -- 000000 (00000)  6  167 003247
    "0000000000000001", -- 000000 (00000)  6  168 003250
    "0000000000000001", -- 000000 (00000)  6  169 003251
    "0000000000000001", -- 000000 (00000)  6  170 003252
    "0000000000000001", -- 000000 (00000)  6  171 003253
    "0000000000000001", -- 000000 (00000)  6  172 003254
    "0000000000000001", -- 000000 (00000)  6  173 003255
    "0000000000000001", -- 000000 (00000)  6  174 003256
    "0000000000000001", -- 000000 (00000)  6  175 003257
    "0000000000000001", -- 000000 (00000)  6  176 003260
    "0000000000000001", -- 000000 (00000)  6  177 003261
    "0000000000000001", -- 000000 (00000)  6  178 003262
    "0000000000000001", -- 000000 (00000)  6  179 003263
    "0000000000000001", -- 000000 (00000)  6  180 003264
    "0000000000000001", -- 000000 (00000)  6  181 003265
    "0000000000000001", -- 000000 (00000)  6  182 003266
    "0000000000000001", -- 000000 (00000)  6  183 003267
    "0000000000000001", -- 000000 (00000)  6  184 003270
    "0000000000000001", -- 000000 (00000)  6  185 003271
    "0000000000000001", -- 000000 (00000)  6  186 003272
    "0000000000000001", -- 000000 (00000)  6  187 003273
    "0000000000000001", -- 000000 (00000)  6  188 003274
    "0000000000000001", -- 000000 (00000)  6  189 003275
    "0000000000000001", -- 000000 (00000)  6  190 003276
    "0000000000000001", -- 000000 (00000)  6  191 003277
    "0000000000000001", -- 000000 (00000)  6  192 003300
    "0000000000000001", -- 000000 (00000)  6  193 003301
    "0000000000000001", -- 000000 (00000)  6  194 003302
    "0000000000000001", -- 000000 (00000)  6  195 003303
    "0000000000000001", -- 000000 (00000)  6  196 003304
    "0000000000000001", -- 000000 (00000)  6  197 003305
    "0000000000000001", -- 000000 (00000)  6  198 003306
    "0000000000000001", -- 000000 (00000)  6  199 003307
    "0000000000000001", -- 000000 (00000)  6  200 003310
    "0000000000000001", -- 000000 (00000)  6  201 003311
    "0000000000000001", -- 000000 (00000)  6  202 003312
    "0000000000000001", -- 000000 (00000)  6  203 003313
    "0000000000000001", -- 000000 (00000)  6  204 003314
    "0000000000000001", -- 000000 (00000)  6  205 003315
    "0000000000000001", -- 000000 (00000)  6  206 003316
    "0000000000000001", -- 000000 (00000)  6  207 003317
    "0000000000000001", -- 000000 (00000)  6  208 003320
    "0000000000000001", -- 000000 (00000)  6  209 003321
    "0000000000000001", -- 000000 (00000)  6  210 003322
    "0000000000000001", -- 000000 (00000)  6  211 003323
    "0000000000000001", -- 000000 (00000)  6  212 003324
    "0000000000000001", -- 000000 (00000)  6  213 003325
    "0000000000000001", -- 000000 (00000)  6  214 003326
    "0000000000000001", -- 000000 (00000)  6  215 003327
    "0000000000000001", -- 000000 (00000)  6  216 003330
    "0000000000000001", -- 000000 (00000)  6  217 003331
    "0000000000000001", -- 000000 (00000)  6  218 003332
    "0000000000000001", -- 000000 (00000)  6  219 003333
    "0000000000000001", -- 000000 (00000)  6  220 003334
    "0000000000000001", -- 000000 (00000)  6  221 003335
    "0000000000000001", -- 000000 (00000)  6  222 003336
    "0000000000000001", -- 000000 (00000)  6  223 003337
    "0000000000000001", -- 000000 (00000)  6  224 003340
    "0000000000000001", -- 000000 (00000)  6  225 003341
    "0000000000000001", -- 000000 (00000)  6  226 003342
    "0000000000000001", -- 000000 (00000)  6  227 003343
    "0000000000000001", -- 000000 (00000)  6  228 003344
    "0000000000000001", -- 000000 (00000)  6  229 003345
    "0000000000000001", -- 000000 (00000)  6  230 003346
    "0000000000000001", -- 000000 (00000)  6  231 003347
    "0000000000000001", -- 000000 (00000)  6  232 003350
    "0000000000000001", -- 000000 (00000)  6  233 003351
    "0000000000000001", -- 000000 (00000)  6  234 003352
    "0000000000000001", -- 000000 (00000)  6  235 003353
    "0000000000000001", -- 000000 (00000)  6  236 003354
    "0000000000000001", -- 000000 (00000)  6  237 003355
    "0000000000000001", -- 000000 (00000)  6  238 003356
    "0000000000000001", -- 000000 (00000)  6  239 003357
    "0000000000000001", -- 000000 (00000)  6  240 003360
    "0000000000000001", -- 000000 (00000)  6  241 003361
    "0000000000000001", -- 000000 (00000)  6  242 003362
    "0000000000000001", -- 000000 (00000)  6  243 003363
    "0000000000000001", -- 000000 (00000)  6  244 003364
    "0000000000000001", -- 000000 (00000)  6  245 003365
    "0000000000000001", -- 000000 (00000)  6  246 003366
    "0000000000000001", -- 000000 (00000)  6  247 003367
    "0000000000000001", -- 000000 (00000)  6  248 003370
    "0000000000000001", -- 000000 (00000)  6  249 003371
    "0000000000000001", -- 000000 (00000)  6  250 003372
    "0000000000000001", -- 000000 (00000)  6  251 003373
    "0000000000000001", -- 000000 (00000)  6  252 003374
    "0000000000000001", -- 000000 (00000)  6  253 003375
    "0000000000000001", -- 000000 (00000)  6  254 003376
    "0000000000000001", -- 000000 (00000)  6  255 003377
    "0000000000000001", -- 000000 (00000)  7    0 003400
    "0000000000000001", -- 000000 (00000)  7    1 003401
    "0000000000000001", -- 000000 (00000)  7    2 003402
    "0000000000000001", -- 000000 (00000)  7    3 003403
    "0000000000000001", -- 000000 (00000)  7    4 003404
    "0000000000000001", -- 000000 (00000)  7    5 003405
    "0000000000000001", -- 000000 (00000)  7    6 003406
    "0000000000000001", -- 000000 (00000)  7    7 003407
    "0000000000000001", -- 000000 (00000)  7    8 003410
    "0000000000000001", -- 000000 (00000)  7    9 003411
    "0000000000000001", -- 000000 (00000)  7   10 003412
    "0000000000000001", -- 000000 (00000)  7   11 003413
    "0000000000000001", -- 000000 (00000)  7   12 003414
    "0000000000000001", -- 000000 (00000)  7   13 003415
    "0000000000000001", -- 000000 (00000)  7   14 003416
    "0000000000000001", -- 000000 (00000)  7   15 003417
    "0000000000000001", -- 000000 (00000)  7   16 003420
    "0000000000000001", -- 000000 (00000)  7   17 003421
    "0000000000000001", -- 000000 (00000)  7   18 003422
    "0000000000000001", -- 000000 (00000)  7   19 003423
    "0000000000000001", -- 000000 (00000)  7   20 003424
    "0000000000000001", -- 000000 (00000)  7   21 003425
    "0000000000000001", -- 000000 (00000)  7   22 003426
    "0000000000000001", -- 000000 (00000)  7   23 003427
    "0000000000000001", -- 000000 (00000)  7   24 003430
    "0000000000000001", -- 000000 (00000)  7   25 003431
    "0000000000000001", -- 000000 (00000)  7   26 003432
    "0000000000000001", -- 000000 (00000)  7   27 003433
    "0000000000000001", -- 000000 (00000)  7   28 003434
    "0000000000000001", -- 000000 (00000)  7   29 003435
    "0000000000000001", -- 000000 (00000)  7   30 003436
    "0000000000000001", -- 000000 (00000)  7   31 003437
    "0000000000000001", -- 000000 (00000)  7   32 003440
    "0000000000000001", -- 000000 (00000)  7   33 003441
    "0000000000000001", -- 000000 (00000)  7   34 003442
    "0000000000000001", -- 000000 (00000)  7   35 003443
    "0000000000000001", -- 000000 (00000)  7   36 003444
    "0000000000000001", -- 000000 (00000)  7   37 003445
    "0000000000000001", -- 000000 (00000)  7   38 003446
    "0000000000000001", -- 000000 (00000)  7   39 003447
    "0000000000000001", -- 000000 (00000)  7   40 003450
    "0000000000000001", -- 000000 (00000)  7   41 003451
    "0000000000000001", -- 000000 (00000)  7   42 003452
    "0000000000000001", -- 000000 (00000)  7   43 003453
    "0000000000000001", -- 000000 (00000)  7   44 003454
    "0000000000000001", -- 000000 (00000)  7   45 003455
    "0000000000000001", -- 000000 (00000)  7   46 003456
    "0000000000000001", -- 000000 (00000)  7   47 003457
    "0000000000000001", -- 000000 (00000)  7   48 003460
    "0000000000000001", -- 000000 (00000)  7   49 003461
    "0000000000000001", -- 000000 (00000)  7   50 003462
    "0000000000000001", -- 000000 (00000)  7   51 003463
    "0000000000000001", -- 000000 (00000)  7   52 003464
    "0000000000000001", -- 000000 (00000)  7   53 003465
    "0000000000000001", -- 000000 (00000)  7   54 003466
    "0000000000000001", -- 000000 (00000)  7   55 003467
    "0000000000000001", -- 000000 (00000)  7   56 003470
    "0000000000000001", -- 000000 (00000)  7   57 003471
    "0000000000000001", -- 000000 (00000)  7   58 003472
    "0000000000000001", -- 000000 (00000)  7   59 003473
    "0000000000000001", -- 000000 (00000)  7   60 003474
    "0000000000000001", -- 000000 (00000)  7   61 003475
    "0000000000000001", -- 000000 (00000)  7   62 003476
    "0000000000000001", -- 000000 (00000)  7   63 003477
    "0000000000000001", -- 000000 (00000)  7   64 003500
    "0000000000000001", -- 000000 (00000)  7   65 003501
    "0000000000000001", -- 000000 (00000)  7   66 003502
    "0000000000000001", -- 000000 (00000)  7   67 003503
    "0000000000000001", -- 000000 (00000)  7   68 003504
    "0000000000000001", -- 000000 (00000)  7   69 003505
    "0000000000000001", -- 000000 (00000)  7   70 003506
    "0000000000000001", -- 000000 (00000)  7   71 003507
    "0000000000000001", -- 000000 (00000)  7   72 003510
    "0000000000000001", -- 000000 (00000)  7   73 003511
    "0000000000000001", -- 000000 (00000)  7   74 003512
    "0000000000000001", -- 000000 (00000)  7   75 003513
    "0000000000000001", -- 000000 (00000)  7   76 003514
    "0000000000000001", -- 000000 (00000)  7   77 003515
    "0000000000000001", -- 000000 (00000)  7   78 003516
    "0000000000000001", -- 000000 (00000)  7   79 003517
    "0000000000000001", -- 000000 (00000)  7   80 003520
    "0000000000000001", -- 000000 (00000)  7   81 003521
    "0000000000000001", -- 000000 (00000)  7   82 003522
    "0000000000000001", -- 000000 (00000)  7   83 003523
    "0000000000000001", -- 000000 (00000)  7   84 003524
    "0000000000000001", -- 000000 (00000)  7   85 003525
    "0000000000000001", -- 000000 (00000)  7   86 003526
    "0000000000000001", -- 000000 (00000)  7   87 003527
    "0000000000000001", -- 000000 (00000)  7   88 003530
    "0000000000000001", -- 000000 (00000)  7   89 003531
    "0000000000000001", -- 000000 (00000)  7   90 003532
    "0000000000000001", -- 000000 (00000)  7   91 003533
    "0000000000000001", -- 000000 (00000)  7   92 003534
    "0000000000000001", -- 000000 (00000)  7   93 003535
    "0000000000000001", -- 000000 (00000)  7   94 003536
    "0000000000000001", -- 000000 (00000)  7   95 003537
    "0000000000000001", -- 000000 (00000)  7   96 003540
    "0000000000000001", -- 000000 (00000)  7   97 003541
    "0000000000000001", -- 000000 (00000)  7   98 003542
    "0000000000000001", -- 000000 (00000)  7   99 003543
    "0000000000000001", -- 000000 (00000)  7  100 003544
    "0000000000000001", -- 000000 (00000)  7  101 003545
    "0000000000000001", -- 000000 (00000)  7  102 003546
    "0000000000000001", -- 000000 (00000)  7  103 003547
    "0000000000000001", -- 000000 (00000)  7  104 003550
    "0000000000000001", -- 000000 (00000)  7  105 003551
    "0000000000000001", -- 000000 (00000)  7  106 003552
    "0000000000000001", -- 000000 (00000)  7  107 003553
    "0000000000000001", -- 000000 (00000)  7  108 003554
    "0000000000000001", -- 000000 (00000)  7  109 003555
    "0000000000000001", -- 000000 (00000)  7  110 003556
    "0000000000000001", -- 000000 (00000)  7  111 003557
    "0000000000000001", -- 000000 (00000)  7  112 003560
    "0000000000000001", -- 000000 (00000)  7  113 003561
    "0000000000000001", -- 000000 (00000)  7  114 003562
    "0000000000000001", -- 000000 (00000)  7  115 003563
    "0000000000000001", -- 000000 (00000)  7  116 003564
    "0000000000000001", -- 000000 (00000)  7  117 003565
    "0000000000000001", -- 000000 (00000)  7  118 003566
    "0000000000000001", -- 000000 (00000)  7  119 003567
    "0000000000000001", -- 000000 (00000)  7  120 003570
    "0000000000000001", -- 000000 (00000)  7  121 003571
    "0000000000000001", -- 000000 (00000)  7  122 003572
    "0000000000000001", -- 000000 (00000)  7  123 003573
    "0000000000000001", -- 000000 (00000)  7  124 003574
    "0000000000000001", -- 000000 (00000)  7  125 003575
    "0000000000000001", -- 000000 (00000)  7  126 003576
    "0000000000000001", -- 000000 (00000)  7  127 003577
    "0000000000000001", -- 000000 (00000)  7  128 003600
    "0000000000000001", -- 000000 (00000)  7  129 003601
    "0000000000000001", -- 000000 (00000)  7  130 003602
    "0000000000000001", -- 000000 (00000)  7  131 003603
    "0000000000000001", -- 000000 (00000)  7  132 003604
    "0000000000000001", -- 000000 (00000)  7  133 003605
    "0000000000000001", -- 000000 (00000)  7  134 003606
    "0000000000000001", -- 000000 (00000)  7  135 003607
    "0000000000000001", -- 000000 (00000)  7  136 003610
    "0000000000000001", -- 000000 (00000)  7  137 003611
    "0000000000000001", -- 000000 (00000)  7  138 003612
    "0000000000000001", -- 000000 (00000)  7  139 003613
    "0000000000000001", -- 000000 (00000)  7  140 003614
    "0000000000000001", -- 000000 (00000)  7  141 003615
    "0000000000000001", -- 000000 (00000)  7  142 003616
    "0000000000000001", -- 000000 (00000)  7  143 003617
    "0000000000000001", -- 000000 (00000)  7  144 003620
    "0000000000000001", -- 000000 (00000)  7  145 003621
    "0000000000000001", -- 000000 (00000)  7  146 003622
    "0000000000000001", -- 000000 (00000)  7  147 003623
    "0000000000000001", -- 000000 (00000)  7  148 003624
    "0000000000000001", -- 000000 (00000)  7  149 003625
    "0000000000000001", -- 000000 (00000)  7  150 003626
    "0000000000000001", -- 000000 (00000)  7  151 003627
    "0000000000000001", -- 000000 (00000)  7  152 003630
    "0000000000000001", -- 000000 (00000)  7  153 003631
    "0000000000000001", -- 000000 (00000)  7  154 003632
    "0000000000000001", -- 000000 (00000)  7  155 003633
    "0000000000000001", -- 000000 (00000)  7  156 003634
    "0000000000000001", -- 000000 (00000)  7  157 003635
    "0000000000000001", -- 000000 (00000)  7  158 003636
    "0000000000000001", -- 000000 (00000)  7  159 003637
    "0000000000000001", -- 000000 (00000)  7  160 003640
    "0000000000000001", -- 000000 (00000)  7  161 003641
    "0000000000000001", -- 000000 (00000)  7  162 003642
    "0000000000000001", -- 000000 (00000)  7  163 003643
    "0000000000000001", -- 000000 (00000)  7  164 003644
    "0000000000000001", -- 000000 (00000)  7  165 003645
    "0000000000000001", -- 000000 (00000)  7  166 003646
    "0000000000000001", -- 000000 (00000)  7  167 003647
    "0000000000000001", -- 000000 (00000)  7  168 003650
    "0000000000000001", -- 000000 (00000)  7  169 003651
    "0000000000000001", -- 000000 (00000)  7  170 003652
    "0000000000000001", -- 000000 (00000)  7  171 003653
    "0000000000000001", -- 000000 (00000)  7  172 003654
    "0000000000000001", -- 000000 (00000)  7  173 003655
    "0000000000000001", -- 000000 (00000)  7  174 003656
    "0000000000000001", -- 000000 (00000)  7  175 003657
    "0000000000000001", -- 000000 (00000)  7  176 003660
    "0000000000000001", -- 000000 (00000)  7  177 003661
    "0000000000000001", -- 000000 (00000)  7  178 003662
    "0000000000000001", -- 000000 (00000)  7  179 003663
    "0000000000000001", -- 000000 (00000)  7  180 003664
    "0000000000000001", -- 000000 (00000)  7  181 003665
    "0000000000000001", -- 000000 (00000)  7  182 003666
    "0000000000000001", -- 000000 (00000)  7  183 003667
    "0000000000000001", -- 000000 (00000)  7  184 003670
    "0000000000000001", -- 000000 (00000)  7  185 003671
    "0000000000000001", -- 000000 (00000)  7  186 003672
    "0000000000000001", -- 000000 (00000)  7  187 003673
    "0000000000000001", -- 000000 (00000)  7  188 003674
    "0000000000000001", -- 000000 (00000)  7  189 003675
    "0000000000000001", -- 000000 (00000)  7  190 003676
    "0000000000000001", -- 000000 (00000)  7  191 003677
    "0000000000000001", -- 000000 (00000)  7  192 003700
    "0000000000000001", -- 000000 (00000)  7  193 003701
    "0000000000000001", -- 000000 (00000)  7  194 003702
    "0000000000000001", -- 000000 (00000)  7  195 003703
    "0000000000000001", -- 000000 (00000)  7  196 003704
    "0000000000000001", -- 000000 (00000)  7  197 003705
    "0000000000000001", -- 000000 (00000)  7  198 003706
    "0000000000000001", -- 000000 (00000)  7  199 003707
    "0000000000000001", -- 000000 (00000)  7  200 003710
    "0000000000000001", -- 000000 (00000)  7  201 003711
    "0000000000000001", -- 000000 (00000)  7  202 003712
    "0000000000000001", -- 000000 (00000)  7  203 003713
    "0000000000000001", -- 000000 (00000)  7  204 003714
    "0000000000000001", -- 000000 (00000)  7  205 003715
    "0000000000000001", -- 000000 (00000)  7  206 003716
    "0000000000000001", -- 000000 (00000)  7  207 003717
    "0000000000000001", -- 000000 (00000)  7  208 003720
    "0000000000000001", -- 000000 (00000)  7  209 003721
    "0000000000000001", -- 000000 (00000)  7  210 003722
    "0000000000000001", -- 000000 (00000)  7  211 003723
    "0000000000000001", -- 000000 (00000)  7  212 003724
    "0000000000000001", -- 000000 (00000)  7  213 003725
    "0000000000000001", -- 000000 (00000)  7  214 003726
    "0000000000000001", -- 000000 (00000)  7  215 003727
    "0000000000000001", -- 000000 (00000)  7  216 003730
    "0000000000000001", -- 000000 (00000)  7  217 003731
    "0000000000000001", -- 000000 (00000)  7  218 003732
    "0000000000000001", -- 000000 (00000)  7  219 003733
    "0000000000000001", -- 000000 (00000)  7  220 003734
    "0000000000000001", -- 000000 (00000)  7  221 003735
    "0000000000000001", -- 000000 (00000)  7  222 003736
    "0000000000000001", -- 000000 (00000)  7  223 003737
    "0000000000000001", -- 000000 (00000)  7  224 003740
    "0000000000000001", -- 000000 (00000)  7  225 003741
    "0000000000000001", -- 000000 (00000)  7  226 003742
    "0000000000000001", -- 000000 (00000)  7  227 003743
    "0000000000000001", -- 000000 (00000)  7  228 003744
    "0000000000000001", -- 000000 (00000)  7  229 003745
    "0000000000000001", -- 000000 (00000)  7  230 003746
    "0000000000000001", -- 000000 (00000)  7  231 003747
    "0000000000000001", -- 000000 (00000)  7  232 003750
    "0000000000000001", -- 000000 (00000)  7  233 003751
    "0000000000000001", -- 000000 (00000)  7  234 003752
    "0000000000000001", -- 000000 (00000)  7  235 003753
    "0000000000000001", -- 000000 (00000)  7  236 003754
    "0000000000000001", -- 000000 (00000)  7  237 003755
    "0000000000000001", -- 000000 (00000)  7  238 003756
    "0000000000000001", -- 000000 (00000)  7  239 003757
    "0000000000000001", -- 000000 (00000)  7  240 003760
    "0000000000000001", -- 000000 (00000)  7  241 003761
    "0000000000000001", -- 000000 (00000)  7  242 003762
    "0000000000000001", -- 000000 (00000)  7  243 003763
    "0000000000000001", -- 000000 (00000)  7  244 003764
    "0000000000000001", -- 000000 (00000)  7  245 003765
    "0000000000000001", -- 000000 (00000)  7  246 003766
    "0000000000000001", -- 000000 (00000)  7  247 003767
    "0000000000000001", -- 000000 (00000)  7  248 003770
    "0000000000000001", -- 000000 (00000)  7  249 003771
    "0000000000000001", -- 000000 (00000)  7  250 003772
    "0000000000000001", -- 000000 (00000)  7  251 003773
    "0000000000000001", -- 000000 (00000)  7  252 003774
    "0000000000000001", -- 000000 (00000)  7  253 003775
    "0000000000000001", -- 000000 (00000)  7  254 003776
    "0000000000000001"  -- 000000 (00000)  7  255 003777
  );

begin

  process( clka, wea, addra, dina ) is
  begin
  
    if rising_edge( clka ) then
	 
      if wea(0) = '1' then

        -- Perform a write.
        CORES( conv_integer(addra) ) <= dina;

      else
      
        -- Perform the read.
        -- doutb <= CORES( conv_integer(addrb) );

      end if; -- wea

    end if; -- clka
	 
  end process;
  
  process( clkb, addrb ) is
  begin

    if rising_edge( clkb ) then
    
      doutb <= CORES( conv_integer(addrb) );
      
    end if; -- clkb
    
  end process;
  
  -- doutb <= CORES( conv_integer(addrb) );

end Rtl;

-- **********************
-- ***                ***
-- ***  END OF FILE.  ***
-- ***                ***
-- **********************


