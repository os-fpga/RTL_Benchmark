`ifdef ATCIIC100_CONFIG_VH
`else
//	`define ATCIIC100_FIFO_DEPTH_2
	`define ATCIIC100_FIFO_DEPTH_4
//	`define ATCIIC100_FIFO_DEPTH_8
//	`define ATCIIC100_FIFO_DEPTH_16
`endif
