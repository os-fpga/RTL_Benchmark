// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: data_output_sequencer.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2016-04-18-EP on Sat Apr 27 13:59:59 2019
//=============================================================================
// Description: Sequencer for data_output
//=============================================================================

`ifndef DATA_OUTPUT_SEQUENCER_SV
`define DATA_OUTPUT_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(output_tx) data_output_sequencer_t;


`endif // DATA_OUTPUT_SEQUENCER_SV

