--
-- crc32_fast512_tab.vhd: A 32-bit CRC (IEEE) table for processing fixed 512 bits in parallel
-- Copyright (C) 2011 CESNET
-- Author(s): Lukas Kekely <xkekel00@stud.fit.vutbr.cz>
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in
--    the documentation and/or other materials provided with the
--    distribution.
-- 3. Neither the name of the Company nor the names of its contributors
--    may be used to endorse or promote products derived from this
--    software without specific prior written permission.
--
-- This software is provided ``as is'', and any express or implied
-- warranties, including, but not limited to, the implied warranties of
-- merchantability and fitness for a particular purpose are disclaimed.
-- In no event shall the company or contributors be liable for any
-- direct, indirect, incidental, special, exemplary, or consequential
-- damages (including, but not limited to, procurement of substitute
-- goods or services; loss of use, data, or profits; or business
-- interruption) however caused and on any theory of liability, whether
-- in contract, strict liability, or tort (including negligence or
-- otherwise) arising in any way out of the use of this software, even
-- if advised of the possibility of such damage.
--
-- $Id$
--
-- TODO:
--
--

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.numeric_std.all;
use WORK.math_pack.all;
-- ----------------------------------------------------------------------------
--                        Entity declaration
-- ----------------------------------------------------------------------------
entity crc32_fast512_tab is
   port(
      DI    : in  std_logic_vector(512-1 downto 0);
      DO    : out std_logic_vector(31 downto 0)
   );
end entity crc32_fast512_tab;

-- ----------------------------------------------------------------------------
--                      Architecture declaration
-- ----------------------------------------------------------------------------
architecture arch of crc32_fast512_tab is
begin
-- 32-bit CRC equations processing 512 bits in parallel (VHDL code)
-- Generator polynomial: 0x104C11DB7
   DO(0) <= DI(64) XOR DI(488) XOR DI(236) XOR DI(75) XOR DI(257) XOR DI(264) XOR DI(394) XOR DI(356) XOR DI(195) XOR DI(76) XOR DI(322) XOR DI(483) XOR DI(285) XOR DI(343) XOR DI(60) XOR DI(467) XOR DI(47) XOR DI(428) XOR DI(413) XOR DI(177) XOR DI(361) XOR DI(63) XOR DI(284) XOR DI(414) XOR DI(326) XOR DI(464) XOR DI(253) XOR DI(222) XOR DI(100) XOR DI(329) XOR DI(484) XOR DI(346) XOR DI(50) XOR DI(457) XOR DI(454) XOR DI(243) XOR DI(319) XOR DI(40) XOR DI(447) XOR DI(444) XOR DI(126) XOR DI(68) XOR DI(192) XOR DI(225) XOR DI(93) XOR DI(136) XOR DI(190) XOR DI(121) XOR DI(398) XOR DI(468) XOR DI(330) XOR DI(174) XOR DI(401) XOR DI(486) XOR DI(286) XOR DI(19) XOR DI(415) XOR DI(78) XOR DI(288) XOR DI(124) XOR DI(465) XOR DI(202) XOR DI(32) XOR DI(429) XOR DI(417) XOR DI(163) XOR DI(502) XOR DI(248) XOR DI(255) XOR DI(385) XOR DI(51) XOR DI(275) XOR DI(244) XOR DI(213) XOR DI(310) XOR DI(31) XOR DI(112) XOR DI(321) XOR DI(10) XOR DI(406) XOR DI(193) XOR DI(154) XOR DI(239) XOR DI(376) XOR DI(235) XOR DI(22) XOR DI(103) XOR DI(1) XOR DI(226) XOR DI(217) XOR DI(368) XOR DI(302) XOR DI(377) XOR DI(215) XOR DI(122) XOR DI(375) XOR DI(146) XOR DI(96) XOR DI(341) XOR DI(399) XOR DI(311) XOR DI(449) XOR DI(35) XOR DI(175) XOR DI(386) XOR DI(487) XOR DI(260) XOR DI(224) XOR DI(200) XOR DI(131) XOR DI(384) XOR DI(416) XOR DI(155) XOR DI(79) XOR DI(105) XOR DI(300) XOR DI(354) XOR DI(33) XOR DI(150) XOR DI(430) XOR DI(104) XOR DI(431) XOR DI(342) XOR DI(2) XOR DI(21) XOR DI(418) XOR DI(170) XOR DI(503) XOR DI(482) XOR DI(251) XOR DI(350) XOR DI(54) XOR DI(171) XOR DI(278) XOR DI(408) XOR DI(320) XOR DI(458) XOR DI(247) XOR DI(216) XOR DI(94) XOR DI(478) XOR DI(340) XOR DI(44) XOR DI(451) XOR DI(313) XOR DI(120) XOR DI(62) XOR DI(184) XOR DI(462) XOR DI(324) XOR DI(168) XOR DI(395) XOR DI(480) XOR DI(409) XOR DI(282) XOR DI(459) XOR DI(26) XOR DI(411) XOR DI(496) XOR DI(269) XOR DI(238) XOR DI(207) XOR DI(304) XOR DI(315) XOR DI(4) XOR DI(233) XOR DI(229) XOR DI(220) XOR DI(296) XOR DI(209) XOR DI(116) XOR DI(369) XOR DI(140) XOR DI(90) XOR DI(393) XOR DI(305) XOR DI(29) XOR DI(380) XOR DI(481) XOR DI(218) XOR DI(194) XOR DI(125) XOR DI(378) XOR DI(149) XOR DI(144) XOR DI(98) XOR DI(425) XOR DI(164) XOR DI(48) XOR DI(165) XOR DI(402) XOR DI(314) XOR DI(452) XOR DI(210) XOR DI(88) XOR DI(445) XOR DI(114) XOR DI(178) XOR DI(318) XOR DI(389) XOR DI(20) XOR DI(298) XOR DI(309) XOR DI(214) XOR DI(203) XOR DI(363) XOR DI(134) XOR DI(387) XOR DI(23) XOR DI(475) XOR DI(212) XOR DI(119) XOR DI(143) XOR DI(138) XOR DI(42) XOR DI(159) XOR DI(396) XOR DI(446) XOR DI(439) XOR DI(108) XOR DI(303) XOR DI(197) XOR DI(357) XOR DI(17) XOR DI(113) XOR DI(36) XOR DI(153) XOR DI(440) XOR DI(433) XOR DI(191) XOR DI(351) XOR DI(11) XOR DI(107) XOR DI(30) XOR DI(427) XOR DI(185) XOR DI(345) XOR DI(5) XOR DI(24) XOR DI(179) XOR DI(18) XOR DI(173) XOR DI(12) XOR DI(167) XOR DI(6) XOR DI(0) XOR DI(500) XOR DI(506);
   DO(1) <= DI(65) XOR DI(489) XOR DI(237) XOR DI(76) XOR DI(258) XOR DI(265) XOR DI(395) XOR DI(357) XOR DI(196) XOR DI(77) XOR DI(323) XOR DI(484) XOR DI(286) XOR DI(344) XOR DI(61) XOR DI(468) XOR DI(48) XOR DI(429) XOR DI(414) XOR DI(178) XOR DI(362) XOR DI(64) XOR DI(285) XOR DI(415) XOR DI(327) XOR DI(465) XOR DI(254) XOR DI(223) XOR DI(101) XOR DI(330) XOR DI(485) XOR DI(347) XOR DI(51) XOR DI(458) XOR DI(455) XOR DI(244) XOR DI(320) XOR DI(41) XOR DI(448) XOR DI(445) XOR DI(127) XOR DI(69) XOR DI(193) XOR DI(226) XOR DI(94) XOR DI(137) XOR DI(191) XOR DI(122) XOR DI(399) XOR DI(469) XOR DI(331) XOR DI(175) XOR DI(402) XOR DI(487) XOR DI(287) XOR DI(20) XOR DI(416) XOR DI(79) XOR DI(289) XOR DI(125) XOR DI(466) XOR DI(203) XOR DI(33) XOR DI(430) XOR DI(418) XOR DI(164) XOR DI(503) XOR DI(249) XOR DI(256) XOR DI(386) XOR DI(52) XOR DI(276) XOR DI(245) XOR DI(214) XOR DI(311) XOR DI(32) XOR DI(113) XOR DI(322) XOR DI(11) XOR DI(407) XOR DI(194) XOR DI(155) XOR DI(240) XOR DI(377) XOR DI(236) XOR DI(23) XOR DI(104) XOR DI(2) XOR DI(227) XOR DI(218) XOR DI(369) XOR DI(303) XOR DI(378) XOR DI(216) XOR DI(123) XOR DI(376) XOR DI(147) XOR DI(97) XOR DI(342) XOR DI(400) XOR DI(312) XOR DI(450) XOR DI(36) XOR DI(176) XOR DI(387) XOR DI(488) XOR DI(261) XOR DI(225) XOR DI(201) XOR DI(132) XOR DI(385) XOR DI(417) XOR DI(156) XOR DI(80) XOR DI(106) XOR DI(301) XOR DI(355) XOR DI(34) XOR DI(151) XOR DI(431) XOR DI(105) XOR DI(432) XOR DI(343) XOR DI(3) XOR DI(22) XOR DI(419) XOR DI(171) XOR DI(504) XOR DI(483) XOR DI(252) XOR DI(351) XOR DI(55) XOR DI(172) XOR DI(279) XOR DI(409) XOR DI(321) XOR DI(459) XOR DI(248) XOR DI(217) XOR DI(95) XOR DI(479) XOR DI(341) XOR DI(45) XOR DI(452) XOR DI(314) XOR DI(121) XOR DI(63) XOR DI(185) XOR DI(463) XOR DI(325) XOR DI(169) XOR DI(396) XOR DI(481) XOR DI(410) XOR DI(283) XOR DI(460) XOR DI(27) XOR DI(412) XOR DI(497) XOR DI(270) XOR DI(239) XOR DI(208) XOR DI(305) XOR DI(316) XOR DI(5) XOR DI(234) XOR DI(230) XOR DI(221) XOR DI(297) XOR DI(210) XOR DI(117) XOR DI(370) XOR DI(141) XOR DI(91) XOR DI(394) XOR DI(306) XOR DI(30) XOR DI(381) XOR DI(482) XOR DI(219) XOR DI(195) XOR DI(126) XOR DI(379) XOR DI(150) XOR DI(145) XOR DI(99) XOR DI(426) XOR DI(165) XOR DI(49) XOR DI(166) XOR DI(403) XOR DI(315) XOR DI(453) XOR DI(211) XOR DI(89) XOR DI(446) XOR DI(115) XOR DI(179) XOR DI(319) XOR DI(390) XOR DI(21) XOR DI(299) XOR DI(310) XOR DI(215) XOR DI(204) XOR DI(364) XOR DI(135) XOR DI(388) XOR DI(24) XOR DI(476) XOR DI(213) XOR DI(120) XOR DI(144) XOR DI(139) XOR DI(43) XOR DI(160) XOR DI(397) XOR DI(447) XOR DI(440) XOR DI(109) XOR DI(304) XOR DI(198) XOR DI(358) XOR DI(18) XOR DI(114) XOR DI(37) XOR DI(154) XOR DI(441) XOR DI(434) XOR DI(192) XOR DI(352) XOR DI(12) XOR DI(108) XOR DI(31) XOR DI(428) XOR DI(186) XOR DI(346) XOR DI(6) XOR DI(25) XOR DI(180) XOR DI(19) XOR DI(174) XOR DI(13) XOR DI(168) XOR DI(7) XOR DI(1) XOR DI(501) XOR DI(507);
   DO(2) <= DI(66) XOR DI(490) XOR DI(238) XOR DI(77) XOR DI(259) XOR DI(266) XOR DI(396) XOR DI(358) XOR DI(197) XOR DI(78) XOR DI(324) XOR DI(485) XOR DI(287) XOR DI(345) XOR DI(62) XOR DI(469) XOR DI(49) XOR DI(430) XOR DI(415) XOR DI(179) XOR DI(363) XOR DI(65) XOR DI(286) XOR DI(416) XOR DI(328) XOR DI(466) XOR DI(255) XOR DI(224) XOR DI(102) XOR DI(331) XOR DI(486) XOR DI(348) XOR DI(52) XOR DI(459) XOR DI(456) XOR DI(245) XOR DI(321) XOR DI(42) XOR DI(449) XOR DI(446) XOR DI(128) XOR DI(70) XOR DI(194) XOR DI(227) XOR DI(95) XOR DI(138) XOR DI(192) XOR DI(123) XOR DI(400) XOR DI(470) XOR DI(332) XOR DI(176) XOR DI(403) XOR DI(488) XOR DI(288) XOR DI(21) XOR DI(417) XOR DI(80) XOR DI(290) XOR DI(126) XOR DI(467) XOR DI(204) XOR DI(34) XOR DI(431) XOR DI(419) XOR DI(165) XOR DI(504) XOR DI(250) XOR DI(257) XOR DI(387) XOR DI(53) XOR DI(277) XOR DI(246) XOR DI(215) XOR DI(312) XOR DI(33) XOR DI(114) XOR DI(323) XOR DI(12) XOR DI(408) XOR DI(195) XOR DI(156) XOR DI(241) XOR DI(378) XOR DI(237) XOR DI(24) XOR DI(105) XOR DI(3) XOR DI(228) XOR DI(219) XOR DI(370) XOR DI(304) XOR DI(379) XOR DI(217) XOR DI(124) XOR DI(377) XOR DI(148) XOR DI(98) XOR DI(343) XOR DI(401) XOR DI(313) XOR DI(451) XOR DI(37) XOR DI(177) XOR DI(388) XOR DI(489) XOR DI(262) XOR DI(226) XOR DI(202) XOR DI(133) XOR DI(386) XOR DI(418) XOR DI(157) XOR DI(81) XOR DI(107) XOR DI(302) XOR DI(356) XOR DI(35) XOR DI(152) XOR DI(432) XOR DI(106) XOR DI(433) XOR DI(344) XOR DI(4) XOR DI(23) XOR DI(420) XOR DI(172) XOR DI(505) XOR DI(484) XOR DI(253) XOR DI(352) XOR DI(56) XOR DI(173) XOR DI(280) XOR DI(410) XOR DI(322) XOR DI(460) XOR DI(249) XOR DI(218) XOR DI(96) XOR DI(480) XOR DI(342) XOR DI(46) XOR DI(453) XOR DI(315) XOR DI(122) XOR DI(64) XOR DI(186) XOR DI(464) XOR DI(326) XOR DI(170) XOR DI(397) XOR DI(482) XOR DI(411) XOR DI(284) XOR DI(461) XOR DI(28) XOR DI(413) XOR DI(498) XOR DI(271) XOR DI(240) XOR DI(209) XOR DI(306) XOR DI(317) XOR DI(6) XOR DI(235) XOR DI(231) XOR DI(222) XOR DI(298) XOR DI(211) XOR DI(118) XOR DI(371) XOR DI(142) XOR DI(92) XOR DI(395) XOR DI(307) XOR DI(31) XOR DI(382) XOR DI(483) XOR DI(220) XOR DI(196) XOR DI(127) XOR DI(380) XOR DI(151) XOR DI(146) XOR DI(100) XOR DI(427) XOR DI(166) XOR DI(50) XOR DI(167) XOR DI(404) XOR DI(316) XOR DI(454) XOR DI(212) XOR DI(90) XOR DI(447) XOR DI(116) XOR DI(180) XOR DI(320) XOR DI(391) XOR DI(22) XOR DI(300) XOR DI(311) XOR DI(0) XOR DI(216) XOR DI(205) XOR DI(365) XOR DI(136) XOR DI(389) XOR DI(25) XOR DI(477) XOR DI(214) XOR DI(121) XOR DI(145) XOR DI(140) XOR DI(44) XOR DI(161) XOR DI(398) XOR DI(448) XOR DI(441) XOR DI(110) XOR DI(305) XOR DI(199) XOR DI(359) XOR DI(19) XOR DI(115) XOR DI(38) XOR DI(155) XOR DI(442) XOR DI(435) XOR DI(193) XOR DI(353) XOR DI(13) XOR DI(109) XOR DI(32) XOR DI(429) XOR DI(187) XOR DI(347) XOR DI(7) XOR DI(26) XOR DI(181) XOR DI(20) XOR DI(175) XOR DI(14) XOR DI(169) XOR DI(8) XOR DI(2) XOR DI(502) XOR DI(508);
   DO(3) <= DI(67) XOR DI(491) XOR DI(239) XOR DI(78) XOR DI(260) XOR DI(267) XOR DI(397) XOR DI(359) XOR DI(198) XOR DI(79) XOR DI(325) XOR DI(486) XOR DI(288) XOR DI(346) XOR DI(63) XOR DI(470) XOR DI(50) XOR DI(431) XOR DI(416) XOR DI(180) XOR DI(364) XOR DI(66) XOR DI(287) XOR DI(417) XOR DI(329) XOR DI(467) XOR DI(256) XOR DI(225) XOR DI(103) XOR DI(332) XOR DI(487) XOR DI(349) XOR DI(53) XOR DI(460) XOR DI(457) XOR DI(246) XOR DI(322) XOR DI(43) XOR DI(450) XOR DI(447) XOR DI(129) XOR DI(71) XOR DI(195) XOR DI(228) XOR DI(96) XOR DI(139) XOR DI(193) XOR DI(124) XOR DI(401) XOR DI(471) XOR DI(333) XOR DI(177) XOR DI(404) XOR DI(489) XOR DI(289) XOR DI(22) XOR DI(418) XOR DI(81) XOR DI(291) XOR DI(127) XOR DI(468) XOR DI(205) XOR DI(35) XOR DI(432) XOR DI(420) XOR DI(166) XOR DI(505) XOR DI(251) XOR DI(258) XOR DI(388) XOR DI(54) XOR DI(278) XOR DI(247) XOR DI(216) XOR DI(313) XOR DI(34) XOR DI(115) XOR DI(324) XOR DI(13) XOR DI(409) XOR DI(196) XOR DI(157) XOR DI(242) XOR DI(379) XOR DI(238) XOR DI(25) XOR DI(106) XOR DI(4) XOR DI(229) XOR DI(220) XOR DI(371) XOR DI(305) XOR DI(380) XOR DI(218) XOR DI(125) XOR DI(378) XOR DI(149) XOR DI(99) XOR DI(344) XOR DI(402) XOR DI(314) XOR DI(452) XOR DI(38) XOR DI(178) XOR DI(389) XOR DI(490) XOR DI(263) XOR DI(227) XOR DI(203) XOR DI(134) XOR DI(387) XOR DI(419) XOR DI(158) XOR DI(82) XOR DI(108) XOR DI(303) XOR DI(357) XOR DI(36) XOR DI(153) XOR DI(433) XOR DI(107) XOR DI(434) XOR DI(345) XOR DI(5) XOR DI(24) XOR DI(421) XOR DI(173) XOR DI(506) XOR DI(485) XOR DI(254) XOR DI(353) XOR DI(57) XOR DI(174) XOR DI(281) XOR DI(411) XOR DI(323) XOR DI(461) XOR DI(250) XOR DI(219) XOR DI(97) XOR DI(481) XOR DI(343) XOR DI(47) XOR DI(454) XOR DI(316) XOR DI(123) XOR DI(65) XOR DI(187) XOR DI(465) XOR DI(327) XOR DI(171) XOR DI(398) XOR DI(483) XOR DI(412) XOR DI(285) XOR DI(462) XOR DI(29) XOR DI(414) XOR DI(499) XOR DI(272) XOR DI(241) XOR DI(210) XOR DI(307) XOR DI(318) XOR DI(7) XOR DI(236) XOR DI(232) XOR DI(223) XOR DI(299) XOR DI(212) XOR DI(119) XOR DI(372) XOR DI(143) XOR DI(93) XOR DI(396) XOR DI(308) XOR DI(32) XOR DI(383) XOR DI(484) XOR DI(221) XOR DI(197) XOR DI(128) XOR DI(381) XOR DI(152) XOR DI(147) XOR DI(101) XOR DI(428) XOR DI(167) XOR DI(51) XOR DI(168) XOR DI(405) XOR DI(317) XOR DI(455) XOR DI(213) XOR DI(91) XOR DI(448) XOR DI(117) XOR DI(181) XOR DI(321) XOR DI(392) XOR DI(23) XOR DI(301) XOR DI(312) XOR DI(1) XOR DI(217) XOR DI(206) XOR DI(366) XOR DI(137) XOR DI(390) XOR DI(26) XOR DI(478) XOR DI(215) XOR DI(122) XOR DI(146) XOR DI(141) XOR DI(45) XOR DI(162) XOR DI(399) XOR DI(449) XOR DI(442) XOR DI(111) XOR DI(306) XOR DI(200) XOR DI(360) XOR DI(20) XOR DI(116) XOR DI(39) XOR DI(156) XOR DI(443) XOR DI(436) XOR DI(194) XOR DI(354) XOR DI(14) XOR DI(110) XOR DI(33) XOR DI(430) XOR DI(188) XOR DI(348) XOR DI(8) XOR DI(27) XOR DI(182) XOR DI(21) XOR DI(176) XOR DI(15) XOR DI(170) XOR DI(9) XOR DI(3) XOR DI(503) XOR DI(509);
   DO(4) <= DI(68) XOR DI(492) XOR DI(240) XOR DI(79) XOR DI(261) XOR DI(268) XOR DI(398) XOR DI(360) XOR DI(199) XOR DI(80) XOR DI(326) XOR DI(487) XOR DI(289) XOR DI(347) XOR DI(64) XOR DI(471) XOR DI(51) XOR DI(432) XOR DI(417) XOR DI(181) XOR DI(365) XOR DI(67) XOR DI(288) XOR DI(418) XOR DI(330) XOR DI(468) XOR DI(257) XOR DI(226) XOR DI(104) XOR DI(333) XOR DI(488) XOR DI(350) XOR DI(54) XOR DI(461) XOR DI(458) XOR DI(247) XOR DI(323) XOR DI(44) XOR DI(451) XOR DI(448) XOR DI(130) XOR DI(72) XOR DI(196) XOR DI(229) XOR DI(97) XOR DI(140) XOR DI(194) XOR DI(125) XOR DI(402) XOR DI(472) XOR DI(334) XOR DI(178) XOR DI(405) XOR DI(490) XOR DI(290) XOR DI(23) XOR DI(419) XOR DI(82) XOR DI(292) XOR DI(128) XOR DI(469) XOR DI(206) XOR DI(36) XOR DI(433) XOR DI(421) XOR DI(167) XOR DI(506) XOR DI(252) XOR DI(259) XOR DI(389) XOR DI(55) XOR DI(279) XOR DI(248) XOR DI(217) XOR DI(314) XOR DI(35) XOR DI(116) XOR DI(325) XOR DI(14) XOR DI(410) XOR DI(197) XOR DI(158) XOR DI(243) XOR DI(380) XOR DI(239) XOR DI(26) XOR DI(107) XOR DI(5) XOR DI(230) XOR DI(221) XOR DI(372) XOR DI(306) XOR DI(381) XOR DI(219) XOR DI(126) XOR DI(379) XOR DI(150) XOR DI(100) XOR DI(345) XOR DI(403) XOR DI(315) XOR DI(453) XOR DI(39) XOR DI(179) XOR DI(390) XOR DI(491) XOR DI(264) XOR DI(228) XOR DI(204) XOR DI(135) XOR DI(388) XOR DI(420) XOR DI(159) XOR DI(83) XOR DI(109) XOR DI(304) XOR DI(358) XOR DI(37) XOR DI(154) XOR DI(434) XOR DI(108) XOR DI(435) XOR DI(346) XOR DI(6) XOR DI(25) XOR DI(422) XOR DI(174) XOR DI(507) XOR DI(486) XOR DI(255) XOR DI(354) XOR DI(58) XOR DI(175) XOR DI(282) XOR DI(412) XOR DI(324) XOR DI(462) XOR DI(251) XOR DI(220) XOR DI(98) XOR DI(482) XOR DI(344) XOR DI(48) XOR DI(455) XOR DI(317) XOR DI(124) XOR DI(66) XOR DI(188) XOR DI(466) XOR DI(328) XOR DI(172) XOR DI(399) XOR DI(484) XOR DI(413) XOR DI(286) XOR DI(463) XOR DI(30) XOR DI(415) XOR DI(500) XOR DI(273) XOR DI(242) XOR DI(211) XOR DI(308) XOR DI(319) XOR DI(8) XOR DI(237) XOR DI(233) XOR DI(224) XOR DI(300) XOR DI(213) XOR DI(120) XOR DI(373) XOR DI(144) XOR DI(94) XOR DI(397) XOR DI(309) XOR DI(33) XOR DI(384) XOR DI(485) XOR DI(222) XOR DI(198) XOR DI(129) XOR DI(382) XOR DI(153) XOR DI(148) XOR DI(102) XOR DI(429) XOR DI(0) XOR DI(168) XOR DI(52) XOR DI(169) XOR DI(406) XOR DI(318) XOR DI(456) XOR DI(214) XOR DI(92) XOR DI(449) XOR DI(118) XOR DI(182) XOR DI(322) XOR DI(393) XOR DI(24) XOR DI(302) XOR DI(313) XOR DI(2) XOR DI(218) XOR DI(207) XOR DI(367) XOR DI(138) XOR DI(391) XOR DI(27) XOR DI(479) XOR DI(216) XOR DI(123) XOR DI(147) XOR DI(142) XOR DI(46) XOR DI(163) XOR DI(400) XOR DI(450) XOR DI(443) XOR DI(112) XOR DI(307) XOR DI(201) XOR DI(361) XOR DI(21) XOR DI(117) XOR DI(40) XOR DI(157) XOR DI(444) XOR DI(437) XOR DI(195) XOR DI(355) XOR DI(15) XOR DI(111) XOR DI(34) XOR DI(431) XOR DI(189) XOR DI(349) XOR DI(9) XOR DI(28) XOR DI(183) XOR DI(22) XOR DI(177) XOR DI(16) XOR DI(171) XOR DI(10) XOR DI(4) XOR DI(504) XOR DI(510);
   DO(5) <= DI(69) XOR DI(493) XOR DI(241) XOR DI(80) XOR DI(262) XOR DI(269) XOR DI(399) XOR DI(361) XOR DI(200) XOR DI(81) XOR DI(327) XOR DI(488) XOR DI(290) XOR DI(348) XOR DI(65) XOR DI(472) XOR DI(52) XOR DI(433) XOR DI(418) XOR DI(182) XOR DI(366) XOR DI(68) XOR DI(289) XOR DI(419) XOR DI(331) XOR DI(469) XOR DI(258) XOR DI(227) XOR DI(105) XOR DI(334) XOR DI(489) XOR DI(351) XOR DI(55) XOR DI(462) XOR DI(459) XOR DI(248) XOR DI(324) XOR DI(45) XOR DI(452) XOR DI(449) XOR DI(131) XOR DI(73) XOR DI(197) XOR DI(230) XOR DI(98) XOR DI(141) XOR DI(195) XOR DI(126) XOR DI(403) XOR DI(473) XOR DI(335) XOR DI(179) XOR DI(406) XOR DI(491) XOR DI(291) XOR DI(24) XOR DI(420) XOR DI(83) XOR DI(293) XOR DI(129) XOR DI(470) XOR DI(207) XOR DI(37) XOR DI(434) XOR DI(422) XOR DI(168) XOR DI(507) XOR DI(253) XOR DI(260) XOR DI(390) XOR DI(56) XOR DI(280) XOR DI(249) XOR DI(218) XOR DI(315) XOR DI(36) XOR DI(117) XOR DI(326) XOR DI(15) XOR DI(411) XOR DI(198) XOR DI(159) XOR DI(244) XOR DI(381) XOR DI(240) XOR DI(27) XOR DI(108) XOR DI(6) XOR DI(231) XOR DI(222) XOR DI(373) XOR DI(307) XOR DI(382) XOR DI(220) XOR DI(127) XOR DI(380) XOR DI(151) XOR DI(101) XOR DI(346) XOR DI(404) XOR DI(316) XOR DI(454) XOR DI(40) XOR DI(180) XOR DI(391) XOR DI(492) XOR DI(265) XOR DI(229) XOR DI(205) XOR DI(136) XOR DI(389) XOR DI(421) XOR DI(160) XOR DI(84) XOR DI(110) XOR DI(305) XOR DI(359) XOR DI(38) XOR DI(155) XOR DI(435) XOR DI(109) XOR DI(436) XOR DI(347) XOR DI(7) XOR DI(26) XOR DI(423) XOR DI(175) XOR DI(508) XOR DI(487) XOR DI(256) XOR DI(355) XOR DI(59) XOR DI(176) XOR DI(283) XOR DI(413) XOR DI(325) XOR DI(463) XOR DI(252) XOR DI(221) XOR DI(99) XOR DI(483) XOR DI(345) XOR DI(49) XOR DI(456) XOR DI(318) XOR DI(125) XOR DI(67) XOR DI(189) XOR DI(467) XOR DI(329) XOR DI(173) XOR DI(400) XOR DI(485) XOR DI(414) XOR DI(287) XOR DI(464) XOR DI(31) XOR DI(416) XOR DI(501) XOR DI(274) XOR DI(243) XOR DI(212) XOR DI(309) XOR DI(320) XOR DI(9) XOR DI(238) XOR DI(234) XOR DI(225) XOR DI(301) XOR DI(214) XOR DI(121) XOR DI(374) XOR DI(145) XOR DI(95) XOR DI(398) XOR DI(310) XOR DI(34) XOR DI(385) XOR DI(486) XOR DI(223) XOR DI(199) XOR DI(130) XOR DI(383) XOR DI(154) XOR DI(149) XOR DI(103) XOR DI(430) XOR DI(1) XOR DI(169) XOR DI(53) XOR DI(170) XOR DI(407) XOR DI(319) XOR DI(457) XOR DI(215) XOR DI(93) XOR DI(450) XOR DI(119) XOR DI(183) XOR DI(323) XOR DI(394) XOR DI(25) XOR DI(303) XOR DI(314) XOR DI(3) XOR DI(219) XOR DI(208) XOR DI(368) XOR DI(139) XOR DI(392) XOR DI(28) XOR DI(480) XOR DI(217) XOR DI(124) XOR DI(148) XOR DI(143) XOR DI(47) XOR DI(164) XOR DI(401) XOR DI(451) XOR DI(444) XOR DI(113) XOR DI(308) XOR DI(202) XOR DI(362) XOR DI(22) XOR DI(118) XOR DI(41) XOR DI(158) XOR DI(445) XOR DI(438) XOR DI(196) XOR DI(356) XOR DI(16) XOR DI(112) XOR DI(35) XOR DI(432) XOR DI(190) XOR DI(350) XOR DI(10) XOR DI(29) XOR DI(184) XOR DI(23) XOR DI(178) XOR DI(17) XOR DI(172) XOR DI(11) XOR DI(5) XOR DI(505) XOR DI(511);
   DO(6) <= DI(70) XOR DI(494) XOR DI(345) XOR DI(313) XOR DI(242) XOR DI(269) XOR DI(63) XOR DI(81) XOR DI(263) XOR DI(378) XOR DI(138) XOR DI(62) XOR DI(329) XOR DI(270) XOR DI(400) XOR DI(178) XOR DI(79) XOR DI(107) XOR DI(387) XOR DI(5) XOR DI(362) XOR DI(201) XOR DI(361) XOR DI(82) XOR DI(416) XOR DI(328) XOR DI(489) XOR DI(264) XOR DI(255) XOR DI(195) XOR DI(291) XOR DI(467) XOR DI(349) XOR DI(66) XOR DI(473) XOR DI(418) XOR DI(53) XOR DI(434) XOR DI(419) XOR DI(153) XOR DI(238) XOR DI(183) XOR DI(367) XOR DI(69) XOR DI(290) XOR DI(420) XOR DI(332) XOR DI(303) XOR DI(470) XOR DI(259) XOR DI(228) XOR DI(286) XOR DI(106) XOR DI(368) XOR DI(88) XOR DI(154) XOR DI(78) XOR DI(124) XOR DI(202) XOR DI(98) XOR DI(335) XOR DI(490) XOR DI(260) XOR DI(352) XOR DI(56) XOR DI(463) XOR DI(409) XOR DI(322) XOR DI(460) XOR DI(249) XOR DI(325) XOR DI(46) XOR DI(453) XOR DI(450) XOR DI(440) XOR DI(64) XOR DI(132) XOR DI(394) XOR DI(482) XOR DI(74) XOR DI(198) XOR DI(251) XOR DI(108) XOR DI(231) XOR DI(99) XOR DI(298) XOR DI(142) XOR DI(31) XOR DI(196) XOR DI(127) XOR DI(380) XOR DI(296) XOR DI(350) XOR DI(247) XOR DI(404) XOR DI(243) XOR DI(474) XOR DI(336) XOR DI(40) XOR DI(447) XOR DI(180) XOR DI(278) XOR DI(22) XOR DI(407) XOR DI(492) XOR DI(229) XOR DI(225) XOR DI(292) XOR DI(112) XOR DI(136) XOR DI(389) XOR DI(25) XOR DI(376) XOR DI(421) XOR DI(84) XOR DI(314) XOR DI(385) XOR DI(294) XOR DI(305) XOR DI(130) XOR DI(471) XOR DI(208) XOR DI(134) XOR DI(38) XOR DI(435) XOR DI(193) XOR DI(429) XOR DI(103) XOR DI(423) XOR DI(341) XOR DI(169) XOR DI(163) XOR DI(496) XOR DI(508) XOR DI(233) XOR DI(254) XOR DI(261) XOR DI(391) XOR DI(192) XOR DI(480) XOR DI(282) XOR DI(340) XOR DI(57) XOR DI(44) XOR DI(425) XOR DI(281) XOR DI(411) XOR DI(250) XOR DI(219) XOR DI(343) XOR DI(47) XOR DI(454) XOR DI(316) XOR DI(37) XOR DI(444) XOR DI(90) XOR DI(118) XOR DI(327) XOR DI(398) XOR DI(483) XOR DI(16) XOR DI(412) XOR DI(75) XOR DI(285) XOR DI(121) XOR DI(462) XOR DI(199) XOR DI(160) XOR DI(245) XOR DI(382) XOR DI(241) XOR DI(210) XOR DI(28) XOR DI(109) XOR DI(318) XOR DI(7) XOR DI(236) XOR DI(232) XOR DI(19) XOR DI(223) XOR DI(214) XOR DI(374) XOR DI(212) XOR DI(143) XOR DI(93) XOR DI(396) XOR DI(308) XOR DI(383) XOR DI(221) XOR DI(128) XOR DI(381) XOR DI(413) XOR DI(152) XOR DI(76) XOR DI(102) XOR DI(427) XOR DI(428) XOR DI(167) XOR DI(500) XOR DI(248) XOR DI(347) XOR DI(51) XOR DI(168) XOR DI(405) XOR DI(317) XOR DI(455) XOR DI(475) XOR DI(41) XOR DI(181) XOR DI(459) XOR DI(392) XOR DI(406) XOR DI(493) XOR DI(266) XOR DI(1) XOR DI(230) XOR DI(217) XOR DI(206) XOR DI(137) XOR DI(390) XOR DI(377) XOR DI(478) XOR DI(422) XOR DI(161) XOR DI(449) XOR DI(207) XOR DI(85) XOR DI(111) XOR DI(175) XOR DI(306) XOR DI(360) XOR DI(20) XOR DI(116) XOR DI(39) XOR DI(156) XOR DI(436) XOR DI(105) XOR DI(300) XOR DI(194) XOR DI(354) XOR DI(110) XOR DI(33) XOR DI(437) XOR DI(430) XOR DI(348) XOR DI(8) XOR DI(27) XOR DI(424) XOR DI(342) XOR DI(21) XOR DI(176) XOR DI(164) XOR DI(503) XOR DI(509);
   DO(7) <= DI(71) XOR DI(495) XOR DI(346) XOR DI(314) XOR DI(243) XOR DI(270) XOR DI(64) XOR DI(82) XOR DI(264) XOR DI(379) XOR DI(139) XOR DI(63) XOR DI(330) XOR DI(271) XOR DI(401) XOR DI(179) XOR DI(80) XOR DI(108) XOR DI(388) XOR DI(6) XOR DI(363) XOR DI(202) XOR DI(362) XOR DI(83) XOR DI(417) XOR DI(329) XOR DI(490) XOR DI(265) XOR DI(256) XOR DI(196) XOR DI(292) XOR DI(468) XOR DI(350) XOR DI(67) XOR DI(474) XOR DI(419) XOR DI(54) XOR DI(435) XOR DI(420) XOR DI(154) XOR DI(239) XOR DI(184) XOR DI(368) XOR DI(70) XOR DI(291) XOR DI(421) XOR DI(333) XOR DI(304) XOR DI(471) XOR DI(260) XOR DI(229) XOR DI(287) XOR DI(107) XOR DI(369) XOR DI(89) XOR DI(155) XOR DI(79) XOR DI(125) XOR DI(203) XOR DI(99) XOR DI(336) XOR DI(491) XOR DI(261) XOR DI(353) XOR DI(57) XOR DI(464) XOR DI(410) XOR DI(323) XOR DI(461) XOR DI(250) XOR DI(326) XOR DI(47) XOR DI(454) XOR DI(451) XOR DI(441) XOR DI(65) XOR DI(133) XOR DI(395) XOR DI(483) XOR DI(75) XOR DI(199) XOR DI(252) XOR DI(109) XOR DI(232) XOR DI(100) XOR DI(299) XOR DI(143) XOR DI(32) XOR DI(197) XOR DI(128) XOR DI(381) XOR DI(297) XOR DI(351) XOR DI(248) XOR DI(405) XOR DI(244) XOR DI(475) XOR DI(337) XOR DI(41) XOR DI(448) XOR DI(181) XOR DI(279) XOR DI(23) XOR DI(408) XOR DI(493) XOR DI(230) XOR DI(226) XOR DI(293) XOR DI(113) XOR DI(137) XOR DI(390) XOR DI(26) XOR DI(377) XOR DI(422) XOR DI(85) XOR DI(315) XOR DI(386) XOR DI(295) XOR DI(306) XOR DI(131) XOR DI(472) XOR DI(209) XOR DI(135) XOR DI(39) XOR DI(436) XOR DI(194) XOR DI(430) XOR DI(104) XOR DI(424) XOR DI(342) XOR DI(170) XOR DI(164) XOR DI(497) XOR DI(509) XOR DI(234) XOR DI(255) XOR DI(262) XOR DI(392) XOR DI(193) XOR DI(481) XOR DI(283) XOR DI(341) XOR DI(58) XOR DI(45) XOR DI(426) XOR DI(282) XOR DI(412) XOR DI(251) XOR DI(220) XOR DI(344) XOR DI(48) XOR DI(455) XOR DI(317) XOR DI(38) XOR DI(445) XOR DI(91) XOR DI(119) XOR DI(328) XOR DI(399) XOR DI(484) XOR DI(17) XOR DI(413) XOR DI(76) XOR DI(286) XOR DI(122) XOR DI(463) XOR DI(200) XOR DI(161) XOR DI(246) XOR DI(383) XOR DI(242) XOR DI(211) XOR DI(29) XOR DI(110) XOR DI(319) XOR DI(8) XOR DI(237) XOR DI(233) XOR DI(20) XOR DI(224) XOR DI(215) XOR DI(375) XOR DI(213) XOR DI(144) XOR DI(94) XOR DI(397) XOR DI(309) XOR DI(384) XOR DI(222) XOR DI(129) XOR DI(382) XOR DI(414) XOR DI(153) XOR DI(77) XOR DI(103) XOR DI(428) XOR DI(429) XOR DI(0) XOR DI(168) XOR DI(501) XOR DI(249) XOR DI(348) XOR DI(52) XOR DI(169) XOR DI(406) XOR DI(318) XOR DI(456) XOR DI(476) XOR DI(42) XOR DI(182) XOR DI(460) XOR DI(393) XOR DI(407) XOR DI(494) XOR DI(267) XOR DI(2) XOR DI(231) XOR DI(218) XOR DI(207) XOR DI(138) XOR DI(391) XOR DI(378) XOR DI(479) XOR DI(423) XOR DI(162) XOR DI(450) XOR DI(208) XOR DI(86) XOR DI(112) XOR DI(176) XOR DI(307) XOR DI(361) XOR DI(21) XOR DI(117) XOR DI(40) XOR DI(157) XOR DI(437) XOR DI(106) XOR DI(301) XOR DI(195) XOR DI(355) XOR DI(111) XOR DI(34) XOR DI(438) XOR DI(431) XOR DI(349) XOR DI(9) XOR DI(28) XOR DI(425) XOR DI(343) XOR DI(22) XOR DI(177) XOR DI(165) XOR DI(504) XOR DI(510);
   DO(8) <= DI(72) XOR DI(496) XOR DI(347) XOR DI(315) XOR DI(244) XOR DI(271) XOR DI(65) XOR DI(83) XOR DI(265) XOR DI(380) XOR DI(140) XOR DI(64) XOR DI(331) XOR DI(272) XOR DI(402) XOR DI(180) XOR DI(81) XOR DI(109) XOR DI(389) XOR DI(7) XOR DI(364) XOR DI(203) XOR DI(363) XOR DI(84) XOR DI(418) XOR DI(330) XOR DI(491) XOR DI(266) XOR DI(257) XOR DI(197) XOR DI(293) XOR DI(469) XOR DI(351) XOR DI(68) XOR DI(475) XOR DI(420) XOR DI(55) XOR DI(436) XOR DI(421) XOR DI(155) XOR DI(240) XOR DI(185) XOR DI(369) XOR DI(71) XOR DI(292) XOR DI(422) XOR DI(334) XOR DI(305) XOR DI(472) XOR DI(261) XOR DI(230) XOR DI(288) XOR DI(108) XOR DI(370) XOR DI(90) XOR DI(156) XOR DI(80) XOR DI(126) XOR DI(204) XOR DI(100) XOR DI(337) XOR DI(492) XOR DI(262) XOR DI(354) XOR DI(58) XOR DI(465) XOR DI(411) XOR DI(324) XOR DI(462) XOR DI(251) XOR DI(327) XOR DI(48) XOR DI(455) XOR DI(452) XOR DI(442) XOR DI(66) XOR DI(134) XOR DI(396) XOR DI(484) XOR DI(76) XOR DI(200) XOR DI(253) XOR DI(110) XOR DI(233) XOR DI(101) XOR DI(300) XOR DI(144) XOR DI(33) XOR DI(198) XOR DI(129) XOR DI(382) XOR DI(298) XOR DI(352) XOR DI(249) XOR DI(406) XOR DI(245) XOR DI(476) XOR DI(338) XOR DI(42) XOR DI(449) XOR DI(182) XOR DI(280) XOR DI(24) XOR DI(409) XOR DI(494) XOR DI(231) XOR DI(227) XOR DI(294) XOR DI(114) XOR DI(138) XOR DI(391) XOR DI(27) XOR DI(378) XOR DI(423) XOR DI(86) XOR DI(316) XOR DI(387) XOR DI(296) XOR DI(307) XOR DI(132) XOR DI(473) XOR DI(210) XOR DI(136) XOR DI(40) XOR DI(437) XOR DI(195) XOR DI(431) XOR DI(105) XOR DI(425) XOR DI(343) XOR DI(171) XOR DI(165) XOR DI(498) XOR DI(510) XOR DI(235) XOR DI(256) XOR DI(263) XOR DI(393) XOR DI(194) XOR DI(482) XOR DI(284) XOR DI(342) XOR DI(59) XOR DI(46) XOR DI(427) XOR DI(283) XOR DI(413) XOR DI(252) XOR DI(221) XOR DI(345) XOR DI(49) XOR DI(456) XOR DI(318) XOR DI(39) XOR DI(446) XOR DI(92) XOR DI(120) XOR DI(329) XOR DI(400) XOR DI(485) XOR DI(18) XOR DI(414) XOR DI(77) XOR DI(287) XOR DI(123) XOR DI(464) XOR DI(201) XOR DI(162) XOR DI(247) XOR DI(384) XOR DI(243) XOR DI(212) XOR DI(30) XOR DI(111) XOR DI(320) XOR DI(9) XOR DI(238) XOR DI(234) XOR DI(21) XOR DI(0) XOR DI(225) XOR DI(216) XOR DI(376) XOR DI(214) XOR DI(145) XOR DI(95) XOR DI(398) XOR DI(310) XOR DI(385) XOR DI(223) XOR DI(130) XOR DI(383) XOR DI(415) XOR DI(154) XOR DI(78) XOR DI(104) XOR DI(429) XOR DI(430) XOR DI(1) XOR DI(169) XOR DI(502) XOR DI(250) XOR DI(349) XOR DI(53) XOR DI(170) XOR DI(407) XOR DI(319) XOR DI(457) XOR DI(477) XOR DI(43) XOR DI(183) XOR DI(461) XOR DI(394) XOR DI(408) XOR DI(495) XOR DI(268) XOR DI(3) XOR DI(232) XOR DI(219) XOR DI(208) XOR DI(139) XOR DI(392) XOR DI(379) XOR DI(480) XOR DI(424) XOR DI(163) XOR DI(451) XOR DI(209) XOR DI(87) XOR DI(113) XOR DI(177) XOR DI(308) XOR DI(362) XOR DI(22) XOR DI(118) XOR DI(41) XOR DI(158) XOR DI(438) XOR DI(107) XOR DI(302) XOR DI(196) XOR DI(356) XOR DI(112) XOR DI(35) XOR DI(439) XOR DI(432) XOR DI(350) XOR DI(10) XOR DI(29) XOR DI(426) XOR DI(344) XOR DI(23) XOR DI(178) XOR DI(166) XOR DI(505) XOR DI(511);
   DO(9) <= DI(255) XOR DI(324) XOR DI(282) XOR DI(459) XOR DI(175) XOR DI(260) XOR DI(326) XOR DI(116) XOR DI(73) XOR DI(497) XOR DI(348) XOR DI(316) XOR DI(150) XOR DI(90) XOR DI(449) XOR DI(305) XOR DI(245) XOR DI(48) XOR DI(165) XOR DI(272) XOR DI(66) XOR DI(134) XOR DI(84) XOR DI(266) XOR DI(396) XOR DI(484) XOR DI(381) XOR DI(76) XOR DI(286) XOR DI(122) XOR DI(126) XOR DI(141) XOR DI(488) XOR DI(500) XOR DI(64) XOR DI(65) XOR DI(332) XOR DI(273) XOR DI(403) XOR DI(181) XOR DI(82) XOR DI(110) XOR DI(390) XOR DI(8) XOR DI(454) XOR DI(365) XOR DI(204) XOR DI(364) XOR DI(85) XOR DI(300) XOR DI(144) XOR DI(94) XOR DI(419) XOR DI(331) XOR DI(492) XOR DI(267) XOR DI(51) XOR DI(258) XOR DI(198) XOR DI(294) XOR DI(470) XOR DI(138) XOR DI(352) XOR DI(6) XOR DI(229) XOR DI(68) XOR DI(387) XOR DI(69) XOR DI(315) XOR DI(476) XOR DI(278) XOR DI(421) XOR DI(406) XOR DI(354) XOR DI(56) XOR DI(322) XOR DI(33) XOR DI(437) XOR DI(185) XOR DI(218) XOR DI(12) XOR DI(422) XOR DI(156) XOR DI(241) XOR DI(378) XOR DI(186) XOR DI(369) XOR DI(361) XOR DI(370) XOR DI(168) XOR DI(72) XOR DI(98) XOR DI(293) XOR DI(26) XOR DI(423) XOR DI(335) XOR DI(411) XOR DI(475) XOR DI(306) XOR DI(473) XOR DI(402) XOR DI(275) XOR DI(262) XOR DI(231) XOR DI(200) XOR DI(289) XOR DI(109) XOR DI(298) XOR DI(371) XOR DI(91) XOR DI(418) XOR DI(157) XOR DI(203) XOR DI(81) XOR DI(207) XOR DI(127) XOR DI(468) XOR DI(205) XOR DI(136) XOR DI(389) XOR DI(101) XOR DI(296) XOR DI(100) XOR DI(338) XOR DI(493) XOR DI(63) XOR DI(487) XOR DI(263) XOR DI(355) XOR DI(194) XOR DI(75) XOR DI(482) XOR DI(342) XOR DI(59) XOR DI(466) XOR DI(412) XOR DI(62) XOR DI(413) XOR DI(325) XOR DI(463) XOR DI(252) XOR DI(328) XOR DI(49) XOR DI(456) XOR DI(453) XOR DI(318) XOR DI(446) XOR DI(443) XOR DI(125) XOR DI(67) XOR DI(191) XOR DI(135) XOR DI(120) XOR DI(397) XOR DI(467) XOR DI(329) XOR DI(173) XOR DI(485) XOR DI(18) XOR DI(77) XOR DI(464) XOR DI(201) XOR DI(247) XOR DI(254) XOR DI(243) XOR DI(212) XOR DI(111) XOR DI(192) XOR DI(153) XOR DI(238) XOR DI(375) XOR DI(234) XOR DI(21) XOR DI(102) XOR DI(225) XOR DI(216) XOR DI(301) XOR DI(376) XOR DI(214) XOR DI(145) XOR DI(340) XOR DI(398) XOR DI(310) XOR DI(34) XOR DI(174) XOR DI(199) XOR DI(130) XOR DI(383) XOR DI(154) XOR DI(104) XOR DI(299) XOR DI(353) XOR DI(32) XOR DI(149) XOR DI(429) XOR DI(103) XOR DI(341) XOR DI(20) XOR DI(417) XOR DI(502) XOR DI(250) XOR DI(407) XOR DI(246) XOR DI(477) XOR DI(339) XOR DI(43) XOR DI(450) XOR DI(183) XOR DI(281) XOR DI(25) XOR DI(410) XOR DI(495) XOR DI(314) XOR DI(232) XOR DI(228) XOR DI(295) XOR DI(115) XOR DI(368) XOR DI(139) XOR DI(392) XOR DI(304) XOR DI(28) XOR DI(379) XOR DI(480) XOR DI(193) XOR DI(143) XOR DI(424) XOR DI(313) XOR DI(451) XOR DI(87) XOR DI(444) XOR DI(177) XOR DI(317) XOR DI(388) XOR DI(297) XOR DI(308) XOR DI(133) XOR DI(474) XOR DI(211) XOR DI(137) XOR DI(41) XOR DI(445) XOR DI(438) XOR DI(107) XOR DI(302) XOR DI(196) XOR DI(356) XOR DI(35) XOR DI(432) XOR DI(190) XOR DI(106) XOR DI(29) XOR DI(426) XOR DI(344) XOR DI(17) XOR DI(172) XOR DI(166) XOR DI(5) XOR DI(499) XOR DI(511);
   DO(10) <= DI(256) XOR DI(321) XOR DI(322) XOR DI(487) XOR DI(260) XOR DI(325) XOR DI(47) XOR DI(75) XOR DI(283) XOR DI(460) XOR DI(176) XOR DI(261) XOR DI(361) XOR DI(327) XOR DI(117) XOR DI(170) XOR DI(74) XOR DI(431) XOR DI(177) XOR DI(498) XOR DI(349) XOR DI(317) XOR DI(151) XOR DI(100) XOR DI(394) XOR DI(91) XOR DI(450) XOR DI(484) XOR DI(257) XOR DI(284) XOR DI(306) XOR DI(122) XOR DI(246) XOR DI(49) XOR DI(166) XOR DI(273) XOR DI(67) XOR DI(224) XOR DI(135) XOR DI(85) XOR DI(267) XOR DI(397) XOR DI(236) XOR DI(51) XOR DI(485) XOR DI(222) XOR DI(285) XOR DI(79) XOR DI(382) XOR DI(77) XOR DI(287) XOR DI(123) XOR DI(127) XOR DI(31) XOR DI(428) XOR DI(142) XOR DI(96) XOR DI(416) XOR DI(489) XOR DI(501) XOR DI(65) XOR DI(346) XOR DI(66) XOR DI(275) XOR DI(333) XOR DI(274) XOR DI(404) XOR DI(243) XOR DI(40) XOR DI(182) XOR DI(83) XOR DI(111) XOR DI(391) XOR DI(9) XOR DI(455) XOR DI(375) XOR DI(366) XOR DI(225) XOR DI(93) XOR DI(205) XOR DI(365) XOR DI(86) XOR DI(301) XOR DI(190) XOR DI(406) XOR DI(145) XOR DI(95) XOR DI(420) XOR DI(332) XOR DI(493) XOR DI(268) XOR DI(310) XOR DI(52) XOR DI(385) XOR DI(449) XOR DI(401) XOR DI(259) XOR DI(286) XOR DI(199) XOR DI(295) XOR DI(471) XOR DI(368) XOR DI(139) XOR DI(415) XOR DI(10) XOR DI(288) XOR DI(353) XOR DI(124) XOR DI(32) XOR DI(386) XOR DI(429) XOR DI(7) XOR DI(1) XOR DI(417) XOR DI(163) XOR DI(2) XOR DI(502) XOR DI(482) XOR DI(230) XOR DI(69) XOR DI(388) XOR DI(350) XOR DI(70) XOR DI(316) XOR DI(477) XOR DI(279) XOR DI(54) XOR DI(422) XOR DI(407) XOR DI(171) XOR DI(355) XOR DI(57) XOR DI(278) XOR DI(320) XOR DI(458) XOR DI(216) XOR DI(94) XOR DI(323) XOR DI(313) XOR DI(34) XOR DI(438) XOR DI(120) XOR DI(62) XOR DI(186) XOR DI(219) XOR DI(462) XOR DI(324) XOR DI(168) XOR DI(395) XOR DI(480) XOR DI(13) XOR DI(409) XOR DI(459) XOR DI(423) XOR DI(157) XOR DI(242) XOR DI(379) XOR DI(269) XOR DI(238) XOR DI(207) XOR DI(304) XOR DI(4) XOR DI(187) XOR DI(370) XOR DI(220) XOR DI(362) XOR DI(371) XOR DI(209) XOR DI(90) XOR DI(169) XOR DI(218) XOR DI(125) XOR DI(378) XOR DI(149) XOR DI(73) XOR DI(99) XOR DI(294) XOR DI(27) XOR DI(424) XOR DI(98) XOR DI(336) XOR DI(412) XOR DI(164) XOR DI(476) XOR DI(48) XOR DI(165) XOR DI(402) XOR DI(210) XOR DI(307) XOR DI(114) XOR DI(474) XOR DI(403) XOR DI(276) XOR DI(20) XOR DI(263) XOR DI(232) XOR DI(201) XOR DI(214) XOR DI(290) XOR DI(203) XOR DI(110) XOR DI(363) XOR DI(387) XOR DI(299) XOR DI(23) XOR DI(119) XOR DI(372) XOR DI(143) XOR DI(92) XOR DI(419) XOR DI(158) XOR DI(159) XOR DI(396) XOR DI(204) XOR DI(82) XOR DI(208) XOR DI(128) XOR DI(17) XOR DI(469) XOR DI(206) XOR DI(113) XOR DI(137) XOR DI(153) XOR DI(390) XOR DI(440) XOR DI(102) XOR DI(297) XOR DI(351) XOR DI(11) XOR DI(185) XOR DI(5) XOR DI(101) XOR DI(24) XOR DI(179) XOR DI(339) XOR DI(12) XOR DI(0) XOR DI(494) XOR DI(506);
   DO(11) <= DI(257) XOR DI(322) XOR DI(323) XOR DI(488) XOR DI(261) XOR DI(326) XOR DI(48) XOR DI(76) XOR DI(284) XOR DI(461) XOR DI(177) XOR DI(262) XOR DI(362) XOR DI(328) XOR DI(118) XOR DI(171) XOR DI(75) XOR DI(432) XOR DI(178) XOR DI(499) XOR DI(350) XOR DI(318) XOR DI(152) XOR DI(101) XOR DI(395) XOR DI(92) XOR DI(451) XOR DI(485) XOR DI(258) XOR DI(285) XOR DI(307) XOR DI(123) XOR DI(247) XOR DI(50) XOR DI(167) XOR DI(274) XOR DI(68) XOR DI(225) XOR DI(136) XOR DI(86) XOR DI(268) XOR DI(398) XOR DI(237) XOR DI(52) XOR DI(486) XOR DI(223) XOR DI(286) XOR DI(80) XOR DI(383) XOR DI(78) XOR DI(288) XOR DI(124) XOR DI(128) XOR DI(32) XOR DI(429) XOR DI(143) XOR DI(97) XOR DI(417) XOR DI(490) XOR DI(502) XOR DI(66) XOR DI(347) XOR DI(67) XOR DI(276) XOR DI(334) XOR DI(275) XOR DI(405) XOR DI(244) XOR DI(41) XOR DI(183) XOR DI(84) XOR DI(112) XOR DI(392) XOR DI(10) XOR DI(456) XOR DI(376) XOR DI(367) XOR DI(226) XOR DI(94) XOR DI(206) XOR DI(366) XOR DI(87) XOR DI(302) XOR DI(191) XOR DI(407) XOR DI(146) XOR DI(96) XOR DI(421) XOR DI(333) XOR DI(494) XOR DI(269) XOR DI(311) XOR DI(53) XOR DI(386) XOR DI(450) XOR DI(402) XOR DI(260) XOR DI(287) XOR DI(200) XOR DI(296) XOR DI(472) XOR DI(369) XOR DI(140) XOR DI(416) XOR DI(11) XOR DI(289) XOR DI(354) XOR DI(125) XOR DI(33) XOR DI(387) XOR DI(430) XOR DI(8) XOR DI(2) XOR DI(418) XOR DI(164) XOR DI(3) XOR DI(503) XOR DI(483) XOR DI(231) XOR DI(70) XOR DI(389) XOR DI(351) XOR DI(71) XOR DI(317) XOR DI(478) XOR DI(280) XOR DI(55) XOR DI(423) XOR DI(408) XOR DI(172) XOR DI(356) XOR DI(58) XOR DI(279) XOR DI(321) XOR DI(459) XOR DI(217) XOR DI(95) XOR DI(324) XOR DI(314) XOR DI(35) XOR DI(439) XOR DI(121) XOR DI(63) XOR DI(187) XOR DI(220) XOR DI(463) XOR DI(325) XOR DI(169) XOR DI(396) XOR DI(481) XOR DI(14) XOR DI(410) XOR DI(460) XOR DI(424) XOR DI(158) XOR DI(243) XOR DI(380) XOR DI(270) XOR DI(239) XOR DI(208) XOR DI(305) XOR DI(5) XOR DI(188) XOR DI(371) XOR DI(221) XOR DI(363) XOR DI(372) XOR DI(210) XOR DI(91) XOR DI(170) XOR DI(219) XOR DI(126) XOR DI(379) XOR DI(150) XOR DI(74) XOR DI(100) XOR DI(295) XOR DI(28) XOR DI(425) XOR DI(99) XOR DI(337) XOR DI(413) XOR DI(165) XOR DI(477) XOR DI(49) XOR DI(166) XOR DI(403) XOR DI(211) XOR DI(308) XOR DI(115) XOR DI(475) XOR DI(404) XOR DI(277) XOR DI(21) XOR DI(264) XOR DI(233) XOR DI(202) XOR DI(215) XOR DI(291) XOR DI(204) XOR DI(111) XOR DI(364) XOR DI(388) XOR DI(300) XOR DI(24) XOR DI(120) XOR DI(373) XOR DI(144) XOR DI(93) XOR DI(420) XOR DI(159) XOR DI(160) XOR DI(397) XOR DI(205) XOR DI(83) XOR DI(209) XOR DI(129) XOR DI(18) XOR DI(470) XOR DI(207) XOR DI(114) XOR DI(138) XOR DI(154) XOR DI(391) XOR DI(441) XOR DI(103) XOR DI(298) XOR DI(352) XOR DI(12) XOR DI(186) XOR DI(6) XOR DI(102) XOR DI(25) XOR DI(180) XOR DI(340) XOR DI(0) XOR DI(13) XOR DI(1) XOR DI(495) XOR DI(507);
   DO(12) <= DI(258) XOR DI(323) XOR DI(324) XOR DI(489) XOR DI(262) XOR DI(327) XOR DI(49) XOR DI(77) XOR DI(285) XOR DI(462) XOR DI(178) XOR DI(263) XOR DI(363) XOR DI(329) XOR DI(119) XOR DI(172) XOR DI(76) XOR DI(433) XOR DI(179) XOR DI(500) XOR DI(351) XOR DI(319) XOR DI(153) XOR DI(102) XOR DI(396) XOR DI(93) XOR DI(452) XOR DI(486) XOR DI(259) XOR DI(286) XOR DI(308) XOR DI(124) XOR DI(248) XOR DI(51) XOR DI(168) XOR DI(275) XOR DI(69) XOR DI(226) XOR DI(137) XOR DI(87) XOR DI(269) XOR DI(399) XOR DI(238) XOR DI(53) XOR DI(487) XOR DI(224) XOR DI(287) XOR DI(81) XOR DI(384) XOR DI(79) XOR DI(289) XOR DI(125) XOR DI(129) XOR DI(33) XOR DI(430) XOR DI(144) XOR DI(98) XOR DI(418) XOR DI(491) XOR DI(503) XOR DI(67) XOR DI(348) XOR DI(68) XOR DI(277) XOR DI(335) XOR DI(276) XOR DI(406) XOR DI(245) XOR DI(42) XOR DI(184) XOR DI(85) XOR DI(113) XOR DI(393) XOR DI(11) XOR DI(457) XOR DI(377) XOR DI(368) XOR DI(227) XOR DI(95) XOR DI(207) XOR DI(367) XOR DI(88) XOR DI(303) XOR DI(192) XOR DI(408) XOR DI(147) XOR DI(97) XOR DI(422) XOR DI(334) XOR DI(495) XOR DI(270) XOR DI(312) XOR DI(54) XOR DI(387) XOR DI(451) XOR DI(403) XOR DI(261) XOR DI(288) XOR DI(201) XOR DI(297) XOR DI(473) XOR DI(370) XOR DI(141) XOR DI(417) XOR DI(12) XOR DI(290) XOR DI(355) XOR DI(126) XOR DI(34) XOR DI(388) XOR DI(431) XOR DI(9) XOR DI(3) XOR DI(419) XOR DI(165) XOR DI(4) XOR DI(504) XOR DI(484) XOR DI(232) XOR DI(71) XOR DI(390) XOR DI(352) XOR DI(72) XOR DI(318) XOR DI(479) XOR DI(281) XOR DI(56) XOR DI(424) XOR DI(409) XOR DI(173) XOR DI(357) XOR DI(59) XOR DI(280) XOR DI(322) XOR DI(460) XOR DI(218) XOR DI(96) XOR DI(325) XOR DI(315) XOR DI(36) XOR DI(440) XOR DI(122) XOR DI(64) XOR DI(188) XOR DI(221) XOR DI(464) XOR DI(326) XOR DI(170) XOR DI(397) XOR DI(482) XOR DI(15) XOR DI(411) XOR DI(461) XOR DI(425) XOR DI(159) XOR DI(244) XOR DI(381) XOR DI(271) XOR DI(240) XOR DI(209) XOR DI(306) XOR DI(6) XOR DI(189) XOR DI(372) XOR DI(222) XOR DI(364) XOR DI(373) XOR DI(211) XOR DI(92) XOR DI(171) XOR DI(220) XOR DI(127) XOR DI(380) XOR DI(151) XOR DI(75) XOR DI(101) XOR DI(296) XOR DI(29) XOR DI(426) XOR DI(100) XOR DI(338) XOR DI(414) XOR DI(166) XOR DI(478) XOR DI(50) XOR DI(167) XOR DI(404) XOR DI(212) XOR DI(309) XOR DI(116) XOR DI(476) XOR DI(405) XOR DI(278) XOR DI(22) XOR DI(265) XOR DI(234) XOR DI(203) XOR DI(216) XOR DI(292) XOR DI(205) XOR DI(112) XOR DI(365) XOR DI(389) XOR DI(301) XOR DI(25) XOR DI(121) XOR DI(374) XOR DI(145) XOR DI(94) XOR DI(421) XOR DI(160) XOR DI(161) XOR DI(398) XOR DI(206) XOR DI(84) XOR DI(210) XOR DI(130) XOR DI(19) XOR DI(471) XOR DI(208) XOR DI(115) XOR DI(139) XOR DI(155) XOR DI(392) XOR DI(442) XOR DI(104) XOR DI(299) XOR DI(353) XOR DI(13) XOR DI(187) XOR DI(7) XOR DI(103) XOR DI(26) XOR DI(181) XOR DI(341) XOR DI(1) XOR DI(14) XOR DI(2) XOR DI(496) XOR DI(508);
   DO(13) <= DI(259) XOR DI(324) XOR DI(325) XOR DI(490) XOR DI(263) XOR DI(328) XOR DI(50) XOR DI(78) XOR DI(286) XOR DI(463) XOR DI(179) XOR DI(264) XOR DI(364) XOR DI(330) XOR DI(120) XOR DI(173) XOR DI(77) XOR DI(434) XOR DI(180) XOR DI(0) XOR DI(501) XOR DI(352) XOR DI(320) XOR DI(154) XOR DI(103) XOR DI(397) XOR DI(94) XOR DI(453) XOR DI(487) XOR DI(260) XOR DI(287) XOR DI(309) XOR DI(125) XOR DI(249) XOR DI(52) XOR DI(169) XOR DI(276) XOR DI(70) XOR DI(227) XOR DI(138) XOR DI(88) XOR DI(270) XOR DI(400) XOR DI(239) XOR DI(54) XOR DI(488) XOR DI(225) XOR DI(288) XOR DI(82) XOR DI(385) XOR DI(80) XOR DI(290) XOR DI(126) XOR DI(130) XOR DI(34) XOR DI(431) XOR DI(145) XOR DI(99) XOR DI(419) XOR DI(492) XOR DI(504) XOR DI(68) XOR DI(349) XOR DI(69) XOR DI(278) XOR DI(336) XOR DI(277) XOR DI(407) XOR DI(246) XOR DI(43) XOR DI(185) XOR DI(86) XOR DI(114) XOR DI(394) XOR DI(12) XOR DI(458) XOR DI(378) XOR DI(369) XOR DI(228) XOR DI(96) XOR DI(208) XOR DI(368) XOR DI(89) XOR DI(304) XOR DI(193) XOR DI(409) XOR DI(148) XOR DI(98) XOR DI(423) XOR DI(335) XOR DI(496) XOR DI(271) XOR DI(313) XOR DI(55) XOR DI(388) XOR DI(452) XOR DI(404) XOR DI(262) XOR DI(289) XOR DI(202) XOR DI(298) XOR DI(474) XOR DI(371) XOR DI(142) XOR DI(418) XOR DI(13) XOR DI(291) XOR DI(356) XOR DI(127) XOR DI(35) XOR DI(389) XOR DI(432) XOR DI(10) XOR DI(4) XOR DI(420) XOR DI(166) XOR DI(5) XOR DI(505) XOR DI(485) XOR DI(233) XOR DI(72) XOR DI(391) XOR DI(353) XOR DI(73) XOR DI(319) XOR DI(480) XOR DI(282) XOR DI(57) XOR DI(425) XOR DI(410) XOR DI(174) XOR DI(358) XOR DI(60) XOR DI(281) XOR DI(323) XOR DI(461) XOR DI(219) XOR DI(97) XOR DI(326) XOR DI(316) XOR DI(37) XOR DI(441) XOR DI(123) XOR DI(65) XOR DI(189) XOR DI(222) XOR DI(465) XOR DI(327) XOR DI(171) XOR DI(398) XOR DI(483) XOR DI(16) XOR DI(412) XOR DI(462) XOR DI(426) XOR DI(160) XOR DI(245) XOR DI(382) XOR DI(272) XOR DI(241) XOR DI(210) XOR DI(307) XOR DI(7) XOR DI(190) XOR DI(373) XOR DI(223) XOR DI(365) XOR DI(374) XOR DI(212) XOR DI(93) XOR DI(172) XOR DI(221) XOR DI(128) XOR DI(381) XOR DI(152) XOR DI(76) XOR DI(102) XOR DI(297) XOR DI(30) XOR DI(427) XOR DI(101) XOR DI(339) XOR DI(415) XOR DI(167) XOR DI(479) XOR DI(51) XOR DI(168) XOR DI(405) XOR DI(213) XOR DI(310) XOR DI(117) XOR DI(477) XOR DI(406) XOR DI(279) XOR DI(23) XOR DI(266) XOR DI(235) XOR DI(204) XOR DI(217) XOR DI(293) XOR DI(206) XOR DI(113) XOR DI(366) XOR DI(390) XOR DI(302) XOR DI(26) XOR DI(122) XOR DI(375) XOR DI(146) XOR DI(95) XOR DI(422) XOR DI(161) XOR DI(162) XOR DI(399) XOR DI(207) XOR DI(85) XOR DI(211) XOR DI(131) XOR DI(20) XOR DI(472) XOR DI(209) XOR DI(116) XOR DI(140) XOR DI(156) XOR DI(393) XOR DI(443) XOR DI(105) XOR DI(300) XOR DI(354) XOR DI(14) XOR DI(188) XOR DI(8) XOR DI(104) XOR DI(27) XOR DI(182) XOR DI(342) XOR DI(2) XOR DI(15) XOR DI(3) XOR DI(497) XOR DI(509);
   DO(14) <= DI(260) XOR DI(325) XOR DI(326) XOR DI(491) XOR DI(264) XOR DI(329) XOR DI(51) XOR DI(79) XOR DI(287) XOR DI(464) XOR DI(180) XOR DI(265) XOR DI(365) XOR DI(331) XOR DI(121) XOR DI(174) XOR DI(78) XOR DI(435) XOR DI(181) XOR DI(1) XOR DI(502) XOR DI(353) XOR DI(321) XOR DI(155) XOR DI(104) XOR DI(398) XOR DI(95) XOR DI(454) XOR DI(488) XOR DI(261) XOR DI(288) XOR DI(310) XOR DI(126) XOR DI(250) XOR DI(53) XOR DI(170) XOR DI(277) XOR DI(71) XOR DI(228) XOR DI(139) XOR DI(89) XOR DI(271) XOR DI(401) XOR DI(240) XOR DI(55) XOR DI(489) XOR DI(226) XOR DI(289) XOR DI(83) XOR DI(386) XOR DI(81) XOR DI(291) XOR DI(127) XOR DI(131) XOR DI(35) XOR DI(432) XOR DI(146) XOR DI(100) XOR DI(420) XOR DI(493) XOR DI(505) XOR DI(69) XOR DI(350) XOR DI(70) XOR DI(279) XOR DI(337) XOR DI(278) XOR DI(408) XOR DI(247) XOR DI(44) XOR DI(186) XOR DI(87) XOR DI(115) XOR DI(395) XOR DI(13) XOR DI(459) XOR DI(379) XOR DI(370) XOR DI(229) XOR DI(97) XOR DI(209) XOR DI(369) XOR DI(90) XOR DI(305) XOR DI(194) XOR DI(410) XOR DI(149) XOR DI(99) XOR DI(424) XOR DI(336) XOR DI(497) XOR DI(272) XOR DI(314) XOR DI(56) XOR DI(389) XOR DI(453) XOR DI(405) XOR DI(263) XOR DI(290) XOR DI(203) XOR DI(299) XOR DI(475) XOR DI(372) XOR DI(143) XOR DI(419) XOR DI(14) XOR DI(292) XOR DI(357) XOR DI(128) XOR DI(36) XOR DI(390) XOR DI(433) XOR DI(11) XOR DI(5) XOR DI(421) XOR DI(167) XOR DI(6) XOR DI(506) XOR DI(486) XOR DI(234) XOR DI(73) XOR DI(392) XOR DI(354) XOR DI(74) XOR DI(320) XOR DI(481) XOR DI(283) XOR DI(58) XOR DI(426) XOR DI(411) XOR DI(175) XOR DI(359) XOR DI(61) XOR DI(282) XOR DI(324) XOR DI(462) XOR DI(220) XOR DI(98) XOR DI(327) XOR DI(317) XOR DI(38) XOR DI(442) XOR DI(124) XOR DI(66) XOR DI(190) XOR DI(223) XOR DI(466) XOR DI(328) XOR DI(172) XOR DI(399) XOR DI(484) XOR DI(17) XOR DI(413) XOR DI(463) XOR DI(427) XOR DI(161) XOR DI(246) XOR DI(383) XOR DI(273) XOR DI(242) XOR DI(211) XOR DI(308) XOR DI(8) XOR DI(191) XOR DI(374) XOR DI(224) XOR DI(366) XOR DI(375) XOR DI(213) XOR DI(94) XOR DI(173) XOR DI(222) XOR DI(129) XOR DI(382) XOR DI(153) XOR DI(77) XOR DI(103) XOR DI(298) XOR DI(31) XOR DI(428) XOR DI(102) XOR DI(340) XOR DI(416) XOR DI(168) XOR DI(480) XOR DI(52) XOR DI(169) XOR DI(406) XOR DI(214) XOR DI(311) XOR DI(118) XOR DI(478) XOR DI(407) XOR DI(280) XOR DI(24) XOR DI(267) XOR DI(236) XOR DI(205) XOR DI(218) XOR DI(294) XOR DI(207) XOR DI(114) XOR DI(367) XOR DI(391) XOR DI(303) XOR DI(27) XOR DI(123) XOR DI(376) XOR DI(147) XOR DI(96) XOR DI(423) XOR DI(162) XOR DI(163) XOR DI(400) XOR DI(208) XOR DI(86) XOR DI(212) XOR DI(132) XOR DI(21) XOR DI(473) XOR DI(210) XOR DI(117) XOR DI(141) XOR DI(157) XOR DI(394) XOR DI(444) XOR DI(106) XOR DI(301) XOR DI(355) XOR DI(15) XOR DI(189) XOR DI(9) XOR DI(105) XOR DI(28) XOR DI(183) XOR DI(343) XOR DI(3) XOR DI(16) XOR DI(4) XOR DI(498) XOR DI(510);
   DO(15) <= DI(261) XOR DI(326) XOR DI(327) XOR DI(492) XOR DI(265) XOR DI(330) XOR DI(52) XOR DI(80) XOR DI(288) XOR DI(465) XOR DI(181) XOR DI(266) XOR DI(366) XOR DI(332) XOR DI(122) XOR DI(175) XOR DI(79) XOR DI(436) XOR DI(182) XOR DI(2) XOR DI(503) XOR DI(354) XOR DI(322) XOR DI(156) XOR DI(105) XOR DI(399) XOR DI(96) XOR DI(455) XOR DI(489) XOR DI(262) XOR DI(289) XOR DI(311) XOR DI(127) XOR DI(251) XOR DI(54) XOR DI(171) XOR DI(278) XOR DI(72) XOR DI(229) XOR DI(140) XOR DI(90) XOR DI(272) XOR DI(402) XOR DI(241) XOR DI(56) XOR DI(490) XOR DI(227) XOR DI(290) XOR DI(84) XOR DI(387) XOR DI(82) XOR DI(292) XOR DI(128) XOR DI(132) XOR DI(36) XOR DI(433) XOR DI(147) XOR DI(101) XOR DI(421) XOR DI(494) XOR DI(506) XOR DI(70) XOR DI(351) XOR DI(71) XOR DI(280) XOR DI(338) XOR DI(279) XOR DI(409) XOR DI(248) XOR DI(45) XOR DI(187) XOR DI(88) XOR DI(116) XOR DI(396) XOR DI(14) XOR DI(460) XOR DI(380) XOR DI(371) XOR DI(230) XOR DI(98) XOR DI(210) XOR DI(370) XOR DI(91) XOR DI(306) XOR DI(195) XOR DI(411) XOR DI(150) XOR DI(100) XOR DI(425) XOR DI(337) XOR DI(498) XOR DI(273) XOR DI(315) XOR DI(57) XOR DI(390) XOR DI(454) XOR DI(406) XOR DI(264) XOR DI(291) XOR DI(204) XOR DI(300) XOR DI(476) XOR DI(373) XOR DI(144) XOR DI(420) XOR DI(15) XOR DI(293) XOR DI(358) XOR DI(129) XOR DI(37) XOR DI(391) XOR DI(434) XOR DI(12) XOR DI(6) XOR DI(422) XOR DI(168) XOR DI(7) XOR DI(507) XOR DI(487) XOR DI(235) XOR DI(74) XOR DI(393) XOR DI(355) XOR DI(75) XOR DI(321) XOR DI(482) XOR DI(284) XOR DI(59) XOR DI(427) XOR DI(412) XOR DI(176) XOR DI(360) XOR DI(62) XOR DI(283) XOR DI(325) XOR DI(463) XOR DI(221) XOR DI(99) XOR DI(328) XOR DI(318) XOR DI(39) XOR DI(443) XOR DI(125) XOR DI(67) XOR DI(191) XOR DI(224) XOR DI(467) XOR DI(329) XOR DI(173) XOR DI(400) XOR DI(485) XOR DI(18) XOR DI(414) XOR DI(464) XOR DI(428) XOR DI(162) XOR DI(247) XOR DI(384) XOR DI(274) XOR DI(243) XOR DI(212) XOR DI(309) XOR DI(9) XOR DI(192) XOR DI(375) XOR DI(225) XOR DI(367) XOR DI(376) XOR DI(214) XOR DI(95) XOR DI(174) XOR DI(223) XOR DI(130) XOR DI(383) XOR DI(154) XOR DI(78) XOR DI(104) XOR DI(299) XOR DI(32) XOR DI(429) XOR DI(103) XOR DI(341) XOR DI(417) XOR DI(169) XOR DI(481) XOR DI(53) XOR DI(170) XOR DI(407) XOR DI(215) XOR DI(312) XOR DI(119) XOR DI(479) XOR DI(408) XOR DI(281) XOR DI(25) XOR DI(268) XOR DI(237) XOR DI(206) XOR DI(219) XOR DI(295) XOR DI(208) XOR DI(115) XOR DI(368) XOR DI(392) XOR DI(304) XOR DI(28) XOR DI(124) XOR DI(377) XOR DI(148) XOR DI(97) XOR DI(424) XOR DI(163) XOR DI(164) XOR DI(401) XOR DI(209) XOR DI(87) XOR DI(213) XOR DI(133) XOR DI(22) XOR DI(474) XOR DI(211) XOR DI(118) XOR DI(142) XOR DI(158) XOR DI(395) XOR DI(445) XOR DI(107) XOR DI(302) XOR DI(356) XOR DI(16) XOR DI(190) XOR DI(10) XOR DI(106) XOR DI(29) XOR DI(184) XOR DI(344) XOR DI(4) XOR DI(17) XOR DI(5) XOR DI(499) XOR DI(511);
   DO(16) <= DI(262) XOR DI(327) XOR DI(124) XOR DI(328) XOR DI(257) XOR DI(78) XOR DI(286) XOR DI(51) XOR DI(493) XOR DI(266) XOR DI(399) XOR DI(331) XOR DI(53) XOR DI(487) XOR DI(200) XOR DI(81) XOR DI(416) XOR DI(289) XOR DI(354) XOR DI(466) XOR DI(503) XOR DI(386) XOR DI(182) XOR DI(267) XOR DI(302) XOR DI(367) XOR DI(333) XOR DI(123) XOR DI(176) XOR DI(288) XOR DI(417) XOR DI(80) XOR DI(437) XOR DI(467) XOR DI(431) XOR DI(183) XOR DI(343) XOR DI(3) XOR DI(504) XOR DI(355) XOR DI(323) XOR DI(451) XOR DI(62) XOR DI(184) XOR DI(157) XOR DI(106) XOR DI(4) XOR DI(400) XOR DI(97) XOR DI(194) XOR DI(48) XOR DI(178) XOR DI(456) XOR DI(490) XOR DI(263) XOR DI(290) XOR DI(387) XOR DI(312) XOR DI(128) XOR DI(113) XOR DI(153) XOR DI(433) XOR DI(506) XOR DI(252) XOR DI(351) XOR DI(55) XOR DI(462) XOR DI(42) XOR DI(172) XOR DI(279) XOR DI(321) XOR DI(459) XOR DI(217) XOR DI(324) XOR DI(452) XOR DI(449) XOR DI(35) XOR DI(439) XOR DI(481) XOR DI(73) XOR DI(197) XOR DI(230) XOR DI(363) XOR DI(141) XOR DI(91) XOR DI(255) XOR DI(195) XOR DI(273) XOR DI(403) XOR DI(242) XOR DI(57) XOR DI(179) XOR DI(457) XOR DI(21) XOR DI(406) XOR DI(491) XOR DI(264) XOR DI(233) XOR DI(202) XOR DI(228) XOR DI(291) XOR DI(85) XOR DI(388) XOR DI(24) XOR DI(375) XOR DI(144) XOR DI(93) XOR DI(83) XOR DI(293) XOR DI(304) XOR DI(129) XOR DI(114) XOR DI(138) XOR DI(133) XOR DI(37) XOR DI(154) XOR DI(434) XOR DI(12) XOR DI(148) XOR DI(102) XOR DI(422) XOR DI(340) XOR DI(168) XOR DI(495) XOR DI(507) XOR DI(484) XOR DI(71) XOR DI(253) XOR DI(260) XOR DI(352) XOR DI(72) XOR DI(318) XOR DI(281) XOR DI(339) XOR DI(173) XOR DI(280) XOR DI(410) XOR DI(249) XOR DI(218) XOR DI(46) XOR DI(239) XOR DI(315) XOR DI(36) XOR DI(440) XOR DI(122) XOR DI(64) XOR DI(188) XOR DI(89) XOR DI(117) XOR DI(397) XOR DI(15) XOR DI(411) XOR DI(461) XOR DI(251) XOR DI(381) XOR DI(47) XOR DI(150) XOR DI(235) XOR DI(372) XOR DI(231) XOR DI(99) XOR DI(298) XOR DI(211) XOR DI(371) XOR DI(92) XOR DI(395) XOR DI(307) XOR DI(445) XOR DI(31) XOR DI(196) XOR DI(380) XOR DI(412) XOR DI(151) XOR DI(101) XOR DI(350) XOR DI(146) XOR DI(426) XOR DI(427) XOR DI(338) XOR DI(414) XOR DI(499) XOR DI(478) XOR DI(247) XOR DI(346) XOR DI(50) XOR DI(167) XOR DI(274) XOR DI(316) XOR DI(454) XOR DI(243) XOR DI(90) XOR DI(447) XOR DI(309) XOR DI(58) XOR DI(458) XOR DI(320) XOR DI(391) XOR DI(278) XOR DI(455) XOR DI(22) XOR DI(407) XOR DI(265) XOR DI(203) XOR DI(311) XOR DI(0) XOR DI(229) XOR DI(292) XOR DI(205) XOR DI(112) XOR DI(136) XOR DI(389) XOR DI(301) XOR DI(477) XOR DI(190) XOR DI(121) XOR DI(374) XOR DI(145) XOR DI(140) XOR DI(94) XOR DI(421) XOR DI(44) XOR DI(398) XOR DI(314) XOR DI(16) XOR DI(294) XOR DI(359) XOR DI(130) XOR DI(38) XOR DI(392) XOR DI(435) XOR DI(13) XOR DI(32) XOR DI(7) XOR DI(103) XOR DI(423) XOR DI(341) XOR DI(1) XOR DI(20) XOR DI(169) XOR DI(8) XOR DI(2) XOR DI(496) XOR DI(502) XOR DI(508);
   DO(17) <= DI(263) XOR DI(328) XOR DI(125) XOR DI(329) XOR DI(258) XOR DI(79) XOR DI(287) XOR DI(52) XOR DI(494) XOR DI(267) XOR DI(400) XOR DI(332) XOR DI(54) XOR DI(488) XOR DI(201) XOR DI(82) XOR DI(417) XOR DI(290) XOR DI(355) XOR DI(467) XOR DI(504) XOR DI(387) XOR DI(183) XOR DI(268) XOR DI(303) XOR DI(368) XOR DI(334) XOR DI(124) XOR DI(177) XOR DI(289) XOR DI(418) XOR DI(81) XOR DI(438) XOR DI(468) XOR DI(432) XOR DI(184) XOR DI(344) XOR DI(4) XOR DI(505) XOR DI(356) XOR DI(324) XOR DI(452) XOR DI(63) XOR DI(185) XOR DI(158) XOR DI(107) XOR DI(5) XOR DI(401) XOR DI(98) XOR DI(195) XOR DI(49) XOR DI(179) XOR DI(457) XOR DI(491) XOR DI(264) XOR DI(291) XOR DI(388) XOR DI(313) XOR DI(129) XOR DI(114) XOR DI(154) XOR DI(434) XOR DI(507) XOR DI(253) XOR DI(352) XOR DI(56) XOR DI(463) XOR DI(43) XOR DI(173) XOR DI(280) XOR DI(322) XOR DI(460) XOR DI(218) XOR DI(325) XOR DI(453) XOR DI(450) XOR DI(36) XOR DI(440) XOR DI(482) XOR DI(74) XOR DI(198) XOR DI(231) XOR DI(364) XOR DI(142) XOR DI(92) XOR DI(256) XOR DI(196) XOR DI(274) XOR DI(404) XOR DI(243) XOR DI(58) XOR DI(180) XOR DI(458) XOR DI(22) XOR DI(407) XOR DI(492) XOR DI(265) XOR DI(234) XOR DI(203) XOR DI(229) XOR DI(292) XOR DI(86) XOR DI(389) XOR DI(25) XOR DI(376) XOR DI(145) XOR DI(94) XOR DI(84) XOR DI(294) XOR DI(305) XOR DI(130) XOR DI(115) XOR DI(139) XOR DI(134) XOR DI(38) XOR DI(155) XOR DI(435) XOR DI(13) XOR DI(149) XOR DI(103) XOR DI(423) XOR DI(341) XOR DI(169) XOR DI(496) XOR DI(508) XOR DI(485) XOR DI(72) XOR DI(254) XOR DI(261) XOR DI(353) XOR DI(73) XOR DI(319) XOR DI(282) XOR DI(340) XOR DI(174) XOR DI(281) XOR DI(411) XOR DI(250) XOR DI(219) XOR DI(47) XOR DI(240) XOR DI(316) XOR DI(37) XOR DI(441) XOR DI(123) XOR DI(65) XOR DI(189) XOR DI(90) XOR DI(118) XOR DI(398) XOR DI(16) XOR DI(412) XOR DI(462) XOR DI(252) XOR DI(382) XOR DI(48) XOR DI(151) XOR DI(236) XOR DI(373) XOR DI(232) XOR DI(100) XOR DI(299) XOR DI(212) XOR DI(372) XOR DI(93) XOR DI(396) XOR DI(308) XOR DI(446) XOR DI(32) XOR DI(197) XOR DI(381) XOR DI(413) XOR DI(152) XOR DI(102) XOR DI(351) XOR DI(147) XOR DI(427) XOR DI(428) XOR DI(339) XOR DI(415) XOR DI(500) XOR DI(479) XOR DI(248) XOR DI(347) XOR DI(51) XOR DI(168) XOR DI(275) XOR DI(317) XOR DI(455) XOR DI(244) XOR DI(91) XOR DI(448) XOR DI(310) XOR DI(59) XOR DI(459) XOR DI(321) XOR DI(392) XOR DI(279) XOR DI(456) XOR DI(23) XOR DI(408) XOR DI(266) XOR DI(204) XOR DI(312) XOR DI(1) XOR DI(230) XOR DI(293) XOR DI(206) XOR DI(113) XOR DI(137) XOR DI(390) XOR DI(302) XOR DI(478) XOR DI(191) XOR DI(122) XOR DI(375) XOR DI(146) XOR DI(141) XOR DI(95) XOR DI(422) XOR DI(45) XOR DI(399) XOR DI(315) XOR DI(17) XOR DI(295) XOR DI(360) XOR DI(131) XOR DI(39) XOR DI(393) XOR DI(436) XOR DI(14) XOR DI(33) XOR DI(8) XOR DI(104) XOR DI(424) XOR DI(342) XOR DI(2) XOR DI(21) XOR DI(170) XOR DI(9) XOR DI(3) XOR DI(497) XOR DI(503) XOR DI(509);
   DO(18) <= DI(264) XOR DI(329) XOR DI(126) XOR DI(330) XOR DI(259) XOR DI(80) XOR DI(288) XOR DI(53) XOR DI(495) XOR DI(268) XOR DI(401) XOR DI(333) XOR DI(55) XOR DI(489) XOR DI(202) XOR DI(83) XOR DI(418) XOR DI(291) XOR DI(356) XOR DI(468) XOR DI(505) XOR DI(388) XOR DI(184) XOR DI(269) XOR DI(304) XOR DI(369) XOR DI(335) XOR DI(125) XOR DI(178) XOR DI(290) XOR DI(419) XOR DI(82) XOR DI(439) XOR DI(469) XOR DI(433) XOR DI(185) XOR DI(345) XOR DI(5) XOR DI(506) XOR DI(357) XOR DI(325) XOR DI(453) XOR DI(64) XOR DI(186) XOR DI(159) XOR DI(108) XOR DI(6) XOR DI(402) XOR DI(99) XOR DI(196) XOR DI(50) XOR DI(180) XOR DI(458) XOR DI(492) XOR DI(265) XOR DI(292) XOR DI(389) XOR DI(314) XOR DI(130) XOR DI(115) XOR DI(155) XOR DI(435) XOR DI(508) XOR DI(254) XOR DI(353) XOR DI(57) XOR DI(464) XOR DI(44) XOR DI(174) XOR DI(281) XOR DI(323) XOR DI(461) XOR DI(219) XOR DI(326) XOR DI(454) XOR DI(451) XOR DI(37) XOR DI(441) XOR DI(483) XOR DI(75) XOR DI(199) XOR DI(232) XOR DI(365) XOR DI(143) XOR DI(93) XOR DI(257) XOR DI(197) XOR DI(275) XOR DI(405) XOR DI(244) XOR DI(59) XOR DI(181) XOR DI(459) XOR DI(23) XOR DI(408) XOR DI(493) XOR DI(266) XOR DI(235) XOR DI(204) XOR DI(230) XOR DI(293) XOR DI(87) XOR DI(390) XOR DI(26) XOR DI(377) XOR DI(146) XOR DI(95) XOR DI(85) XOR DI(295) XOR DI(306) XOR DI(131) XOR DI(116) XOR DI(140) XOR DI(135) XOR DI(39) XOR DI(156) XOR DI(436) XOR DI(14) XOR DI(150) XOR DI(104) XOR DI(424) XOR DI(342) XOR DI(170) XOR DI(497) XOR DI(509) XOR DI(486) XOR DI(73) XOR DI(255) XOR DI(262) XOR DI(354) XOR DI(74) XOR DI(320) XOR DI(283) XOR DI(341) XOR DI(175) XOR DI(282) XOR DI(412) XOR DI(251) XOR DI(220) XOR DI(48) XOR DI(241) XOR DI(317) XOR DI(38) XOR DI(442) XOR DI(124) XOR DI(66) XOR DI(190) XOR DI(91) XOR DI(119) XOR DI(399) XOR DI(17) XOR DI(413) XOR DI(463) XOR DI(253) XOR DI(383) XOR DI(49) XOR DI(152) XOR DI(237) XOR DI(374) XOR DI(233) XOR DI(101) XOR DI(300) XOR DI(213) XOR DI(373) XOR DI(94) XOR DI(397) XOR DI(309) XOR DI(447) XOR DI(33) XOR DI(198) XOR DI(382) XOR DI(414) XOR DI(153) XOR DI(103) XOR DI(352) XOR DI(148) XOR DI(428) XOR DI(429) XOR DI(340) XOR DI(0) XOR DI(416) XOR DI(501) XOR DI(480) XOR DI(249) XOR DI(348) XOR DI(52) XOR DI(169) XOR DI(276) XOR DI(318) XOR DI(456) XOR DI(245) XOR DI(92) XOR DI(449) XOR DI(311) XOR DI(60) XOR DI(460) XOR DI(322) XOR DI(393) XOR DI(280) XOR DI(457) XOR DI(24) XOR DI(409) XOR DI(267) XOR DI(205) XOR DI(313) XOR DI(2) XOR DI(231) XOR DI(294) XOR DI(207) XOR DI(114) XOR DI(138) XOR DI(391) XOR DI(303) XOR DI(479) XOR DI(192) XOR DI(123) XOR DI(376) XOR DI(147) XOR DI(142) XOR DI(96) XOR DI(423) XOR DI(46) XOR DI(400) XOR DI(316) XOR DI(18) XOR DI(296) XOR DI(361) XOR DI(132) XOR DI(40) XOR DI(394) XOR DI(437) XOR DI(15) XOR DI(34) XOR DI(9) XOR DI(105) XOR DI(425) XOR DI(343) XOR DI(3) XOR DI(22) XOR DI(171) XOR DI(10) XOR DI(4) XOR DI(498) XOR DI(504) XOR DI(510);
   DO(19) <= DI(265) XOR DI(330) XOR DI(127) XOR DI(331) XOR DI(260) XOR DI(81) XOR DI(289) XOR DI(54) XOR DI(496) XOR DI(269) XOR DI(402) XOR DI(334) XOR DI(56) XOR DI(490) XOR DI(203) XOR DI(84) XOR DI(419) XOR DI(292) XOR DI(357) XOR DI(469) XOR DI(506) XOR DI(389) XOR DI(185) XOR DI(270) XOR DI(305) XOR DI(370) XOR DI(336) XOR DI(126) XOR DI(179) XOR DI(291) XOR DI(420) XOR DI(83) XOR DI(440) XOR DI(470) XOR DI(434) XOR DI(186) XOR DI(346) XOR DI(6) XOR DI(507) XOR DI(358) XOR DI(326) XOR DI(454) XOR DI(65) XOR DI(187) XOR DI(160) XOR DI(109) XOR DI(7) XOR DI(403) XOR DI(100) XOR DI(197) XOR DI(51) XOR DI(181) XOR DI(459) XOR DI(493) XOR DI(266) XOR DI(293) XOR DI(390) XOR DI(315) XOR DI(131) XOR DI(116) XOR DI(156) XOR DI(436) XOR DI(509) XOR DI(255) XOR DI(354) XOR DI(58) XOR DI(465) XOR DI(45) XOR DI(175) XOR DI(282) XOR DI(324) XOR DI(462) XOR DI(220) XOR DI(327) XOR DI(455) XOR DI(452) XOR DI(38) XOR DI(442) XOR DI(484) XOR DI(76) XOR DI(200) XOR DI(233) XOR DI(366) XOR DI(144) XOR DI(94) XOR DI(258) XOR DI(198) XOR DI(276) XOR DI(406) XOR DI(245) XOR DI(60) XOR DI(182) XOR DI(460) XOR DI(24) XOR DI(409) XOR DI(494) XOR DI(267) XOR DI(236) XOR DI(205) XOR DI(231) XOR DI(294) XOR DI(88) XOR DI(391) XOR DI(27) XOR DI(378) XOR DI(147) XOR DI(96) XOR DI(86) XOR DI(296) XOR DI(307) XOR DI(132) XOR DI(117) XOR DI(141) XOR DI(136) XOR DI(40) XOR DI(157) XOR DI(437) XOR DI(15) XOR DI(151) XOR DI(105) XOR DI(425) XOR DI(343) XOR DI(171) XOR DI(498) XOR DI(510) XOR DI(487) XOR DI(74) XOR DI(256) XOR DI(263) XOR DI(355) XOR DI(75) XOR DI(321) XOR DI(284) XOR DI(342) XOR DI(176) XOR DI(283) XOR DI(413) XOR DI(252) XOR DI(221) XOR DI(49) XOR DI(242) XOR DI(318) XOR DI(39) XOR DI(443) XOR DI(125) XOR DI(67) XOR DI(191) XOR DI(92) XOR DI(120) XOR DI(400) XOR DI(18) XOR DI(414) XOR DI(464) XOR DI(254) XOR DI(384) XOR DI(50) XOR DI(153) XOR DI(238) XOR DI(375) XOR DI(234) XOR DI(102) XOR DI(301) XOR DI(214) XOR DI(374) XOR DI(95) XOR DI(398) XOR DI(310) XOR DI(448) XOR DI(34) XOR DI(199) XOR DI(383) XOR DI(415) XOR DI(154) XOR DI(104) XOR DI(353) XOR DI(149) XOR DI(429) XOR DI(430) XOR DI(341) XOR DI(1) XOR DI(417) XOR DI(502) XOR DI(481) XOR DI(250) XOR DI(349) XOR DI(53) XOR DI(170) XOR DI(277) XOR DI(319) XOR DI(457) XOR DI(246) XOR DI(93) XOR DI(450) XOR DI(312) XOR DI(61) XOR DI(461) XOR DI(323) XOR DI(394) XOR DI(281) XOR DI(458) XOR DI(25) XOR DI(410) XOR DI(268) XOR DI(206) XOR DI(314) XOR DI(3) XOR DI(232) XOR DI(295) XOR DI(208) XOR DI(115) XOR DI(139) XOR DI(392) XOR DI(304) XOR DI(480) XOR DI(193) XOR DI(124) XOR DI(377) XOR DI(148) XOR DI(143) XOR DI(97) XOR DI(424) XOR DI(47) XOR DI(401) XOR DI(317) XOR DI(19) XOR DI(297) XOR DI(362) XOR DI(133) XOR DI(41) XOR DI(395) XOR DI(438) XOR DI(16) XOR DI(35) XOR DI(10) XOR DI(106) XOR DI(426) XOR DI(344) XOR DI(4) XOR DI(23) XOR DI(172) XOR DI(11) XOR DI(5) XOR DI(499) XOR DI(505) XOR DI(511);
   DO(20) <= DI(266) XOR DI(79) XOR DI(331) XOR DI(330) XOR DI(128) XOR DI(332) XOR DI(261) XOR DI(288) XOR DI(82) XOR DI(290) XOR DI(369) XOR DI(275) XOR DI(226) XOR DI(468) XOR DI(433) XOR DI(351) XOR DI(55) XOR DI(248) XOR DI(131) XOR DI(185) XOR DI(197) XOR DI(497) XOR DI(270) XOR DI(403) XOR DI(335) XOR DI(57) XOR DI(179) XOR DI(475) XOR DI(491) XOR DI(204) XOR DI(85) XOR DI(420) XOR DI(293) XOR DI(358) XOR DI(470) XOR DI(507) XOR DI(260) XOR DI(390) XOR DI(357) XOR DI(440) XOR DI(64) XOR DI(186) XOR DI(326) XOR DI(159) XOR DI(244) XOR DI(271) XOR DI(306) XOR DI(108) XOR DI(371) XOR DI(337) XOR DI(127) XOR DI(380) XOR DI(146) XOR DI(100) XOR DI(346) XOR DI(454) XOR DI(90) XOR DI(180) XOR DI(203) XOR DI(229) XOR DI(292) XOR DI(389) XOR DI(421) XOR DI(44) XOR DI(84) XOR DI(441) XOR DI(471) XOR DI(435) XOR DI(187) XOR DI(347) XOR DI(7) XOR DI(496) XOR DI(508) XOR DI(175) XOR DI(359) XOR DI(220) XOR DI(327) XOR DI(455) XOR DI(452) XOR DI(66) XOR DI(188) XOR DI(484) XOR DI(286) XOR DI(122) XOR DI(161) XOR DI(110) XOR DI(8) XOR DI(404) XOR DI(101) XOR DI(300) XOR DI(447) XOR DI(33) XOR DI(198) XOR DI(168) XOR DI(52) XOR DI(406) XOR DI(60) XOR DI(182) XOR DI(460) XOR DI(478) XOR DI(409) XOR DI(494) XOR DI(267) XOR DI(236) XOR DI(218) XOR DI(294) XOR DI(114) XOR DI(138) XOR DI(88) XOR DI(391) XOR DI(316) XOR DI(387) XOR DI(361) XOR DI(132) XOR DI(210) XOR DI(117) XOR DI(136) XOR DI(157) XOR DI(437) XOR DI(195) XOR DI(165) XOR DI(510) XOR DI(63) XOR DI(487) XOR DI(256) XOR DI(355) XOR DI(321) XOR DI(59) XOR DI(466) XOR DI(46) XOR DI(176) XOR DI(283) XOR DI(413) XOR DI(325) XOR DI(463) XOR DI(221) XOR DI(328) XOR DI(483) XOR DI(456) XOR DI(453) XOR DI(39) XOR DI(446) XOR DI(443) XOR DI(191) XOR DI(224) XOR DI(120) XOR DI(467) XOR DI(329) XOR DI(485) XOR DI(18) XOR DI(77) XOR DI(464) XOR DI(201) XOR DI(31) XOR DI(428) XOR DI(212) XOR DI(309) XOR DI(30) XOR DI(153) XOR DI(238) XOR DI(234) XOR DI(21) XOR DI(0) XOR DI(225) XOR DI(216) XOR DI(367) XOR DI(214) XOR DI(145) XOR DI(95) XOR DI(340) XOR DI(398) XOR DI(310) XOR DI(174) XOR DI(486) XOR DI(259) XOR DI(199) XOR DI(78) XOR DI(104) XOR DI(32) XOR DI(429) XOR DI(341) XOR DI(1) XOR DI(417) XOR DI(502) XOR DI(170) XOR DI(277) XOR DI(407) XOR DI(457) XOR DI(246) XOR DI(119) XOR DI(61) XOR DI(183) XOR DI(461) XOR DI(167) XOR DI(394) XOR DI(408) XOR DI(25) XOR DI(410) XOR DI(495) XOR DI(268) XOR DI(237) XOR DI(206) XOR DI(303) XOR DI(314) XOR DI(232) XOR DI(295) XOR DI(368) XOR DI(89) XOR DI(392) XOR DI(304) XOR DI(28) XOR DI(379) XOR DI(480) XOR DI(217) XOR DI(193) XOR DI(124) XOR DI(377) XOR DI(148) XOR DI(143) XOR DI(97) XOR DI(163) XOR DI(47) XOR DI(164) XOR DI(87) XOR DI(113) XOR DI(297) XOR DI(308) XOR DI(213) XOR DI(202) XOR DI(133) XOR DI(386) XOR DI(22) XOR DI(118) XOR DI(142) XOR DI(137) XOR DI(41) XOR DI(158) XOR DI(445) XOR DI(438) XOR DI(16) XOR DI(112) XOR DI(152) XOR DI(190) XOR DI(10) XOR DI(106) XOR DI(29) XOR DI(426) XOR DI(184) XOR DI(344) XOR DI(23) XOR DI(178) XOR DI(172) XOR DI(499) XOR DI(511);
   DO(21) <= DI(264) XOR DI(267) XOR DI(126) XOR DI(286) XOR DI(80) XOR DI(288) XOR DI(255) XOR DI(332) XOR DI(331) XOR DI(431) XOR DI(68) XOR DI(129) XOR DI(195) XOR DI(361) XOR DI(333) XOR DI(262) XOR DI(289) XOR DI(83) XOR DI(291) XOR DI(54) XOR DI(324) XOR DI(370) XOR DI(452) XOR DI(276) XOR DI(227) XOR DI(363) XOR DI(469) XOR DI(433) XOR DI(434) XOR DI(12) XOR DI(506) XOR DI(253) XOR DI(352) XOR DI(56) XOR DI(357) XOR DI(249) XOR DI(36) XOR DI(440) XOR DI(132) XOR DI(186) XOR DI(198) XOR DI(498) XOR DI(251) XOR DI(271) XOR DI(108) XOR DI(6) XOR DI(402) XOR DI(220) XOR DI(346) XOR DI(404) XOR DI(336) XOR DI(58) XOR DI(180) XOR DI(476) XOR DI(492) XOR DI(229) XOR DI(205) XOR DI(136) XOR DI(86) XOR DI(389) XOR DI(94) XOR DI(421) XOR DI(294) XOR DI(359) XOR DI(471) XOR DI(155) XOR DI(508) XOR DI(261) XOR DI(391) XOR DI(282) XOR DI(44) XOR DI(425) XOR DI(358) XOR DI(343) XOR DI(441) XOR DI(65) XOR DI(187) XOR DI(327) XOR DI(160) XOR DI(245) XOR DI(272) XOR DI(210) XOR DI(307) XOR DI(109) XOR DI(236) XOR DI(100) XOR DI(372) XOR DI(338) XOR DI(396) XOR DI(197) XOR DI(128) XOR DI(381) XOR DI(76) XOR DI(351) XOR DI(147) XOR DI(101) XOR DI(248) XOR DI(347) XOR DI(51) XOR DI(275) XOR DI(455) XOR DI(244) XOR DI(91) XOR DI(475) XOR DI(181) XOR DI(459) XOR DI(406) XOR DI(204) XOR DI(230) XOR DI(293) XOR DI(390) XOR DI(478) XOR DI(122) XOR DI(422) XOR DI(45) XOR DI(449) XOR DI(85) XOR DI(442) XOR DI(131) XOR DI(472) XOR DI(116) XOR DI(140) XOR DI(436) XOR DI(300) XOR DI(354) XOR DI(150) XOR DI(188) XOR DI(348) XOR DI(8) XOR DI(497) XOR DI(509) XOR DI(63) XOR DI(75) XOR DI(321) XOR DI(482) XOR DI(176) XOR DI(360) XOR DI(413) XOR DI(221) XOR DI(328) XOR DI(483) XOR DI(456) XOR DI(453) XOR DI(318) XOR DI(67) XOR DI(224) XOR DI(189) XOR DI(485) XOR DI(285) XOR DI(18) XOR DI(287) XOR DI(123) XOR DI(428) XOR DI(416) XOR DI(162) XOR DI(384) XOR DI(50) XOR DI(243) XOR DI(212) XOR DI(111) XOR DI(320) XOR DI(9) XOR DI(405) XOR DI(375) XOR DI(21) XOR DI(102) XOR DI(0) XOR DI(216) XOR DI(301) XOR DI(376) XOR DI(340) XOR DI(398) XOR DI(448) XOR DI(34) XOR DI(174) XOR DI(385) XOR DI(199) XOR DI(415) XOR DI(104) XOR DI(103) XOR DI(20) XOR DI(417) XOR DI(169) XOR DI(502) XOR DI(53) XOR DI(170) XOR DI(407) XOR DI(319) XOR DI(93) XOR DI(61) XOR DI(183) XOR DI(461) XOR DI(167) XOR DI(394) XOR DI(479) XOR DI(410) XOR DI(495) XOR DI(268) XOR DI(237) XOR DI(303) XOR DI(314) XOR DI(219) XOR DI(295) XOR DI(115) XOR DI(139) XOR DI(89) XOR DI(392) XOR DI(480) XOR DI(193) XOR DI(124) XOR DI(377) XOR DI(163) XOR DI(401) XOR DI(313) XOR DI(451) XOR DI(209) XOR DI(317) XOR DI(388) XOR DI(362) XOR DI(133) XOR DI(386) XOR DI(211) XOR DI(118) XOR DI(137) XOR DI(158) XOR DI(445) XOR DI(438) XOR DI(302) XOR DI(196) XOR DI(112) XOR DI(35) XOR DI(190) XOR DI(350) XOR DI(10) XOR DI(4) XOR DI(178) XOR DI(166) XOR DI(5) XOR DI(511);
   DO(22) <= DI(50) XOR DI(265) XOR DI(268) XOR DI(468) XOR DI(330) XOR DI(78) XOR DI(502) XOR DI(127) XOR DI(487) XOR DI(260) XOR DI(287) XOR DI(81) XOR DI(79) XOR DI(289) XOR DI(256) XOR DI(155) XOR DI(368) XOR DI(333) XOR DI(332) XOR DI(488) XOR DI(467) XOR DI(432) XOR DI(69) XOR DI(350) XOR DI(278) XOR DI(458) XOR DI(247) XOR DI(130) XOR DI(196) XOR DI(229) XOR DI(362) XOR DI(369) XOR DI(334) XOR DI(178) XOR DI(263) XOR DI(290) XOR DI(203) XOR DI(84) XOR DI(292) XOR DI(357) XOR DI(433) XOR DI(506) XOR DI(55) XOR DI(356) XOR DI(63) XOR DI(185) XOR DI(325) XOR DI(243) XOR DI(380) XOR DI(239) XOR DI(305) XOR DI(107) XOR DI(401) XOR DI(149) XOR DI(371) XOR DI(126) XOR DI(345) XOR DI(453) XOR DI(277) XOR DI(264) XOR DI(202) XOR DI(228) XOR DI(364) XOR DI(440) XOR DI(470) XOR DI(154) XOR DI(434) XOR DI(12) XOR DI(108) XOR DI(435) XOR DI(346) XOR DI(13) XOR DI(507) XOR DI(254) XOR DI(353) XOR DI(57) XOR DI(464) XOR DI(44) XOR DI(174) XOR DI(358) XOR DI(250) XOR DI(326) XOR DI(47) XOR DI(451) XOR DI(37) XOR DI(441) XOR DI(133) XOR DI(187) XOR DI(398) XOR DI(75) XOR DI(285) XOR DI(121) XOR DI(199) XOR DI(499) XOR DI(252) XOR DI(272) XOR DI(109) XOR DI(7) XOR DI(403) XOR DI(100) XOR DI(143) XOR DI(93) XOR DI(32) XOR DI(257) XOR DI(221) XOR DI(248) XOR DI(347) XOR DI(275) XOR DI(405) XOR DI(475) XOR DI(337) XOR DI(310) XOR DI(59) XOR DI(181) XOR DI(459) XOR DI(477) XOR DI(23) XOR DI(493) XOR DI(235) XOR DI(230) XOR DI(226) XOR DI(206) XOR DI(137) XOR DI(87) XOR DI(390) XOR DI(26) XOR DI(146) XOR DI(95) XOR DI(422) XOR DI(295) XOR DI(360) XOR DI(131) XOR DI(472) XOR DI(209) XOR DI(156) XOR DI(150) XOR DI(430) XOR DI(342) XOR DI(509) XOR DI(255) XOR DI(262) XOR DI(392) XOR DI(354) XOR DI(193) XOR DI(283) XOR DI(465) XOR DI(45) XOR DI(426) XOR DI(359) XOR DI(282) XOR DI(324) XOR DI(251) XOR DI(98) XOR DI(482) XOR DI(344) XOR DI(48) XOR DI(445) XOR DI(442) XOR DI(66) XOR DI(188) XOR DI(396) XOR DI(328) XOR DI(284) XOR DI(17) XOR DI(413) XOR DI(122) XOR DI(30) XOR DI(427) XOR DI(415) XOR DI(161) XOR DI(500) XOR DI(246) XOR DI(253) XOR DI(273) XOR DI(211) XOR DI(308) XOR DI(29) XOR DI(110) XOR DI(237) XOR DI(233) XOR DI(20) XOR DI(101) XOR DI(224) XOR DI(215) XOR DI(300) XOR DI(375) XOR DI(120) XOR DI(373) XOR DI(144) XOR DI(339) XOR DI(397) XOR DI(309) XOR DI(447) XOR DI(33) XOR DI(173) XOR DI(384) XOR DI(198) XOR DI(129) XOR DI(382) XOR DI(153) XOR DI(77) XOR DI(298) XOR DI(352) XOR DI(31) XOR DI(148) XOR DI(428) XOR DI(102) XOR DI(340) XOR DI(249) XOR DI(348) XOR DI(52) XOR DI(276) XOR DI(456) XOR DI(245) XOR DI(214) XOR DI(92) XOR DI(476) XOR DI(42) XOR DI(311) XOR DI(60) XOR DI(182) XOR DI(460) XOR DI(478) XOR DI(407) XOR DI(24) XOR DI(409) XOR DI(236) XOR DI(205) XOR DI(313) XOR DI(2) XOR DI(231) XOR DI(218) XOR DI(294) XOR DI(207) XOR DI(114) XOR DI(88) XOR DI(391) XOR DI(479) XOR DI(216) XOR DI(192) XOR DI(123) XOR DI(96) XOR DI(423) XOR DI(46) XOR DI(450) XOR DI(86) XOR DI(443) XOR DI(18) XOR DI(132) XOR DI(473) XOR DI(117) XOR DI(141) XOR DI(136) XOR DI(40) XOR DI(394) XOR DI(444) XOR DI(437) XOR DI(301) XOR DI(195) XOR DI(355) XOR DI(151) XOR DI(431) XOR DI(189) XOR DI(349) XOR DI(9) XOR DI(425) XOR DI(343) XOR DI(165) XOR DI(4) XOR DI(498) XOR DI(510);
   DO(23) <= DI(51) XOR DI(266) XOR DI(269) XOR DI(469) XOR DI(331) XOR DI(79) XOR DI(503) XOR DI(128) XOR DI(488) XOR DI(261) XOR DI(288) XOR DI(82) XOR DI(80) XOR DI(290) XOR DI(257) XOR DI(156) XOR DI(369) XOR DI(334) XOR DI(333) XOR DI(489) XOR DI(468) XOR DI(433) XOR DI(70) XOR DI(351) XOR DI(279) XOR DI(459) XOR DI(248) XOR DI(131) XOR DI(197) XOR DI(230) XOR DI(363) XOR DI(370) XOR DI(335) XOR DI(179) XOR DI(264) XOR DI(291) XOR DI(204) XOR DI(85) XOR DI(293) XOR DI(358) XOR DI(434) XOR DI(507) XOR DI(56) XOR DI(357) XOR DI(64) XOR DI(186) XOR DI(326) XOR DI(244) XOR DI(381) XOR DI(240) XOR DI(306) XOR DI(108) XOR DI(402) XOR DI(150) XOR DI(372) XOR DI(127) XOR DI(346) XOR DI(454) XOR DI(278) XOR DI(265) XOR DI(203) XOR DI(229) XOR DI(365) XOR DI(441) XOR DI(471) XOR DI(155) XOR DI(435) XOR DI(13) XOR DI(109) XOR DI(436) XOR DI(347) XOR DI(14) XOR DI(508) XOR DI(255) XOR DI(354) XOR DI(58) XOR DI(465) XOR DI(45) XOR DI(175) XOR DI(359) XOR DI(251) XOR DI(327) XOR DI(48) XOR DI(452) XOR DI(38) XOR DI(442) XOR DI(134) XOR DI(188) XOR DI(399) XOR DI(76) XOR DI(286) XOR DI(122) XOR DI(200) XOR DI(500) XOR DI(253) XOR DI(273) XOR DI(110) XOR DI(8) XOR DI(404) XOR DI(101) XOR DI(144) XOR DI(94) XOR DI(33) XOR DI(258) XOR DI(222) XOR DI(249) XOR DI(348) XOR DI(276) XOR DI(406) XOR DI(476) XOR DI(338) XOR DI(311) XOR DI(60) XOR DI(182) XOR DI(460) XOR DI(478) XOR DI(24) XOR DI(494) XOR DI(236) XOR DI(231) XOR DI(227) XOR DI(207) XOR DI(138) XOR DI(88) XOR DI(391) XOR DI(27) XOR DI(147) XOR DI(96) XOR DI(423) XOR DI(296) XOR DI(361) XOR DI(132) XOR DI(473) XOR DI(210) XOR DI(157) XOR DI(151) XOR DI(431) XOR DI(343) XOR DI(510) XOR DI(256) XOR DI(263) XOR DI(393) XOR DI(355) XOR DI(194) XOR DI(284) XOR DI(466) XOR DI(46) XOR DI(427) XOR DI(360) XOR DI(283) XOR DI(325) XOR DI(252) XOR DI(99) XOR DI(483) XOR DI(345) XOR DI(49) XOR DI(446) XOR DI(443) XOR DI(67) XOR DI(189) XOR DI(397) XOR DI(329) XOR DI(285) XOR DI(18) XOR DI(414) XOR DI(123) XOR DI(31) XOR DI(428) XOR DI(416) XOR DI(162) XOR DI(501) XOR DI(247) XOR DI(254) XOR DI(274) XOR DI(212) XOR DI(309) XOR DI(30) XOR DI(111) XOR DI(238) XOR DI(234) XOR DI(21) XOR DI(102) XOR DI(225) XOR DI(216) XOR DI(301) XOR DI(376) XOR DI(121) XOR DI(374) XOR DI(145) XOR DI(340) XOR DI(398) XOR DI(310) XOR DI(448) XOR DI(34) XOR DI(174) XOR DI(385) XOR DI(199) XOR DI(130) XOR DI(383) XOR DI(154) XOR DI(78) XOR DI(299) XOR DI(353) XOR DI(32) XOR DI(149) XOR DI(429) XOR DI(103) XOR DI(341) XOR DI(250) XOR DI(349) XOR DI(53) XOR DI(277) XOR DI(457) XOR DI(246) XOR DI(215) XOR DI(93) XOR DI(477) XOR DI(43) XOR DI(312) XOR DI(61) XOR DI(183) XOR DI(461) XOR DI(479) XOR DI(408) XOR DI(25) XOR DI(410) XOR DI(237) XOR DI(206) XOR DI(314) XOR DI(3) XOR DI(232) XOR DI(219) XOR DI(295) XOR DI(208) XOR DI(115) XOR DI(89) XOR DI(392) XOR DI(480) XOR DI(217) XOR DI(193) XOR DI(124) XOR DI(97) XOR DI(424) XOR DI(47) XOR DI(451) XOR DI(87) XOR DI(444) XOR DI(19) XOR DI(133) XOR DI(474) XOR DI(118) XOR DI(142) XOR DI(137) XOR DI(41) XOR DI(395) XOR DI(445) XOR DI(438) XOR DI(302) XOR DI(196) XOR DI(356) XOR DI(152) XOR DI(432) XOR DI(190) XOR DI(350) XOR DI(10) XOR DI(426) XOR DI(344) XOR DI(166) XOR DI(5) XOR DI(499) XOR DI(511);
   DO(24) <= DI(52) XOR DI(267) XOR DI(270) XOR DI(470) XOR DI(332) XOR DI(488) XOR DI(288) XOR DI(80) XOR DI(126) XOR DI(431) XOR DI(504) XOR DI(129) XOR DI(489) XOR DI(262) XOR DI(289) XOR DI(83) XOR DI(418) XOR DI(81) XOR DI(291) XOR DI(468) XOR DI(258) XOR DI(324) XOR DI(157) XOR DI(269) XOR DI(370) XOR DI(369) XOR DI(335) XOR DI(378) XOR DI(144) XOR DI(334) XOR DI(114) XOR DI(490) XOR DI(363) XOR DI(387) XOR DI(469) XOR DI(434) XOR DI(185) XOR DI(24) XOR DI(179) XOR DI(12) XOR DI(506) XOR DI(71) XOR DI(260) XOR DI(352) XOR DI(280) XOR DI(322) XOR DI(460) XOR DI(249) XOR DI(96) XOR DI(36) XOR DI(440) XOR DI(64) XOR DI(132) XOR DI(198) XOR DI(159) XOR DI(108) XOR DI(402) XOR DI(231) XOR DI(364) XOR DI(298) XOR DI(371) XOR DI(380) XOR DI(336) XOR DI(40) XOR DI(180) XOR DI(265) XOR DI(203) XOR DI(229) XOR DI(292) XOR DI(205) XOR DI(136) XOR DI(86) XOR DI(389) XOR DI(294) XOR DI(305) XOR DI(359) XOR DI(435) XOR DI(496) XOR DI(508) XOR DI(282) XOR DI(57) XOR DI(358) XOR DI(60) XOR DI(343) XOR DI(454) XOR DI(65) XOR DI(222) XOR DI(187) XOR DI(465) XOR DI(327) XOR DI(171) XOR DI(245) XOR DI(382) XOR DI(241) XOR DI(210) XOR DI(307) XOR DI(109) XOR DI(403) XOR DI(151) XOR DI(236) XOR DI(373) XOR DI(128) XOR DI(76) XOR DI(347) XOR DI(51) XOR DI(168) XOR DI(455) XOR DI(244) XOR DI(459) XOR DI(165) XOR DI(406) XOR DI(279) XOR DI(266) XOR DI(204) XOR DI(230) XOR DI(366) XOR DI(442) XOR DI(472) XOR DI(140) XOR DI(156) XOR DI(436) XOR DI(105) XOR DI(14) XOR DI(110) XOR DI(437) XOR DI(348) XOR DI(2) XOR DI(15) XOR DI(503) XOR DI(509) XOR DI(63) XOR DI(487) XOR DI(256) XOR DI(355) XOR DI(75) XOR DI(321) XOR DI(482) XOR DI(59) XOR DI(466) XOR DI(46) XOR DI(176) XOR DI(360) XOR DI(413) XOR DI(252) XOR DI(328) XOR DI(483) XOR DI(49) XOR DI(453) XOR DI(318) XOR DI(39) XOR DI(443) XOR DI(224) XOR DI(135) XOR DI(189) XOR DI(120) XOR DI(329) XOR DI(173) XOR DI(400) XOR DI(18) XOR DI(414) XOR DI(77) XOR DI(287) XOR DI(123) XOR DI(464) XOR DI(201) XOR DI(416) XOR DI(501) XOR DI(254) XOR DI(274) XOR DI(243) XOR DI(212) XOR DI(309) XOR DI(30) XOR DI(111) XOR DI(320) XOR DI(9) XOR DI(405) XOR DI(192) XOR DI(21) XOR DI(102) XOR DI(0) XOR DI(225) XOR DI(376) XOR DI(214) XOR DI(121) XOR DI(145) XOR DI(95) XOR DI(340) XOR DI(34) XOR DI(174) XOR DI(385) XOR DI(486) XOR DI(259) XOR DI(223) XOR DI(154) XOR DI(78) XOR DI(149) XOR DI(1) XOR DI(250) XOR DI(349) XOR DI(170) XOR DI(277) XOR DI(407) XOR DI(319) XOR DI(457) XOR DI(215) XOR DI(93) XOR DI(477) XOR DI(339) XOR DI(312) XOR DI(61) XOR DI(183) XOR DI(461) XOR DI(479) XOR DI(408) XOR DI(25) XOR DI(495) XOR DI(237) XOR DI(314) XOR DI(232) XOR DI(228) XOR DI(208) XOR DI(368) XOR DI(139) XOR DI(89) XOR DI(392) XOR DI(304) XOR DI(28) XOR DI(193) XOR DI(148) XOR DI(97) XOR DI(424) XOR DI(164) XOR DI(401) XOR DI(451) XOR DI(113) XOR DI(177) XOR DI(297) XOR DI(202) XOR DI(362) XOR DI(133) XOR DI(474) XOR DI(211) XOR DI(158) XOR DI(395) XOR DI(107) XOR DI(152) XOR DI(432) XOR DI(10) XOR DI(29) XOR DI(344) XOR DI(23) XOR DI(178) XOR DI(17) XOR DI(5) XOR DI(511);
   DO(25) <= DI(68) XOR DI(53) XOR DI(268) XOR DI(368) XOR DI(271) XOR DI(471) XOR DI(333) XOR DI(489) XOR DI(289) XOR DI(418) XOR DI(81) XOR DI(127) XOR DI(468) XOR DI(432) XOR DI(505) XOR DI(54) XOR DI(247) XOR DI(130) XOR DI(269) XOR DI(125) XOR DI(490) XOR DI(263) XOR DI(290) XOR DI(84) XOR DI(419) XOR DI(82) XOR DI(292) XOR DI(357) XOR DI(469) XOR DI(36) XOR DI(506) XOR DI(259) XOR DI(389) XOR DI(314) XOR DI(439) XOR DI(63) XOR DI(185) XOR DI(325) XOR DI(158) XOR DI(243) XOR DI(380) XOR DI(270) XOR DI(239) XOR DI(107) XOR DI(5) XOR DI(371) XOR DI(370) XOR DI(336) XOR DI(126) XOR DI(379) XOR DI(145) XOR DI(335) XOR DI(115) XOR DI(491) XOR DI(264) XOR DI(364) XOR DI(388) XOR DI(440) XOR DI(304) XOR DI(470) XOR DI(154) XOR DI(12) XOR DI(435) XOR DI(186) XOR DI(346) XOR DI(25) XOR DI(180) XOR DI(13) XOR DI(507) XOR DI(72) XOR DI(261) XOR DI(353) XOR DI(464) XOR DI(44) XOR DI(281) XOR DI(323) XOR DI(461) XOR DI(250) XOR DI(97) XOR DI(326) XOR DI(451) XOR DI(37) XOR DI(441) XOR DI(65) XOR DI(133) XOR DI(395) XOR DI(398) XOR DI(75) XOR DI(285) XOR DI(199) XOR DI(160) XOR DI(109) XOR DI(403) XOR DI(232) XOR DI(100) XOR DI(365) XOR DI(299) XOR DI(372) XOR DI(143) XOR DI(93) XOR DI(446) XOR DI(32) XOR DI(197) XOR DI(381) XOR DI(351) XOR DI(167) XOR DI(248) XOR DI(51) XOR DI(337) XOR DI(41) XOR DI(181) XOR DI(459) XOR DI(23) XOR DI(266) XOR DI(235) XOR DI(204) XOR DI(230) XOR DI(217) XOR DI(293) XOR DI(206) XOR DI(113) XOR DI(137) XOR DI(87) XOR DI(390) XOR DI(295) XOR DI(306) XOR DI(360) XOR DI(131) XOR DI(116) XOR DI(436) XOR DI(430) XOR DI(104) XOR DI(342) XOR DI(170) XOR DI(164) XOR DI(497) XOR DI(503) XOR DI(509) XOR DI(486) XOR DI(354) XOR DI(481) XOR DI(283) XOR DI(58) XOR DI(411) XOR DI(359) XOR DI(61) XOR DI(282) XOR DI(324) XOR DI(220) XOR DI(482) XOR DI(344) XOR DI(48) XOR DI(455) XOR DI(445) XOR DI(66) XOR DI(223) XOR DI(188) XOR DI(119) XOR DI(466) XOR DI(328) XOR DI(172) XOR DI(399) XOR DI(284) XOR DI(17) XOR DI(413) XOR DI(286) XOR DI(200) XOR DI(427) XOR DI(500) XOR DI(246) XOR DI(383) XOR DI(242) XOR DI(211) XOR DI(308) XOR DI(110) XOR DI(404) XOR DI(191) XOR DI(152) XOR DI(237) XOR DI(374) XOR DI(20) XOR DI(300) XOR DI(375) XOR DI(120) XOR DI(144) XOR DI(309) XOR DI(447) XOR DI(33) XOR DI(173) XOR DI(384) XOR DI(222) XOR DI(129) XOR DI(77) XOR DI(428) XOR DI(429) XOR DI(0) XOR DI(416) XOR DI(168) XOR DI(348) XOR DI(52) XOR DI(169) XOR DI(318) XOR DI(456) XOR DI(245) XOR DI(214) XOR DI(42) XOR DI(449) XOR DI(311) XOR DI(460) XOR DI(166) XOR DI(407) XOR DI(280) XOR DI(457) XOR DI(267) XOR DI(236) XOR DI(205) XOR DI(302) XOR DI(231) XOR DI(218) XOR DI(207) XOR DI(367) XOR DI(138) XOR DI(88) XOR DI(303) XOR DI(378) XOR DI(192) XOR DI(376) XOR DI(163) XOR DI(443) XOR DI(387) XOR DI(296) XOR DI(385) XOR DI(21) XOR DI(473) XOR DI(210) XOR DI(141) XOR DI(157) XOR DI(394) XOR DI(437) XOR DI(106) XOR DI(195) XOR DI(15) XOR DI(111) XOR DI(438) XOR DI(431) XOR DI(349) XOR DI(105) XOR DI(343) XOR DI(3) XOR DI(16) XOR DI(4) XOR DI(504) XOR DI(510);
   DO(26) <= DI(69) XOR DI(54) XOR DI(269) XOR DI(369) XOR DI(272) XOR DI(472) XOR DI(334) XOR DI(490) XOR DI(290) XOR DI(419) XOR DI(82) XOR DI(128) XOR DI(469) XOR DI(433) XOR DI(506) XOR DI(55) XOR DI(248) XOR DI(131) XOR DI(270) XOR DI(126) XOR DI(491) XOR DI(264) XOR DI(291) XOR DI(85) XOR DI(420) XOR DI(83) XOR DI(293) XOR DI(358) XOR DI(470) XOR DI(37) XOR DI(507) XOR DI(260) XOR DI(390) XOR DI(315) XOR DI(440) XOR DI(64) XOR DI(186) XOR DI(326) XOR DI(159) XOR DI(244) XOR DI(381) XOR DI(271) XOR DI(240) XOR DI(108) XOR DI(6) XOR DI(372) XOR DI(371) XOR DI(337) XOR DI(127) XOR DI(380) XOR DI(146) XOR DI(336) XOR DI(116) XOR DI(492) XOR DI(265) XOR DI(365) XOR DI(389) XOR DI(441) XOR DI(305) XOR DI(471) XOR DI(155) XOR DI(13) XOR DI(436) XOR DI(187) XOR DI(347) XOR DI(26) XOR DI(181) XOR DI(14) XOR DI(508) XOR DI(73) XOR DI(262) XOR DI(354) XOR DI(465) XOR DI(45) XOR DI(282) XOR DI(324) XOR DI(462) XOR DI(251) XOR DI(98) XOR DI(327) XOR DI(452) XOR DI(38) XOR DI(442) XOR DI(66) XOR DI(134) XOR DI(396) XOR DI(399) XOR DI(76) XOR DI(286) XOR DI(200) XOR DI(161) XOR DI(110) XOR DI(404) XOR DI(233) XOR DI(101) XOR DI(366) XOR DI(300) XOR DI(373) XOR DI(144) XOR DI(94) XOR DI(447) XOR DI(33) XOR DI(198) XOR DI(382) XOR DI(352) XOR DI(168) XOR DI(249) XOR DI(52) XOR DI(338) XOR DI(42) XOR DI(182) XOR DI(460) XOR DI(24) XOR DI(267) XOR DI(236) XOR DI(205) XOR DI(231) XOR DI(218) XOR DI(294) XOR DI(207) XOR DI(114) XOR DI(138) XOR DI(88) XOR DI(391) XOR DI(296) XOR DI(307) XOR DI(361) XOR DI(132) XOR DI(117) XOR DI(437) XOR DI(431) XOR DI(105) XOR DI(343) XOR DI(171) XOR DI(165) XOR DI(498) XOR DI(504) XOR DI(510) XOR DI(487) XOR DI(355) XOR DI(482) XOR DI(284) XOR DI(59) XOR DI(412) XOR DI(360) XOR DI(62) XOR DI(283) XOR DI(325) XOR DI(221) XOR DI(483) XOR DI(345) XOR DI(49) XOR DI(456) XOR DI(446) XOR DI(67) XOR DI(224) XOR DI(189) XOR DI(120) XOR DI(467) XOR DI(329) XOR DI(173) XOR DI(400) XOR DI(285) XOR DI(18) XOR DI(414) XOR DI(287) XOR DI(201) XOR DI(428) XOR DI(501) XOR DI(247) XOR DI(384) XOR DI(243) XOR DI(212) XOR DI(309) XOR DI(111) XOR DI(405) XOR DI(192) XOR DI(153) XOR DI(238) XOR DI(375) XOR DI(21) XOR DI(0) XOR DI(301) XOR DI(376) XOR DI(121) XOR DI(145) XOR DI(310) XOR DI(448) XOR DI(34) XOR DI(174) XOR DI(385) XOR DI(223) XOR DI(130) XOR DI(78) XOR DI(429) XOR DI(430) XOR DI(1) XOR DI(417) XOR DI(169) XOR DI(349) XOR DI(53) XOR DI(170) XOR DI(319) XOR DI(457) XOR DI(246) XOR DI(215) XOR DI(43) XOR DI(450) XOR DI(312) XOR DI(461) XOR DI(167) XOR DI(408) XOR DI(281) XOR DI(458) XOR DI(268) XOR DI(237) XOR DI(206) XOR DI(303) XOR DI(232) XOR DI(219) XOR DI(208) XOR DI(368) XOR DI(139) XOR DI(89) XOR DI(304) XOR DI(379) XOR DI(193) XOR DI(377) XOR DI(164) XOR DI(444) XOR DI(388) XOR DI(297) XOR DI(386) XOR DI(22) XOR DI(474) XOR DI(211) XOR DI(142) XOR DI(158) XOR DI(395) XOR DI(438) XOR DI(107) XOR DI(196) XOR DI(16) XOR DI(112) XOR DI(439) XOR DI(432) XOR DI(350) XOR DI(106) XOR DI(344) XOR DI(4) XOR DI(17) XOR DI(5) XOR DI(505) XOR DI(511);
   DO(27) <= DI(70) XOR DI(55) XOR DI(42) XOR DI(324) XOR DI(452) XOR DI(88) XOR DI(185) XOR DI(270) XOR DI(98) XOR DI(363) XOR DI(370) XOR DI(255) XOR DI(195) XOR DI(126) XOR DI(273) XOR DI(473) XOR DI(335) XOR DI(179) XOR DI(491) XOR DI(264) XOR DI(291) XOR DI(24) XOR DI(144) XOR DI(420) XOR DI(83) XOR DI(129) XOR DI(470) XOR DI(114) XOR DI(138) XOR DI(434) XOR DI(12) XOR DI(507) XOR DI(253) XOR DI(260) XOR DI(56) XOR DI(357) XOR DI(322) XOR DI(249) XOR DI(218) XOR DI(96) XOR DI(36) XOR DI(64) XOR DI(132) XOR DI(251) XOR DI(271) XOR DI(402) XOR DI(127) XOR DI(296) XOR DI(40) XOR DI(278) XOR DI(492) XOR DI(265) XOR DI(203) XOR DI(229) XOR DI(292) XOR DI(136) XOR DI(86) XOR DI(94) XOR DI(421) XOR DI(84) XOR DI(294) XOR DI(359) XOR DI(471) XOR DI(134) XOR DI(38) XOR DI(155) XOR DI(496) XOR DI(508) XOR DI(261) XOR DI(391) XOR DI(425) XOR DI(411) XOR DI(343) XOR DI(454) XOR DI(316) XOR DI(441) XOR DI(65) XOR DI(187) XOR DI(465) XOR DI(327) XOR DI(160) XOR DI(245) XOR DI(382) XOR DI(48) XOR DI(272) XOR DI(241) XOR DI(210) XOR DI(109) XOR DI(7) XOR DI(236) XOR DI(373) XOR DI(100) XOR DI(372) XOR DI(338) XOR DI(257) XOR DI(128) XOR DI(381) XOR DI(76) XOR DI(147) XOR DI(500) XOR DI(51) XOR DI(275) XOR DI(337) XOR DI(117) XOR DI(493) XOR DI(266) XOR DI(226) XOR DI(366) XOR DI(390) XOR DI(26) XOR DI(478) XOR DI(399) XOR DI(442) XOR DI(315) XOR DI(306) XOR DI(200) XOR DI(472) XOR DI(116) XOR DI(156) XOR DI(105) XOR DI(300) XOR DI(354) XOR DI(14) XOR DI(33) XOR DI(150) XOR DI(437) XOR DI(188) XOR DI(348) XOR DI(27) XOR DI(182) XOR DI(15) XOR DI(503) XOR DI(509) XOR DI(487) XOR DI(235) XOR DI(74) XOR DI(263) XOR DI(393) XOR DI(355) XOR DI(75) XOR DI(321) XOR DI(482) XOR DI(342) XOR DI(466) XOR DI(46) XOR DI(427) XOR DI(62) XOR DI(283) XOR DI(325) XOR DI(463) XOR DI(252) XOR DI(99) XOR DI(328) XOR DI(453) XOR DI(318) XOR DI(39) XOR DI(446) XOR DI(443) XOR DI(125) XOR DI(67) XOR DI(191) XOR DI(135) XOR DI(120) XOR DI(397) XOR DI(467) XOR DI(329) XOR DI(173) XOR DI(400) XOR DI(414) XOR DI(77) XOR DI(287) XOR DI(464) XOR DI(201) XOR DI(31) XOR DI(428) XOR DI(416) XOR DI(162) XOR DI(384) XOR DI(243) XOR DI(309) XOR DI(30) XOR DI(111) XOR DI(405) XOR DI(192) XOR DI(153) XOR DI(375) XOR DI(234) XOR DI(21) XOR DI(102) XOR DI(0) XOR DI(367) XOR DI(301) XOR DI(214) XOR DI(374) XOR DI(145) XOR DI(95) XOR DI(340) XOR DI(398) XOR DI(448) XOR DI(34) XOR DI(486) XOR DI(199) XOR DI(383) XOR DI(78) XOR DI(104) XOR DI(353) XOR DI(32) XOR DI(149) XOR DI(103) XOR DI(341) XOR DI(20) XOR DI(417) XOR DI(169) XOR DI(481) XOR DI(250) XOR DI(53) XOR DI(319) XOR DI(215) XOR DI(93) XOR DI(339) XOR DI(43) XOR DI(119) XOR DI(183) XOR DI(461) XOR DI(167) XOR DI(394) XOR DI(408) XOR DI(25) XOR DI(268) XOR DI(237) XOR DI(206) XOR DI(303) XOR DI(314) XOR DI(232) XOR DI(219) XOR DI(295) XOR DI(208) XOR DI(115) XOR DI(368) XOR DI(139) XOR DI(89) XOR DI(392) XOR DI(480) XOR DI(217) XOR DI(124) XOR DI(163) XOR DI(47) XOR DI(164) XOR DI(444) XOR DI(177) XOR DI(297) XOR DI(308) XOR DI(362) XOR DI(133) XOR DI(118) XOR DI(395) XOR DI(438) XOR DI(432) XOR DI(10) XOR DI(106) XOR DI(29) XOR DI(184) XOR DI(344) XOR DI(4) XOR DI(178) XOR DI(172) XOR DI(11) XOR DI(166) XOR DI(499) XOR DI(505) XOR DI(511);
   DO(28) <= DI(71) XOR DI(260) XOR DI(56) XOR DI(43) XOR DI(357) XOR DI(325) XOR DI(453) XOR DI(239) XOR DI(36) XOR DI(440) XOR DI(64) XOR DI(89) XOR DI(186) XOR DI(159) XOR DI(271) XOR DI(108) XOR DI(6) XOR DI(402) XOR DI(99) XOR DI(364) XOR DI(371) XOR DI(256) XOR DI(196) XOR DI(127) XOR DI(380) XOR DI(350) XOR DI(247) XOR DI(346) XOR DI(50) XOR DI(274) XOR DI(243) XOR DI(474) XOR DI(336) XOR DI(180) XOR DI(458) XOR DI(278) XOR DI(492) XOR DI(265) XOR DI(203) XOR DI(229) XOR DI(225) XOR DI(292) XOR DI(389) XOR DI(25) XOR DI(145) XOR DI(421) XOR DI(84) XOR DI(314) XOR DI(305) XOR DI(130) XOR DI(471) XOR DI(115) XOR DI(139) XOR DI(155) XOR DI(435) XOR DI(13) XOR DI(149) XOR DI(496) XOR DI(502) XOR DI(508) XOR DI(254) XOR DI(261) XOR DI(57) XOR DI(358) XOR DI(323) XOR DI(250) XOR DI(219) XOR DI(97) XOR DI(451) XOR DI(37) XOR DI(65) XOR DI(133) XOR DI(285) XOR DI(252) XOR DI(272) XOR DI(403) XOR DI(143) XOR DI(93) XOR DI(446) XOR DI(257) XOR DI(197) XOR DI(128) XOR DI(297) XOR DI(351) XOR DI(248) XOR DI(51) XOR DI(275) XOR DI(475) XOR DI(41) XOR DI(459) XOR DI(321) XOR DI(279) XOR DI(23) XOR DI(408) XOR DI(493) XOR DI(266) XOR DI(204) XOR DI(230) XOR DI(226) XOR DI(217) XOR DI(293) XOR DI(113) XOR DI(137) XOR DI(87) XOR DI(377) XOR DI(95) XOR DI(422) XOR DI(85) XOR DI(386) XOR DI(295) XOR DI(360) XOR DI(131) XOR DI(472) XOR DI(135) XOR DI(39) XOR DI(156) XOR DI(194) XOR DI(430) XOR DI(497) XOR DI(503) XOR DI(509) XOR DI(62) XOR DI(486) XOR DI(255) XOR DI(262) XOR DI(392) XOR DI(426) XOR DI(411) XOR DI(175) XOR DI(282) XOR DI(412) XOR DI(324) XOR DI(98) XOR DI(344) XOR DI(455) XOR DI(452) XOR DI(317) XOR DI(442) XOR DI(124) XOR DI(66) XOR DI(190) XOR DI(188) XOR DI(466) XOR DI(328) XOR DI(484) XOR DI(17) XOR DI(413) XOR DI(286) XOR DI(122) XOR DI(427) XOR DI(161) XOR DI(246) XOR DI(383) XOR DI(49) XOR DI(273) XOR DI(242) XOR DI(211) XOR DI(29) XOR DI(110) XOR DI(8) XOR DI(191) XOR DI(237) XOR DI(374) XOR DI(20) XOR DI(101) XOR DI(224) XOR DI(300) XOR DI(213) XOR DI(373) XOR DI(144) XOR DI(339) XOR DI(258) XOR DI(222) XOR DI(129) XOR DI(382) XOR DI(414) XOR DI(153) XOR DI(77) XOR DI(148) XOR DI(19) XOR DI(416) XOR DI(501) XOR DI(480) XOR DI(52) XOR DI(276) XOR DI(318) XOR DI(214) XOR DI(338) XOR DI(42) XOR DI(311) XOR DI(118) XOR DI(60) XOR DI(478) XOR DI(457) XOR DI(24) XOR DI(494) XOR DI(267) XOR DI(313) XOR DI(2) XOR DI(227) XOR DI(114) XOR DI(367) XOR DI(138) XOR DI(88) XOR DI(391) XOR DI(303) XOR DI(27) XOR DI(378) XOR DI(479) XOR DI(400) XOR DI(443) XOR DI(316) XOR DI(387) XOR DI(18) XOR DI(307) XOR DI(212) XOR DI(201) XOR DI(361) XOR DI(473) XOR DI(210) XOR DI(117) XOR DI(157) XOR DI(106) XOR DI(301) XOR DI(195) XOR DI(355) XOR DI(15) XOR DI(34) XOR DI(151) XOR DI(438) XOR DI(431) XOR DI(189) XOR DI(349) XOR DI(28) XOR DI(425) XOR DI(183) XOR DI(177) XOR DI(16) XOR DI(171) XOR DI(10) XOR DI(4) XOR DI(504) XOR DI(510);
   DO(29) <= DI(72) XOR DI(261) XOR DI(57) XOR DI(44) XOR DI(358) XOR DI(326) XOR DI(454) XOR DI(240) XOR DI(37) XOR DI(441) XOR DI(65) XOR DI(90) XOR DI(187) XOR DI(160) XOR DI(272) XOR DI(109) XOR DI(7) XOR DI(403) XOR DI(100) XOR DI(365) XOR DI(372) XOR DI(257) XOR DI(197) XOR DI(128) XOR DI(381) XOR DI(351) XOR DI(248) XOR DI(347) XOR DI(51) XOR DI(275) XOR DI(244) XOR DI(475) XOR DI(337) XOR DI(181) XOR DI(459) XOR DI(279) XOR DI(493) XOR DI(266) XOR DI(204) XOR DI(230) XOR DI(226) XOR DI(293) XOR DI(390) XOR DI(26) XOR DI(146) XOR DI(422) XOR DI(85) XOR DI(315) XOR DI(306) XOR DI(131) XOR DI(472) XOR DI(116) XOR DI(140) XOR DI(156) XOR DI(436) XOR DI(14) XOR DI(150) XOR DI(497) XOR DI(503) XOR DI(509) XOR DI(255) XOR DI(262) XOR DI(58) XOR DI(359) XOR DI(324) XOR DI(251) XOR DI(220) XOR DI(98) XOR DI(452) XOR DI(38) XOR DI(66) XOR DI(134) XOR DI(286) XOR DI(253) XOR DI(273) XOR DI(404) XOR DI(144) XOR DI(94) XOR DI(447) XOR DI(258) XOR DI(198) XOR DI(129) XOR DI(298) XOR DI(352) XOR DI(249) XOR DI(52) XOR DI(276) XOR DI(476) XOR DI(42) XOR DI(460) XOR DI(322) XOR DI(280) XOR DI(24) XOR DI(409) XOR DI(494) XOR DI(267) XOR DI(205) XOR DI(231) XOR DI(227) XOR DI(218) XOR DI(294) XOR DI(114) XOR DI(138) XOR DI(88) XOR DI(378) XOR DI(96) XOR DI(423) XOR DI(86) XOR DI(387) XOR DI(296) XOR DI(361) XOR DI(132) XOR DI(473) XOR DI(136) XOR DI(40) XOR DI(157) XOR DI(195) XOR DI(431) XOR DI(498) XOR DI(504) XOR DI(510) XOR DI(63) XOR DI(487) XOR DI(256) XOR DI(263) XOR DI(393) XOR DI(427) XOR DI(412) XOR DI(176) XOR DI(283) XOR DI(413) XOR DI(325) XOR DI(99) XOR DI(345) XOR DI(456) XOR DI(453) XOR DI(318) XOR DI(443) XOR DI(125) XOR DI(67) XOR DI(191) XOR DI(189) XOR DI(467) XOR DI(329) XOR DI(485) XOR DI(18) XOR DI(414) XOR DI(287) XOR DI(123) XOR DI(428) XOR DI(162) XOR DI(247) XOR DI(384) XOR DI(50) XOR DI(274) XOR DI(243) XOR DI(212) XOR DI(30) XOR DI(111) XOR DI(9) XOR DI(192) XOR DI(238) XOR DI(375) XOR DI(21) XOR DI(102) XOR DI(225) XOR DI(301) XOR DI(214) XOR DI(374) XOR DI(145) XOR DI(340) XOR DI(259) XOR DI(223) XOR DI(130) XOR DI(383) XOR DI(415) XOR DI(154) XOR DI(78) XOR DI(149) XOR DI(20) XOR DI(417) XOR DI(502) XOR DI(481) XOR DI(53) XOR DI(277) XOR DI(319) XOR DI(215) XOR DI(339) XOR DI(43) XOR DI(312) XOR DI(119) XOR DI(61) XOR DI(479) XOR DI(458) XOR DI(25) XOR DI(495) XOR DI(268) XOR DI(314) XOR DI(3) XOR DI(228) XOR DI(115) XOR DI(368) XOR DI(139) XOR DI(89) XOR DI(392) XOR DI(304) XOR DI(28) XOR DI(379) XOR DI(480) XOR DI(401) XOR DI(444) XOR DI(317) XOR DI(388) XOR DI(19) XOR DI(308) XOR DI(213) XOR DI(202) XOR DI(362) XOR DI(474) XOR DI(211) XOR DI(118) XOR DI(158) XOR DI(107) XOR DI(302) XOR DI(196) XOR DI(356) XOR DI(16) XOR DI(35) XOR DI(152) XOR DI(439) XOR DI(432) XOR DI(190) XOR DI(350) XOR DI(29) XOR DI(426) XOR DI(184) XOR DI(178) XOR DI(17) XOR DI(172) XOR DI(11) XOR DI(5) XOR DI(505) XOR DI(511);
   DO(30) <= DI(73) XOR DI(255) XOR DI(262) XOR DI(354) XOR DI(58) XOR DI(465) XOR DI(45) XOR DI(411) XOR DI(175) XOR DI(359) XOR DI(282) XOR DI(324) XOR DI(462) XOR DI(251) XOR DI(220) XOR DI(98) XOR DI(327) XOR DI(48) XOR DI(455) XOR DI(452) XOR DI(241) XOR DI(38) XOR DI(442) XOR DI(66) XOR DI(91) XOR DI(134) XOR DI(188) XOR DI(396) XOR DI(399) XOR DI(484) XOR DI(76) XOR DI(286) XOR DI(122) XOR DI(200) XOR DI(161) XOR DI(500) XOR DI(253) XOR DI(273) XOR DI(110) XOR DI(8) XOR DI(404) XOR DI(233) XOR DI(101) XOR DI(366) XOR DI(300) XOR DI(373) XOR DI(144) XOR DI(94) XOR DI(447) XOR DI(33) XOR DI(258) XOR DI(222) XOR DI(198) XOR DI(129) XOR DI(382) XOR DI(298) XOR DI(352) XOR DI(168) XOR DI(249) XOR DI(348) XOR DI(52) XOR DI(276) XOR DI(406) XOR DI(245) XOR DI(476) XOR DI(338) XOR DI(42) XOR DI(449) XOR DI(311) XOR DI(60) XOR DI(182) XOR DI(460) XOR DI(322) XOR DI(478) XOR DI(280) XOR DI(24) XOR DI(409) XOR DI(494) XOR DI(267) XOR DI(236) XOR DI(205) XOR DI(2) XOR DI(231) XOR DI(227) XOR DI(218) XOR DI(294) XOR DI(207) XOR DI(114) XOR DI(138) XOR DI(88) XOR DI(391) XOR DI(27) XOR DI(378) XOR DI(147) XOR DI(96) XOR DI(423) XOR DI(86) XOR DI(316) XOR DI(387) XOR DI(296) XOR DI(307) XOR DI(361) XOR DI(132) XOR DI(473) XOR DI(210) XOR DI(117) XOR DI(141) XOR DI(136) XOR DI(40) XOR DI(157) XOR DI(437) XOR DI(195) XOR DI(15) XOR DI(151) XOR DI(431) XOR DI(105) XOR DI(425) XOR DI(343) XOR DI(171) XOR DI(165) XOR DI(498) XOR DI(504) XOR DI(510) XOR DI(63) XOR DI(487) XOR DI(235) XOR DI(256) XOR DI(263) XOR DI(194) XOR DI(75) XOR DI(321) XOR DI(342) XOR DI(59) XOR DI(360) XOR DI(325) XOR DI(252) XOR DI(221) XOR DI(99) XOR DI(483) XOR DI(345) XOR DI(453) XOR DI(39) XOR DI(446) XOR DI(125) XOR DI(67) XOR DI(135) XOR DI(467) XOR DI(329) XOR DI(285) XOR DI(287) XOR DI(464) XOR DI(247) XOR DI(254) XOR DI(50) XOR DI(274) XOR DI(243) XOR DI(405) XOR DI(238) XOR DI(225) XOR DI(121) XOR DI(145) XOR DI(95) XOR DI(398) XOR DI(310) XOR DI(448) XOR DI(174) XOR DI(259) XOR DI(199) XOR DI(130) XOR DI(154) XOR DI(78) XOR DI(104) XOR DI(299) XOR DI(353) XOR DI(32) XOR DI(149) XOR DI(430) XOR DI(1) XOR DI(417) XOR DI(502) XOR DI(250) XOR DI(53) XOR DI(170) XOR DI(277) XOR DI(93) XOR DI(477) XOR DI(43) XOR DI(461) XOR DI(323) XOR DI(167) XOR DI(408) XOR DI(281) XOR DI(458) XOR DI(25) XOR DI(410) XOR DI(495) XOR DI(268) XOR DI(206) XOR DI(314) XOR DI(232) XOR DI(228) XOR DI(219) XOR DI(295) XOR DI(115) XOR DI(368) XOR DI(139) XOR DI(89) XOR DI(304) XOR DI(379) XOR DI(217) XOR DI(377) XOR DI(143) XOR DI(97) XOR DI(424) XOR DI(47) XOR DI(164) XOR DI(401) XOR DI(451) XOR DI(209) XOR DI(87) XOR DI(113) XOR DI(388) XOR DI(297) XOR DI(202) XOR DI(362) XOR DI(133) XOR DI(386) XOR DI(474) XOR DI(137) XOR DI(41) XOR DI(158) XOR DI(395) XOR DI(107) XOR DI(196) XOR DI(356) XOR DI(35) XOR DI(439) XOR DI(432) XOR DI(350) XOR DI(184) XOR DI(23) XOR DI(178) XOR DI(11) XOR DI(5) XOR DI(499) XOR DI(505) XOR DI(511);
   DO(31) <= DI(63) XOR DI(487) XOR DI(235) XOR DI(74) XOR DI(256) XOR DI(263) XOR DI(393) XOR DI(355) XOR DI(194) XOR DI(75) XOR DI(321) XOR DI(482) XOR DI(284) XOR DI(342) XOR DI(59) XOR DI(466) XOR DI(46) XOR DI(427) XOR DI(412) XOR DI(176) XOR DI(360) XOR DI(62) XOR DI(283) XOR DI(413) XOR DI(325) XOR DI(463) XOR DI(252) XOR DI(221) XOR DI(99) XOR DI(328) XOR DI(483) XOR DI(345) XOR DI(49) XOR DI(456) XOR DI(453) XOR DI(242) XOR DI(318) XOR DI(39) XOR DI(446) XOR DI(443) XOR DI(125) XOR DI(67) XOR DI(191) XOR DI(224) XOR DI(92) XOR DI(135) XOR DI(189) XOR DI(120) XOR DI(397) XOR DI(467) XOR DI(329) XOR DI(173) XOR DI(400) XOR DI(485) XOR DI(285) XOR DI(18) XOR DI(414) XOR DI(77) XOR DI(287) XOR DI(123) XOR DI(464) XOR DI(201) XOR DI(31) XOR DI(428) XOR DI(416) XOR DI(162) XOR DI(501) XOR DI(247) XOR DI(254) XOR DI(384) XOR DI(50) XOR DI(274) XOR DI(243) XOR DI(212) XOR DI(309) XOR DI(30) XOR DI(111) XOR DI(320) XOR DI(9) XOR DI(405) XOR DI(192) XOR DI(153) XOR DI(238) XOR DI(375) XOR DI(234) XOR DI(21) XOR DI(102) XOR DI(0) XOR DI(225) XOR DI(216) XOR DI(367) XOR DI(301) XOR DI(376) XOR DI(214) XOR DI(121) XOR DI(374) XOR DI(145) XOR DI(95) XOR DI(340) XOR DI(398) XOR DI(310) XOR DI(448) XOR DI(34) XOR DI(174) XOR DI(385) XOR DI(486) XOR DI(259) XOR DI(223) XOR DI(199) XOR DI(130) XOR DI(383) XOR DI(415) XOR DI(154) XOR DI(78) XOR DI(104) XOR DI(299) XOR DI(353) XOR DI(32) XOR DI(149) XOR DI(429) XOR DI(103) XOR DI(430) XOR DI(341) XOR DI(1) XOR DI(20) XOR DI(417) XOR DI(169) XOR DI(502) XOR DI(481) XOR DI(250) XOR DI(349) XOR DI(53) XOR DI(170) XOR DI(277) XOR DI(407) XOR DI(319) XOR DI(457) XOR DI(246) XOR DI(215) XOR DI(93) XOR DI(477) XOR DI(339) XOR DI(43) XOR DI(450) XOR DI(312) XOR DI(119) XOR DI(61) XOR DI(183) XOR DI(461) XOR DI(323) XOR DI(167) XOR DI(394) XOR DI(479) XOR DI(408) XOR DI(281) XOR DI(458) XOR DI(25) XOR DI(410) XOR DI(495) XOR DI(268) XOR DI(237) XOR DI(206) XOR DI(303) XOR DI(314) XOR DI(3) XOR DI(232) XOR DI(228) XOR DI(219) XOR DI(295) XOR DI(208) XOR DI(115) XOR DI(368) XOR DI(139) XOR DI(89) XOR DI(392) XOR DI(304) XOR DI(28) XOR DI(379) XOR DI(480) XOR DI(217) XOR DI(193) XOR DI(124) XOR DI(377) XOR DI(148) XOR DI(143) XOR DI(97) XOR DI(424) XOR DI(163) XOR DI(47) XOR DI(164) XOR DI(401) XOR DI(313) XOR DI(451) XOR DI(209) XOR DI(87) XOR DI(444) XOR DI(113) XOR DI(177) XOR DI(317) XOR DI(388) XOR DI(19) XOR DI(297) XOR DI(308) XOR DI(213) XOR DI(202) XOR DI(362) XOR DI(133) XOR DI(386) XOR DI(22) XOR DI(474) XOR DI(211) XOR DI(118) XOR DI(142) XOR DI(137) XOR DI(41) XOR DI(158) XOR DI(395) XOR DI(445) XOR DI(438) XOR DI(107) XOR DI(302) XOR DI(196) XOR DI(356) XOR DI(16) XOR DI(112) XOR DI(35) XOR DI(152) XOR DI(439) XOR DI(432) XOR DI(190) XOR DI(350) XOR DI(10) XOR DI(106) XOR DI(29) XOR DI(426) XOR DI(184) XOR DI(344) XOR DI(4) XOR DI(23) XOR DI(178) XOR DI(17) XOR DI(172) XOR DI(11) XOR DI(166) XOR DI(5) XOR DI(499) XOR DI(505) XOR DI(511);
end architecture;