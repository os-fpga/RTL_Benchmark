LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
ENTITY FinalBalancedFIR IS PORT (
	Load : IN std_logic;
	Ct0 : OUT std_logic;
	Ct1 : OUT std_logic;
	nRST : IN std_logic;
	Ct2 : OUT std_logic;
	Ct3 : OUT std_logic;
	Total10 : OUT std_logic;
	Total11 : OUT std_logic;
	Total12 : OUT std_logic;
	Total13 : OUT std_logic;
	Total14 : OUT std_logic;
	Total15 : OUT std_logic;
	Qco0 : OUT std_logic;
	Qco1 : OUT std_logic;
	Qco2 : OUT std_logic;
	Qco3 : OUT std_logic;
	Qco4 : OUT std_logic;
	Qco5 : OUT std_logic;
	Qco6 : OUT std_logic;
	Qco7 : OUT std_logic;
	Dsg0 : IN std_logic;
	Dsg1 : IN std_logic;
	Dsg2 : IN std_logic;
	Dsg3 : IN std_logic;
	Dsg4 : IN std_logic;
	Dsg5 : IN std_logic;
	Dsg6 : IN std_logic;
	Dsg7 : IN std_logic;
	Total0 : OUT std_logic;
	Total1 : OUT std_logic;
	Total2 : OUT std_logic;
	Total3 : OUT std_logic;
	Total4 : OUT std_logic;
	Total5 : OUT std_logic;
	Total6 : OUT std_logic;
	Total7 : OUT std_logic;
	Total8 : OUT std_logic;
	Total9 : OUT std_logic;
	Clk : IN std_logic;
	nCt0 : OUT std_logic;
	nCt1 : OUT std_logic;
	nCt2 : OUT std_logic;
	nCt3 : OUT std_logic;
	Qsg0 : OUT std_logic;
	Qsg1 : OUT std_logic;
	Qsg2 : OUT std_logic;
	Qsg3 : OUT std_logic;
	Qsg4 : OUT std_logic;
	Qsg5 : OUT std_logic;
	Qsg6 : OUT std_logic;
	Qsg7 : OUT std_logic;
	Dco0 : IN std_logic;
	Dco1 : IN std_logic;
	Dco2 : IN std_logic;
	Dco3 : IN std_logic;
	Dco4 : IN std_logic;
	Dco5 : IN std_logic;
	Dco6 : IN std_logic;
	Dco7 : IN std_logic
); 

END FinalBalancedFIR;



ARCHITECTURE STRUCTURE OF FinalBalancedFIR IS

-- COMPONENTS

COMPONENT NEWSLICE
	PORT (
	CLK : IN std_logic;
	DCO0 : IN std_logic;
	DCO1 : IN std_logic;
	DCO2 : IN std_logic;
	DCO3 : IN std_logic;
	DCO4 : IN std_logic;
	DCO5 : IN std_logic;
	DCO6 : IN std_logic;
	DCO7 : IN std_logic;
	DSG0 : IN std_logic;
	DSG1 : IN std_logic;
	DSG2 : IN std_logic;
	DSG3 : IN std_logic;
	DSG4 : IN std_logic;
	DSG5 : IN std_logic;
	DSG6 : IN std_logic;
	DSG7 : IN std_logic;
	ENABLE : IN std_logic;
	LOAD : IN std_logic;
	NRST : IN std_logic;
	QCO0 : OUT std_logic;
	QCO1 : OUT std_logic;
	QCO2 : OUT std_logic;
	QCO3 : OUT std_logic;
	QCO4 : OUT std_logic;
	QCO5 : OUT std_logic;
	QCO6 : OUT std_logic;
	QCO7 : OUT std_logic;
	QSG0 : OUT std_logic;
	QSG1 : OUT std_logic;
	QSG2 : OUT std_logic;
	QSG3 : OUT std_logic;
	QSG4 : OUT std_logic;
	QSG5 : OUT std_logic;
	QSG6 : OUT std_logic;
	QSG7 : OUT std_logic;
	S0 : OUT std_logic;
	S1 : OUT std_logic;
	S2 : OUT std_logic;
	S3 : OUT std_logic;
	S4 : OUT std_logic;
	S5 : OUT std_logic;
	S6 : OUT std_logic;
	S7 : OUT std_logic;
	S8 : OUT std_logic;
	S9 : OUT std_logic;
	S10 : OUT std_logic;
	S11 : OUT std_logic;
	S12 : OUT std_logic;
	S13 : OUT std_logic;
	S14 : OUT std_logic;
	S15 : OUT std_logic;
	SIGNED : OUT std_logic
	); END COMPONENT;

COMPONENT EIGHTBITREG
	PORT (
	CLK : IN std_logic;
	D0 : IN std_logic;
	D1 : IN std_logic;
	D2 : IN std_logic;
	D3 : IN std_logic;
	D4 : IN std_logic;
	D5 : IN std_logic;
	D6 : IN std_logic;
	D7 : IN std_logic;
	NPRESET : IN std_logic;
	NRESET : IN std_logic;
	Q0 : OUT std_logic;
	Q1 : OUT std_logic;
	Q2 : OUT std_logic;
	Q3 : OUT std_logic;
	Q4 : OUT std_logic;
	Q5 : OUT std_logic;
	Q6 : OUT std_logic;
	Q7 : OUT std_logic
	); END COMPONENT;

COMPONENT ADDERDELAY
	PORT (
	DIN0 : IN std_logic;
	DIN1 : IN std_logic;
	DIN2 : IN std_logic;
	DIN3 : IN std_logic;
	DIN4 : IN std_logic;
	DIN5 : IN std_logic;
	DIN6 : IN std_logic;
	DIN7 : IN std_logic;
	DIN8 : IN std_logic;
	DIN9 : IN std_logic;
	DIN10 : IN std_logic;
	DIN11 : IN std_logic;
	DIN12 : IN std_logic;
	DIN13 : IN std_logic;
	DIN14 : IN std_logic;
	DIN15 : IN std_logic;
	DOUT0 : OUT std_logic;
	DOUT1 : OUT std_logic;
	DOUT2 : OUT std_logic;
	DOUT3 : OUT std_logic;
	DOUT4 : OUT std_logic;
	DOUT5 : OUT std_logic;
	DOUT6 : OUT std_logic;
	DOUT7 : OUT std_logic;
	DOUT8 : OUT std_logic;
	DOUT9 : OUT std_logic;
	DOUT10 : OUT std_logic;
	DOUT11 : OUT std_logic;
	DOUT12 : OUT std_logic;
	DOUT13 : OUT std_logic;
	DOUT14 : OUT std_logic;
	DOUT15 : OUT std_logic;
	SIGNEDIN : IN std_logic;
	SIGNEDOUT : OUT std_logic
	); END COMPONENT;

COMPONENT \16adderBalanced\
	PORT (
	A0 : IN std_logic;
	A1 : IN std_logic;
	A2 : IN std_logic;
	A3 : IN std_logic;
	A4 : IN std_logic;
	A5 : IN std_logic;
	A6 : IN std_logic;
	A7 : IN std_logic;
	A8 : IN std_logic;
	A9 : IN std_logic;
	A10 : IN std_logic;
	A11 : IN std_logic;
	A12 : IN std_logic;
	A13 : IN std_logic;
	A14 : IN std_logic;
	A15 : IN std_logic;
	B0 : IN std_logic;
	B1 : IN std_logic;
	B2 : IN std_logic;
	B3 : IN std_logic;
	B4 : IN std_logic;
	B5 : IN std_logic;
	B6 : IN std_logic;
	B7 : IN std_logic;
	B8 : IN std_logic;
	B9 : IN std_logic;
	B10 : IN std_logic;
	B11 : IN std_logic;
	B12 : IN std_logic;
	B13 : IN std_logic;
	B14 : IN std_logic;
	B15 : IN std_logic;
	CIN : IN std_logic;
	COUT : OUT std_logic;
	Y0 : OUT std_logic;
	Y1 : OUT std_logic;
	Y2 : OUT std_logic;
	Y3 : OUT std_logic;
	Y4 : OUT std_logic;
	Y5 : OUT std_logic;
	Y6 : OUT std_logic;
	Y7 : OUT std_logic;
	Y8 : OUT std_logic;
	Y9 : OUT std_logic;
	Y10 : OUT std_logic;
	Y11 : OUT std_logic;
	Y12 : OUT std_logic;
	Y13 : OUT std_logic;
	Y14 : OUT std_logic;
	Y15 : OUT std_logic
	); END COMPONENT;

COMPONENT TAPADDER
	PORT (
	A0 : IN std_logic;
	A1 : IN std_logic;
	A2 : IN std_logic;
	A3 : IN std_logic;
	A4 : IN std_logic;
	A5 : IN std_logic;
	A6 : IN std_logic;
	A7 : IN std_logic;
	A8 : IN std_logic;
	A9 : IN std_logic;
	A10 : IN std_logic;
	A11 : IN std_logic;
	A12 : IN std_logic;
	A13 : IN std_logic;
	A14 : IN std_logic;
	A15 : IN std_logic;
	AND1 : IN std_logic;
	AND2 : IN std_logic;
	AND3 : IN std_logic;
	B0 : IN std_logic;
	B1 : IN std_logic;
	B2 : IN std_logic;
	B3 : IN std_logic;
	B4 : IN std_logic;
	B5 : IN std_logic;
	B6 : IN std_logic;
	B7 : IN std_logic;
	B8 : IN std_logic;
	B9 : IN std_logic;
	B10 : IN std_logic;
	B11 : IN std_logic;
	B12 : IN std_logic;
	B13 : IN std_logic;
	B14 : IN std_logic;
	B15 : IN std_logic;
	CIN : IN std_logic;
	COUT : OUT std_logic;
	O0 : OUT std_logic;
	O1 : OUT std_logic;
	O2 : OUT std_logic;
	O3 : OUT std_logic;
	O4 : OUT std_logic;
	O5 : OUT std_logic;
	O6 : OUT std_logic;
	O7 : OUT std_logic;
	O8 : OUT std_logic;
	O9 : OUT std_logic;
	O10 : OUT std_logic;
	O11 : OUT std_logic;
	O12 : OUT std_logic;
	O13 : OUT std_logic;
	O14 : OUT std_logic;
	O15 : OUT std_logic;
	OR1 : IN std_logic;
	OR2 : IN std_logic;
	OR3 : IN std_logic;
	Y0 : OUT std_logic;
	Y1 : OUT std_logic;
	Y2 : OUT std_logic;
	Y3 : OUT std_logic;
	Y4 : OUT std_logic;
	Y5 : OUT std_logic;
	Y6 : OUT std_logic;
	Y7 : OUT std_logic;
	Y8 : OUT std_logic;
	Y9 : OUT std_logic;
	Y10 : OUT std_logic;
	Y11 : OUT std_logic;
	Y12 : OUT std_logic;
	Y13 : OUT std_logic;
	Y14 : OUT std_logic;
	Y15 : OUT std_logic
	); END COMPONENT;

COMPONENT COUNTER
	PORT (
	CLK : IN std_logic;
	NCLR : IN std_logic;
	NPRE : IN std_logic;
	NQ0 : OUT std_logic;
	NQ1 : OUT std_logic;
	NQ2 : OUT std_logic;
	NQ3 : OUT std_logic;
	Q0 : OUT std_logic;
	Q1 : OUT std_logic;
	Q2 : OUT std_logic;
	Q3 : OUT std_logic
	); END COMPONENT;

COMPONENT ORBLOCK
	PORT (
	A0 : INOUT std_logic;
	A1 : INOUT std_logic;
	A2 : INOUT std_logic;
	A3 : INOUT std_logic;
	A4 : INOUT std_logic;
	A5 : INOUT std_logic;
	A6 : INOUT std_logic;
	A7 : INOUT std_logic;
	A8 : INOUT std_logic;
	A9 : INOUT std_logic;
	A10 : INOUT std_logic;
	A11 : INOUT std_logic;
	A12 : INOUT std_logic;
	A13 : INOUT std_logic;
	A14 : INOUT std_logic;
	A15 : INOUT std_logic;
	B0 : INOUT std_logic;
	B1 : INOUT std_logic;
	B2 : INOUT std_logic;
	B3 : INOUT std_logic;
	B4 : INOUT std_logic;
	B5 : INOUT std_logic;
	B6 : INOUT std_logic;
	B7 : INOUT std_logic;
	B8 : INOUT std_logic;
	B9 : INOUT std_logic;
	B10 : INOUT std_logic;
	B11 : INOUT std_logic;
	B12 : INOUT std_logic;
	B13 : INOUT std_logic;
	B14 : INOUT std_logic;
	B15 : INOUT std_logic;
	C0 : INOUT std_logic;
	C1 : INOUT std_logic;
	C2 : INOUT std_logic;
	C3 : INOUT std_logic;
	C4 : INOUT std_logic;
	C5 : INOUT std_logic;
	C6 : INOUT std_logic;
	C7 : INOUT std_logic;
	C8 : INOUT std_logic;
	C9 : INOUT std_logic;
	C10 : INOUT std_logic;
	C11 : INOUT std_logic;
	C12 : INOUT std_logic;
	C13 : INOUT std_logic;
	C14 : INOUT std_logic;
	C15 : INOUT std_logic;
	D0 : INOUT std_logic;
	D1 : INOUT std_logic;
	D2 : INOUT std_logic;
	D3 : INOUT std_logic;
	D4 : INOUT std_logic;
	D5 : INOUT std_logic;
	D6 : INOUT std_logic;
	D7 : INOUT std_logic;
	D8 : INOUT std_logic;
	D9 : INOUT std_logic;
	D10 : INOUT std_logic;
	D11 : INOUT std_logic;
	D12 : INOUT std_logic;
	D13 : INOUT std_logic;
	D14 : INOUT std_logic;
	D15 : INOUT std_logic;
	E0 : INOUT std_logic;
	E1 : INOUT std_logic;
	E2 : INOUT std_logic;
	E3 : INOUT std_logic;
	E4 : INOUT std_logic;
	E5 : INOUT std_logic;
	E6 : INOUT std_logic;
	E7 : INOUT std_logic;
	E8 : INOUT std_logic;
	E9 : INOUT std_logic;
	E10 : INOUT std_logic;
	E11 : INOUT std_logic;
	E12 : INOUT std_logic;
	E13 : INOUT std_logic;
	E14 : INOUT std_logic;
	E15 : INOUT std_logic;
	F0 : INOUT std_logic;
	F1 : INOUT std_logic;
	F2 : INOUT std_logic;
	F3 : INOUT std_logic;
	F4 : INOUT std_logic;
	F5 : INOUT std_logic;
	F6 : INOUT std_logic;
	F7 : INOUT std_logic;
	F8 : INOUT std_logic;
	F9 : INOUT std_logic;
	F10 : INOUT std_logic;
	F11 : INOUT std_logic;
	F12 : INOUT std_logic;
	F13 : INOUT std_logic;
	F14 : INOUT std_logic;
	F15 : INOUT std_logic;
	G0 : INOUT std_logic;
	G1 : INOUT std_logic;
	G2 : INOUT std_logic;
	G3 : INOUT std_logic;
	G4 : INOUT std_logic;
	G5 : INOUT std_logic;
	G6 : INOUT std_logic;
	G7 : INOUT std_logic;
	G8 : INOUT std_logic;
	G9 : INOUT std_logic;
	G10 : INOUT std_logic;
	G11 : INOUT std_logic;
	G12 : INOUT std_logic;
	G13 : INOUT std_logic;
	G14 : INOUT std_logic;
	G15 : INOUT std_logic;
	H0 : INOUT std_logic;
	H1 : INOUT std_logic;
	H2 : INOUT std_logic;
	H3 : INOUT std_logic;
	H4 : INOUT std_logic;
	H5 : INOUT std_logic;
	H6 : INOUT std_logic;
	H7 : INOUT std_logic;
	H8 : INOUT std_logic;
	H9 : INOUT std_logic;
	H10 : INOUT std_logic;
	H11 : INOUT std_logic;
	H12 : INOUT std_logic;
	H13 : INOUT std_logic;
	H14 : INOUT std_logic;
	H15 : INOUT std_logic;
	OUTPUT0 : INOUT std_logic;
	OUTPUT1 : INOUT std_logic;
	OUTPUT2 : INOUT std_logic;
	OUTPUT3 : INOUT std_logic;
	OUTPUT4 : INOUT std_logic;
	OUTPUT5 : INOUT std_logic;
	OUTPUT6 : INOUT std_logic;
	OUTPUT7 : INOUT std_logic;
	OUTPUT8 : INOUT std_logic;
	OUTPUT9 : INOUT std_logic;
	OUTPUT10 : INOUT std_logic;
	OUTPUT11 : INOUT std_logic;
	OUTPUT12 : INOUT std_logic;
	OUTPUT13 : INOUT std_logic;
	OUTPUT14 : INOUT std_logic;
	OUTPUT15 : INOUT std_logic
	); END COMPONENT;

COMPONENT \7404\
	PORT (
	A_A : IN std_logic;
	Y_A : OUT std_logic;
	GND : IN std_logic;
	VCC : IN std_logic;
	A_B : IN std_logic;
	Y_B : OUT std_logic;
	A_C : IN std_logic;
	Y_C : OUT std_logic;
	A_D : IN std_logic;
	Y_D : OUT std_logic;
	A_E : IN std_logic;
	Y_E : OUT std_logic;
	A_F : IN std_logic;
	Y_F : OUT std_logic
	); END COMPONENT;

COMPONENT \7408\
	PORT (
	A_A : IN std_logic;
	B_A : IN std_logic;
	Y_A : OUT std_logic;
	VCC : IN std_logic;
	GND : IN std_logic;
	A_B : IN std_logic;
	B_B : IN std_logic;
	Y_B : OUT std_logic;
	A_C : IN std_logic;
	B_C : IN std_logic;
	Y_C : OUT std_logic;
	A_D : IN std_logic;
	B_D : IN std_logic;
	Y_D : OUT std_logic
	); END COMPONENT;

COMPONENT ENABLEALL
	PORT (
	C0 : IN std_logic;
	C1 : IN std_logic;
	C2 : IN std_logic;
	C3 : IN std_logic;
	ENABLEELEVEN : OUT std_logic;
	ENABLEFIFTEEN : OUT std_logic;
	ENABLEFIVE : OUT std_logic;
	ENABLEFOUR : OUT std_logic;
	ENABLEFOURTEEN : OUT std_logic;
	ENABLENINE : OUT std_logic;
	ENABLEONE : OUT std_logic;
	ENABLESEVEN : OUT std_logic;
	ENABLESIX : OUT std_logic;
	ENABLETEN : OUT std_logic;
	ENABLETHIRTEEN : OUT std_logic;
	ENABLETHREE : OUT std_logic;
	ENABLETWELVE : OUT std_logic;
	ENABLETWO : OUT std_logic;
	NC0 : IN std_logic;
	NC1 : IN std_logic;
	NC2 : IN std_logic
	); END COMPONENT;

-- SIGNALS

SIGNAL N107814 : std_logic;
SIGNAL N112080923 : std_logic;
SIGNAL N112178123 : std_logic;
SIGNAL N84208 : std_logic;
SIGNAL N108274 : std_logic;
SIGNAL N112080916 : std_logic;
SIGNAL N112615518 : std_logic;
SIGNAL N83415 : std_logic;
SIGNAL N107818 : std_logic;
SIGNAL N111716427 : std_logic;
SIGNAL N110807428 : std_logic;
SIGNAL N83423 : std_logic;
SIGNAL N110985131 : std_logic;
SIGNAL N111886530 : std_logic;
SIGNAL N1147618 : std_logic;
SIGNAL N06027 : std_logic;
SIGNAL N108266 : std_logic;
SIGNAL N11085609 : std_logic;
SIGNAL N112251024 : std_logic;
SIGNAL N06035 : std_logic;
SIGNAL N107826 : std_logic;
SIGNAL N110678325 : std_logic;
SIGNAL COTEST6 : std_logic;
SIGNAL TF9 : std_logic;
SIGNAL N112712724 : std_logic;
SIGNAL N110985133 : std_logic;
SIGNAL COTEST7 : std_logic;
SIGNAL N108282 : std_logic;
SIGNAL N112518330 : std_logic;
SIGNAL N111716420 : std_logic;
SIGNAL ENABLE12 : std_logic;
SIGNAL N108254 : std_logic;
SIGNAL N110985124 : std_logic;
SIGNAL ENABLE3 : std_logic;
SIGNAL N110960826 : std_logic;
SIGNAL N1147650 : std_logic;
SIGNAL N1143318 : std_logic;
SIGNAL N111424833 : std_logic;
SIGNAL N113729323 : std_logic;
SIGNAL N1147602 : std_logic;
SIGNAL B15 : std_logic;
SIGNAL N11054923 : std_logic;
SIGNAL N112712716 : std_logic;
SIGNAL N1147626 : std_logic;
SIGNAL N78511 : std_logic;
SIGNAL N11077939 : std_logic;
SIGNAL N110960818 : std_logic;
SIGNAL N1147594 : std_logic;
SIGNAL N78513 : std_logic;
SIGNAL N110960817 : std_logic;
SIGNAL N111449127 : std_logic;
SIGNAL N1147598 : std_logic;
SIGNAL N78525 : std_logic;
SIGNAL TF1 : std_logic;
SIGNAL N110625912 : std_logic;
SIGNAL N111424830 : std_logic;
SIGNAL C9 : std_logic;
SIGNAL N11062593 : std_logic;
SIGNAL N111424818 : std_logic;
SIGNAL N1147606 : std_logic;
SIGNAL N1146797 : std_logic;
SIGNAL N112494016 : std_logic;
SIGNAL N110549215 : std_logic;
SIGNAL N1147630 : std_logic;
SIGNAL N1146825 : std_logic;
SIGNAL N112469725 : std_logic;
SIGNAL N110960827 : std_logic;
SIGNAL N1147658 : std_logic;
SIGNAL N1146837 : std_logic;
SIGNAL N111983733 : std_logic;
SIGNAL N110932726 : std_logic;
SIGNAL N1147610 : std_logic;
SIGNAL N1146801 : std_logic;
SIGNAL TF4 : std_logic;
SIGNAL N111959418 : std_logic;
SIGNAL N111983728 : std_logic;
SIGNAL TEST0 : std_logic;
SIGNAL TF12 : std_logic;
SIGNAL N111959427 : std_logic;
SIGNAL N111959431 : std_logic;
SIGNAL TF14 : std_logic;
SIGNAL N111959420 : std_logic;
SIGNAL N112105223 : std_logic;
SIGNAL N107806 : std_logic;
SIGNAL N112372531 : std_logic;
SIGNAL N111473419 : std_logic;
SIGNAL N108286 : std_logic;
SIGNAL N112348230 : std_logic;
SIGNAL N110347225 : std_logic;
SIGNAL B2 : std_logic;
SIGNAL TF10 : std_logic;
SIGNAL N112348221 : std_logic;
SIGNAL N111009433 : std_logic;
SIGNAL C2 : std_logic;
SIGNAL TF11 : std_logic;
SIGNAL N111473431 : std_logic;
SIGNAL N111037523 : std_logic;
SIGNAL D6 : std_logic;
SIGNAL TF7 : std_logic;
SIGNAL N111473416 : std_logic;
SIGNAL N111009425 : std_logic;
SIGNAL E14 : std_logic;
SIGNAL F12 : std_logic;
SIGNAL N110347216 : std_logic;
SIGNAL N111594933 : std_logic;
SIGNAL N1057701 : std_logic;
SIGNAL F15 : std_logic;
SIGNAL N111009430 : std_logic;
SIGNAL N111619218 : std_logic;
SIGNAL N1147646 : std_logic;
SIGNAL G2 : std_logic;
SIGNAL N111009416 : std_logic;
SIGNAL N112566927 : std_logic;
SIGNAL N1147638 : std_logic;
SIGNAL G12 : std_logic;
SIGNAL N112032325 : std_logic;
SIGNAL N112566920 : std_logic;
SIGNAL N1147642 : std_logic;
SIGNAL TF3 : std_logic;
SIGNAL H11 : std_logic;
SIGNAL N112032316 : std_logic;
SIGNAL N112542621 : std_logic;
SIGNAL N108258 : std_logic;
SIGNAL N11047252 : std_logic;
SIGNAL N111215229 : std_logic;
SIGNAL N80159 : std_logic;
SIGNAL N110500625 : std_logic;
SIGNAL N111215220 : std_logic;
SIGNAL N1147336 : std_logic;
SIGNAL N79348 : std_logic;
SIGNAL N110500620 : std_logic;
SIGNAL N110779331 : std_logic;
SIGNAL N1147292 : std_logic;
SIGNAL N77700 : std_logic;
SIGNAL N110472527 : std_logic;
SIGNAL N110779322 : std_logic;
SIGNAL TE11 : std_logic;
SIGNAL N77718 : std_logic;
SIGNAL N103471 : std_logic;
SIGNAL N110472520 : std_logic;
SIGNAL N111162831 : std_logic;
SIGNAL N77720 : std_logic;
SIGNAL H14 : std_logic;
SIGNAL N111594925 : std_logic;
SIGNAL N11116287 : std_logic;
SIGNAL N1147288 : std_logic;
SIGNAL MONITOR4 : std_logic;
SIGNAL N111594916 : std_logic;
SIGNAL N111910826 : std_logic;
SIGNAL N1147308 : std_logic;
SIGNAL MONITOR8 : std_logic;
SIGNAL N111813630 : std_logic;
SIGNAL N111570622 : std_logic;
SIGNAL TE5 : std_logic;
SIGNAL MONITOR11 : std_logic;
SIGNAL N111813620 : std_logic;
SIGNAL N110831729 : std_logic;
SIGNAL TE8 : std_logic;
SIGNAL N103475 : std_logic;
SIGNAL N1131487 : std_logic;
SIGNAL N111813616 : std_logic;
SIGNAL N110831724 : std_logic;
SIGNAL N103927 : std_logic;
SIGNAL N1130640 : std_logic;
SIGNAL N110472526 : std_logic;
SIGNAL N110932712 : std_logic;
SIGNAL N103903 : std_logic;
SIGNAL N1129254 : std_logic;
SIGNAL N11047259 : std_logic;
SIGNAL N110831721 : std_logic;
SIGNAL N1128792 : std_logic;
SIGNAL N111935131 : std_logic;
SIGNAL N111594926 : std_logic;
SIGNAL N1147324 : std_logic;
SIGNAL N103459 : std_logic;
SIGNAL G14 : std_logic;
SIGNAL N111935121 : std_logic;
SIGNAL N111594917 : std_logic;
SIGNAL N103907 : std_logic;
SIGNAL N111215228 : std_logic;
SIGNAL N111570619 : std_logic;
SIGNAL N1078491 : std_logic;
SIGNAL N110779330 : std_logic;
SIGNAL N111765019 : std_logic;
SIGNAL N1059428 : std_logic;
SIGNAL TE0 : std_logic;
SIGNAL N111162812 : std_logic;
SIGNAL N112080931 : std_logic;
SIGNAL A1 : std_logic;
SIGNAL TE14 : std_logic;
SIGNAL N103931 : std_logic;
SIGNAL N11116289 : std_logic;
SIGNAL N112712729 : std_logic;
SIGNAL N84216 : std_logic;
SIGNAL N103911 : std_logic;
SIGNAL N112445429 : std_logic;
SIGNAL N112712722 : std_logic;
SIGNAL COTEST5 : std_logic;
SIGNAL N110625911 : std_logic;
SIGNAL CHECK2 : std_logic;
SIGNAL TE13 : std_logic;
SIGNAL N103455 : std_logic;
SIGNAL N111570630 : std_logic;
SIGNAL N112542620 : std_logic;
SIGNAL ENABLE13 : std_logic;
SIGNAL N110831716 : std_logic;
SIGNAL N111983727 : std_logic;
SIGNAL N1147328 : std_logic;
SIGNAL N80960 : std_logic;
SIGNAL N111692125 : std_logic;
SIGNAL N111086114 : std_logic;
SIGNAL TE9 : std_logic;
SIGNAL N80980 : std_logic;
SIGNAL N111570629 : std_logic;
SIGNAL N11108610 : std_logic;
SIGNAL N1147332 : std_logic;
SIGNAL N1143354 : std_logic;
SIGNAL N111570616 : std_logic;
SIGNAL N111138527 : std_logic;
SIGNAL B4 : std_logic;
SIGNAL TE12 : std_logic;
SIGNAL TE15 : std_logic;
SIGNAL N112251025 : std_logic;
SIGNAL N112032328 : std_logic;
SIGNAL N78535 : std_logic;
SIGNAL N103915 : std_logic;
SIGNAL N112251016 : std_logic;
SIGNAL N111546331 : std_logic;
SIGNAL N111765027 : std_logic;
SIGNAL N10716208 : std_logic;
SIGNAL N1147312 : std_logic;
SIGNAL N1146829 : std_logic;
SIGNAL N111765018 : std_logic;
SIGNAL N111643519 : std_logic;
SIGNAL N1147272 : std_logic;
SIGNAL D9 : std_logic;
SIGNAL N111361025 : std_logic;
SIGNAL N112275331 : std_logic;
SIGNAL N91226 : std_logic;
SIGNAL TE3 : std_logic;
SIGNAL E15 : std_logic;
SIGNAL N111361016 : std_logic;
SIGNAL N111789317 : std_logic;
SIGNAL TE4 : std_logic;
SIGNAL N110856030 : std_logic;
SIGNAL N112664123 : std_logic;
SIGNAL TE6 : std_logic;
SIGNAL N110856016 : std_logic;
SIGNAL N112323928 : std_logic;
SIGNAL N1147280 : std_logic;
SIGNAL N94155 : std_logic;
SIGNAL N11085601 : std_logic;
SIGNAL N112323921 : std_logic;
SIGNAL N1147300 : std_logic;
SIGNAL B7 : std_logic;
SIGNAL N112105226 : std_logic;
SIGNAL N111473422 : std_logic;
SIGNAL N1147276 : std_logic;
SIGNAL C6 : std_logic;
SIGNAL N103467 : std_logic;
SIGNAL N112105216 : std_logic;
SIGNAL N110755031 : std_logic;
SIGNAL C15 : std_logic;
SIGNAL N112080927 : std_logic;
SIGNAL N110755017 : std_logic;
SIGNAL N1147316 : std_logic;
SIGNAL D4 : std_logic;
SIGNAL N103923 : std_logic;
SIGNAL N112080918 : std_logic;
SIGNAL N110730724 : std_logic;
SIGNAL D14 : std_logic;
SIGNAL E2 : std_logic;
SIGNAL N103479 : std_logic;
SIGNAL N112323933 : std_logic;
SIGNAL N112396829 : std_logic;
SIGNAL N112323927 : std_logic;
SIGNAL N111215231 : std_logic;
SIGNAL CHECK4 : std_logic;
SIGNAL TE1 : std_logic;
SIGNAL N112323918 : std_logic;
SIGNAL N111190924 : std_logic;
SIGNAL N1058015 : std_logic;
SIGNAL CHECK10 : std_logic;
SIGNAL N103463 : std_logic;
SIGNAL N112737018 : std_logic;
SIGNAL N111061823 : std_logic;
SIGNAL N79334 : std_logic;
SIGNAL N112712717 : std_logic;
SIGNAL N110395811 : std_logic;
SIGNAL N1147320 : std_logic;
SIGNAL N93236 : std_logic;
SIGNAL N112785628 : std_logic;
SIGNAL N110908416 : std_logic;
SIGNAL N1145381 : std_logic;
SIGNAL TE7 : std_logic;
SIGNAL N103935 : std_logic;
SIGNAL N112761330 : std_logic;
SIGNAL N110884117 : std_logic;
SIGNAL N1145365 : std_logic;
SIGNAL N103919 : std_logic;
SIGNAL N112542628 : std_logic;
SIGNAL N112591217 : std_logic;
SIGNAL N1145389 : std_logic;
SIGNAL N110319128 : std_logic;
SIGNAL N112566919 : std_logic;
SIGNAL N1147296 : std_logic;
SIGNAL N1145357 : std_logic;
SIGNAL N110319114 : std_logic;
SIGNAL N110448224 : std_logic;
SIGNAL H10 : std_logic;
SIGNAL N1147304 : std_logic;
SIGNAL MONITOR7 : std_logic;
SIGNAL N111138519 : std_logic;
SIGNAL N111361030 : std_logic;
SIGNAL TE2 : std_logic;
SIGNAL N112032333 : std_logic;
SIGNAL N110448223 : std_logic;
SIGNAL MONITOR9 : std_logic;
SIGNAL TE10 : std_logic;
SIGNAL N110577328 : std_logic;
SIGNAL N111667823 : std_logic;
SIGNAL MONITOR13 : std_logic;
SIGNAL N1147284 : std_logic;
SIGNAL G3 : std_logic;
SIGNAL N110577323 : std_logic;
SIGNAL N110423930 : std_logic;
SIGNAL N1146958 : std_logic;
SIGNAL G11 : std_logic;
SIGNAL N110549229 : std_logic;
SIGNAL N110423925 : std_logic;
SIGNAL N1146994 : std_logic;
SIGNAL N10716203 : std_logic;
SIGNAL N112664133 : std_logic;
SIGNAL N1078481 : std_logic;
SIGNAL TD5 : std_logic;
SIGNAL N110908433 : std_logic;
SIGNAL N112421118 : std_logic;
SIGNAL N1078483 : std_logic;
SIGNAL TD13 : std_logic;
SIGNAL N102889 : std_logic;
SIGNAL N110908417 : std_logic;
SIGNAL N112348220 : std_logic;
SIGNAL A11 : std_logic;
SIGNAL N112275333 : std_logic;
SIGNAL N111546325 : std_logic;
SIGNAL COONETEST5 : std_logic;
SIGNAL N102425 : std_logic;
SIGNAL N112299623 : std_logic;
SIGNAL N110654031 : std_logic;
SIGNAL N1146986 : std_logic;
SIGNAL N06033 : std_logic;
SIGNAL N111789333 : std_logic;
SIGNAL N111497716 : std_logic;
SIGNAL COTEST0 : std_logic;
SIGNAL N102885 : std_logic;
SIGNAL N111813623 : std_logic;
SIGNAL N112202430 : std_logic;
SIGNAL TD2 : std_logic;
SIGNAL ENABLE2 : std_logic;
SIGNAL N111789325 : std_logic;
SIGNAL N112202416 : std_logic;
SIGNAL N1146990 : std_logic;
SIGNAL N1143338 : std_logic;
SIGNAL N112664125 : std_logic;
SIGNAL N112396828 : std_logic;
SIGNAL TD10 : std_logic;
SIGNAL N78517 : std_logic;
SIGNAL N112469727 : std_logic;
SIGNAL N112396821 : std_logic;
SIGNAL N78527 : std_logic;
SIGNAL N102441 : std_logic;
SIGNAL N102433 : std_logic;
SIGNAL N112469718 : std_logic;
SIGNAL N112372530 : std_logic;
SIGNAL C4 : std_logic;
SIGNAL N110266718 : std_logic;
SIGNAL N110755023 : std_logic;
SIGNAL N1146974 : std_logic;
SIGNAL ENABLE10 : std_logic;
SIGNAL N11026674 : std_logic;
SIGNAL N110755016 : std_logic;
SIGNAL N1146978 : std_logic;
SIGNAL N1146809 : std_logic;
SIGNAL N112323930 : std_logic;
SIGNAL N112785616 : std_logic;
SIGNAL N1146950 : std_logic;
SIGNAL N1146789 : std_logic;
SIGNAL N112299622 : std_logic;
SIGNAL N110500624 : std_logic;
SIGNAL N91244 : std_logic;
SIGNAL N102421 : std_logic;
SIGNAL N111009419 : std_logic;
SIGNAL N111765030 : std_logic;
SIGNAL TEST5 : std_logic;
SIGNAL N102881 : std_logic;
SIGNAL N11100949 : std_logic;
SIGNAL N111740720 : std_logic;
SIGNAL SGTEST5 : std_logic;
SIGNAL N102877 : std_logic;
SIGNAL N11100944 : std_logic;
SIGNAL N110577325 : std_logic;
SIGNAL N1146970 : std_logic;
SIGNAL E8 : std_logic;
SIGNAL N111449129 : std_logic;
SIGNAL N110577316 : std_logic;
SIGNAL TD12 : std_logic;
SIGNAL N110755030 : std_logic;
SIGNAL N110678318 : std_logic;
SIGNAL TD0 : std_logic;
SIGNAL N112396833 : std_logic;
SIGNAL N110654028 : std_logic;
SIGNAL TD8 : std_logic;
SIGNAL N81769 : std_logic;
SIGNAL N112421131 : std_logic;
SIGNAL N110654021 : std_logic;
SIGNAL A2 : std_logic;
SIGNAL N102869 : std_logic;
SIGNAL N112421119 : std_logic;
SIGNAL N110654018 : std_logic;
SIGNAL N1147014 : std_logic;
SIGNAL B8 : std_logic;
SIGNAL N111263829 : std_logic;
SIGNAL N111667824 : std_logic;
SIGNAL N1146982 : std_logic;
SIGNAL B10 : std_logic;
SIGNAL N110347228 : std_logic;
SIGNAL N111643528 : std_logic;
SIGNAL C7 : std_logic;
SIGNAL TD7 : std_logic;
SIGNAL N111215221 : std_logic;
SIGNAL N111643521 : std_logic;
SIGNAL N1146962 : std_logic;
SIGNAL D11 : std_logic;
SIGNAL N111886518 : std_logic;
SIGNAL N111138530 : std_logic;
SIGNAL N1146998 : std_logic;
SIGNAL E6 : std_logic;
SIGNAL N111061825 : std_logic;
SIGNAL N111138516 : std_logic;
SIGNAL N1146954 : std_logic;
SIGNAL N79330 : std_logic;
SIGNAL N111037520 : std_logic;
SIGNAL N112615520 : std_logic;
SIGNAL TD6 : std_logic;
SIGNAL N79338 : std_logic;
SIGNAL N110395832 : std_logic;
SIGNAL N111336731 : std_logic;
SIGNAL N1147006 : std_logic;
SIGNAL N79352 : std_logic;
SIGNAL N110908418 : std_logic;
SIGNAL N111336721 : std_logic;
SIGNAL N1147002 : std_logic;
SIGNAL N1145329 : std_logic;
SIGNAL N110884122 : std_logic;
SIGNAL N110730733 : std_logic;
SIGNAL N1145341 : std_logic;
SIGNAL TD3 : std_logic;
SIGNAL N111162830 : std_logic;
SIGNAL N110730719 : std_logic;
SIGNAL TD4 : std_logic;
SIGNAL N77694 : std_logic;
SIGNAL N111162827 : std_logic;
SIGNAL N111716423 : std_logic;
SIGNAL N77724 : std_logic;
SIGNAL N102893 : std_logic;
SIGNAL N102429 : std_logic;
SIGNAL N11070268 : std_logic;
SIGNAL N112518326 : std_logic;
SIGNAL N75904 : std_logic;
SIGNAL N1130871 : std_logic;
SIGNAL N11070266 : std_logic;
SIGNAL N112494023 : std_logic;
SIGNAL N102901 : std_logic;
SIGNAL G1 : std_logic;
SIGNAL N112566924 : std_logic;
SIGNAL N111114231 : std_logic;
SIGNAL TD1 : std_logic;
SIGNAL G9 : std_logic;
SIGNAL N110423919 : std_logic;
SIGNAL N111086130 : std_logic;
SIGNAL N102445 : std_logic;
SIGNAL N111263816 : std_logic;
SIGNAL N1078487 : std_logic;
SIGNAL TD11 : std_logic;
SIGNAL N110448231 : std_logic;
SIGNAL N110524923 : std_logic;
SIGNAL A8 : std_logic;
SIGNAL N102437 : std_logic;
SIGNAL VCC : std_logic;
SIGNAL N112178125 : std_logic;
SIGNAL TD9 : std_logic;
SIGNAL CHECK8 : std_logic;
SIGNAL N110702616 : std_logic;
SIGNAL N112615526 : std_logic;
SIGNAL TD15 : std_logic;
SIGNAL N1147127 : std_logic;
SIGNAL N111692116 : std_logic;
SIGNAL N110779329 : std_logic;
SIGNAL N1058329 : std_logic;
SIGNAL N1147131 : std_logic;
SIGNAL N102897 : std_logic;
SIGNAL N1147139 : std_logic;
SIGNAL N110549220 : std_logic;
SIGNAL N111886525 : std_logic;
SIGNAL N11054926 : std_logic;
SIGNAL N111886516 : std_logic;
SIGNAL N93230 : std_logic;
SIGNAL N102873 : std_logic;
SIGNAL N111789328 : std_logic;
SIGNAL N111862218 : std_logic;
SIGNAL N1146966 : std_logic;
SIGNAL N93244 : std_logic;
SIGNAL N110395831 : std_logic;
SIGNAL N110884129 : std_logic;
SIGNAL N1147010 : std_logic;
SIGNAL ENABLE5 : std_logic;
SIGNAL N110395817 : std_logic;
SIGNAL N110856022 : std_logic;
SIGNAL TD14 : std_logic;
SIGNAL ENABLE4 : std_logic;
SIGNAL N112737022 : std_logic;
SIGNAL N112251026 : std_logic;
SIGNAL N1146636 : std_logic;
SIGNAL N1143334 : std_logic;
SIGNAL N112737017 : std_logic;
SIGNAL N111619227 : std_logic;
SIGNAL TC1 : std_logic;
SIGNAL N78519 : std_logic;
SIGNAL N112664124 : std_logic;
SIGNAL N111619217 : std_logic;
SIGNAL N78529 : std_logic;
SIGNAL N101361 : std_logic;
SIGNAL N112421126 : std_logic;
SIGNAL N111716422 : std_logic;
SIGNAL C5 : std_logic;
SIGNAL N101357 : std_logic;
SIGNAL N111837926 : std_logic;
SIGNAL N110856013 : std_logic;
SIGNAL N1146644 : std_logic;
SIGNAL TEST4 : std_logic;
SIGNAL N111837917 : std_logic;
SIGNAL N1146632 : std_logic;
SIGNAL N91240 : std_logic;
SIGNAL N110932728 : std_logic;
SIGNAL N113729327 : std_logic;
SIGNAL N94149 : std_logic;
SIGNAL TC8 : std_logic;
SIGNAL N110932719 : std_logic;
SIGNAL N113729318 : std_logic;
SIGNAL TC3 : std_logic;
SIGNAL N82580 : std_logic;
SIGNAL N111522033 : std_logic;
SIGNAL N112712728 : std_logic;
SIGNAL TC9 : std_logic;
SIGNAL N81773 : std_logic;
SIGNAL N111522022 : std_logic;
SIGNAL N110985128 : std_logic;
SIGNAL N1146676 : std_logic;
SIGNAL C0 : std_logic;
SIGNAL N110654022 : std_logic;
SIGNAL N110960830 : std_logic;
SIGNAL TC5 : std_logic;
SIGNAL C13 : std_logic;
SIGNAL N110625924 : std_logic;
SIGNAL N111424825 : std_logic;
SIGNAL D8 : std_logic;
SIGNAL N101349 : std_logic;
SIGNAL N10716204 : std_logic;
SIGNAL N110779313 : std_logic;
SIGNAL TC4 : std_logic;
SIGNAL D13 : std_logic;
SIGNAL N111086122 : std_logic;
SIGNAL N110960829 : std_logic;
SIGNAL N1058643 : std_logic;
SIGNAL E10 : std_logic;
SIGNAL F0 : std_logic;
SIGNAL N112372527 : std_logic;
SIGNAL N110960822 : std_logic;
SIGNAL N1146656 : std_logic;
SIGNAL F5 : std_logic;
SIGNAL N112372517 : std_logic;
SIGNAL N112494033 : std_logic;
SIGNAL TC14 : std_logic;
SIGNAL N110755018 : std_logic;
SIGNAL N111959433 : std_logic;
SIGNAL G0 : std_logic;
SIGNAL N100893 : std_logic;
SIGNAL N113729333 : std_logic;
SIGNAL N112372518 : std_logic;
SIGNAL G13 : std_logic;
SIGNAL N1146660 : std_logic;
SIGNAL N112785619 : std_logic;
SIGNAL N112348225 : std_logic;
SIGNAL H13 : std_logic;
SIGNAL N101341 : std_logic;
SIGNAL N112785617 : std_logic;
SIGNAL N111473426 : std_logic;
SIGNAL N101337 : std_logic;
SIGNAL CHECK5 : std_logic;
SIGNAL N11039588 : std_logic;
SIGNAL N111473421 : std_logic;
SIGNAL N1146664 : std_logic;
SIGNAL N80161 : std_logic;
SIGNAL N110500631 : std_logic;
SIGNAL N110347229 : std_logic;
SIGNAL N1146648 : std_logic;
SIGNAL N79346 : std_logic;
SIGNAL F2 : std_logic;
SIGNAL N111740728 : std_logic;
SIGNAL N110347220 : std_logic;
SIGNAL TC10 : std_logic;
SIGNAL N110601617 : std_logic;
SIGNAL N111037518 : std_logic;
SIGNAL N1146680 : std_logic;
SIGNAL N955599 : std_logic;
SIGNAL N110678326 : std_logic;
SIGNAL N111009429 : std_logic;
SIGNAL TC15 : std_logic;
SIGNAL N75862 : std_logic;
SIGNAL N111667829 : std_logic;
SIGNAL N111009420 : std_logic;
SIGNAL MONITOR16 : std_logic;
SIGNAL N1146684 : std_logic;
SIGNAL N111114223 : std_logic;
SIGNAL N112032329 : std_logic;
SIGNAL H6 : std_logic;
SIGNAL TC0 : std_logic;
SIGNAL N112178129 : std_logic;
SIGNAL N112032320 : std_logic;
SIGNAL N1129716 : std_logic;
SIGNAL TC6 : std_logic;
SIGNAL N112761331 : std_logic;
SIGNAL N1128099 : std_logic;
SIGNAL N110472522 : std_logic;
SIGNAL TC7 : std_logic;
SIGNAL N112615528 : std_logic;
SIGNAL N111594929 : std_logic;
SIGNAL N1078475 : std_logic;
SIGNAL N100909 : std_logic;
SIGNAL N11116286 : std_logic;
SIGNAL N111594920 : std_logic;
SIGNAL N1146668 : std_logic;
SIGNAL CHECK15 : std_logic;
SIGNAL N111336716 : std_logic;
SIGNAL N112566922 : std_logic;
SIGNAL TC11 : std_logic;
SIGNAL N06041 : std_logic;
SIGNAL N110730723 : std_logic;
SIGNAL N111813627 : std_logic;
SIGNAL N101365 : std_logic;
SIGNAL N80964 : std_logic;
SIGNAL N110702622 : std_logic;
SIGNAL N110472530 : std_logic;
SIGNAL N1146652 : std_logic;
SIGNAL N80970 : std_logic;
SIGNAL N111740717 : std_logic;
SIGNAL N111935125 : std_logic;
SIGNAL N1146688 : std_logic;
SIGNAL N78509 : std_logic;
SIGNAL N111716431 : std_logic;
SIGNAL N110779317 : std_logic;
SIGNAL TC12 : std_logic;
SIGNAL C8 : std_logic;
SIGNAL N112518318 : std_logic;
SIGNAL N111162833 : std_logic;
SIGNAL N101345 : std_logic;
SIGNAL N1146845 : std_logic;
SIGNAL N111114233 : std_logic;
SIGNAL N111162817 : std_logic;
SIGNAL N1146841 : std_logic;
SIGNAL N100889 : std_logic;
SIGNAL N110266733 : std_logic;
SIGNAL N110625915 : std_logic;
SIGNAL N1146833 : std_logic;
SIGNAL N100905 : std_logic;
SIGNAL N110266725 : std_logic;
SIGNAL N110831719 : std_logic;
SIGNAL N1146692 : std_logic;
SIGNAL D10 : std_logic;
SIGNAL N111263818 : std_logic;
SIGNAL N110831723 : std_logic;
SIGNAL N91246 : std_logic;
SIGNAL N100897 : std_logic;
SIGNAL N112615523 : std_logic;
SIGNAL N111692120 : std_logic;
SIGNAL N101353 : std_logic;
SIGNAL E9 : std_logic;
SIGNAL N112591231 : std_logic;
SIGNAL N111594928 : std_logic;
SIGNAL N1146672 : std_logic;
SIGNAL N112591224 : std_logic;
SIGNAL N111594919 : std_logic;
SIGNAL N82586 : std_logic;
SIGNAL N101369 : std_logic;
SIGNAL N110779323 : std_logic;
SIGNAL N111570631 : std_logic;
SIGNAL N100913 : std_logic;
SIGNAL N82596 : std_logic;
SIGNAL N110779321 : std_logic;
SIGNAL N111570624 : std_logic;
SIGNAL N100901 : std_logic;
SIGNAL N82600 : std_logic;
SIGNAL N111862223 : std_logic;
SIGNAL N1146628 : std_logic;
SIGNAL N82602 : std_logic;
SIGNAL N112275319 : std_logic;
SIGNAL N112251029 : std_logic;
SIGNAL TC2 : std_logic;
SIGNAL N81775 : std_logic;
SIGNAL N111424821 : std_logic;
SIGNAL N112251020 : std_logic;
SIGNAL TC13 : std_logic;
SIGNAL N81779 : std_logic;
SIGNAL N110678323 : std_logic;
SIGNAL N111765031 : std_logic;
SIGNAL N1146640 : std_logic;
SIGNAL N81783 : std_logic;
SIGNAL F8 : std_logic;
SIGNAL N112080925 : std_logic;
SIGNAL N111361029 : std_logic;
SIGNAL N91214 : std_logic;
SIGNAL N11085604 : std_logic;
SIGNAL N112323931 : std_logic;
SIGNAL N1145079 : std_logic;
SIGNAL CHECK12 : std_logic;
SIGNAL N112761317 : std_logic;
SIGNAL TB4 : std_logic;
SIGNAL N80139 : std_logic;
SIGNAL N111983731 : std_logic;
SIGNAL N1145139 : std_logic;
SIGNAL N80167 : std_logic;
SIGNAL N113729316 : std_logic;
SIGNAL F4 : std_logic;
SIGNAL N111983722 : std_logic;
SIGNAL N91190 : std_logic;
SIGNAL N112712719 : std_logic;
SIGNAL N111983717 : std_logic;
SIGNAL N91210 : std_logic;
SIGNAL N80972 : std_logic;
SIGNAL N112518327 : std_logic;
SIGNAL N11108619 : std_logic;
SIGNAL N1145111 : std_logic;
SIGNAL N1145369 : std_logic;
SIGNAL N110960821 : std_logic;
SIGNAL N110319132 : std_logic;
SIGNAL TB1 : std_logic;
SIGNAL N75820 : std_logic;
SIGNAL N110549212 : std_logic;
SIGNAL N11031911 : std_logic;
SIGNAL N1129023 : std_logic;
SIGNAL TB11 : std_logic;
SIGNAL N11054925 : std_logic;
SIGNAL N111138529 : std_logic;
SIGNAL N1145131 : std_logic;
SIGNAL N1078489 : std_logic;
SIGNAL N11077934 : std_logic;
SIGNAL N111546326 : std_logic;
SIGNAL N1145127 : std_logic;
SIGNAL N1078495 : std_logic;
SIGNAL N110960819 : std_logic;
SIGNAL N111546317 : std_logic;
SIGNAL TB9 : std_logic;
SIGNAL CHECK14 : std_logic;
SIGNAL N110932718 : std_logic;
SIGNAL N107162010 : std_logic;
SIGNAL N1145087 : std_logic;
SIGNAL N84210 : std_logic;
SIGNAL N110625919 : std_logic;
SIGNAL N110908421 : std_logic;
SIGNAL N1066581 : std_logic;
SIGNAL N83409 : std_logic;
SIGNAL N110625914 : std_logic;
SIGNAL N112275326 : std_logic;
SIGNAL N91200 : std_logic;
SIGNAL N83421 : std_logic;
SIGNAL N11062595 : std_logic;
SIGNAL N112469731 : std_logic;
SIGNAL N91206 : std_logic;
SIGNAL COTEST4 : std_logic;
SIGNAL N112494018 : std_logic;
SIGNAL N112469722 : std_logic;
SIGNAL N1145103 : std_logic;
SIGNAL N93234 : std_logic;
SIGNAL N112469717 : std_logic;
SIGNAL N112445421 : std_logic;
SIGNAL N1143362 : std_logic;
SIGNAL N91220 : std_logic;
SIGNAL N111959430 : std_logic;
SIGNAL N110266731 : std_logic;
SIGNAL N1143366 : std_logic;
SIGNAL N91216 : std_logic;
SIGNAL N111959429 : std_logic;
SIGNAL N110266722 : std_logic;
SIGNAL TB7 : std_logic;
SIGNAL C10 : std_logic;
SIGNAL N111959422 : std_logic;
SIGNAL N112323923 : std_logic;
SIGNAL N91196 : std_logic;
SIGNAL D3 : std_logic;
SIGNAL N111935118 : std_logic;
SIGNAL N112299617 : std_logic;
SIGNAL N1145115 : std_logic;
SIGNAL N94157 : std_logic;
SIGNAL N112372526 : std_logic;
SIGNAL N111009426 : std_logic;
SIGNAL N91218 : std_logic;
SIGNAL N111037526 : std_logic;
SIGNAL N111473417 : std_logic;
SIGNAL N91202 : std_logic;
SIGNAL N82588 : std_logic;
SIGNAL N111009428 : std_logic;
SIGNAL N111449119 : std_logic;
SIGNAL N1145099 : std_logic;
SIGNAL N81777 : std_logic;
SIGNAL N110472511 : std_logic;
SIGNAL N110730728 : std_logic;
SIGNAL N1145075 : std_logic;
SIGNAL A3 : std_logic;
SIGNAL N11047254 : std_logic;
SIGNAL N111263819 : std_logic;
SIGNAL TB2 : std_logic;
SIGNAL B6 : std_logic;
SIGNAL N110472529 : std_logic;
SIGNAL N111190919 : std_logic;
SIGNAL TB13 : std_logic;
SIGNAL D15 : std_logic;
SIGNAL N111619221 : std_logic;
SIGNAL N110395815 : std_logic;
SIGNAL F14 : std_logic;
SIGNAL N91208 : std_logic;
SIGNAL N111837933 : std_logic;
SIGNAL N110395813 : std_logic;
SIGNAL G4 : std_logic;
SIGNAL N1145119 : std_logic;
SIGNAL N111837921 : std_logic;
SIGNAL N111190931 : std_logic;
SIGNAL H7 : std_logic;
SIGNAL TB3 : std_logic;
SIGNAL N111837916 : std_logic;
SIGNAL N11070265 : std_logic;
SIGNAL H9 : std_logic;
SIGNAL TB6 : std_logic;
SIGNAL N111813622 : std_logic;
SIGNAL N112566928 : std_logic;
SIGNAL H15 : std_logic;
SIGNAL TB12 : std_logic;
SIGNAL N110472521 : std_logic;
SIGNAL N110423928 : std_logic;
SIGNAL N91212 : std_logic;
SIGNAL N80141 : std_logic;
SIGNAL N111935116 : std_logic;
SIGNAL N111692129 : std_logic;
SIGNAL N1145083 : std_logic;
SIGNAL N80153 : std_logic;
SIGNAL N1147489 : std_logic;
SIGNAL N111215223 : std_logic;
SIGNAL N110549224 : std_logic;
SIGNAL N1145135 : std_logic;
SIGNAL N1147485 : std_logic;
SIGNAL N110779325 : std_logic;
SIGNAL N110549210 : std_logic;
SIGNAL TB10 : std_logic;
SIGNAL N111162825 : std_logic;
SIGNAL N111789318 : std_logic;
SIGNAL N1147445 : std_logic;
SIGNAL N1145107 : std_logic;
SIGNAL N112445431 : std_logic;
SIGNAL N110423927 : std_logic;
SIGNAL N955836 : std_logic;
SIGNAL TB0 : std_logic;
SIGNAL N11062596 : std_logic;
SIGNAL N110395826 : std_logic;
SIGNAL TB8 : std_logic;
SIGNAL N1145333 : std_logic;
SIGNAL N111570625 : std_logic;
SIGNAL N112664128 : std_logic;
SIGNAL TB15 : std_logic;
SIGNAL N77698 : std_logic;
SIGNAL N110831727 : std_logic;
SIGNAL N111837930 : std_logic;
SIGNAL N1145091 : std_logic;
SIGNAL N77710 : std_logic;
SIGNAL N110932715 : std_logic;
SIGNAL N110932732 : std_logic;
SIGNAL N1145123 : std_logic;
SIGNAL N75814 : std_logic;
SIGNAL N11093271 : std_logic;
SIGNAL N110625928 : std_logic;
SIGNAL MONITOR6 : std_logic;
SIGNAL TB5 : std_logic;
SIGNAL N110831718 : std_logic;
SIGNAL N111086131 : std_logic;
SIGNAL N1132733 : std_logic;
SIGNAL TB14 : std_logic;
SIGNAL N110807427 : std_logic;
SIGNAL N112202420 : std_logic;
SIGNAL N1132502 : std_logic;
SIGNAL N1145095 : std_logic;
SIGNAL N112153828 : std_logic;
SIGNAL N112396830 : std_logic;
SIGNAL N1131102 : std_logic;
SIGNAL N91198 : std_logic;
SIGNAL N112153821 : std_logic;
SIGNAL N112396823 : std_logic;
SIGNAL N91204 : std_logic;
SIGNAL N84212 : std_logic;
SIGNAL N112153816 : std_logic;
SIGNAL N112396816 : std_logic;
SIGNAL N91192 : std_logic;
SIGNAL N84218 : std_logic;
SIGNAL N111765022 : std_logic;
SIGNAL N110755033 : std_logic;
SIGNAL N91194 : std_logic;
SIGNAL N84228 : std_logic;
SIGNAL N111361020 : std_logic;
SIGNAL N111497724 : std_logic;
SIGNAL N1141961 : std_logic;
SIGNAL N84236 : std_logic;
SIGNAL N111336727 : std_logic;
SIGNAL N110395821 : std_logic;
SIGNAL TA10 : std_logic;
SIGNAL COONETEST4 : std_logic;
SIGNAL N112105233 : std_logic;
SIGNAL N111740733 : std_logic;
SIGNAL N1142672 : std_logic;
SIGNAL COTEST2 : std_logic;
SIGNAL N112105218 : std_logic;
SIGNAL N111765020 : std_logic;
SIGNAL N1142514 : std_logic;
SIGNAL ENABLE11 : std_logic;
SIGNAL N112080922 : std_logic;
SIGNAL N111765016 : std_logic;
SIGNAL N1142356 : std_logic;
SIGNAL N80952 : std_logic;
SIGNAL N112323922 : std_logic;
SIGNAL N110601621 : std_logic;
SIGNAL TA15 : std_logic;
SIGNAL N1143322 : std_logic;
SIGNAL N112737020 : std_logic;
SIGNAL N110678330 : std_logic;
SIGNAL N1143358 : std_logic;
SIGNAL N100400 : std_logic;
SIGNAL N112785623 : std_logic;
SIGNAL N110654030 : std_logic;
SIGNAL N99948 : std_logic;
SIGNAL N1143310 : std_logic;
SIGNAL N112785618 : std_logic;
SIGNAL N110654023 : std_logic;
SIGNAL N1142988 : std_logic;
SIGNAL N1058800 : std_logic;
SIGNAL N112761325 : std_logic;
SIGNAL N111643530 : std_logic;
SIGNAL N99936 : std_logic;
SIGNAL ENABLE7 : std_logic;
SIGNAL N112542623 : std_logic;
SIGNAL N111643523 : std_logic;
SIGNAL N1142593 : std_logic;
SIGNAL E5 : std_logic;
SIGNAL N111983730 : std_logic;
SIGNAL N111114218 : std_logic;
SIGNAL N1142435 : std_logic;
SIGNAL N11108613 : std_logic;
SIGNAL N112153818 : std_logic;
SIGNAL TA7 : std_logic;
SIGNAL N110319118 : std_logic;
SIGNAL N112761316 : std_logic;
SIGNAL TA9 : std_logic;
SIGNAL N11031919 : std_logic;
SIGNAL N111162810 : std_logic;
SIGNAL N100384 : std_logic;
SIGNAL N94151 : std_logic;
SIGNAL N112032327 : std_logic;
SIGNAL N111336723 : std_logic;
SIGNAL N1143146 : std_logic;
SIGNAL N82594 : std_logic;
SIGNAL N110577330 : std_logic;
SIGNAL N110601625 : std_logic;
SIGNAL TA2 : std_logic;
SIGNAL N82598 : std_logic;
SIGNAL N110549231 : std_logic;
SIGNAL N110702617 : std_logic;
SIGNAL N1063489 : std_logic;
SIGNAL B1 : std_logic;
SIGNAL N10716205 : std_logic;
SIGNAL N111740729 : std_logic;
SIGNAL TA6 : std_logic;
SIGNAL B13 : std_logic;
SIGNAL N111643527 : std_logic;
SIGNAL N112518333 : std_logic;
SIGNAL N100396 : std_logic;
SIGNAL C11 : std_logic;
SIGNAL N111643522 : std_logic;
SIGNAL N111086125 : std_logic;
SIGNAL N1268884 : std_logic;
SIGNAL N100392 : std_logic;
SIGNAL N110908429 : std_logic;
SIGNAL N110524918 : std_logic;
SIGNAL F10 : std_logic;
SIGNAL N1142040 : std_logic;
SIGNAL N112299618 : std_logic;
SIGNAL N111862227 : std_logic;
SIGNAL N99928 : std_logic;
SIGNAL N77702 : std_logic;
SIGNAL N112275325 : std_logic;
SIGNAL N110856024 : std_logic;
SIGNAL N100388 : std_logic;
SIGNAL N75826 : std_logic;
SIGNAL N112275320 : std_logic;
SIGNAL N110856017 : std_logic;
SIGNAL N100376 : std_logic;
SIGNAL N75850 : std_logic;
SIGNAL N110678327 : std_logic;
SIGNAL MONITOR5 : std_logic;
SIGNAL N1142751 : std_logic;
SIGNAL N111789329 : std_logic;
SIGNAL N111619229 : std_logic;
SIGNAL MONITOR12 : std_logic;
SIGNAL TA5 : std_logic;
SIGNAL N111789320 : std_logic;
SIGNAL N111619219 : std_logic;
SIGNAL N1078493 : std_logic;
SIGNAL N99944 : std_logic;
SIGNAL N112664127 : std_logic;
SIGNAL N110985118 : std_logic;
SIGNAL N1078499 : std_logic;
SIGNAL TA8 : std_logic;
SIGNAL N110266713 : std_logic;
SIGNAL N11085608 : std_logic;
SIGNAL A7 : std_logic;
SIGNAL TA12 : std_logic;
SIGNAL N11026678 : std_logic;
SIGNAL N1142830 : std_logic;
SIGNAL N84220 : std_logic;
SIGNAL N112299633 : std_logic;
SIGNAL N1142119 : std_logic;
SIGNAL N84230 : std_logic;
SIGNAL N112299624 : std_logic;
SIGNAL TA0 : std_logic;
SIGNAL N83393 : std_logic;
SIGNAL N111009411 : std_logic;
SIGNAL N112712723 : std_logic;
SIGNAL TA1 : std_logic;
SIGNAL N83413 : std_logic;
SIGNAL N11100946 : std_logic;
SIGNAL N110985123 : std_logic;
SIGNAL N99940 : std_logic;
SIGNAL COONETEST2 : std_logic;
SIGNAL N111473425 : std_logic;
SIGNAL N1143067 : std_logic;
SIGNAL N80966 : std_logic;
SIGNAL N111449124 : std_logic;
SIGNAL N11054922 : std_logic;
SIGNAL N1142909 : std_logic;
SIGNAL N78521 : std_logic;
SIGNAL N110755025 : std_logic;
SIGNAL N11077938 : std_logic;
SIGNAL N1142277 : std_logic;
SIGNAL N78533 : std_logic;
SIGNAL N110755020 : std_logic;
SIGNAL N110960824 : std_logic;
SIGNAL N1142198 : std_logic;
SIGNAL ENABLE15 : std_logic;
SIGNAL N112421121 : std_logic;
SIGNAL N11062599 : std_logic;
SIGNAL TA11 : std_logic;
SIGNAL C1 : std_logic;
SIGNAL N111263824 : std_logic;
SIGNAL N11026672 : std_logic;
SIGNAL TA13 : std_logic;
SIGNAL N1146793 : std_logic;
SIGNAL N110319127 : std_logic;
SIGNAL N112494030 : std_logic;
SIGNAL N99932 : std_logic;
SIGNAL SGTEST0 : std_logic;
SIGNAL N111190927 : std_logic;
SIGNAL N111959417 : std_logic;
SIGNAL N100372 : std_logic;
SIGNAL SGTEST4 : std_logic;
SIGNAL N111910825 : std_logic;
SIGNAL N112348229 : std_logic;
SIGNAL N1141882 : std_logic;
SIGNAL N91236 : std_logic;
SIGNAL N111061827 : std_logic;
SIGNAL N111473428 : std_logic;
SIGNAL N99924 : std_logic;
SIGNAL E1 : std_logic;
SIGNAL N111037527 : std_logic;
SIGNAL N111037530 : std_logic;
SIGNAL N100404 : std_logic;
SIGNAL N111037522 : std_logic;
SIGNAL N112032324 : std_logic;
SIGNAL E11 : std_logic;
SIGNAL N100380 : std_logic;
SIGNAL N110908420 : std_logic;
SIGNAL N110472524 : std_logic;
SIGNAL TA3 : std_logic;
SIGNAL N110884124 : std_logic;
SIGNAL N110472517 : std_logic;
SIGNAL TA4 : std_logic;
SIGNAL N111190916 : std_logic;
SIGNAL N111813617 : std_logic;
SIGNAL TA14 : std_logic;
SIGNAL N111162822 : std_logic;
SIGNAL N111215227 : std_logic;
SIGNAL N110779333 : std_logic;
SIGNAL N81771 : std_logic;
SIGNAL N11093275 : std_logic;
SIGNAL B5 : std_logic;
SIGNAL N11070263 : std_logic;
SIGNAL N111692122 : std_logic;
SIGNAL B9 : std_logic;
SIGNAL N112591220 : std_logic;
SIGNAL N111570626 : std_logic;
SIGNAL N1147457 : std_logic;
SIGNAL N111361027 : std_logic;
SIGNAL N111765017 : std_logic;
SIGNAL N1147477 : std_logic;
SIGNAL N111009410 : std_logic;
SIGNAL N112080926 : std_logic;
SIGNAL N77704 : std_logic;
SIGNAL N11100945 : std_logic;
SIGNAL N112785627 : std_logic;
SIGNAL N77706 : std_logic;
SIGNAL N110448226 : std_logic;
SIGNAL N112542627 : std_logic;
SIGNAL N77712 : std_logic;
SIGNAL N110448217 : std_logic;
SIGNAL N110319122 : std_logic;
SIGNAL N75886 : std_logic;
SIGNAL N110702628 : std_logic;
SIGNAL N110319113 : std_logic;
SIGNAL N75892 : std_logic;
SIGNAL N111667817 : std_logic;
SIGNAL N111546333 : std_logic;
SIGNAL H4 : std_logic;
SIGNAL N110549232 : std_logic;
SIGNAL N110577320 : std_logic;
SIGNAL MONITOR14 : std_logic;
SIGNAL N110549218 : std_logic;
SIGNAL N112299631 : std_logic;
SIGNAL G15 : std_logic;
SIGNAL N11054921 : std_logic;
SIGNAL N112664116 : std_logic;
SIGNAL A0 : std_logic;
SIGNAL N111789330 : std_logic;
SIGNAL N112469726 : std_logic;
SIGNAL A5 : std_logic;
SIGNAL N111061831 : std_logic;
SIGNAL N110266717 : std_logic;
SIGNAL N84214 : std_logic;
SIGNAL N111061826 : std_logic;
SIGNAL N110266712 : std_logic;
SIGNAL N83399 : std_logic;
SIGNAL N111061817 : std_logic;
SIGNAL N112323925 : std_logic;
SIGNAL N83405 : std_logic;
SIGNAL N110319111 : std_logic;
SIGNAL N112299619 : std_logic;
SIGNAL COONETEST0 : std_logic;
SIGNAL N11031914 : std_logic;
SIGNAL N11100941 : std_logic;
SIGNAL CHECK1 : std_logic;
SIGNAL N11031910 : std_logic;
SIGNAL N111449128 : std_logic;
SIGNAL N80962 : std_logic;
SIGNAL N110423917 : std_logic;
SIGNAL N111449123 : std_logic;
SIGNAL N80978 : std_logic;
SIGNAL N110395819 : std_logic;
SIGNAL N111263828 : std_logic;
SIGNAL N1059114 : std_logic;
SIGNAL N112664119 : std_logic;
SIGNAL N111215233 : std_logic;
SIGNAL C12 : std_logic;
SIGNAL N110932723 : std_logic;
SIGNAL N111886520 : std_logic;
SIGNAL D1 : std_logic;
SIGNAL N11093278 : std_logic;
SIGNAL N110884119 : std_logic;
SIGNAL TEST6 : std_logic;
SIGNAL N111546322 : std_logic;
SIGNAL N111162819 : std_logic;
SIGNAL TEST7 : std_logic;
SIGNAL N110654017 : std_logic;
SIGNAL N112566923 : std_logic;
SIGNAL N111522026 : std_logic;
SIGNAL N110448233 : std_logic;
SIGNAL E12 : std_logic;
SIGNAL N111522017 : std_logic;
SIGNAL N110423918 : std_logic;
SIGNAL G6 : std_logic;
SIGNAL N111497728 : std_logic;
SIGNAL N111361033 : std_logic;
SIGNAL CHECK3 : std_logic;
SIGNAL N111497719 : std_logic;
SIGNAL N110448230 : std_logic;
SIGNAL CHECK9 : std_logic;
SIGNAL N107162013 : std_logic;
SIGNAL N111692124 : std_logic;
SIGNAL N80163 : std_logic;
SIGNAL N111086117 : std_logic;
SIGNAL N110549219 : std_logic;
SIGNAL N80165 : std_logic;
SIGNAL N11108612 : std_logic;
SIGNAL N111061830 : std_logic;
SIGNAL N1147449 : std_logic;
SIGNAL N110395812 : std_logic;
SIGNAL N110395828 : std_logic;
SIGNAL N1147461 : std_logic;
SIGNAL N11039583 : std_logic;
SIGNAL N112737021 : std_logic;
SIGNAL N1145345 : std_logic;
SIGNAL N110524926 : std_logic;
SIGNAL N112737016 : std_logic;
SIGNAL N77722 : std_logic;
SIGNAL N110500626 : std_logic;
SIGNAL N112421130 : std_logic;
SIGNAL N75856 : std_logic;
SIGNAL N111740723 : std_logic;
SIGNAL N112421125 : std_logic;
SIGNAL N75898 : std_logic;
SIGNAL N110577319 : std_logic;
SIGNAL N112348222 : std_logic;
SIGNAL H3 : std_logic;
SIGNAL N111667831 : std_logic;
SIGNAL N111837925 : std_logic;
SIGNAL H8 : std_logic;
SIGNAL N111643520 : std_logic;
SIGNAL N111522030 : std_logic;
SIGNAL MONITOR10 : std_logic;
SIGNAL N111138533 : std_logic;
SIGNAL N111522016 : std_logic;
SIGNAL N1128330 : std_logic;
SIGNAL N111138524 : std_logic;
SIGNAL N111522021 : std_logic;
SIGNAL N1078473 : std_logic;
SIGNAL N112178133 : std_logic;
SIGNAL N112396818 : std_logic;
SIGNAL N1078485 : std_logic;
SIGNAL N112178124 : std_logic;
SIGNAL N110395816 : std_logic;
SIGNAL A13 : std_logic;
SIGNAL N112178119 : std_logic;
SIGNAL N110500628 : std_logic;
SIGNAL N112153826 : std_logic;
SIGNAL N111740727 : std_logic;
SIGNAL N1147159 : std_logic;
SIGNAL N83395 : std_logic;
SIGNAL N112761326 : std_logic;
SIGNAL N111740718 : std_logic;
SIGNAL ENABLE6 : std_logic;
SIGNAL N110730725 : std_logic;
SIGNAL N110654025 : std_logic;
SIGNAL N1143314 : std_logic;
SIGNAL N111740719 : std_logic;
SIGNAL N111667816 : std_logic;
SIGNAL N1143350 : std_logic;
SIGNAL N111716426 : std_logic;
SIGNAL N111643525 : std_logic;
SIGNAL N112518320 : std_logic;
SIGNAL N112761328 : std_logic;
SIGNAL N1146813 : std_logic;
SIGNAL N112494026 : std_logic;
SIGNAL N111336725 : std_logic;
SIGNAL D0 : std_logic;
SIGNAL N110266727 : std_logic;
SIGNAL N110601629 : std_logic;
SIGNAL D2 : std_logic;
SIGNAL N91238 : std_logic;
SIGNAL N111263833 : std_logic;
SIGNAL N110702619 : std_logic;
SIGNAL N112615525 : std_logic;
SIGNAL N111740731 : std_logic;
SIGNAL E4 : std_logic;
SIGNAL N112591226 : std_logic;
SIGNAL N110266724 : std_logic;
SIGNAL E13 : std_logic;
SIGNAL N94153 : std_logic;
SIGNAL N110807433 : std_logic;
SIGNAL N112615531 : std_logic;
SIGNAL N110807429 : std_logic;
SIGNAL N112591228 : std_logic;
SIGNAL N110807422 : std_logic;
SIGNAL N110807417 : std_logic;
SIGNAL N82590 : std_logic;
SIGNAL N111886528 : std_logic;
SIGNAL N111862233 : std_logic;
SIGNAL N82608 : std_logic;
SIGNAL N111886519 : std_logic;
SIGNAL N111862222 : std_logic;
SIGNAL C3 : std_logic;
SIGNAL N110856033 : std_logic;
SIGNAL N110856031 : std_logic;
SIGNAL N110856029 : std_logic;
SIGNAL N110856026 : std_logic;
SIGNAL D5 : std_logic;
SIGNAL F6 : std_logic;
SIGNAL N111424823 : std_logic;
SIGNAL N110856019 : std_logic;
SIGNAL N80157 : std_logic;
SIGNAL N111619233 : std_logic;
SIGNAL N112275316 : std_logic;
SIGNAL N1147441 : std_logic;
SIGNAL N110678320 : std_logic;
SIGNAL N1147497 : std_logic;
SIGNAL N111619231 : std_logic;
SIGNAL N78531 : std_logic;
SIGNAL N113729330 : std_logic;
SIGNAL N110985130 : std_logic;
SIGNAL N75880 : std_logic;
SIGNAL N113729321 : std_logic;
SIGNAL N110985120 : std_logic;
SIGNAL H2 : std_logic;
SIGNAL N112518322 : std_logic;
SIGNAL N112518321 : std_logic;
SIGNAL H12 : std_logic;
SIGNAL N110960816 : std_logic;
SIGNAL N110960820 : std_logic;
SIGNAL N1128561 : std_logic;
SIGNAL N111424828 : std_logic;
SIGNAL N111449116 : std_logic;
SIGNAL N1057544 : std_logic;
SIGNAL N111424816 : std_logic;
SIGNAL N111424820 : std_logic;
SIGNAL N1078479 : std_logic;
SIGNAL N11054927 : std_logic;
SIGNAL N110960833 : std_logic;
SIGNAL A14 : std_logic;
SIGNAL N110779332 : std_logic;
SIGNAL N11062592 : std_logic;
SIGNAL N83401 : std_logic;
SIGNAL N110932727 : std_logic;
SIGNAL N111983719 : std_logic;
SIGNAL N83419 : std_logic;
SIGNAL N110932720 : std_logic;
SIGNAL N111959419 : std_logic;
SIGNAL N06029 : std_logic;
SIGNAL N110932716 : std_logic;
SIGNAL N112105225 : std_logic;
SIGNAL CHECK0 : std_logic;
SIGNAL N110625931 : std_logic;
SIGNAL N111473430 : std_logic;
SIGNAL N1143330 : std_logic;
SIGNAL N110625921 : std_logic;
SIGNAL N111037525 : std_logic;
SIGNAL N1143342 : std_logic;
SIGNAL N110625916 : std_logic;
SIGNAL N111009427 : std_logic;
SIGNAL B12 : std_logic;
SIGNAL N11062597 : std_logic;
SIGNAL N11047251 : std_logic;
SIGNAL N112494020 : std_logic;
SIGNAL N110472519 : std_logic;
SIGNAL N78537 : std_logic;
SIGNAL N112469716 : std_logic;
SIGNAL N111813629 : std_logic;
SIGNAL SGTEST1 : std_logic;
SIGNAL N111959425 : std_logic;
SIGNAL N111813619 : std_logic;
SIGNAL SGTEST6 : std_logic;
SIGNAL N111959424 : std_logic;
SIGNAL N91248 : std_logic;
SIGNAL N111935127 : std_logic;
SIGNAL N11047250 : std_logic;
SIGNAL ENABLE1 : std_logic;
SIGNAL N111935120 : std_logic;
SIGNAL N111215222 : std_logic;
SIGNAL N112372521 : std_logic;
SIGNAL N110779324 : std_logic;
SIGNAL N112105230 : std_logic;
SIGNAL N112445428 : std_logic;
SIGNAL N112105221 : std_logic;
SIGNAL N110831731 : std_logic;
SIGNAL N111473423 : std_logic;
SIGNAL N110831726 : std_logic;
SIGNAL N82578 : std_logic;
SIGNAL N110347223 : std_logic;
SIGNAL N111570628 : std_logic;
SIGNAL N82592 : std_logic;
SIGNAL N111037521 : std_logic;
SIGNAL N111361019 : std_logic;
SIGNAL N82604 : std_logic;
SIGNAL N111009423 : std_logic;
SIGNAL N112080933 : std_logic;
SIGNAL N81787 : std_logic;
SIGNAL N110472513 : std_logic;
SIGNAL N112785622 : std_logic;
SIGNAL G10 : std_logic;
SIGNAL N11047256 : std_logic;
SIGNAL N112542622 : std_logic;
SIGNAL CHECK6 : std_logic;
SIGNAL N110472533 : std_logic;
SIGNAL N111983729 : std_logic;
SIGNAL N79326 : std_logic;
SIGNAL N110500618 : std_logic;
SIGNAL N111086132 : std_logic;
SIGNAL N1147493 : std_logic;
SIGNAL N111619225 : std_logic;
SIGNAL N110319117 : std_logic;
SIGNAL N1147465 : std_logic;
SIGNAL N111619216 : std_logic;
SIGNAL N111862217 : std_logic;
SIGNAL F11 : std_logic;
SIGNAL N112566931 : std_logic;
SIGNAL N110577327 : std_logic;
SIGNAL N1145385 : std_logic;
SIGNAL N112542630 : std_logic;
SIGNAL N110577322 : std_logic;
SIGNAL N1145349 : std_logic;
SIGNAL N112542625 : std_logic;
SIGNAL N110549226 : std_logic;
SIGNAL N75832 : std_logic;
SIGNAL N111837923 : std_logic;
SIGNAL N110549216 : std_logic;
SIGNAL N75838 : std_logic;
SIGNAL N111813624 : std_logic;
SIGNAL N10716202 : std_logic;
SIGNAL H0 : std_logic;
SIGNAL N110472516 : std_logic;
SIGNAL N110908428 : std_logic;
SIGNAL MONITOR2 : std_logic;
SIGNAL N111935129 : std_logic;
SIGNAL N112275324 : std_logic;
SIGNAL MONITOR3 : std_logic;
SIGNAL N111215218 : std_logic;
SIGNAL N111789319 : std_logic;
SIGNAL N1130178 : std_logic;
SIGNAL N110779320 : std_logic;
SIGNAL N112299621 : std_logic;
SIGNAL N1129947 : std_logic;
SIGNAL N11077931 : std_logic;
SIGNAL N11100943 : std_logic;
SIGNAL N1078469 : std_logic;
SIGNAL N111162829 : std_logic;
SIGNAL N111473433 : std_logic;
SIGNAL A12 : std_logic;
SIGNAL N11116281 : std_logic;
SIGNAL N111473424 : std_logic;
SIGNAL N84224 : std_logic;
SIGNAL N112445426 : std_logic;
SIGNAL N110755019 : std_logic;
SIGNAL N93242 : std_logic;
SIGNAL N112445418 : std_logic;
SIGNAL N110730726 : std_logic;
SIGNAL ENABLE14 : std_logic;
SIGNAL N111910817 : std_logic;
SIGNAL N111190926 : std_logic;
SIGNAL N78523 : std_logic;
SIGNAL N111570620 : std_logic;
SIGNAL N111910833 : std_logic;
SIGNAL N110831722 : std_logic;
SIGNAL N111886522 : std_logic;
SIGNAL D7 : std_logic;
SIGNAL TEST1 : std_logic;
SIGNAL N112153830 : std_logic;
SIGNAL N110884128 : std_logic;
SIGNAL TEST2 : std_logic;
SIGNAL N112153823 : std_logic;
SIGNAL N110884121 : std_logic;
SIGNAL N91234 : std_logic;
SIGNAL N111594922 : std_logic;
SIGNAL N112591219 : std_logic;
SIGNAL N91250 : std_logic;
SIGNAL N111336722 : std_logic;
SIGNAL N110448225 : std_logic;
SIGNAL N110856023 : std_logic;
SIGNAL N110448216 : std_logic;
SIGNAL E0 : std_logic;
SIGNAL N94147 : std_logic;
SIGNAL N112105220 : std_logic;
SIGNAL N111667825 : std_logic;
SIGNAL N112737029 : std_logic;
SIGNAL N110549217 : std_logic;
SIGNAL N94145 : std_logic;
SIGNAL N112712731 : std_logic;
SIGNAL N11054920 : std_logic;
SIGNAL N112761320 : std_logic;
SIGNAL N111061816 : std_logic;
SIGNAL N112542618 : std_logic;
SIGNAL N112421120 : std_logic;
SIGNAL N111983725 : std_logic;
SIGNAL N112348224 : std_logic;
SIGNAL N82606 : std_logic;
SIGNAL N111983720 : std_logic;
SIGNAL N11093277 : std_logic;
SIGNAL N81795 : std_logic;
SIGNAL N111086112 : std_logic;
SIGNAL N111546316 : std_logic;
SIGNAL A6 : std_logic;
SIGNAL N111138521 : std_logic;
SIGNAL N110654033 : std_logic;
SIGNAL F3 : std_logic;
SIGNAL N112032317 : std_logic;
SIGNAL N110625918 : std_logic;
SIGNAL N80137 : std_logic;
SIGNAL N111546329 : std_logic;
SIGNAL N111522025 : std_logic;
SIGNAL N80149 : std_logic;
SIGNAL N111546320 : std_logic;
SIGNAL N111497718 : std_logic;
SIGNAL N79322 : std_logic;
SIGNAL N110549233 : std_logic;
SIGNAL N112202433 : std_logic;
SIGNAL N79324 : std_logic;
SIGNAL N107162012 : std_logic;
SIGNAL N11039582 : std_logic;
SIGNAL N79342 : std_logic;
SIGNAL N110908424 : std_logic;
SIGNAL N111740722 : std_logic;
SIGNAL F9 : std_logic;
SIGNAL N112275329 : std_logic;
SIGNAL N110577318 : std_logic;
SIGNAL N112664117 : std_logic;
SIGNAL N1145377 : std_logic;
SIGNAL N111667828 : std_logic;
SIGNAL H5 : std_logic;
SIGNAL N112445424 : std_logic;
SIGNAL N112615522 : std_logic;
SIGNAL MONITOR0 : std_logic;
SIGNAL N112445419 : std_logic;
SIGNAL N111716425 : std_logic;
SIGNAL N1078471 : std_logic;
SIGNAL N112299626 : std_logic;
SIGNAL N112494025 : std_logic;
SIGNAL N1078477 : std_logic;
SIGNAL N111009413 : std_logic;
SIGNAL N111114220 : std_logic;
SIGNAL N1147119 : std_logic;
SIGNAL N11100948 : std_logic;
SIGNAL N110266719 : std_logic;
SIGNAL N110524925 : std_logic;
SIGNAL N1147175 : std_logic;
SIGNAL N84206 : std_logic;
SIGNAL N111473420 : std_logic;
SIGNAL N112615533 : std_logic;
SIGNAL N84222 : std_logic;
SIGNAL N111449122 : std_logic;
SIGNAL N112591230 : std_logic;
SIGNAL N83411 : std_logic;
SIGNAL N110730731 : std_logic;
SIGNAL N112591223 : std_logic;
SIGNAL COTEST1 : std_logic;
SIGNAL N110730722 : std_logic;
SIGNAL N110807419 : std_logic;
SIGNAL COTEST3 : std_logic;
SIGNAL N112421123 : std_logic;
SIGNAL N111886527 : std_logic;
SIGNAL N93232 : std_logic;
SIGNAL N112396827 : std_logic;
SIGNAL N110884131 : std_logic;
SIGNAL N80956 : std_logic;
SIGNAL N112396822 : std_logic;
SIGNAL N110856028 : std_logic;
SIGNAL N80968 : std_logic;
SIGNAL N111263822 : std_logic;
SIGNAL N112275318 : std_logic;
SIGNAL N1143326 : std_logic;
SIGNAL N111190922 : std_logic;
SIGNAL N110678322 : std_logic;
SIGNAL N1143306 : std_logic;
SIGNAL N111910820 : std_logic;
SIGNAL N111061829 : std_logic;
SIGNAL N113729320 : std_logic;
SIGNAL N1146817 : std_logic;
SIGNAL N111037529 : std_logic;
SIGNAL N111424827 : std_logic;
SIGNAL D12 : std_logic;
SIGNAL TEST3 : std_logic;
SIGNAL N111037524 : std_logic;
SIGNAL N11054924 : std_logic;
SIGNAL N111037517 : std_logic;
SIGNAL N110932717 : std_logic;
SIGNAL N82582 : std_logic;
SIGNAL N11039585 : std_logic;
SIGNAL N11062594 : std_logic;
SIGNAL N81793 : std_logic;
SIGNAL N110884126 : std_logic;
SIGNAL N112469733 : std_logic;
SIGNAL A10 : std_logic;
SIGNAL N111190933 : std_logic;
SIGNAL N112494017 : std_logic;
SIGNAL G7 : std_logic;
SIGNAL N111190925 : std_logic;
SIGNAL N111959428 : std_logic;
SIGNAL N80155 : std_logic;
SIGNAL N111190918 : std_logic;
SIGNAL N111959421 : std_logic;
SIGNAL N1129485 : std_logic;
SIGNAL N111162824 : std_logic;
SIGNAL N111935117 : std_logic;
SIGNAL G5 : std_logic;
SIGNAL N11070260 : std_logic;
SIGNAL CHECK11 : std_logic;
SIGNAL N112566921 : std_logic;
SIGNAL N112566917 : std_logic;
SIGNAL N112372520 : std_logic;
SIGNAL N1147163 : std_logic;
SIGNAL N110423931 : std_logic;
SIGNAL N110347231 : std_logic;
SIGNAL N1147135 : std_logic;
SIGNAL N110423926 : std_logic;
SIGNAL N110347222 : std_logic;
SIGNAL N1147143 : std_logic;
SIGNAL N1147151 : std_logic;
SIGNAL N111009414 : std_logic;
SIGNAL N111009422 : std_logic;
SIGNAL N11100940 : std_logic;
SIGNAL N112032331 : std_logic;
SIGNAL N1147115 : std_logic;
SIGNAL N83417 : std_logic;
SIGNAL N110448221 : std_logic;
SIGNAL N11047253 : std_logic;
SIGNAL COONETEST6 : std_logic;
SIGNAL N110702623 : std_logic;
SIGNAL N110500617 : std_logic;
SIGNAL N06031 : std_logic;
SIGNAL N110702610 : std_logic;
SIGNAL N110472528 : std_logic;
SIGNAL N93238 : std_logic;
SIGNAL N111667833 : std_logic;
SIGNAL N111813633 : std_logic;
SIGNAL N80950 : std_logic;
SIGNAL N111667821 : std_logic;
SIGNAL N111813631 : std_logic;
SIGNAL N80954 : std_logic;
SIGNAL N110549227 : std_logic;
SIGNAL N111813621 : std_logic;
SIGNAL N80974 : std_logic;
SIGNAL N110549213 : std_logic;
SIGNAL N110472532 : std_logic;
SIGNAL N111061833 : std_logic;
SIGNAL N111935128 : std_logic;
SIGNAL N1143370 : std_logic;
SIGNAL N111061821 : std_logic;
SIGNAL N111215217 : std_logic;
SIGNAL N1146853 : std_logic;
SIGNAL N91224 : std_logic;
SIGNAL N11031916 : std_logic;
SIGNAL N110779319 : std_logic;
SIGNAL N91230 : std_logic;
SIGNAL N112664131 : std_logic;
SIGNAL N110779310 : std_logic;
SIGNAL N112421116 : std_logic;
SIGNAL N112445430 : std_logic;
SIGNAL N111837924 : std_logic;
SIGNAL N110807421 : std_logic;
SIGNAL N81791 : std_logic;
SIGNAL N110932710 : std_logic;
SIGNAL N112153827 : std_logic;
SIGNAL B11 : std_logic;
SIGNAL N11093270 : std_logic;
SIGNAL N111692131 : std_logic;
SIGNAL CHECK13 : std_logic;
SIGNAL N110654029 : std_logic;
SIGNAL N111692126 : std_logic;
SIGNAL N80143 : std_logic;
SIGNAL N111497730 : std_logic;
SIGNAL N110856010 : std_logic;
SIGNAL N79332 : std_logic;
SIGNAL N111497723 : std_logic;
SIGNAL N11085602 : std_logic;
SIGNAL N79350 : std_logic;
SIGNAL N11108614 : std_logic;
SIGNAL N112105227 : std_logic;
SIGNAL N1147469 : std_logic;
SIGNAL N112202428 : std_logic;
SIGNAL N112105217 : std_logic;
SIGNAL N112202423 : std_logic;
SIGNAL N112761319 : std_logic;
SIGNAL N1145353 : std_logic;
SIGNAL N110755022 : std_logic;
SIGNAL N111983724 : std_logic;
SIGNAL N1145337 : std_logic;
SIGNAL N77696 : std_logic;
SIGNAL N110601633 : std_logic;
SIGNAL N111086111 : std_logic;
SIGNAL N75874 : std_logic;
SIGNAL N110601624 : std_logic;
SIGNAL N11031913 : std_logic;
SIGNAL A9 : std_logic;
SIGNAL N110678333 : std_logic;
SIGNAL N112032326 : std_logic;
SIGNAL N110678316 : std_logic;
SIGNAL N111546328 : std_logic;
SIGNAL N1147155 : std_logic;
SIGNAL N84226 : std_logic;
SIGNAL N111667826 : std_logic;
SIGNAL N111546319 : std_logic;
SIGNAL N83403 : std_logic;
SIGNAL N111667818 : std_logic;
SIGNAL N110577329 : std_logic;
SIGNAL N06037 : std_logic;
SIGNAL N111643517 : std_logic;
SIGNAL N110549230 : std_logic;
SIGNAL ENABLE9 : std_logic;
SIGNAL N111138528 : std_logic;
SIGNAL N110908423 : std_logic;
SIGNAL N111114230 : std_logic;
SIGNAL N112299629 : std_logic;
SIGNAL N1143346 : std_logic;
SIGNAL N78539 : std_logic;
SIGNAL N111114221 : std_logic;
SIGNAL N112275328 : std_logic;
SIGNAL N112761333 : std_logic;
SIGNAL N112445423 : std_logic;
SIGNAL C14 : std_logic;
SIGNAL SGTEST7 : std_logic;
SIGNAL N112615516 : std_logic;
SIGNAL N111449121 : std_logic;
SIGNAL N91222 : std_logic;
SIGNAL N111162813 : std_logic;
SIGNAL N110730730 : std_logic;
SIGNAL N91232 : std_logic;
SIGNAL N110730727 : std_logic;
SIGNAL N110730721 : std_logic;
SIGNAL N110702629 : std_logic;
SIGNAL N112421133 : std_logic;
SIGNAL N111716421 : std_logic;
SIGNAL N111263821 : std_logic;
SIGNAL N82584 : std_logic;
SIGNAL N112494021 : std_logic;
SIGNAL N111190921 : std_logic;
SIGNAL N81765 : std_logic;
SIGNAL N111114225 : std_logic;
SIGNAL N111910819 : std_logic;
SIGNAL N81785 : std_logic;
SIGNAL N111086119 : std_logic;
SIGNAL N110884123 : std_logic;
SIGNAL N81789 : std_logic;
SIGNAL N110266729 : std_logic;
SIGNAL N111162828 : std_logic;
SIGNAL N111263827 : std_logic;
SIGNAL N111162821 : std_logic;
SIGNAL E3 : std_logic;
SIGNAL N80147 : std_logic;
SIGNAL N110524930 : std_logic;
SIGNAL N110702615 : std_logic;
SIGNAL N1147453 : std_logic;
SIGNAL N110524921 : std_logic;
SIGNAL N112566930 : std_logic;
SIGNAL N77716 : std_logic;
SIGNAL N112202425 : std_logic;
SIGNAL N110448220 : std_logic;
SIGNAL N75844 : std_logic;
SIGNAL N112615527 : std_logic;
SIGNAL N11070267 : std_logic;
SIGNAL N75868 : std_logic;
SIGNAL N112591218 : std_logic;
SIGNAL N111061820 : std_logic;
SIGNAL N1130409 : std_logic;
SIGNAL N110807431 : std_logic;
SIGNAL N110395818 : std_logic;
SIGNAL N1078467 : std_logic;
SIGNAL N110807424 : std_logic;
SIGNAL N112737028 : std_logic;
SIGNAL GND : std_logic;
SIGNAL N111886523 : std_logic;
SIGNAL N112664130 : std_logic;
SIGNAL N111862230 : std_logic;
SIGNAL N112348231 : std_logic;
SIGNAL N1147123 : std_logic;
SIGNAL N83397 : std_logic;
SIGNAL N110884118 : std_logic;
SIGNAL N111546321 : std_logic;
SIGNAL N83407 : std_logic;
SIGNAL N112275321 : std_logic;
SIGNAL N110625930 : std_logic;
SIGNAL COONETEST1 : std_logic;
SIGNAL N112251027 : std_logic;
SIGNAL N111497722 : std_logic;
SIGNAL COONETEST3 : std_logic;
SIGNAL N110678329 : std_logic;
SIGNAL N112202422 : std_logic;
SIGNAL N06039 : std_logic;
SIGNAL N112080917 : std_logic;
SIGNAL N110577333 : std_logic;
SIGNAL N80958 : std_logic;
SIGNAL N110985127 : std_logic;
SIGNAL N110601623 : std_logic;
SIGNAL N78515 : std_logic;
SIGNAL N110985116 : std_logic;
SIGNAL N111667830 : std_logic;
SIGNAL N110856011 : std_logic;
SIGNAL N112153829 : std_logic;
SIGNAL N1146805 : std_logic;
SIGNAL N112153820 : std_logic;
SIGNAL N1146849 : std_logic;
SIGNAL N113729325 : std_logic;
SIGNAL N110266726 : std_logic;
SIGNAL N1058486 : std_logic;
SIGNAL SGTEST2 : std_logic;
SIGNAL N112712726 : std_logic;
SIGNAL N110524920 : std_logic;
SIGNAL N91228 : std_logic;
SIGNAL N112518319 : std_logic;
SIGNAL N112615524 : std_logic;
SIGNAL N94143 : std_logic;
SIGNAL N112518316 : std_logic;
SIGNAL N112591225 : std_logic;
SIGNAL N81781 : std_logic;
SIGNAL N110985126 : std_logic;
SIGNAL N111862229 : std_logic;
SIGNAL N79336 : std_logic;
SIGNAL N110960828 : std_logic;
SIGNAL N111424822 : std_logic;
SIGNAL SGTEST3 : std_logic;
SIGNAL N111449118 : std_logic;
SIGNAL N110678324 : std_logic;
SIGNAL MONITOR1 : std_logic;
SIGNAL N11054929 : std_logic;
SIGNAL N112712725 : std_logic;
SIGNAL N110779311 : std_logic;
SIGNAL N110985125 : std_logic;
SIGNAL N1147167 : std_logic;
SIGNAL N110932722 : std_logic;
SIGNAL N111449133 : std_logic;
SIGNAL N1147147 : std_logic;
SIGNAL N110625923 : std_logic;
SIGNAL N110625920 : std_logic;
SIGNAL N1147171 : std_logic;
SIGNAL N1147111 : std_logic;
SIGNAL N110266711 : std_logic;
SIGNAL N84232 : std_logic;
SIGNAL N111959426 : std_logic;
SIGNAL N111935119 : std_logic;
SIGNAL N84234 : std_logic;
SIGNAL N111935122 : std_logic;
SIGNAL N111009431 : std_logic;
SIGNAL COONETEST7 : std_logic;
SIGNAL N112372516 : std_logic;
SIGNAL N111009417 : std_logic;
SIGNAL N93240 : std_logic;
SIGNAL N110347227 : std_logic;
SIGNAL N110472512 : std_logic;
SIGNAL N80976 : std_logic;
SIGNAL N110347218 : std_logic;
SIGNAL N112542629 : std_logic;
SIGNAL N111037516 : std_logic;
SIGNAL N112445425 : std_logic;
SIGNAL N1146821 : std_logic;
SIGNAL N91242 : std_logic;
SIGNAL N111009418 : std_logic;
SIGNAL N112153822 : std_logic;
SIGNAL N91252 : std_logic;
SIGNAL N112032318 : std_logic;
SIGNAL N111594923 : std_logic;
SIGNAL N110472515 : std_logic;
SIGNAL N111594921 : std_logic;
SIGNAL N1058172 : std_logic;
SIGNAL N110625933 : std_logic;
SIGNAL N11047258 : std_logic;
SIGNAL N112251017 : std_logic;
SIGNAL N110625917 : std_logic;
SIGNAL N111594927 : std_logic;
SIGNAL N111765028 : std_logic;
SIGNAL N111497731 : std_logic;
SIGNAL N111594918 : std_logic;
SIGNAL N111361031 : std_logic;
SIGNAL N111497726 : std_logic;
SIGNAL N112566933 : std_logic;
SIGNAL N111361017 : std_logic;
SIGNAL N111497717 : std_logic;
SIGNAL N112566916 : std_logic;
SIGNAL N112080928 : std_logic;
SIGNAL N111086113 : std_logic;
SIGNAL N112542617 : std_logic;
SIGNAL N112785629 : std_logic;
SIGNAL N112202431 : std_logic;
SIGNAL N111935123 : std_logic;
SIGNAL N110319129 : std_logic;
SIGNAL N112396831 : std_logic;
SIGNAL N11077933 : std_logic;
SIGNAL N110319115 : std_logic;
SIGNAL N112396824 : std_logic;
SIGNAL N11116283 : std_logic;
SIGNAL N111138520 : std_logic;
SIGNAL N112396817 : std_logic;
SIGNAL N112445420 : std_logic;
SIGNAL N110577331 : std_logic;
SIGNAL N112372525 : std_logic;
SIGNAL N111910829 : std_logic;
SIGNAL N110577324 : std_logic;
SIGNAL N111497725 : std_logic;
SIGNAL N111910822 : std_logic;
SIGNAL N111643533 : std_logic;
SIGNAL N110755024 : std_logic;
SIGNAL N110625913 : std_logic;
SIGNAL N112469728 : std_logic;
SIGNAL N113729329 : std_logic;
SIGNAL N110831733 : std_logic;
SIGNAL N112469719 : std_logic;
SIGNAL N113729324 : std_logic;
SIGNAL N110831717 : std_logic;
SIGNAL N110266728 : std_logic;
SIGNAL N11039581 : std_logic;
SIGNAL N110831725 : std_logic;
SIGNAL N11026675 : std_logic;
SIGNAL N110524927 : std_logic;
SIGNAL N111692133 : std_logic;
SIGNAL N111449130 : std_logic;
SIGNAL N110524922 : std_logic;
SIGNAL N112153825 : std_logic;
SIGNAL N110730716 : std_logic;
SIGNAL N110500627 : std_logic;
SIGNAL N112251018 : std_logic;
SIGNAL N112421122 : std_logic;
SIGNAL N111765021 : std_logic;
SIGNAL N111765029 : std_logic;
SIGNAL N111263830 : std_logic;
SIGNAL N111740721 : std_logic;
SIGNAL N111336733 : std_logic;
SIGNAL N111215224 : std_logic;
SIGNAL N110601627 : std_logic;
SIGNAL N111361018 : std_logic;
SIGNAL N111910828 : std_logic;
SIGNAL N110577326 : std_logic;
SIGNAL N111336717 : std_logic;
SIGNAL N111162823 : std_logic;
SIGNAL N110577317 : std_logic;
SIGNAL N110856032 : std_logic;
SIGNAL N111162816 : std_logic;
SIGNAL N110678319 : std_logic;
SIGNAL N11085605 : std_logic;
SIGNAL N110423920 : std_logic;
SIGNAL N110654024 : std_logic;
SIGNAL N112105222 : std_logic;
SIGNAL N111361028 : std_logic;
SIGNAL N111643531 : std_logic;
SIGNAL N112080929 : std_logic;
SIGNAL N11070269 : std_logic;
SIGNAL N111643524 : std_logic;
SIGNAL N112323929 : std_logic;
SIGNAL N111692117 : std_logic;
SIGNAL N111643518 : std_logic;
SIGNAL N112737031 : std_logic;
SIGNAL N110549221 : std_logic;
SIGNAL N111138531 : std_logic;
SIGNAL N112737024 : std_logic;
SIGNAL N11031915 : std_logic;
SIGNAL N111138522 : std_logic;
SIGNAL N112712718 : std_logic;
SIGNAL N110395820 : std_logic;
SIGNAL N111138517 : std_logic;
SIGNAL N112785630 : std_logic;
SIGNAL N112737023 : std_logic;
SIGNAL N112178122 : std_logic;
SIGNAL N11108617 : std_logic;
SIGNAL N112421127 : std_logic;
SIGNAL N112178117 : std_logic;
SIGNAL N110319130 : std_logic;
SIGNAL N111837927 : std_logic;
SIGNAL N112153824 : std_logic;
SIGNAL N110319116 : std_logic;
SIGNAL N111837918 : std_logic;
SIGNAL N112761327 : std_logic;
SIGNAL N111862219 : std_logic;
SIGNAL N110932729 : std_logic;
SIGNAL N112615521 : std_logic;
SIGNAL N111138523 : std_logic;
SIGNAL N11093279 : std_logic;
SIGNAL N111336728 : std_logic;
SIGNAL N111138518 : std_logic;
SIGNAL N110625925 : std_logic;
SIGNAL N111336724 : std_logic;
SIGNAL N112032319 : std_logic;
SIGNAL N111522023 : std_logic;
SIGNAL N110601626 : std_logic;
SIGNAL N111546324 : std_logic;
SIGNAL N111497720 : std_logic;
SIGNAL N110601618 : std_logic;
SIGNAL N107162014 : std_logic;
SIGNAL N110755021 : std_logic;
SIGNAL N110702618 : std_logic;
SIGNAL N110908419 : std_logic;
SIGNAL N110395823 : std_logic;
SIGNAL N111740730 : std_logic;
SIGNAL N112299625 : std_logic;
SIGNAL N111114224 : std_logic;
SIGNAL N111716424 : std_logic;
SIGNAL N111813625 : std_logic;
SIGNAL N111086118 : std_logic;
SIGNAL N112494024 : std_logic;
SIGNAL N111789327 : std_logic;
SIGNAL N112202424 : std_logic;
SIGNAL N111114217 : std_logic;
SIGNAL N110807430 : std_logic;
SIGNAL N111086126 : std_logic;
SIGNAL N112469729 : std_logic;
SIGNAL N110807423 : std_logic;
SIGNAL N110266723 : std_logic;
SIGNAL N112469720 : std_logic;
SIGNAL N111862224 : std_logic;
SIGNAL N110524924 : std_logic;
SIGNAL N110266720 : std_logic;
SIGNAL N110884133 : std_logic;
SIGNAL N112202417 : std_logic;
SIGNAL N11026676 : std_logic;
SIGNAL N111424824 : std_logic;
SIGNAL N112178118 : std_logic;
SIGNAL N112323917 : std_logic;
SIGNAL N112615530 : std_logic;
SIGNAL N112299630 : std_logic;
SIGNAL N11077935 : std_logic;
SIGNAL N112615519 : std_logic;
SIGNAL N111009415 : std_logic;
SIGNAL N110932721 : std_logic;
SIGNAL N112591227 : std_logic;
SIGNAL N111449131 : std_logic;
SIGNAL N110625922 : std_logic;
SIGNAL N111886526 : std_logic;
SIGNAL N111449117 : std_logic;
SIGNAL N112348217 : std_logic;
SIGNAL N111886517 : std_logic;
SIGNAL N110730717 : std_logic;
SIGNAL N11047257 : std_logic;
SIGNAL N110884130 : std_logic;
SIGNAL N111263831 : std_logic;
SIGNAL N110500621 : std_logic;
SIGNAL N110856025 : std_logic;
SIGNAL N111263817 : std_logic;
SIGNAL N111619222 : std_logic;
SIGNAL N110856018 : std_logic;
SIGNAL N110347217 : std_logic;
SIGNAL N112542631 : std_logic;
SIGNAL N112275330 : std_logic;
SIGNAL N110319124 : std_logic;
SIGNAL N110779326 : std_logic;
SIGNAL N112251031 : std_logic;
SIGNAL N111215225 : std_logic;
SIGNAL N11077932 : std_logic;
SIGNAL N112251019 : std_logic;
SIGNAL N111190917 : std_logic;
SIGNAL N112445427 : std_logic;
SIGNAL N111424829 : std_logic;
SIGNAL N111886529 : std_logic;
SIGNAL N111910821 : std_logic;
SIGNAL N111424817 : std_logic;
SIGNAL N111037531 : std_logic;
SIGNAL N11093272 : std_logic;
SIGNAL N110678328 : std_logic;
SIGNAL N11039587 : std_logic;
SIGNAL N112153831 : std_logic;
SIGNAL N112080921 : std_logic;
SIGNAL N11039580 : std_logic;
SIGNAL N111765023 : std_logic;
SIGNAL N111619230 : std_logic;
SIGNAL N111162826 : std_logic;
SIGNAL N111361021 : std_logic;
SIGNAL N111619220 : std_logic;
SIGNAL N110702632 : std_logic;
SIGNAL N112737030 : std_logic;
SIGNAL N110985119 : std_logic;
SIGNAL N112566926 : std_logic;
SIGNAL N112785624 : std_logic;
SIGNAL N110856014 : std_logic;
SIGNAL N110423921 : std_logic;
SIGNAL N112542624 : std_logic;
SIGNAL N111361024 : std_logic;
SIGNAL N110319119 : std_logic;
SIGNAL N110702612 : std_logic;
SIGNAL N110908430 : std_logic;
SIGNAL N11070262 : std_logic;
SIGNAL N112664118 : std_logic;
SIGNAL N113729328 : std_logic;
SIGNAL N111692127 : std_logic;
SIGNAL N112445416 : std_logic;
SIGNAL N113729319 : std_logic;
SIGNAL N111692118 : std_logic;
SIGNAL N110266714 : std_logic;
SIGNAL N112712733 : std_logic;
SIGNAL N110549222 : std_logic;
SIGNAL N11026679 : std_logic;
SIGNAL N110985129 : std_logic;
SIGNAL N11054928 : std_logic;
SIGNAL N11026670 : std_logic;
SIGNAL N110960831 : std_logic;
SIGNAL N11031918 : std_logic;
SIGNAL N112299616 : std_logic;
SIGNAL N111424826 : std_logic;
SIGNAL N110395830 : std_logic;
SIGNAL N111009424 : std_logic;
SIGNAL N110779314 : std_logic;
SIGNAL N112737019 : std_logic;
SIGNAL N110755026 : std_logic;
SIGNAL N110932733 : std_logic;
SIGNAL N112664126 : std_logic;
SIGNAL N112421124 : std_logic;
SIGNAL N110932731 : std_logic;
SIGNAL N112421128 : std_logic;
SIGNAL N111263825 : std_logic;
SIGNAL N110625927 : std_logic;
SIGNAL N111837928 : std_logic;
SIGNAL N111190928 : std_logic;
SIGNAL N110625910 : std_logic;
SIGNAL N111837919 : std_logic;
SIGNAL N111061818 : std_logic;
SIGNAL N11062591 : std_logic;
SIGNAL N110932730 : std_logic;
SIGNAL N11039586 : std_logic;
SIGNAL N11026673 : std_logic;
SIGNAL N110932714 : std_logic;
SIGNAL N112591221 : std_logic;
SIGNAL N112494031 : std_logic;
SIGNAL N110625926 : std_logic;
SIGNAL N111361023 : std_logic;
SIGNAL N112469730 : std_logic;
SIGNAL N111522024 : std_logic;
SIGNAL N110448227 : std_logic;
SIGNAL N112469723 : std_logic;
SIGNAL N107162011 : std_logic;
SIGNAL N110448218 : std_logic;
SIGNAL N111983726 : std_logic;
SIGNAL N10716206 : std_logic;
SIGNAL N11070261 : std_logic;
SIGNAL N111983718 : std_logic;
SIGNAL N111086133 : std_logic;
SIGNAL N111789316 : std_logic;
SIGNAL N111959423 : std_logic;
SIGNAL N111086129 : std_logic;
SIGNAL N11031917 : std_logic;
SIGNAL N111959416 : std_logic;
SIGNAL N111086124 : std_logic;
SIGNAL N112664120 : std_logic;
SIGNAL N112372533 : std_logic;
SIGNAL N11108616 : std_logic;
SIGNAL N110932713 : std_logic;
SIGNAL N112372519 : std_logic;
SIGNAL N112202418 : std_logic;
SIGNAL N111522027 : std_logic;
SIGNAL N112348226 : std_logic;
SIGNAL N112372523 : std_logic;
SIGNAL N111522018 : std_logic;
SIGNAL N112348216 : std_logic;
SIGNAL N111497733 : std_logic;
SIGNAL N111497729 : std_logic;
SIGNAL N112105219 : std_logic;
SIGNAL N110755027 : std_logic;
SIGNAL N10716200 : std_logic;
SIGNAL N111473429 : std_logic;
SIGNAL N113729317 : std_logic;
SIGNAL N11108615 : std_logic;
SIGNAL N110347230 : std_logic;
SIGNAL N112785621 : std_logic;
SIGNAL N112372522 : std_logic;
SIGNAL N110347221 : std_logic;
SIGNAL N110395833 : std_logic;
SIGNAL N110500619 : std_logic;
SIGNAL N111037519 : std_logic;
SIGNAL N110395824 : std_logic;
SIGNAL N111740724 : std_logic;
SIGNAL N111009421 : std_logic;
SIGNAL N110395810 : std_logic;
SIGNAL N112178120 : std_logic;
SIGNAL N112032330 : std_logic;
SIGNAL N111765024 : std_logic;
SIGNAL N112761321 : std_logic;
SIGNAL N112032321 : std_logic;
SIGNAL N110601628 : std_logic;
SIGNAL N112518328 : std_logic;
SIGNAL N110500630 : std_logic;
SIGNAL N110601619 : std_logic;
SIGNAL N112494027 : std_logic;
SIGNAL N110500616 : std_logic;
SIGNAL N111667820 : std_logic;
SIGNAL N111114226 : std_logic;
SIGNAL N110472525 : std_logic;
SIGNAL N111114216 : std_logic;
SIGNAL N111086120 : std_logic;
SIGNAL N113753628 : std_logic;
SIGNAL N110472518 : std_logic;
SIGNAL N112178131 : std_logic;
SIGNAL N111263823 : std_logic;
SIGNAL N113753619 : std_logic;
SIGNAL N111619228 : std_logic;
SIGNAL N112761322 : std_logic;
SIGNAL N112178127 : std_logic;
SIGNAL N113753626 : std_logic;
SIGNAL N111594930 : std_logic;
SIGNAL N11116288 : std_logic;
SIGNAL N110807425 : std_logic;
SIGNAL N113753630 : std_logic;
SIGNAL N111837929 : std_logic;
SIGNAL N110601616 : std_logic;
SIGNAL N112251028 : std_logic;
SIGNAL N113753621 : std_logic;
SIGNAL N111813618 : std_logic;
SIGNAL N110702631 : std_logic;
SIGNAL N111716429 : std_logic;
SIGNAL N113753627 : std_logic;
SIGNAL N110472531 : std_logic;
SIGNAL N111716416 : std_logic;
SIGNAL N111716417 : std_logic;
SIGNAL N113753623 : std_logic;
SIGNAL N110472514 : std_logic;
SIGNAL N112518329 : std_logic;
SIGNAL N11085600 : std_logic;
SIGNAL N113753633 : std_logic;
SIGNAL N11047255 : std_logic;
SIGNAL N111114227 : std_logic;
SIGNAL N113729322 : std_logic;
SIGNAL N113753620 : std_logic;
SIGNAL N111935126 : std_logic;
SIGNAL N111086121 : std_logic;
SIGNAL N110347224 : std_logic;
SIGNAL N113753625 : std_logic;
SIGNAL N111215216 : std_logic;
SIGNAL N111086116 : std_logic;
SIGNAL N112542626 : std_logic;
SIGNAL N113753617 : std_logic;
SIGNAL N110779318 : std_logic;
SIGNAL N110266716 : std_logic;
SIGNAL N111935130 : std_logic;
SIGNAL N113753624 : std_logic;
SIGNAL N11077937 : std_logic;
SIGNAL N110524916 : std_logic;
SIGNAL N111162814 : std_logic;
SIGNAL N113753629 : std_logic;
SIGNAL N11077930 : std_logic;
SIGNAL N112202427 : std_logic;
SIGNAL N11116284 : std_logic;
SIGNAL N113753616 : std_logic;
SIGNAL N111162818 : std_logic;
SIGNAL N112178128 : std_logic;
SIGNAL N111910830 : std_logic;
SIGNAL N113753618 : std_logic;
SIGNAL N11116280 : std_logic;
SIGNAL N112178121 : std_logic;
SIGNAL N111910823 : std_logic;
SIGNAL N113753622 : std_logic;
SIGNAL N112445417 : std_logic;
SIGNAL N112178116 : std_logic;
SIGNAL N111570621 : std_logic;
SIGNAL N113753631 : std_logic;
SIGNAL N111910816 : std_logic;
SIGNAL N112615529 : std_logic;
SIGNAL N110831728 : std_logic;
SIGNAL N110625932 : std_logic;
SIGNAL N112591216 : std_logic;
SIGNAL N112153833 : std_logic;
SIGNAL N110831720 : std_logic;
SIGNAL N110807426 : std_logic;
SIGNAL N112737025 : std_logic;
SIGNAL N110807420 : std_logic;
SIGNAL N110807416 : std_logic;
SIGNAL N107162032 : std_logic;
SIGNAL N111692123 : std_logic;
SIGNAL N110779316 : std_logic;
SIGNAL N110908425 : std_logic;
SIGNAL N111570627 : std_logic;
SIGNAL N111862225 : std_logic;
SIGNAL N111215226 : std_logic;
SIGNAL N112251030 : std_logic;
SIGNAL N111862220 : std_logic;
SIGNAL N111190923 : std_logic;
SIGNAL N112251021 : std_logic;
SIGNAL N112275323 : std_logic;
SIGNAL N110702624 : std_logic;
SIGNAL N111336720 : std_logic;
SIGNAL N112251022 : std_logic;
SIGNAL N110549228 : std_logic;
SIGNAL N110856021 : std_logic;
SIGNAL N112080919 : std_logic;
SIGNAL N110549214 : std_logic;
SIGNAL N11085607 : std_logic;
SIGNAL N111619223 : std_logic;
SIGNAL N111789323 : std_logic;
SIGNAL N11085603 : std_logic;
SIGNAL N111716430 : std_logic;
SIGNAL N111061822 : std_logic;
SIGNAL N112105231 : std_logic;
SIGNAL N111716418 : std_logic;
SIGNAL N110423922 : std_logic;
SIGNAL N112105224 : std_logic;
SIGNAL N110985122 : std_logic;
SIGNAL N112372524 : std_logic;
SIGNAL N112712727 : std_logic;
SIGNAL N110856015 : std_logic;
SIGNAL N110755028 : std_logic;
SIGNAL N112785633 : std_logic;
SIGNAL N11085606 : std_logic;
SIGNAL N110524931 : std_logic;
SIGNAL N112761318 : std_logic;
SIGNAL N111765025 : std_logic;
SIGNAL N112542633 : std_logic;
SIGNAL N112712730 : std_logic;
SIGNAL N110678317 : std_logic;
SIGNAL N112542616 : std_logic;
SIGNAL N112712721 : std_logic;
SIGNAL N111983723 : std_logic;
SIGNAL N110985121 : std_logic;
SIGNAL N112761323 : std_logic;
SIGNAL N111086110 : std_logic;
SIGNAL N110960823 : std_logic;
SIGNAL N111336718 : std_logic;
SIGNAL N110319133 : std_logic;
SIGNAL N111449125 : std_logic;
SIGNAL N112518323 : std_logic;
SIGNAL N11031912 : std_logic;
SIGNAL N11077936 : std_logic;
SIGNAL N112494022 : std_logic;
SIGNAL N111862216 : std_logic;
SIGNAL N110960825 : std_logic;
SIGNAL N111862231 : std_logic;
SIGNAL N112032323 : std_logic;
SIGNAL N110932724 : std_logic;
SIGNAL N112251023 : std_logic;
SIGNAL N111546327 : std_logic;
SIGNAL N11062590 : std_logic;
SIGNAL N112080930 : std_logic;
SIGNAL N111546318 : std_logic;
SIGNAL N111983721 : std_logic;
SIGNAL N112080920 : std_logic;
SIGNAL N110577321 : std_logic;
SIGNAL N111983716 : std_logic;
SIGNAL N111619224 : std_logic;
SIGNAL N110549225 : std_logic;
SIGNAL N111935124 : std_logic;
SIGNAL N110856012 : std_logic;
SIGNAL N10716201 : std_logic;
SIGNAL N112348233 : std_logic;
SIGNAL N112518325 : std_logic;
SIGNAL N110908422 : std_logic;
SIGNAL N112372528 : std_logic;
SIGNAL N11026677 : std_logic;
SIGNAL N112299628 : std_logic;
SIGNAL N112348227 : std_logic;
SIGNAL N111619226 : std_logic;
SIGNAL N112275327 : std_logic;
SIGNAL N112348218 : std_logic;
SIGNAL N111570633 : std_logic;
SIGNAL N111813628 : std_logic;
SIGNAL N112105228 : std_logic;
SIGNAL N112785631 : std_logic;
SIGNAL N112445433 : std_logic;
SIGNAL N111037528 : std_logic;
SIGNAL N110319131 : std_logic;
SIGNAL N112445422 : std_logic;
SIGNAL N112032322 : std_logic;
SIGNAL N111862226 : std_logic;
SIGNAL N110266732 : std_logic;
SIGNAL N110472510 : std_logic;
SIGNAL N10716207 : std_logic;
SIGNAL N112323926 : std_logic;
SIGNAL N110500622 : std_logic;
SIGNAL N111813626 : std_logic;
SIGNAL N112299627 : std_logic;
SIGNAL N112566925 : std_logic;
SIGNAL N112664122 : std_logic;
SIGNAL N112299620 : std_logic;
SIGNAL N112566918 : std_logic;
SIGNAL N112469721 : std_logic;
SIGNAL N11100942 : std_logic;
SIGNAL N112542619 : std_logic;
SIGNAL N110266721 : std_logic;
SIGNAL N111473427 : std_logic;
SIGNAL N110472523 : std_logic;
SIGNAL N112323920 : std_logic;
SIGNAL N111473418 : std_logic;
SIGNAL N110779327 : std_logic;
SIGNAL N110730718 : std_logic;
SIGNAL N111449120 : std_logic;
SIGNAL N110779315 : std_logic;
SIGNAL N111215230 : std_logic;
SIGNAL N110730729 : std_logic;
SIGNAL N110779312 : std_logic;
SIGNAL N111037533 : std_logic;
SIGNAL N110730720 : std_logic;
SIGNAL N111162815 : std_logic;
SIGNAL N111692128 : std_logic;
SIGNAL N112421129 : std_logic;
SIGNAL N11116285 : std_logic;
SIGNAL N111692119 : std_logic;
SIGNAL N112421117 : std_logic;
SIGNAL N111910831 : std_logic;
SIGNAL N110549223 : std_logic;
SIGNAL N112396825 : std_logic;
SIGNAL N111910824 : std_logic;
SIGNAL N112348219 : std_logic;
SIGNAL N112396820 : std_logic;
SIGNAL N11062598 : std_logic;
SIGNAL N111837920 : std_logic;
SIGNAL N111263820 : std_logic;
SIGNAL N111570618 : std_logic;
SIGNAL N112372529 : std_logic;
SIGNAL N110347233 : std_logic;
SIGNAL N11093273 : std_logic;
SIGNAL N110395825 : std_logic;
SIGNAL N110319123 : std_logic;
SIGNAL N112153817 : std_logic;
SIGNAL N110500623 : std_logic;
SIGNAL N111215219 : std_logic;
SIGNAL N111594931 : std_logic;
SIGNAL N111190920 : std_logic;
SIGNAL N111594924 : std_logic;
SIGNAL N111886533 : std_logic;
SIGNAL N111570617 : std_logic;
SIGNAL N110654020 : std_logic;
SIGNAL N111910827 : std_logic;
SIGNAL N111361022 : std_logic;
SIGNAL N111336730 : std_logic;
SIGNAL N111910818 : std_logic;
SIGNAL N111336729 : std_logic;
SIGNAL N110702626 : std_logic;
SIGNAL N111886521 : std_logic;
SIGNAL N112080924 : std_logic;
SIGNAL N112615517 : std_logic;
SIGNAL N11039584 : std_logic;
SIGNAL N112323924 : std_logic;
SIGNAL N110779328 : std_logic;
SIGNAL N110884127 : std_logic;
SIGNAL N112737033 : std_logic;
SIGNAL N110985117 : std_logic;
SIGNAL N110884120 : std_logic;
SIGNAL N112737026 : std_logic;
SIGNAL N111935133 : std_logic;
SIGNAL N111162820 : std_logic;
SIGNAL N112712720 : std_logic;
SIGNAL N112105229 : std_logic;
SIGNAL N110702611 : std_logic;
SIGNAL N112785625 : std_logic;
SIGNAL N11093274 : std_logic;
SIGNAL N112566929 : std_logic;
SIGNAL N112785620 : std_logic;
SIGNAL N110831730 : std_logic;
SIGNAL N110448229 : std_logic;
SIGNAL N110319125 : std_logic;
SIGNAL N111570623 : std_logic;
SIGNAL N110423929 : std_logic;
SIGNAL N110319120 : std_logic;
SIGNAL N112785626 : std_logic;
SIGNAL N110423924 : std_logic;
SIGNAL N111862221 : std_logic;
SIGNAL N110319121 : std_logic;
SIGNAL N111009412 : std_logic;
SIGNAL N111138525 : std_logic;
SIGNAL N111190930 : std_logic;
SIGNAL N110448219 : std_logic;
SIGNAL N111643529 : std_logic;
SIGNAL N111061824 : std_logic;
SIGNAL N110702621 : std_logic;
SIGNAL N110908431 : std_logic;
SIGNAL N110423933 : std_logic;
SIGNAL N111692130 : std_logic;
SIGNAL N112275322 : std_logic;
SIGNAL N111692121 : std_logic;
SIGNAL N111789331 : std_logic;
SIGNAL N111522029 : std_logic;
SIGNAL N110549211 : std_logic;
SIGNAL N111789322 : std_logic;
SIGNAL N11108611 : std_logic;
SIGNAL N111789326 : std_logic;
SIGNAL N112664121 : std_logic;
SIGNAL N111740726 : std_logic;
SIGNAL N111789321 : std_logic;
SIGNAL N112469724 : std_logic;
SIGNAL N112518317 : std_logic;
SIGNAL N111061819 : std_logic;
SIGNAL N110266715 : std_logic;
SIGNAL N112494029 : std_logic;
SIGNAL TG5 : std_logic;
SIGNAL N110319112 : std_logic;
SIGNAL N110266710 : std_logic;
SIGNAL TG6 : std_logic;
SIGNAL N110395829 : std_logic;
SIGNAL N11026671 : std_logic;
SIGNAL N112737027 : std_logic;
SIGNAL N112323919 : std_logic;
SIGNAL N1056495 : std_logic;
SIGNAL TG0 : std_logic;
SIGNAL N112664129 : std_logic;
SIGNAL N112323916 : std_logic;
SIGNAL TG14 : std_logic;
SIGNAL N112348223 : std_logic;
SIGNAL N111009432 : std_logic;
SIGNAL TG15 : std_logic;
SIGNAL N111837931 : std_logic;
SIGNAL N111449126 : std_logic;
SIGNAL N109348 : std_logic;
SIGNAL N111837922 : std_logic;
SIGNAL N111263826 : std_logic;
SIGNAL N110932711 : std_logic;
SIGNAL N110347226 : std_logic;
SIGNAL N1260508 : std_logic;
SIGNAL N11093276 : std_logic;
SIGNAL N110347219 : std_logic;
SIGNAL N1263850 : std_logic;
SIGNAL N111546330 : std_logic;
SIGNAL N110319126 : std_logic;
SIGNAL N1267774 : std_logic;
SIGNAL TG1 : std_logic;
SIGNAL N111522031 : std_logic;
SIGNAL N111190929 : std_logic;
SIGNAL TG3 : std_logic;
SIGNAL N111522020 : std_logic;
SIGNAL N111886531 : std_logic;
SIGNAL TG12 : std_logic;
SIGNAL N110654027 : std_logic;
SIGNAL N111886524 : std_logic;
SIGNAL N110625929 : std_logic;
SIGNAL N11039589 : std_logic;
SIGNAL N1256014 : std_logic;
SIGNAL N108996 : std_logic;
SIGNAL N111497721 : std_logic;
SIGNAL N110908427 : std_logic;
SIGNAL N10716209 : std_logic;
SIGNAL N110908426 : std_logic;
SIGNAL N1262264 : std_logic;
SIGNAL TG8 : std_logic;
SIGNAL N111086127 : std_logic;
SIGNAL N110702613 : std_logic;
SIGNAL N109008 : std_logic;
SIGNAL N111086115 : std_logic;
SIGNAL N110448222 : std_logic;
SIGNAL N109324 : std_logic;
SIGNAL N112202426 : std_logic;
SIGNAL N110423916 : std_logic;
SIGNAL N112202421 : std_logic;
SIGNAL N111361026 : std_logic;
SIGNAL N1251498 : std_logic;
SIGNAL N112396826 : std_logic;
SIGNAL N11100947 : std_logic;
SIGNAL N1254680 : std_logic;
SIGNAL TG7 : std_logic;
SIGNAL N111497727 : std_logic;
SIGNAL N110448228 : std_logic;
SIGNAL N108992 : std_logic;
SIGNAL N113729331 : std_logic;
SIGNAL N110702633 : std_logic;
SIGNAL N109352 : std_logic;
SIGNAL N113729326 : std_logic;
SIGNAL N110702630 : std_logic;
SIGNAL TG9 : std_logic;
SIGNAL N110395827 : std_logic;
SIGNAL N110702614 : std_logic;
SIGNAL TG2 : std_logic;
SIGNAL N110395822 : std_logic;
SIGNAL N11070264 : std_logic;
SIGNAL TG10 : std_logic;
SIGNAL N110524933 : std_logic;
SIGNAL N111667819 : std_logic;
SIGNAL N109356 : std_logic;
SIGNAL N110524929 : std_logic;
SIGNAL N111789324 : std_logic;
SIGNAL N109340 : std_logic;
SIGNAL N110500629 : std_logic;
SIGNAL N111061828 : std_logic;
SIGNAL N111765033 : std_logic;
SIGNAL N110319110 : std_logic;
SIGNAL N1258106 : std_logic;
SIGNAL N110601631 : std_logic;
SIGNAL N110423923 : std_logic;
SIGNAL N1250090 : std_logic;
SIGNAL TG4 : std_logic;
SIGNAL N110601622 : std_logic;
SIGNAL N112348228 : std_logic;
SIGNAL TG11 : std_logic;
SIGNAL N110678331 : std_logic;
SIGNAL N110932725 : std_logic;
SIGNAL N109004 : std_logic;
SIGNAL N111667827 : std_logic;
SIGNAL N111546323 : std_logic;
SIGNAL N111643526 : std_logic;
SIGNAL N110654019 : std_logic;
SIGNAL N1257374 : std_logic;
SIGNAL N111114228 : std_logic;
SIGNAL N111522028 : std_logic;
SIGNAL N1261526 : std_logic;
SIGNAL N111114219 : std_logic;
SIGNAL N111522019 : std_logic;
SIGNAL N1244642 : std_logic;
SIGNAL N112153819 : std_logic;
SIGNAL N107162015 : std_logic;
SIGNAL N1263768 : std_logic;
SIGNAL N81767 : std_logic;
SIGNAL N112761329 : std_logic;
SIGNAL N11108618 : std_logic;
SIGNAL N1248836 : std_logic;
SIGNAL N112761324 : std_logic;
SIGNAL N112396819 : std_logic;
SIGNAL N1265342 : std_logic;
SIGNAL A4 : std_logic;
SIGNAL N109344 : std_logic;
SIGNAL N111162832 : std_logic;
SIGNAL N110755029 : std_logic;
SIGNAL B0 : std_logic;
SIGNAL N109332 : std_logic;
SIGNAL N111162811 : std_logic;
SIGNAL N110395814 : std_logic;
SIGNAL B3 : std_logic;
SIGNAL N109328 : std_logic;
SIGNAL N11116282 : std_logic;
SIGNAL N110500633 : std_logic;
SIGNAL B14 : std_logic;
SIGNAL TG13 : std_logic;
SIGNAL N111336726 : std_logic;
SIGNAL N110524917 : std_logic;
SIGNAL E7 : std_logic;
SIGNAL F7 : std_logic;
SIGNAL N109336 : std_logic;
SIGNAL N110601630 : std_logic;
SIGNAL N111765026 : std_logic;
SIGNAL F13 : std_logic;
SIGNAL N109016 : std_logic;
SIGNAL N110601620 : std_logic;
SIGNAL N111740725 : std_logic;
SIGNAL N110702620 : std_logic;
SIGNAL N111740716 : std_logic;
SIGNAL N1268390 : std_logic;
SIGNAL CHECK7 : std_logic;
SIGNAL N111716433 : std_logic;
SIGNAL N110654026 : std_logic;
SIGNAL N1257164 : std_logic;
SIGNAL N80145 : std_logic;
SIGNAL N109000 : std_logic;
SIGNAL N111716419 : std_logic;
SIGNAL N110654016 : std_logic;
SIGNAL N80151 : std_logic;
SIGNAL N109012 : std_logic;
SIGNAL N112494019 : std_logic;
SIGNAL N111667822 : std_logic;
SIGNAL N79328 : std_logic;
SIGNAL N110266730 : std_logic;
SIGNAL N111643516 : std_logic;
SIGNAL N1147622 : std_logic;
SIGNAL N79340 : std_logic;
SIGNAL TF5 : std_logic;
SIGNAL N110524919 : std_logic;
SIGNAL N111138526 : std_logic;
SIGNAL N79344 : std_logic;
SIGNAL N1257378 : std_logic;
SIGNAL N108278 : std_logic;
SIGNAL N112202419 : std_logic;
SIGNAL N112178126 : std_logic;
SIGNAL N1147433 : std_logic;
SIGNAL N107830 : std_logic;
SIGNAL N112591233 : std_logic;
SIGNAL N111336719 : std_logic;
SIGNAL N1147437 : std_logic;
SIGNAL N112591229 : std_logic;
SIGNAL N110702627 : std_logic;
SIGNAL N1147634 : std_logic;
SIGNAL N1057858 : std_logic;
SIGNAL TF6 : std_logic;
SIGNAL N112591222 : std_logic;
SIGNAL N110702625 : std_logic;
SIGNAL TF8 : std_logic;
SIGNAL F1 : std_logic;
SIGNAL N110807418 : std_logic;
SIGNAL N111716428 : std_logic;
SIGNAL N111862228 : std_logic;
SIGNAL N112518331 : std_logic;
SIGNAL N1147614 : std_logic;
SIGNAL N1145393 : std_logic;
SIGNAL TF15 : std_logic;
SIGNAL N110884125 : std_logic;
SIGNAL N112518324 : std_logic;
SIGNAL N1145373 : std_logic;
SIGNAL N108270 : std_logic;
SIGNAL N110884116 : std_logic;
SIGNAL N112494028 : std_logic;
SIGNAL N1145361 : std_logic;
SIGNAL TF0 : std_logic;
SIGNAL N110856027 : std_logic;
SIGNAL N111114229 : std_logic;
SIGNAL N77708 : std_logic;
SIGNAL TF2 : std_logic;
SIGNAL N110856020 : std_logic;
SIGNAL N111114222 : std_logic;
SIGNAL N77714 : std_logic;
SIGNAL N107810 : std_logic;
SIGNAL H1 : std_logic;
SIGNAL N112251033 : std_logic;
SIGNAL N111086128 : std_logic;
SIGNAL MONITOR15 : std_logic;
SIGNAL N112275317 : std_logic;
SIGNAL N111086123 : std_logic;
SIGNAL N1147654 : std_logic;
SIGNAL TF13 : std_logic;
SIGNAL G8 : std_logic;
SIGNAL N111424831 : std_logic;
SIGNAL N110524928 : std_logic;
SIGNAL N107822 : std_logic;
SIGNAL N111424819 : std_logic;
SIGNAL N112202429 : std_logic;
SIGNAL N1078497 : std_logic;
SIGNAL N108262 : std_logic;
SIGNAL N110678321 : std_logic;
SIGNAL N112178130 : std_logic;
SIGNAL A15 : std_logic;

-- GATE INSTANCES

BEGIN
VCC <= '1';
GND <= '0';
CT3<=N94157;
NCT0<=N94143;
NCT1<=N94145;
NCT2<=N94147;
NCT3<=N94149;
CT0<=N94151;
CT1<=N94153;
CT2<=N94155;
U45 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => N77694, 
	DCO1 => N77696, 
	DCO2 => N77698, 
	DCO3 => N77700, 
	DCO4 => N77702, 
	DCO5 => N77704, 
	DCO6 => N77706, 
	DCO7 => N77708, 
	DSG0 => N77710, 
	DSG1 => N77712, 
	DSG2 => N77714, 
	DSG3 => N77716, 
	DSG4 => N77718, 
	DSG5 => N77720, 
	DSG6 => N77722, 
	DSG7 => N77724, 
	ENABLE => ENABLE14, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => N75814, 
	QCO1 => N75820, 
	QCO2 => N75826, 
	QCO3 => N75832, 
	QCO4 => N75838, 
	QCO5 => N75844, 
	QCO6 => N75850, 
	QCO7 => N75856, 
	QSG0 => N75862, 
	QSG1 => N75868, 
	QSG2 => N75874, 
	QSG3 => N75880, 
	QSG4 => N75886, 
	QSG5 => N75892, 
	QSG6 => N75898, 
	QSG7 => N75904, 
	S0 => N11108610, 
	S1 => N11108611, 
	S2 => N11108612, 
	S3 => N11108613, 
	S4 => N11108614, 
	S5 => N11108615, 
	S6 => N11108616, 
	S7 => N11108617, 
	S8 => N11108618, 
	S9 => N11108619, 
	S10 => N111086110, 
	S11 => N111086111, 
	S12 => N111086112, 
	S13 => N111086113, 
	S14 => N111086114, 
	S15 => N111086115, 
	SIGNED => N111086132
);
U46 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => N75814, 
	DCO1 => N75820, 
	DCO2 => N75826, 
	DCO3 => N75832, 
	DCO4 => N75838, 
	DCO5 => N75844, 
	DCO6 => N75850, 
	DCO7 => N75856, 
	DSG0 => N75862, 
	DSG1 => N75868, 
	DSG2 => N75874, 
	DSG3 => N75880, 
	DSG4 => N75886, 
	DSG5 => N75892, 
	DSG6 => N75898, 
	DSG7 => N75904, 
	ENABLE => ENABLE15, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => QCO0, 
	QCO1 => QCO1, 
	QCO2 => QCO2, 
	QCO3 => QCO3, 
	QCO4 => QCO4, 
	QCO5 => QCO5, 
	QCO6 => QCO6, 
	QCO7 => QCO7, 
	QSG0 => QSG0, 
	QSG1 => QSG1, 
	QSG2 => QSG2, 
	QSG3 => QSG3, 
	QSG4 => QSG4, 
	QSG5 => QSG5, 
	QSG6 => QSG6, 
	QSG7 => QSG7, 
	S0 => N11116280, 
	S1 => N11116281, 
	S2 => N11116282, 
	S3 => N11116283, 
	S4 => N11116284, 
	S5 => N11116285, 
	S6 => N11116286, 
	S7 => N11116287, 
	S8 => N11116288, 
	S9 => N11116289, 
	S10 => N111162810, 
	S11 => N111162811, 
	S12 => N111162812, 
	S13 => N111162813, 
	S14 => N111162814, 
	S15 => N111162815, 
	SIGNED => N111162832
);
U47 : EIGHTBITREG	PORT MAP(
	CLK => CLK, 
	D0 => CHECK0, 
	D1 => CHECK1, 
	D2 => CHECK2, 
	D3 => CHECK3, 
	D4 => CHECK4, 
	D5 => CHECK5, 
	D6 => CHECK6, 
	D7 => CHECK7, 
	NPRESET => VCC, 
	NRESET => NRST, 
	Q0 => TOTAL0, 
	Q1 => TOTAL1, 
	Q2 => TOTAL2, 
	Q3 => TOTAL3, 
	Q4 => TOTAL4, 
	Q5 => TOTAL5, 
	Q6 => TOTAL6, 
	Q7 => TOTAL7
);
U48 : EIGHTBITREG	PORT MAP(
	CLK => CLK, 
	D0 => CHECK8, 
	D1 => CHECK9, 
	D2 => CHECK10, 
	D3 => CHECK11, 
	D4 => CHECK12, 
	D5 => CHECK13, 
	D6 => CHECK14, 
	D7 => CHECK15, 
	NPRESET => VCC, 
	NRESET => NRST, 
	Q0 => TOTAL8, 
	Q1 => TOTAL9, 
	Q2 => TOTAL10, 
	Q3 => TOTAL11, 
	Q4 => TOTAL12, 
	Q5 => TOTAL13, 
	Q6 => TOTAL14, 
	Q7 => TOTAL15
);
U180 : ADDERDELAY	PORT MAP(
	DIN0 => N112542616, 
	DIN1 => N112542617, 
	DIN2 => N112542618, 
	DIN3 => N112542619, 
	DIN4 => N112542620, 
	DIN5 => N112542621, 
	DIN6 => N112542622, 
	DIN7 => N112542623, 
	DIN8 => N112542624, 
	DIN9 => N112542625, 
	DIN10 => N112542626, 
	DIN11 => N112542627, 
	DIN12 => N112542628, 
	DIN13 => N112542629, 
	DIN14 => N112542630, 
	DIN15 => N112542631, 
	DOUT0 => N112566916, 
	DOUT1 => N112566917, 
	DOUT2 => N112566918, 
	DOUT3 => N112566919, 
	DOUT4 => N112566920, 
	DOUT5 => N112566921, 
	DOUT6 => N112566922, 
	DOUT7 => N112566923, 
	DOUT8 => N112566924, 
	DOUT9 => N112566925, 
	DOUT10 => N112566926, 
	DOUT11 => N112566927, 
	DOUT12 => N112566928, 
	DOUT13 => N112566929, 
	DOUT14 => N112566930, 
	DOUT15 => N112566931, 
	SIGNEDIN => N112542633, 
	SIGNEDOUT => N112566933
);
U181 : ADDERDELAY	PORT MAP(
	DIN0 => N112566916, 
	DIN1 => N112566917, 
	DIN2 => N112566918, 
	DIN3 => N112566919, 
	DIN4 => N112566920, 
	DIN5 => N112566921, 
	DIN6 => N112566922, 
	DIN7 => N112566923, 
	DIN8 => N112566924, 
	DIN9 => N112566925, 
	DIN10 => N112566926, 
	DIN11 => N112566927, 
	DIN12 => N112566928, 
	DIN13 => N112566929, 
	DIN14 => N112566930, 
	DIN15 => N112566931, 
	DOUT0 => N112591216, 
	DOUT1 => N112591217, 
	DOUT2 => N112591218, 
	DOUT3 => N112591219, 
	DOUT4 => N112591220, 
	DOUT5 => N112591221, 
	DOUT6 => N112591222, 
	DOUT7 => N112591223, 
	DOUT8 => N112591224, 
	DOUT9 => N112591225, 
	DOUT10 => N112591226, 
	DOUT11 => N112591227, 
	DOUT12 => N112591228, 
	DOUT13 => N112591229, 
	DOUT14 => N112591230, 
	DOUT15 => N112591231, 
	SIGNEDIN => N112566933, 
	SIGNEDOUT => N112591233
);
U182 : ADDERDELAY	PORT MAP(
	DIN0 => N112591216, 
	DIN1 => N112591217, 
	DIN2 => N112591218, 
	DIN3 => N112591219, 
	DIN4 => N112591220, 
	DIN5 => N112591221, 
	DIN6 => N112591222, 
	DIN7 => N112591223, 
	DIN8 => N112591224, 
	DIN9 => N112591225, 
	DIN10 => N112591226, 
	DIN11 => N112591227, 
	DIN12 => N112591228, 
	DIN13 => N112591229, 
	DIN14 => N112591230, 
	DIN15 => N112591231, 
	DOUT0 => N112615516, 
	DOUT1 => N112615517, 
	DOUT2 => N112615518, 
	DOUT3 => N112615519, 
	DOUT4 => N112615520, 
	DOUT5 => N112615521, 
	DOUT6 => N112615522, 
	DOUT7 => N112615523, 
	DOUT8 => N112615524, 
	DOUT9 => N112615525, 
	DOUT10 => N112615526, 
	DOUT11 => N112615527, 
	DOUT12 => N112615528, 
	DOUT13 => N112615529, 
	DOUT14 => N112615530, 
	DOUT15 => N112615531, 
	SIGNEDIN => N112591233, 
	SIGNEDOUT => N112615533
);
U150 : ADDERDELAY	PORT MAP(
	DIN0 => N111813616, 
	DIN1 => N111813617, 
	DIN2 => N111813618, 
	DIN3 => N111813619, 
	DIN4 => N111813620, 
	DIN5 => N111813621, 
	DIN6 => N111813622, 
	DIN7 => N111813623, 
	DIN8 => N111813624, 
	DIN9 => N111813625, 
	DIN10 => N111813626, 
	DIN11 => N111813627, 
	DIN12 => N111813628, 
	DIN13 => N111813629, 
	DIN14 => N111813630, 
	DIN15 => N111813631, 
	DOUT0 => N111837916, 
	DOUT1 => N111837917, 
	DOUT2 => N111837918, 
	DOUT3 => N111837919, 
	DOUT4 => N111837920, 
	DOUT5 => N111837921, 
	DOUT6 => N111837922, 
	DOUT7 => N111837923, 
	DOUT8 => N111837924, 
	DOUT9 => N111837925, 
	DOUT10 => N111837926, 
	DOUT11 => N111837927, 
	DOUT12 => N111837928, 
	DOUT13 => N111837929, 
	DOUT14 => N111837930, 
	DOUT15 => N111837931, 
	SIGNEDIN => N111813633, 
	SIGNEDOUT => N111837933
);
U183 : ADDERDELAY	PORT MAP(
	DIN0 => N112323916, 
	DIN1 => N112323917, 
	DIN2 => N112323918, 
	DIN3 => N112323919, 
	DIN4 => N112323920, 
	DIN5 => N112323921, 
	DIN6 => N112323922, 
	DIN7 => N112323923, 
	DIN8 => N112323924, 
	DIN9 => N112323925, 
	DIN10 => N112323926, 
	DIN11 => N112323927, 
	DIN12 => N112323928, 
	DIN13 => N112323929, 
	DIN14 => N112323930, 
	DIN15 => N112323931, 
	DOUT0 => N1147650, 
	DOUT1 => N1147610, 
	DOUT2 => N1147646, 
	DOUT3 => N1147618, 
	DOUT4 => N1147602, 
	DOUT5 => N1147630, 
	DOUT6 => N1147658, 
	DOUT7 => N1147654, 
	DOUT8 => N1147638, 
	DOUT9 => N1147626, 
	DOUT10 => N1147642, 
	DOUT11 => N1147634, 
	DOUT12 => N1147614, 
	DOUT13 => N1147622, 
	DOUT14 => N1147594, 
	DOUT15 => N1147598, 
	SIGNEDIN => N112323933, 
	SIGNEDOUT => N1147606
);
U151 : ADDERDELAY	PORT MAP(
	DIN0 => N111138516, 
	DIN1 => N111138517, 
	DIN2 => N111138518, 
	DIN3 => N111138519, 
	DIN4 => N111138520, 
	DIN5 => N111138521, 
	DIN6 => N111138522, 
	DIN7 => N111138523, 
	DIN8 => N111138524, 
	DIN9 => N111138525, 
	DIN10 => N111138526, 
	DIN11 => N111138527, 
	DIN12 => N111138528, 
	DIN13 => N111138529, 
	DIN14 => N111138530, 
	DIN15 => N111138531, 
	DOUT0 => N111862216, 
	DOUT1 => N111862217, 
	DOUT2 => N111862218, 
	DOUT3 => N111862219, 
	DOUT4 => N111862220, 
	DOUT5 => N111862221, 
	DOUT6 => N111862222, 
	DOUT7 => N111862223, 
	DOUT8 => N111862224, 
	DOUT9 => N111862225, 
	DOUT10 => N111862226, 
	DOUT11 => N111862227, 
	DOUT12 => N111862228, 
	DOUT13 => N111862229, 
	DOUT14 => N111862230, 
	DOUT15 => N111862231, 
	SIGNEDIN => N111138533, 
	SIGNEDOUT => N111862233
);
U184 : ADDERDELAY	PORT MAP(
	DIN0 => N112421116, 
	DIN1 => N112421117, 
	DIN2 => N112421118, 
	DIN3 => N112421119, 
	DIN4 => N112421120, 
	DIN5 => N112421121, 
	DIN6 => N112421122, 
	DIN7 => N112421123, 
	DIN8 => N112421124, 
	DIN9 => N112421125, 
	DIN10 => N112421126, 
	DIN11 => N112421127, 
	DIN12 => N112421128, 
	DIN13 => N112421129, 
	DIN14 => N112421130, 
	DIN15 => N112421131, 
	DOUT0 => N112664116, 
	DOUT1 => N112664117, 
	DOUT2 => N112664118, 
	DOUT3 => N112664119, 
	DOUT4 => N112664120, 
	DOUT5 => N112664121, 
	DOUT6 => N112664122, 
	DOUT7 => N112664123, 
	DOUT8 => N112664124, 
	DOUT9 => N112664125, 
	DOUT10 => N112664126, 
	DOUT11 => N112664127, 
	DOUT12 => N112664128, 
	DOUT13 => N112664129, 
	DOUT14 => N112664130, 
	DOUT15 => N112664131, 
	SIGNEDIN => N112421133, 
	SIGNEDOUT => N112664133
);
U152 : ADDERDELAY	PORT MAP(
	DIN0 => N111862216, 
	DIN1 => N111862217, 
	DIN2 => N111862218, 
	DIN3 => N111862219, 
	DIN4 => N111862220, 
	DIN5 => N111862221, 
	DIN6 => N111862222, 
	DIN7 => N111862223, 
	DIN8 => N111862224, 
	DIN9 => N111862225, 
	DIN10 => N111862226, 
	DIN11 => N111862227, 
	DIN12 => N111862228, 
	DIN13 => N111862229, 
	DIN14 => N111862230, 
	DIN15 => N111862231, 
	DOUT0 => N111886516, 
	DOUT1 => N111886517, 
	DOUT2 => N111886518, 
	DOUT3 => N111886519, 
	DOUT4 => N111886520, 
	DOUT5 => N111886521, 
	DOUT6 => N111886522, 
	DOUT7 => N111886523, 
	DOUT8 => N111886524, 
	DOUT9 => N111886525, 
	DOUT10 => N111886526, 
	DOUT11 => N111886527, 
	DOUT12 => N111886528, 
	DOUT13 => N111886529, 
	DOUT14 => N111886530, 
	DOUT15 => N111886531, 
	SIGNEDIN => N111862233, 
	SIGNEDOUT => N111886533
);
U120 : ADDERDELAY	PORT MAP(
	DIN0 => N11108610, 
	DIN1 => N11108611, 
	DIN2 => N11108612, 
	DIN3 => N11108613, 
	DIN4 => N11108614, 
	DIN5 => N11108615, 
	DIN6 => N11108616, 
	DIN7 => N11108617, 
	DIN8 => N11108618, 
	DIN9 => N11108619, 
	DIN10 => N111086110, 
	DIN11 => N111086111, 
	DIN12 => N111086112, 
	DIN13 => N111086113, 
	DIN14 => N111086114, 
	DIN15 => N111086115, 
	DOUT0 => N111086116, 
	DOUT1 => N111086117, 
	DOUT2 => N111086118, 
	DOUT3 => N111086119, 
	DOUT4 => N111086120, 
	DOUT5 => N111086121, 
	DOUT6 => N111086122, 
	DOUT7 => N111086123, 
	DOUT8 => N111086124, 
	DOUT9 => N111086125, 
	DOUT10 => N111086126, 
	DOUT11 => N111086127, 
	DOUT12 => N111086128, 
	DOUT13 => N111086129, 
	DOUT14 => N111086130, 
	DOUT15 => N111086131, 
	SIGNEDIN => N111086132, 
	SIGNEDOUT => N111086133
);
U185 : ADDERDELAY	PORT MAP(
	DIN0 => N112664116, 
	DIN1 => N112664117, 
	DIN2 => N112664118, 
	DIN3 => N112664119, 
	DIN4 => N112664120, 
	DIN5 => N112664121, 
	DIN6 => N112664122, 
	DIN7 => N112664123, 
	DIN8 => N112664124, 
	DIN9 => N112664125, 
	DIN10 => N112664126, 
	DIN11 => N112664127, 
	DIN12 => N112664128, 
	DIN13 => N112664129, 
	DIN14 => N112664130, 
	DIN15 => N112664131, 
	DOUT0 => N1132733, 
	DOUT1 => N1132502, 
	DOUT2 => N1131487, 
	DOUT3 => N1131102, 
	DOUT4 => N1130871, 
	DOUT5 => N1130640, 
	DOUT6 => N1130409, 
	DOUT7 => N1130178, 
	DOUT8 => N1129947, 
	DOUT9 => N1129716, 
	DOUT10 => N1129485, 
	DOUT11 => N1129254, 
	DOUT12 => N1129023, 
	DOUT13 => N1128792, 
	DOUT14 => N1128561, 
	DOUT15 => N1128330, 
	SIGNEDIN => N112664133, 
	SIGNEDOUT => N1128099
);
U153 : ADDERDELAY	PORT MAP(
	DIN0 => N111886516, 
	DIN1 => N111886517, 
	DIN2 => N111886518, 
	DIN3 => N111886519, 
	DIN4 => N111886520, 
	DIN5 => N111886521, 
	DIN6 => N111886522, 
	DIN7 => N111886523, 
	DIN8 => N111886524, 
	DIN9 => N111886525, 
	DIN10 => N111886526, 
	DIN11 => N111886527, 
	DIN12 => N111886528, 
	DIN13 => N111886529, 
	DIN14 => N111886530, 
	DIN15 => N111886531, 
	DOUT0 => N111910816, 
	DOUT1 => N111910817, 
	DOUT2 => N111910818, 
	DOUT3 => N111910819, 
	DOUT4 => N111910820, 
	DOUT5 => N111910821, 
	DOUT6 => N111910822, 
	DOUT7 => N111910823, 
	DOUT8 => N111910824, 
	DOUT9 => N111910825, 
	DOUT10 => N111910826, 
	DOUT11 => N111910827, 
	DOUT12 => N111910828, 
	DOUT13 => N111910829, 
	DOUT14 => N111910830, 
	DOUT15 => N111910831, 
	SIGNEDIN => N111886533, 
	SIGNEDOUT => N111910833
);
U121 : ADDERDELAY	PORT MAP(
	DIN0 => N111086116, 
	DIN1 => N111086117, 
	DIN2 => N111086118, 
	DIN3 => N111086119, 
	DIN4 => N111086120, 
	DIN5 => N111086121, 
	DIN6 => N111086122, 
	DIN7 => N111086123, 
	DIN8 => N111086124, 
	DIN9 => N111086125, 
	DIN10 => N111086126, 
	DIN11 => N111086127, 
	DIN12 => N111086128, 
	DIN13 => N111086129, 
	DIN14 => N111086130, 
	DIN15 => N111086131, 
	DOUT0 => N111114216, 
	DOUT1 => N111114217, 
	DOUT2 => N111114218, 
	DOUT3 => N111114219, 
	DOUT4 => N111114220, 
	DOUT5 => N111114221, 
	DOUT6 => N111114222, 
	DOUT7 => N111114223, 
	DOUT8 => N111114224, 
	DOUT9 => N111114225, 
	DOUT10 => N111114226, 
	DOUT11 => N111114227, 
	DOUT12 => N111114228, 
	DOUT13 => N111114229, 
	DOUT14 => N111114230, 
	DOUT15 => N111114231, 
	SIGNEDIN => N111086133, 
	SIGNEDOUT => N111114233
);
U186 : ADDERDELAY	PORT MAP(
	DIN0 => N112518316, 
	DIN1 => N112518317, 
	DIN2 => N112518318, 
	DIN3 => N112518319, 
	DIN4 => N112518320, 
	DIN5 => N112518321, 
	DIN6 => N112518322, 
	DIN7 => N112518323, 
	DIN8 => N112518324, 
	DIN9 => N112518325, 
	DIN10 => N112518326, 
	DIN11 => N112518327, 
	DIN12 => N112518328, 
	DIN13 => N112518329, 
	DIN14 => N112518330, 
	DIN15 => N112518331, 
	DOUT0 => N112712716, 
	DOUT1 => N112712717, 
	DOUT2 => N112712718, 
	DOUT3 => N112712719, 
	DOUT4 => N112712720, 
	DOUT5 => N112712721, 
	DOUT6 => N112712722, 
	DOUT7 => N112712723, 
	DOUT8 => N112712724, 
	DOUT9 => N112712725, 
	DOUT10 => N112712726, 
	DOUT11 => N112712727, 
	DOUT12 => N112712728, 
	DOUT13 => N112712729, 
	DOUT14 => N112712730, 
	DOUT15 => N112712731, 
	SIGNEDIN => N112518333, 
	SIGNEDOUT => N112712733
);
U154 : ADDERDELAY	PORT MAP(
	DIN0 => N111215216, 
	DIN1 => N111215217, 
	DIN2 => N111215218, 
	DIN3 => N111215219, 
	DIN4 => N111215220, 
	DIN5 => N111215221, 
	DIN6 => N111215222, 
	DIN7 => N111215223, 
	DIN8 => N111215224, 
	DIN9 => N111215225, 
	DIN10 => N111215226, 
	DIN11 => N111215227, 
	DIN12 => N111215228, 
	DIN13 => N111215229, 
	DIN14 => N111215230, 
	DIN15 => N111215231, 
	DOUT0 => N111935116, 
	DOUT1 => N111935117, 
	DOUT2 => N111935118, 
	DOUT3 => N111935119, 
	DOUT4 => N111935120, 
	DOUT5 => N111935121, 
	DOUT6 => N111935122, 
	DOUT7 => N111935123, 
	DOUT8 => N111935124, 
	DOUT9 => N111935125, 
	DOUT10 => N111935126, 
	DOUT11 => N111935127, 
	DOUT12 => N111935128, 
	DOUT13 => N111935129, 
	DOUT14 => N111935130, 
	DOUT15 => N111935131, 
	SIGNEDIN => N111215233, 
	SIGNEDOUT => N111935133
);
U122 : ADDERDELAY	PORT MAP(
	DIN0 => N111114216, 
	DIN1 => N111114217, 
	DIN2 => N111114218, 
	DIN3 => N111114219, 
	DIN4 => N111114220, 
	DIN5 => N111114221, 
	DIN6 => N111114222, 
	DIN7 => N111114223, 
	DIN8 => N111114224, 
	DIN9 => N111114225, 
	DIN10 => N111114226, 
	DIN11 => N111114227, 
	DIN12 => N111114228, 
	DIN13 => N111114229, 
	DIN14 => N111114230, 
	DIN15 => N111114231, 
	DOUT0 => N111138516, 
	DOUT1 => N111138517, 
	DOUT2 => N111138518, 
	DOUT3 => N111138519, 
	DOUT4 => N111138520, 
	DOUT5 => N111138521, 
	DOUT6 => N111138522, 
	DOUT7 => N111138523, 
	DOUT8 => N111138524, 
	DOUT9 => N111138525, 
	DOUT10 => N111138526, 
	DOUT11 => N111138527, 
	DOUT12 => N111138528, 
	DOUT13 => N111138529, 
	DOUT14 => N111138530, 
	DOUT15 => N111138531, 
	SIGNEDIN => N111114233, 
	SIGNEDOUT => N111138533
);
U187 : ADDERDELAY	PORT MAP(
	DIN0 => N112712716, 
	DIN1 => N112712717, 
	DIN2 => N112712718, 
	DIN3 => N112712719, 
	DIN4 => N112712720, 
	DIN5 => N112712721, 
	DIN6 => N112712722, 
	DIN7 => N112712723, 
	DIN8 => N112712724, 
	DIN9 => N112712725, 
	DIN10 => N112712726, 
	DIN11 => N112712727, 
	DIN12 => N112712728, 
	DIN13 => N112712729, 
	DIN14 => N112712730, 
	DIN15 => N112712731, 
	DOUT0 => N112737016, 
	DOUT1 => N112737017, 
	DOUT2 => N112737018, 
	DOUT3 => N112737019, 
	DOUT4 => N112737020, 
	DOUT5 => N112737021, 
	DOUT6 => N112737022, 
	DOUT7 => N112737023, 
	DOUT8 => N112737024, 
	DOUT9 => N112737025, 
	DOUT10 => N112737026, 
	DOUT11 => N112737027, 
	DOUT12 => N112737028, 
	DOUT13 => N112737029, 
	DOUT14 => N112737030, 
	DOUT15 => N112737031, 
	SIGNEDIN => N112712733, 
	SIGNEDOUT => N112737033
);
U155 : ADDERDELAY	PORT MAP(
	DIN0 => N111935116, 
	DIN1 => N111935117, 
	DIN2 => N111935118, 
	DIN3 => N111935119, 
	DIN4 => N111935120, 
	DIN5 => N111935121, 
	DIN6 => N111935122, 
	DIN7 => N111935123, 
	DIN8 => N111935124, 
	DIN9 => N111935125, 
	DIN10 => N111935126, 
	DIN11 => N111935127, 
	DIN12 => N111935128, 
	DIN13 => N111935129, 
	DIN14 => N111935130, 
	DIN15 => N111935131, 
	DOUT0 => N111959416, 
	DOUT1 => N111959417, 
	DOUT2 => N111959418, 
	DOUT3 => N111959419, 
	DOUT4 => N111959420, 
	DOUT5 => N111959421, 
	DOUT6 => N111959422, 
	DOUT7 => N111959423, 
	DOUT8 => N111959424, 
	DOUT9 => N111959425, 
	DOUT10 => N111959426, 
	DOUT11 => N111959427, 
	DOUT12 => N111959428, 
	DOUT13 => N111959429, 
	DOUT14 => N111959430, 
	DOUT15 => N111959431, 
	SIGNEDIN => N111935133, 
	SIGNEDOUT => N111959433
);
U123 : ADDERDELAY	PORT MAP(
	DIN0 => N11116280, 
	DIN1 => N11116281, 
	DIN2 => N11116282, 
	DIN3 => N11116283, 
	DIN4 => N11116284, 
	DIN5 => N11116285, 
	DIN6 => N11116286, 
	DIN7 => N11116287, 
	DIN8 => N11116288, 
	DIN9 => N11116289, 
	DIN10 => N111162810, 
	DIN11 => N111162811, 
	DIN12 => N111162812, 
	DIN13 => N111162813, 
	DIN14 => N111162814, 
	DIN15 => N111162815, 
	DOUT0 => N111162816, 
	DOUT1 => N111162817, 
	DOUT2 => N111162818, 
	DOUT3 => N111162819, 
	DOUT4 => N111162820, 
	DOUT5 => N111162821, 
	DOUT6 => N111162822, 
	DOUT7 => N111162823, 
	DOUT8 => N111162824, 
	DOUT9 => N111162825, 
	DOUT10 => N111162826, 
	DOUT11 => N111162827, 
	DOUT12 => N111162828, 
	DOUT13 => N111162829, 
	DOUT14 => N111162830, 
	DOUT15 => N111162831, 
	SIGNEDIN => N111162832, 
	SIGNEDOUT => N111162833
);
U188 : ADDERDELAY	PORT MAP(
	DIN0 => N112615516, 
	DIN1 => N112615517, 
	DIN2 => N112615518, 
	DIN3 => N112615519, 
	DIN4 => N112615520, 
	DIN5 => N112615521, 
	DIN6 => N112615522, 
	DIN7 => N112615523, 
	DIN8 => N112615524, 
	DIN9 => N112615525, 
	DIN10 => N112615526, 
	DIN11 => N112615527, 
	DIN12 => N112615528, 
	DIN13 => N112615529, 
	DIN14 => N112615530, 
	DIN15 => N112615531, 
	DOUT0 => N112761316, 
	DOUT1 => N112761317, 
	DOUT2 => N112761318, 
	DOUT3 => N112761319, 
	DOUT4 => N112761320, 
	DOUT5 => N112761321, 
	DOUT6 => N112761322, 
	DOUT7 => N112761323, 
	DOUT8 => N112761324, 
	DOUT9 => N112761325, 
	DOUT10 => N112761326, 
	DOUT11 => N112761327, 
	DOUT12 => N112761328, 
	DOUT13 => N112761329, 
	DOUT14 => N112761330, 
	DOUT15 => N112761331, 
	SIGNEDIN => N112615533, 
	SIGNEDOUT => N112761333
);
U124 : ADDERDELAY	PORT MAP(
	DIN0 => N111162816, 
	DIN1 => N111162817, 
	DIN2 => N111162818, 
	DIN3 => N111162819, 
	DIN4 => N111162820, 
	DIN5 => N111162821, 
	DIN6 => N111162822, 
	DIN7 => N111162823, 
	DIN8 => N111162824, 
	DIN9 => N111162825, 
	DIN10 => N111162826, 
	DIN11 => N111162827, 
	DIN12 => N111162828, 
	DIN13 => N111162829, 
	DIN14 => N111162830, 
	DIN15 => N111162831, 
	DOUT0 => N111190916, 
	DOUT1 => N111190917, 
	DOUT2 => N111190918, 
	DOUT3 => N111190919, 
	DOUT4 => N111190920, 
	DOUT5 => N111190921, 
	DOUT6 => N111190922, 
	DOUT7 => N111190923, 
	DOUT8 => N111190924, 
	DOUT9 => N111190925, 
	DOUT10 => N111190926, 
	DOUT11 => N111190927, 
	DOUT12 => N111190928, 
	DOUT13 => N111190929, 
	DOUT14 => N111190930, 
	DOUT15 => N111190931, 
	SIGNEDIN => N111162833, 
	SIGNEDOUT => N111190933
);
U156 : ADDERDELAY	PORT MAP(
	DIN0 => N111959416, 
	DIN1 => N111959417, 
	DIN2 => N111959418, 
	DIN3 => N111959419, 
	DIN4 => N111959420, 
	DIN5 => N111959421, 
	DIN6 => N111959422, 
	DIN7 => N111959423, 
	DIN8 => N111959424, 
	DIN9 => N111959425, 
	DIN10 => N111959426, 
	DIN11 => N111959427, 
	DIN12 => N111959428, 
	DIN13 => N111959429, 
	DIN14 => N111959430, 
	DIN15 => N111959431, 
	DOUT0 => N111983716, 
	DOUT1 => N111983717, 
	DOUT2 => N111983718, 
	DOUT3 => N111983719, 
	DOUT4 => N111983720, 
	DOUT5 => N111983721, 
	DOUT6 => N111983722, 
	DOUT7 => N111983723, 
	DOUT8 => N111983724, 
	DOUT9 => N111983725, 
	DOUT10 => N111983726, 
	DOUT11 => N111983727, 
	DOUT12 => N111983728, 
	DOUT13 => N111983729, 
	DOUT14 => N111983730, 
	DOUT15 => N111983731, 
	SIGNEDIN => N111959433, 
	SIGNEDOUT => N111983733
);
U189 : ADDERDELAY	PORT MAP(
	DIN0 => N112761316, 
	DIN1 => N112761317, 
	DIN2 => N112761318, 
	DIN3 => N112761319, 
	DIN4 => N112761320, 
	DIN5 => N112761321, 
	DIN6 => N112761322, 
	DIN7 => N112761323, 
	DIN8 => N112761324, 
	DIN9 => N112761325, 
	DIN10 => N112761326, 
	DIN11 => N112761327, 
	DIN12 => N112761328, 
	DIN13 => N112761329, 
	DIN14 => N112761330, 
	DIN15 => N112761331, 
	DOUT0 => N112785616, 
	DOUT1 => N112785617, 
	DOUT2 => N112785618, 
	DOUT3 => N112785619, 
	DOUT4 => N112785620, 
	DOUT5 => N112785621, 
	DOUT6 => N112785622, 
	DOUT7 => N112785623, 
	DOUT8 => N112785624, 
	DOUT9 => N112785625, 
	DOUT10 => N112785626, 
	DOUT11 => N112785627, 
	DOUT12 => N112785628, 
	DOUT13 => N112785629, 
	DOUT14 => N112785630, 
	DOUT15 => N112785631, 
	SIGNEDIN => N112761333, 
	SIGNEDOUT => N112785633
);
U125 : ADDERDELAY	PORT MAP(
	DIN0 => N111190916, 
	DIN1 => N111190917, 
	DIN2 => N111190918, 
	DIN3 => N111190919, 
	DIN4 => N111190920, 
	DIN5 => N111190921, 
	DIN6 => N111190922, 
	DIN7 => N111190923, 
	DIN8 => N111190924, 
	DIN9 => N111190925, 
	DIN10 => N111190926, 
	DIN11 => N111190927, 
	DIN12 => N111190928, 
	DIN13 => N111190929, 
	DIN14 => N111190930, 
	DIN15 => N111190931, 
	DOUT0 => N111215216, 
	DOUT1 => N111215217, 
	DOUT2 => N111215218, 
	DOUT3 => N111215219, 
	DOUT4 => N111215220, 
	DOUT5 => N111215221, 
	DOUT6 => N111215222, 
	DOUT7 => N111215223, 
	DOUT8 => N111215224, 
	DOUT9 => N111215225, 
	DOUT10 => N111215226, 
	DOUT11 => N111215227, 
	DOUT12 => N111215228, 
	DOUT13 => N111215229, 
	DOUT14 => N111215230, 
	DOUT15 => N111215231, 
	SIGNEDIN => N111190933, 
	SIGNEDOUT => N111215233
);
U157 : ADDERDELAY	PORT MAP(
	DIN0 => N111473416, 
	DIN1 => N111473417, 
	DIN2 => N111473418, 
	DIN3 => N111473419, 
	DIN4 => N111473420, 
	DIN5 => N111473421, 
	DIN6 => N111473422, 
	DIN7 => N111473423, 
	DIN8 => N111473424, 
	DIN9 => N111473425, 
	DIN10 => N111473426, 
	DIN11 => N111473427, 
	DIN12 => N111473428, 
	DIN13 => N111473429, 
	DIN14 => N111473430, 
	DIN15 => N111473431, 
	DOUT0 => N1147006, 
	DOUT1 => N1146966, 
	DOUT2 => N1147002, 
	DOUT3 => N1146974, 
	DOUT4 => N1146958, 
	DOUT5 => N1146986, 
	DOUT6 => N1147014, 
	DOUT7 => N1147010, 
	DOUT8 => N1146994, 
	DOUT9 => N1146982, 
	DOUT10 => N1146998, 
	DOUT11 => N1146990, 
	DOUT12 => N1146970, 
	DOUT13 => N1146978, 
	DOUT14 => N1146950, 
	DOUT15 => N1146954, 
	SIGNEDIN => N111473433, 
	SIGNEDOUT => N1146962
);
U126 : ADDERDELAY	PORT MAP(
	DIN0 => N110448216, 
	DIN1 => N110448217, 
	DIN2 => N110448218, 
	DIN3 => N110448219, 
	DIN4 => N110448220, 
	DIN5 => N110448221, 
	DIN6 => N110448222, 
	DIN7 => N110448223, 
	DIN8 => N110448224, 
	DIN9 => N110448225, 
	DIN10 => N110448226, 
	DIN11 => N110448227, 
	DIN12 => N110448228, 
	DIN13 => N110448229, 
	DIN14 => N110448230, 
	DIN15 => N110448231, 
	DOUT0 => N1145385, 
	DOUT1 => N1145345, 
	DOUT2 => N1145381, 
	DOUT3 => N1145353, 
	DOUT4 => N1145337, 
	DOUT5 => N1145365, 
	DOUT6 => N1145393, 
	DOUT7 => N1145389, 
	DOUT8 => N1145373, 
	DOUT9 => N1145361, 
	DOUT10 => N1145377, 
	DOUT11 => N1145369, 
	DOUT12 => N1145349, 
	DOUT13 => N1145357, 
	DOUT14 => N1145329, 
	DOUT15 => N1145333, 
	SIGNEDIN => N110448233, 
	SIGNEDOUT => N1145341
);
U158 : ADDERDELAY	PORT MAP(
	DIN0 => N111546316, 
	DIN1 => N111546317, 
	DIN2 => N111546318, 
	DIN3 => N111546319, 
	DIN4 => N111546320, 
	DIN5 => N111546321, 
	DIN6 => N111546322, 
	DIN7 => N111546323, 
	DIN8 => N111546324, 
	DIN9 => N111546325, 
	DIN10 => N111546326, 
	DIN11 => N111546327, 
	DIN12 => N111546328, 
	DIN13 => N111546329, 
	DIN14 => N111546330, 
	DIN15 => N111546331, 
	DOUT0 => N112032316, 
	DOUT1 => N112032317, 
	DOUT2 => N112032318, 
	DOUT3 => N112032319, 
	DOUT4 => N112032320, 
	DOUT5 => N112032321, 
	DOUT6 => N112032322, 
	DOUT7 => N112032323, 
	DOUT8 => N112032324, 
	DOUT9 => N112032325, 
	DOUT10 => N112032326, 
	DOUT11 => N112032327, 
	DOUT12 => N112032328, 
	DOUT13 => N112032329, 
	DOUT14 => N112032330, 
	DOUT15 => N112032331, 
	SIGNEDIN => N111546333, 
	SIGNEDOUT => N112032333
);
U127 : ADDERDELAY	PORT MAP(
	DIN0 => N110524916, 
	DIN1 => N110524917, 
	DIN2 => N110524918, 
	DIN3 => N110524919, 
	DIN4 => N110524920, 
	DIN5 => N110524921, 
	DIN6 => N110524922, 
	DIN7 => N110524923, 
	DIN8 => N110524924, 
	DIN9 => N110524925, 
	DIN10 => N110524926, 
	DIN11 => N110524927, 
	DIN12 => N110524928, 
	DIN13 => N110524929, 
	DIN14 => N110524930, 
	DIN15 => N110524931, 
	DOUT0 => N111263816, 
	DOUT1 => N111263817, 
	DOUT2 => N111263818, 
	DOUT3 => N111263819, 
	DOUT4 => N111263820, 
	DOUT5 => N111263821, 
	DOUT6 => N111263822, 
	DOUT7 => N111263823, 
	DOUT8 => N111263824, 
	DOUT9 => N111263825, 
	DOUT10 => N111263826, 
	DOUT11 => N111263827, 
	DOUT12 => N111263828, 
	DOUT13 => N111263829, 
	DOUT14 => N111263830, 
	DOUT15 => N111263831, 
	SIGNEDIN => N110524933, 
	SIGNEDOUT => N111263833
);
U159 : ADDERDELAY	PORT MAP(
	DIN0 => N112032316, 
	DIN1 => N112032317, 
	DIN2 => N112032318, 
	DIN3 => N112032319, 
	DIN4 => N112032320, 
	DIN5 => N112032321, 
	DIN6 => N112032322, 
	DIN7 => N112032323, 
	DIN8 => N112032324, 
	DIN9 => N112032325, 
	DIN10 => N112032326, 
	DIN11 => N112032327, 
	DIN12 => N112032328, 
	DIN13 => N112032329, 
	DIN14 => N112032330, 
	DIN15 => N112032331, 
	DOUT0 => N1147167, 
	DOUT1 => N1147127, 
	DOUT2 => N1147163, 
	DOUT3 => N1147135, 
	DOUT4 => N1147119, 
	DOUT5 => N1147147, 
	DOUT6 => N1147175, 
	DOUT7 => N1147171, 
	DOUT8 => N1147155, 
	DOUT9 => N1147143, 
	DOUT10 => N1147159, 
	DOUT11 => N1147151, 
	DOUT12 => N1147131, 
	DOUT13 => N1147139, 
	DOUT14 => N1147111, 
	DOUT15 => N1147115, 
	SIGNEDIN => N112032333, 
	SIGNEDOUT => N1147123
);
U128 : ADDERDELAY	PORT MAP(
	DIN0 => N111263816, 
	DIN1 => N111263817, 
	DIN2 => N111263818, 
	DIN3 => N111263819, 
	DIN4 => N111263820, 
	DIN5 => N111263821, 
	DIN6 => N111263822, 
	DIN7 => N111263823, 
	DIN8 => N111263824, 
	DIN9 => N111263825, 
	DIN10 => N111263826, 
	DIN11 => N111263827, 
	DIN12 => N111263828, 
	DIN13 => N111263829, 
	DIN14 => N111263830, 
	DIN15 => N111263831, 
	DOUT0 => N1146684, 
	DOUT1 => N1146644, 
	DOUT2 => N1146680, 
	DOUT3 => N1146652, 
	DOUT4 => N1146636, 
	DOUT5 => N1146664, 
	DOUT6 => N1146692, 
	DOUT7 => N1146688, 
	DOUT8 => N1146672, 
	DOUT9 => N1146660, 
	DOUT10 => N1146676, 
	DOUT11 => N1146668, 
	DOUT12 => N1146648, 
	DOUT13 => N1146656, 
	DOUT14 => N1146628, 
	DOUT15 => N1146632, 
	SIGNEDIN => N111263833, 
	SIGNEDOUT => N1146640
);
U129 : \16adderBalanced\	PORT MAP(
	A0 => N1263850, 
	A1 => N1251498, 
	A2 => N1268390, 
	A3 => N1244642, 
	A4 => N1258106, 
	A5 => N1260508, 
	A6 => N1257374, 
	A7 => N1261526, 
	A8 => N1254680, 
	A9 => N1263768, 
	A10 => N1250090, 
	A11 => N1257164, 
	A12 => N1248836, 
	A13 => N1267774, 
	A14 => N1265342, 
	A15 => N1262264, 
	B0 => TG0, 
	B1 => TG1, 
	B2 => TG2, 
	B3 => TG3, 
	B4 => TG4, 
	B5 => TG5, 
	B6 => TG6, 
	B7 => TG7, 
	B8 => TG8, 
	B9 => TG9, 
	B10 => TG10, 
	B11 => TG11, 
	B12 => TG12, 
	B13 => TG13, 
	B14 => TG14, 
	B15 => TG15, 
	CIN => N1256014, 
	COUT => N1056495, 
	Y0 => N108992, 
	Y1 => N109348, 
	Y2 => N109000, 
	Y3 => N109356, 
	Y4 => N109344, 
	Y5 => N109008, 
	Y6 => N108996, 
	Y7 => N109352, 
	Y8 => N109340, 
	Y9 => N109336, 
	Y10 => N109332, 
	Y11 => N109328, 
	Y12 => N109324, 
	Y13 => N109012, 
	Y14 => N109016, 
	Y15 => N109004
);
U200 : TAPADDER	PORT MAP(
	A0 => N1132733, 
	A1 => N1132502, 
	A2 => N1131487, 
	A3 => N1131102, 
	A4 => N1130871, 
	A5 => N1130640, 
	A6 => N1130409, 
	A7 => N1130178, 
	A8 => N1129947, 
	A9 => N1129716, 
	A10 => N1129485, 
	A11 => N1129254, 
	A12 => N1129023, 
	A13 => N1128792, 
	A14 => N1128561, 
	A15 => N1128330, 
	AND1 => N94153, 
	AND2 => N94147, 
	AND3 => N94157, 
	B0 => N107806, 
	B1 => N108278, 
	B2 => N107814, 
	B3 => N108286, 
	B4 => N108274, 
	B5 => N107822, 
	B6 => N107810, 
	B7 => N108282, 
	B8 => N108270, 
	B9 => N108266, 
	B10 => N108262, 
	B11 => N108258, 
	B12 => N108254, 
	B13 => N107826, 
	B14 => N107830, 
	B15 => N107818, 
	CIN => N1128099, 
	COUT => N1057544, 
	O0 => G0, 
	O1 => G1, 
	O2 => G2, 
	O3 => G3, 
	O4 => G4, 
	O5 => G5, 
	O6 => G6, 
	O7 => G7, 
	O8 => G8, 
	O9 => G9, 
	O10 => G10, 
	O11 => G11, 
	O12 => G12, 
	O13 => G13, 
	O14 => G14, 
	O15 => G15, 
	OR1 => N94145, 
	OR2 => N94155, 
	OR3 => N94149, 
	Y0 => TG0, 
	Y1 => TG1, 
	Y2 => TG2, 
	Y3 => TG3, 
	Y4 => TG4, 
	Y5 => TG5, 
	Y6 => TG6, 
	Y7 => TG7, 
	Y8 => TG8, 
	Y9 => TG9, 
	Y10 => TG10, 
	Y11 => TG11, 
	Y12 => TG12, 
	Y13 => TG13, 
	Y14 => TG14, 
	Y15 => TG15
);
U201 : TAPADDER	PORT MAP(
	A0 => N1147489, 
	A1 => N1147449, 
	A2 => N1147485, 
	A3 => N1147457, 
	A4 => N1147441, 
	A5 => N1147469, 
	A6 => N1147497, 
	A7 => N1147493, 
	A8 => N1147477, 
	A9 => N1147465, 
	A10 => N1268884, 
	A11 => N1257378, 
	A12 => N1147453, 
	A13 => N1147461, 
	A14 => N1147433, 
	A15 => N1147437, 
	AND1 => N94153, 
	AND2 => N94155, 
	AND3 => N94157, 
	B0 => N103455, 
	B1 => N103927, 
	B2 => N103463, 
	B3 => N103935, 
	B4 => N103923, 
	B5 => N103471, 
	B6 => N103459, 
	B7 => N103931, 
	B8 => N103919, 
	B9 => N103915, 
	B10 => N103911, 
	B11 => N103907, 
	B12 => N103903, 
	B13 => N103475, 
	B14 => N103479, 
	B15 => N103467, 
	CIN => N1147445, 
	COUT => N1057858, 
	O0 => F0, 
	O1 => F1, 
	O2 => F2, 
	O3 => F3, 
	O4 => F4, 
	O5 => F5, 
	O6 => F6, 
	O7 => F7, 
	O8 => F8, 
	O9 => F9, 
	O10 => F10, 
	O11 => F11, 
	O12 => F12, 
	O13 => F13, 
	O14 => F14, 
	O15 => F15, 
	OR1 => N94145, 
	OR2 => N94147, 
	OR3 => N94149, 
	Y0 => TF0, 
	Y1 => TF1, 
	Y2 => TF2, 
	Y3 => TF3, 
	Y4 => TF4, 
	Y5 => TF5, 
	Y6 => TF6, 
	Y7 => TF7, 
	Y8 => TF8, 
	Y9 => TF9, 
	Y10 => TF10, 
	Y11 => TF11, 
	Y12 => TF12, 
	Y13 => TF13, 
	Y14 => TF14, 
	Y15 => TF15
);
U202 : TAPADDER	PORT MAP(
	A0 => N1147167, 
	A1 => N1147127, 
	A2 => N1147163, 
	A3 => N1147135, 
	A4 => N1147119, 
	A5 => N1147147, 
	A6 => N1147175, 
	A7 => N1147171, 
	A8 => N1147155, 
	A9 => N1147143, 
	A10 => N1147159, 
	A11 => N1147151, 
	A12 => N1147131, 
	A13 => N1147139, 
	A14 => N1147111, 
	A15 => N1147115, 
	AND1 => N94145, 
	AND2 => N94155, 
	AND3 => N94157, 
	B0 => N102421, 
	B1 => N102893, 
	B2 => N102429, 
	B3 => N102901, 
	B4 => N102889, 
	B5 => N102437, 
	B6 => N102425, 
	B7 => N102897, 
	B8 => N102885, 
	B9 => N102881, 
	B10 => N102877, 
	B11 => N102873, 
	B12 => N102869, 
	B13 => N102441, 
	B14 => N102445, 
	B15 => N102433, 
	CIN => N1147123, 
	COUT => N1058172, 
	O0 => E0, 
	O1 => E1, 
	O2 => E2, 
	O3 => E3, 
	O4 => E4, 
	O5 => E5, 
	O6 => E6, 
	O7 => E7, 
	O8 => E8, 
	O9 => E9, 
	O10 => E10, 
	O11 => E11, 
	O12 => E12, 
	O13 => E13, 
	O14 => E14, 
	O15 => E15, 
	OR1 => N94153, 
	OR2 => N94147, 
	OR3 => N94149, 
	Y0 => TE0, 
	Y1 => TE1, 
	Y2 => TE2, 
	Y3 => TE3, 
	Y4 => TE4, 
	Y5 => TE5, 
	Y6 => TE6, 
	Y7 => TE7, 
	Y8 => TE8, 
	Y9 => TE9, 
	Y10 => TE10, 
	Y11 => TE11, 
	Y12 => TE12, 
	Y13 => TE13, 
	Y14 => TE14, 
	Y15 => TE15
);
U203 : TAPADDER	PORT MAP(
	A0 => N1146845, 
	A1 => N1146805, 
	A2 => N1146841, 
	A3 => N1146813, 
	A4 => N1146797, 
	A5 => N1146825, 
	A6 => N1146853, 
	A7 => N1146849, 
	A8 => N1146833, 
	A9 => N1146821, 
	A10 => N1146837, 
	A11 => N1146829, 
	A12 => N1146809, 
	A13 => N1146817, 
	A14 => N1146789, 
	A15 => N1146793, 
	AND1 => N94145, 
	AND2 => N94155, 
	AND3 => N94149, 
	B0 => N100889, 
	B1 => N101361, 
	B2 => N100897, 
	B3 => N101369, 
	B4 => N101357, 
	B5 => N100905, 
	B6 => N100893, 
	B7 => N101365, 
	B8 => N101353, 
	B9 => N101349, 
	B10 => N101345, 
	B11 => N101341, 
	B12 => N101337, 
	B13 => N100909, 
	B14 => N100913, 
	B15 => N100901, 
	CIN => N1146801, 
	COUT => N1058486, 
	O0 => D0, 
	O1 => D1, 
	O2 => D2, 
	O3 => D3, 
	O4 => D4, 
	O5 => D5, 
	O6 => D6, 
	O7 => D7, 
	O8 => D8, 
	O9 => D9, 
	O10 => D10, 
	O11 => D11, 
	O12 => D12, 
	O13 => D13, 
	O14 => D14, 
	O15 => D15, 
	OR1 => N94153, 
	OR2 => N94147, 
	OR3 => N94157, 
	Y0 => TD0, 
	Y1 => TD1, 
	Y2 => TD2, 
	Y3 => TD3, 
	Y4 => TD4, 
	Y5 => TD5, 
	Y6 => TD6, 
	Y7 => TD7, 
	Y8 => TD8, 
	Y9 => TD9, 
	Y10 => TD10, 
	Y11 => TD11, 
	Y12 => TD12, 
	Y13 => TD13, 
	Y14 => TD14, 
	Y15 => TD15
);
U204 : TAPADDER	PORT MAP(
	A0 => N1145385, 
	A1 => N1145345, 
	A2 => N1145381, 
	A3 => N1145353, 
	A4 => N1145337, 
	A5 => N1145365, 
	A6 => N1145393, 
	A7 => N1145389, 
	A8 => N1145373, 
	A9 => N1145361, 
	A10 => N1145377, 
	A11 => N1145369, 
	A12 => N1145349, 
	A13 => N1145357, 
	A14 => N1145329, 
	A15 => N1145333, 
	AND1 => N94153, 
	AND2 => N94155, 
	AND3 => N94149, 
	B0 => N91218, 
	B1 => N91220, 
	B2 => N91190, 
	B3 => N91192, 
	B4 => N91194, 
	B5 => N91196, 
	B6 => N91198, 
	B7 => N91200, 
	B8 => N91202, 
	B9 => N91204, 
	B10 => N91206, 
	B11 => N91208, 
	B12 => N91210, 
	B13 => N91212, 
	B14 => N91214, 
	B15 => N91216, 
	CIN => N1145341, 
	COUT => N1058800, 
	O0 => C0, 
	O1 => C1, 
	O2 => C2, 
	O3 => C3, 
	O4 => C4, 
	O5 => C5, 
	O6 => C6, 
	O7 => C7, 
	O8 => C8, 
	O9 => C9, 
	O10 => C10, 
	O11 => C11, 
	O12 => C12, 
	O13 => C13, 
	O14 => C14, 
	O15 => C15, 
	OR1 => N94145, 
	OR2 => N94147, 
	OR3 => N94157, 
	Y0 => TC0, 
	Y1 => TC1, 
	Y2 => TC2, 
	Y3 => TC3, 
	Y4 => TC4, 
	Y5 => TC5, 
	Y6 => TC6, 
	Y7 => TC7, 
	Y8 => TC8, 
	Y9 => TC9, 
	Y10 => TC10, 
	Y11 => TC11, 
	Y12 => TC12, 
	Y13 => TC13, 
	Y14 => TC14, 
	Y15 => TC15
);
U205 : TAPADDER	PORT MAP(
	A0 => N1143362, 
	A1 => N1143322, 
	A2 => N1143358, 
	A3 => N1143330, 
	A4 => N1143314, 
	A5 => N1143342, 
	A6 => N1143370, 
	A7 => N1143366, 
	A8 => N1143350, 
	A9 => N1143338, 
	A10 => N1143354, 
	A11 => N1143346, 
	A12 => N1143326, 
	A13 => N1143334, 
	A14 => N1143306, 
	A15 => N1143310, 
	AND1 => N94153, 
	AND2 => N94147, 
	AND3 => N94149, 
	B0 => N99924, 
	B1 => N100396, 
	B2 => N99932, 
	B3 => N100404, 
	B4 => N100392, 
	B5 => N99940, 
	B6 => N99928, 
	B7 => N100400, 
	B8 => N100388, 
	B9 => N100384, 
	B10 => N100380, 
	B11 => N100376, 
	B12 => N100372, 
	B13 => N99944, 
	B14 => N99948, 
	B15 => N99936, 
	CIN => N1143318, 
	COUT => N1059114, 
	O0 => B0, 
	O1 => B1, 
	O2 => B2, 
	O3 => B3, 
	O4 => B4, 
	O5 => B5, 
	O6 => B6, 
	O7 => B7, 
	O8 => B8, 
	O9 => B9, 
	O10 => B10, 
	O11 => B11, 
	O12 => B12, 
	O13 => B13, 
	O14 => B14, 
	O15 => B15, 
	OR1 => N94155, 
	OR2 => N94157, 
	OR3 => N94145, 
	Y0 => TB0, 
	Y1 => TB1, 
	Y2 => TB2, 
	Y3 => TB3, 
	Y4 => TB4, 
	Y5 => TB5, 
	Y6 => TB6, 
	Y7 => TB7, 
	Y8 => TB8, 
	Y9 => TB9, 
	Y10 => TB10, 
	Y11 => TB11, 
	Y12 => TB12, 
	Y13 => TB13, 
	Y14 => TB14, 
	Y15 => TB15
);
U206 : TAPADDER	PORT MAP(
	A0 => N1078467, 
	A1 => N1078469, 
	A2 => N1078471, 
	A3 => N1078473, 
	A4 => N1078475, 
	A5 => N1078477, 
	A6 => N1078479, 
	A7 => N1078481, 
	A8 => N1078483, 
	A9 => N1078485, 
	A10 => N1078487, 
	A11 => N1078489, 
	A12 => N1078491, 
	A13 => N1078493, 
	A14 => N1078495, 
	A15 => N1078497, 
	AND1 => N955836, 
	AND2 => N94147, 
	AND3 => N94149, 
	B0 => GND, 
	B1 => GND, 
	B2 => GND, 
	B3 => GND, 
	B4 => GND, 
	B5 => GND, 
	B6 => GND, 
	B7 => GND, 
	B8 => GND, 
	B9 => GND, 
	B10 => GND, 
	B11 => GND, 
	B12 => GND, 
	B13 => GND, 
	B14 => GND, 
	B15 => GND, 
	CIN => N1078499, 
	COUT => N1059428, 
	O0 => A0, 
	O1 => A1, 
	O2 => A2, 
	O3 => A3, 
	O4 => A4, 
	O5 => A5, 
	O6 => A6, 
	O7 => A7, 
	O8 => A8, 
	O9 => A9, 
	O10 => A10, 
	O11 => A11, 
	O12 => A12, 
	O13 => A13, 
	O14 => A14, 
	O15 => A15, 
	OR1 => N94155, 
	OR2 => N94157, 
	OR3 => N955599, 
	Y0 => TA0, 
	Y1 => TA1, 
	Y2 => TA2, 
	Y3 => TA3, 
	Y4 => TA4, 
	Y5 => TA5, 
	Y6 => TA6, 
	Y7 => TA7, 
	Y8 => TA8, 
	Y9 => TA9, 
	Y10 => TA10, 
	Y11 => TA11, 
	Y12 => TA12, 
	Y13 => TA13, 
	Y14 => TA14, 
	Y15 => TA15
);
U88 : ADDERDELAY	PORT MAP(
	DIN0 => N11026670, 
	DIN1 => N11026671, 
	DIN2 => N11026672, 
	DIN3 => N11026673, 
	DIN4 => N11026674, 
	DIN5 => N11026675, 
	DIN6 => N11026676, 
	DIN7 => N11026677, 
	DIN8 => N11026678, 
	DIN9 => N11026679, 
	DIN10 => N110266710, 
	DIN11 => N110266711, 
	DIN12 => N110266712, 
	DIN13 => N110266713, 
	DIN14 => N110266714, 
	DIN15 => N110266715, 
	DOUT0 => N110266716, 
	DOUT1 => N110266717, 
	DOUT2 => N110266718, 
	DOUT3 => N110266719, 
	DOUT4 => N110266720, 
	DOUT5 => N110266721, 
	DOUT6 => N110266722, 
	DOUT7 => N110266723, 
	DOUT8 => N110266724, 
	DOUT9 => N110266725, 
	DOUT10 => N110266726, 
	DOUT11 => N110266727, 
	DOUT12 => N110266728, 
	DOUT13 => N110266729, 
	DOUT14 => N110266730, 
	DOUT15 => N110266731, 
	SIGNEDIN => N110266732, 
	SIGNEDOUT => N110266733
);
U89 : ADDERDELAY	PORT MAP(
	DIN0 => N110266716, 
	DIN1 => N110266717, 
	DIN2 => N110266718, 
	DIN3 => N110266719, 
	DIN4 => N110266720, 
	DIN5 => N110266721, 
	DIN6 => N110266722, 
	DIN7 => N110266723, 
	DIN8 => N110266724, 
	DIN9 => N110266725, 
	DIN10 => N110266726, 
	DIN11 => N110266727, 
	DIN12 => N110266728, 
	DIN13 => N110266729, 
	DIN14 => N110266730, 
	DIN15 => N110266731, 
	DOUT0 => N1143362, 
	DOUT1 => N1143322, 
	DOUT2 => N1143358, 
	DOUT3 => N1143330, 
	DOUT4 => N1143314, 
	DOUT5 => N1143342, 
	DOUT6 => N1143370, 
	DOUT7 => N1143366, 
	DOUT8 => N1143350, 
	DOUT9 => N1143338, 
	DOUT10 => N1143354, 
	DOUT11 => N1143346, 
	DOUT12 => N1143326, 
	DOUT13 => N1143334, 
	DOUT14 => N1143306, 
	DOUT15 => N1143310, 
	SIGNEDIN => N110266733, 
	SIGNEDOUT => N1143318
);
U190 : ADDERDELAY	PORT MAP(
	DIN0 => N112737016, 
	DIN1 => N112737017, 
	DIN2 => N112737018, 
	DIN3 => N112737019, 
	DIN4 => N112737020, 
	DIN5 => N112737021, 
	DIN6 => N112737022, 
	DIN7 => N112737023, 
	DIN8 => N112737024, 
	DIN9 => N112737025, 
	DIN10 => N112737026, 
	DIN11 => N112737027, 
	DIN12 => N112737028, 
	DIN13 => N112737029, 
	DIN14 => N112737030, 
	DIN15 => N112737031, 
	DOUT0 => N1263850, 
	DOUT1 => N1251498, 
	DOUT2 => N1268390, 
	DOUT3 => N1244642, 
	DOUT4 => N1258106, 
	DOUT5 => N1260508, 
	DOUT6 => N1257374, 
	DOUT7 => N1261526, 
	DOUT8 => N1254680, 
	DOUT9 => N1263768, 
	DOUT10 => N1250090, 
	DOUT11 => N1257164, 
	DOUT12 => N1248836, 
	DOUT13 => N1267774, 
	DOUT14 => N1265342, 
	DOUT15 => N1262264, 
	SIGNEDIN => N112737033, 
	SIGNEDOUT => N1256014
);
U191 : ADDERDELAY	PORT MAP(
	DIN0 => N112785616, 
	DIN1 => N112785617, 
	DIN2 => N112785618, 
	DIN3 => N112785619, 
	DIN4 => N112785620, 
	DIN5 => N112785621, 
	DIN6 => N112785622, 
	DIN7 => N112785623, 
	DIN8 => N112785624, 
	DIN9 => N112785625, 
	DIN10 => N112785626, 
	DIN11 => N112785627, 
	DIN12 => N112785628, 
	DIN13 => N112785629, 
	DIN14 => N112785630, 
	DIN15 => N112785631, 
	DOUT0 => N113729316, 
	DOUT1 => N113729317, 
	DOUT2 => N113729318, 
	DOUT3 => N113729319, 
	DOUT4 => N113729320, 
	DOUT5 => N113729321, 
	DOUT6 => N113729322, 
	DOUT7 => N113729323, 
	DOUT8 => N113729324, 
	DOUT9 => N113729325, 
	DOUT10 => N113729326, 
	DOUT11 => N113729327, 
	DOUT12 => N113729328, 
	DOUT13 => N113729329, 
	DOUT14 => N113729330, 
	DOUT15 => N113729331, 
	SIGNEDIN => N112785633, 
	SIGNEDOUT => N113729333
);
U160 : ADDERDELAY	PORT MAP(
	DIN0 => N111619216, 
	DIN1 => N111619217, 
	DIN2 => N111619218, 
	DIN3 => N111619219, 
	DIN4 => N111619220, 
	DIN5 => N111619221, 
	DIN6 => N111619222, 
	DIN7 => N111619223, 
	DIN8 => N111619224, 
	DIN9 => N111619225, 
	DIN10 => N111619226, 
	DIN11 => N111619227, 
	DIN12 => N111619228, 
	DIN13 => N111619229, 
	DIN14 => N111619230, 
	DIN15 => N111619231, 
	DOUT0 => N112080916, 
	DOUT1 => N112080917, 
	DOUT2 => N112080918, 
	DOUT3 => N112080919, 
	DOUT4 => N112080920, 
	DOUT5 => N112080921, 
	DOUT6 => N112080922, 
	DOUT7 => N112080923, 
	DOUT8 => N112080924, 
	DOUT9 => N112080925, 
	DOUT10 => N112080926, 
	DOUT11 => N112080927, 
	DOUT12 => N112080928, 
	DOUT13 => N112080929, 
	DOUT14 => N112080930, 
	DOUT15 => N112080931, 
	SIGNEDIN => N111619233, 
	SIGNEDOUT => N112080933
);
U192 : ADDERDELAY	PORT MAP(
	DIN0 => N113729316, 
	DIN1 => N113729317, 
	DIN2 => N113729318, 
	DIN3 => N113729319, 
	DIN4 => N113729320, 
	DIN5 => N113729321, 
	DIN6 => N113729322, 
	DIN7 => N113729323, 
	DIN8 => N113729324, 
	DIN9 => N113729325, 
	DIN10 => N113729326, 
	DIN11 => N113729327, 
	DIN12 => N113729328, 
	DIN13 => N113729329, 
	DIN14 => N113729330, 
	DIN15 => N113729331, 
	DOUT0 => N113753616, 
	DOUT1 => N113753617, 
	DOUT2 => N113753618, 
	DOUT3 => N113753619, 
	DOUT4 => N113753620, 
	DOUT5 => N113753621, 
	DOUT6 => N113753622, 
	DOUT7 => N113753623, 
	DOUT8 => N113753624, 
	DOUT9 => N113753625, 
	DOUT10 => N113753626, 
	DOUT11 => N113753627, 
	DOUT12 => N113753628, 
	DOUT13 => N113753629, 
	DOUT14 => N113753630, 
	DOUT15 => N113753631, 
	SIGNEDIN => N113729333, 
	SIGNEDOUT => N113753633
);
U161 : ADDERDELAY	PORT MAP(
	DIN0 => N112080916, 
	DIN1 => N112080917, 
	DIN2 => N112080918, 
	DIN3 => N112080919, 
	DIN4 => N112080920, 
	DIN5 => N112080921, 
	DIN6 => N112080922, 
	DIN7 => N112080923, 
	DIN8 => N112080924, 
	DIN9 => N112080925, 
	DIN10 => N112080926, 
	DIN11 => N112080927, 
	DIN12 => N112080928, 
	DIN13 => N112080929, 
	DIN14 => N112080930, 
	DIN15 => N112080931, 
	DOUT0 => N112105216, 
	DOUT1 => N112105217, 
	DOUT2 => N112105218, 
	DOUT3 => N112105219, 
	DOUT4 => N112105220, 
	DOUT5 => N112105221, 
	DOUT6 => N112105222, 
	DOUT7 => N112105223, 
	DOUT8 => N112105224, 
	DOUT9 => N112105225, 
	DOUT10 => N112105226, 
	DOUT11 => N112105227, 
	DOUT12 => N112105228, 
	DOUT13 => N112105229, 
	DOUT14 => N112105230, 
	DOUT15 => N112105231, 
	SIGNEDIN => N112080933, 
	SIGNEDOUT => N112105233
);
U193 : \16adderBalanced\	PORT MAP(
	A0 => N1147650, 
	A1 => N1147610, 
	A2 => N1147646, 
	A3 => N1147618, 
	A4 => N1147602, 
	A5 => N1147630, 
	A6 => N1147658, 
	A7 => N1147654, 
	A8 => N1147638, 
	A9 => N1147626, 
	A10 => N1147642, 
	A11 => N1147634, 
	A12 => N1147614, 
	A13 => N1147622, 
	A14 => N1147594, 
	A15 => N1147598, 
	B0 => TF0, 
	B1 => TF1, 
	B2 => TF2, 
	B3 => TF3, 
	B4 => TF4, 
	B5 => TF5, 
	B6 => TF6, 
	B7 => TF7, 
	B8 => TF8, 
	B9 => TF9, 
	B10 => TF10, 
	B11 => TF11, 
	B12 => TF12, 
	B13 => TF13, 
	B14 => TF14, 
	B15 => TF15, 
	CIN => N1147606, 
	COUT => N1057701, 
	Y0 => N107806, 
	Y1 => N108278, 
	Y2 => N107814, 
	Y3 => N108286, 
	Y4 => N108274, 
	Y5 => N107822, 
	Y6 => N107810, 
	Y7 => N108282, 
	Y8 => N108270, 
	Y9 => N108266, 
	Y10 => N108262, 
	Y11 => N108258, 
	Y12 => N108254, 
	Y13 => N107826, 
	Y14 => N107830, 
	Y15 => N107818
);
U194 : \16adderBalanced\	PORT MAP(
	A0 => N1147328, 
	A1 => N1147288, 
	A2 => N1147324, 
	A3 => N1147296, 
	A4 => N1147280, 
	A5 => N1147308, 
	A6 => N1147336, 
	A7 => N1147332, 
	A8 => N1147316, 
	A9 => N1147304, 
	A10 => N1147320, 
	A11 => N1147312, 
	A12 => N1147292, 
	A13 => N1147300, 
	A14 => N1147272, 
	A15 => N1147276, 
	B0 => TE0, 
	B1 => TE1, 
	B2 => TE2, 
	B3 => TE3, 
	B4 => TE4, 
	B5 => TE5, 
	B6 => TE6, 
	B7 => TE7, 
	B8 => TE8, 
	B9 => TE9, 
	B10 => TE10, 
	B11 => TE11, 
	B12 => TE12, 
	B13 => TE13, 
	B14 => TE14, 
	B15 => TE15, 
	CIN => N1147284, 
	COUT => N1058015, 
	Y0 => N103455, 
	Y1 => N103927, 
	Y2 => N103463, 
	Y3 => N103935, 
	Y4 => N103923, 
	Y5 => N103471, 
	Y6 => N103459, 
	Y7 => N103931, 
	Y8 => N103919, 
	Y9 => N103915, 
	Y10 => N103911, 
	Y11 => N103907, 
	Y12 => N103903, 
	Y13 => N103475, 
	Y14 => N103479, 
	Y15 => N103467
);
U130 : ADDERDELAY	PORT MAP(
	DIN0 => N110601616, 
	DIN1 => N110601617, 
	DIN2 => N110601618, 
	DIN3 => N110601619, 
	DIN4 => N110601620, 
	DIN5 => N110601621, 
	DIN6 => N110601622, 
	DIN7 => N110601623, 
	DIN8 => N110601624, 
	DIN9 => N110601625, 
	DIN10 => N110601626, 
	DIN11 => N110601627, 
	DIN12 => N110601628, 
	DIN13 => N110601629, 
	DIN14 => N110601630, 
	DIN15 => N110601631, 
	DOUT0 => N111336716, 
	DOUT1 => N111336717, 
	DOUT2 => N111336718, 
	DOUT3 => N111336719, 
	DOUT4 => N111336720, 
	DOUT5 => N111336721, 
	DOUT6 => N111336722, 
	DOUT7 => N111336723, 
	DOUT8 => N111336724, 
	DOUT9 => N111336725, 
	DOUT10 => N111336726, 
	DOUT11 => N111336727, 
	DOUT12 => N111336728, 
	DOUT13 => N111336729, 
	DOUT14 => N111336730, 
	DOUT15 => N111336731, 
	SIGNEDIN => N110601633, 
	SIGNEDOUT => N111336733
);
U162 : ADDERDELAY	PORT MAP(
	DIN0 => N112105216, 
	DIN1 => N112105217, 
	DIN2 => N112105218, 
	DIN3 => N112105219, 
	DIN4 => N112105220, 
	DIN5 => N112105221, 
	DIN6 => N112105222, 
	DIN7 => N112105223, 
	DIN8 => N112105224, 
	DIN9 => N112105225, 
	DIN10 => N112105226, 
	DIN11 => N112105227, 
	DIN12 => N112105228, 
	DIN13 => N112105229, 
	DIN14 => N112105230, 
	DIN15 => N112105231, 
	DOUT0 => N1147328, 
	DOUT1 => N1147288, 
	DOUT2 => N1147324, 
	DOUT3 => N1147296, 
	DOUT4 => N1147280, 
	DOUT5 => N1147308, 
	DOUT6 => N1147336, 
	DOUT7 => N1147332, 
	DOUT8 => N1147316, 
	DOUT9 => N1147304, 
	DOUT10 => N1147320, 
	DOUT11 => N1147312, 
	DOUT12 => N1147292, 
	DOUT13 => N1147300, 
	DOUT14 => N1147272, 
	DOUT15 => N1147276, 
	SIGNEDIN => N112105233, 
	SIGNEDOUT => N1147284
);
U131 : ADDERDELAY	PORT MAP(
	DIN0 => N111336716, 
	DIN1 => N111336717, 
	DIN2 => N111336718, 
	DIN3 => N111336719, 
	DIN4 => N111336720, 
	DIN5 => N111336721, 
	DIN6 => N111336722, 
	DIN7 => N111336723, 
	DIN8 => N111336724, 
	DIN9 => N111336725, 
	DIN10 => N111336726, 
	DIN11 => N111336727, 
	DIN12 => N111336728, 
	DIN13 => N111336729, 
	DIN14 => N111336730, 
	DIN15 => N111336731, 
	DOUT0 => N111361016, 
	DOUT1 => N111361017, 
	DOUT2 => N111361018, 
	DOUT3 => N111361019, 
	DOUT4 => N111361020, 
	DOUT5 => N111361021, 
	DOUT6 => N111361022, 
	DOUT7 => N111361023, 
	DOUT8 => N111361024, 
	DOUT9 => N111361025, 
	DOUT10 => N111361026, 
	DOUT11 => N111361027, 
	DOUT12 => N111361028, 
	DOUT13 => N111361029, 
	DOUT14 => N111361030, 
	DOUT15 => N111361031, 
	SIGNEDIN => N111336733, 
	SIGNEDOUT => N111361033
);
U163 : ADDERDELAY	PORT MAP(
	DIN0 => N111692116, 
	DIN1 => N111692117, 
	DIN2 => N111692118, 
	DIN3 => N111692119, 
	DIN4 => N111692120, 
	DIN5 => N111692121, 
	DIN6 => N111692122, 
	DIN7 => N111692123, 
	DIN8 => N111692124, 
	DIN9 => N111692125, 
	DIN10 => N111692126, 
	DIN11 => N111692127, 
	DIN12 => N111692128, 
	DIN13 => N111692129, 
	DIN14 => N111692130, 
	DIN15 => N111692131, 
	DOUT0 => N112153816, 
	DOUT1 => N112153817, 
	DOUT2 => N112153818, 
	DOUT3 => N112153819, 
	DOUT4 => N112153820, 
	DOUT5 => N112153821, 
	DOUT6 => N112153822, 
	DOUT7 => N112153823, 
	DOUT8 => N112153824, 
	DOUT9 => N112153825, 
	DOUT10 => N112153826, 
	DOUT11 => N112153827, 
	DOUT12 => N112153828, 
	DOUT13 => N112153829, 
	DOUT14 => N112153830, 
	DOUT15 => N112153831, 
	SIGNEDIN => N111692133, 
	SIGNEDOUT => N112153833
);
U195 : \16adderBalanced\	PORT MAP(
	A0 => N1147006, 
	A1 => N1146966, 
	A2 => N1147002, 
	A3 => N1146974, 
	A4 => N1146958, 
	A5 => N1146986, 
	A6 => N1147014, 
	A7 => N1147010, 
	A8 => N1146994, 
	A9 => N1146982, 
	A10 => N1146998, 
	A11 => N1146990, 
	A12 => N1146970, 
	A13 => N1146978, 
	A14 => N1146950, 
	A15 => N1146954, 
	B0 => TD0, 
	B1 => TD1, 
	B2 => TD2, 
	B3 => TD3, 
	B4 => TD4, 
	B5 => TD5, 
	B6 => TD6, 
	B7 => TD7, 
	B8 => TD8, 
	B9 => TD9, 
	B10 => TD10, 
	B11 => TD11, 
	B12 => TD12, 
	B13 => TD13, 
	B14 => TD14, 
	B15 => TD15, 
	CIN => N1146962, 
	COUT => N1058329, 
	Y0 => N102421, 
	Y1 => N102893, 
	Y2 => N102429, 
	Y3 => N102901, 
	Y4 => N102889, 
	Y5 => N102437, 
	Y6 => N102425, 
	Y7 => N102897, 
	Y8 => N102885, 
	Y9 => N102881, 
	Y10 => N102877, 
	Y11 => N102873, 
	Y12 => N102869, 
	Y13 => N102441, 
	Y14 => N102445, 
	Y15 => N102433
);
U132 : ADDERDELAY	PORT MAP(
	DIN0 => N111361016, 
	DIN1 => N111361017, 
	DIN2 => N111361018, 
	DIN3 => N111361019, 
	DIN4 => N111361020, 
	DIN5 => N111361021, 
	DIN6 => N111361022, 
	DIN7 => N111361023, 
	DIN8 => N111361024, 
	DIN9 => N111361025, 
	DIN10 => N111361026, 
	DIN11 => N111361027, 
	DIN12 => N111361028, 
	DIN13 => N111361029, 
	DIN14 => N111361030, 
	DIN15 => N111361031, 
	DOUT0 => N1146845, 
	DOUT1 => N1146805, 
	DOUT2 => N1146841, 
	DOUT3 => N1146813, 
	DOUT4 => N1146797, 
	DOUT5 => N1146825, 
	DOUT6 => N1146853, 
	DOUT7 => N1146849, 
	DOUT8 => N1146833, 
	DOUT9 => N1146821, 
	DOUT10 => N1146837, 
	DOUT11 => N1146829, 
	DOUT12 => N1146809, 
	DOUT13 => N1146817, 
	DOUT14 => N1146789, 
	DOUT15 => N1146793, 
	SIGNEDIN => N111361033, 
	SIGNEDOUT => N1146801
);
U164 : ADDERDELAY	PORT MAP(
	DIN0 => N112153816, 
	DIN1 => N112153817, 
	DIN2 => N112153818, 
	DIN3 => N112153819, 
	DIN4 => N112153820, 
	DIN5 => N112153821, 
	DIN6 => N112153822, 
	DIN7 => N112153823, 
	DIN8 => N112153824, 
	DIN9 => N112153825, 
	DIN10 => N112153826, 
	DIN11 => N112153827, 
	DIN12 => N112153828, 
	DIN13 => N112153829, 
	DIN14 => N112153830, 
	DIN15 => N112153831, 
	DOUT0 => N112178116, 
	DOUT1 => N112178117, 
	DOUT2 => N112178118, 
	DOUT3 => N112178119, 
	DOUT4 => N112178120, 
	DOUT5 => N112178121, 
	DOUT6 => N112178122, 
	DOUT7 => N112178123, 
	DOUT8 => N112178124, 
	DOUT9 => N112178125, 
	DOUT10 => N112178126, 
	DOUT11 => N112178127, 
	DOUT12 => N112178128, 
	DOUT13 => N112178129, 
	DOUT14 => N112178130, 
	DOUT15 => N112178131, 
	SIGNEDIN => N112153833, 
	SIGNEDOUT => N112178133
);
U100 : ADDERDELAY	PORT MAP(
	DIN0 => N110549216, 
	DIN1 => N110549217, 
	DIN2 => N110549218, 
	DIN3 => N110549219, 
	DIN4 => N110549220, 
	DIN5 => N110549221, 
	DIN6 => N110549222, 
	DIN7 => N110549223, 
	DIN8 => N110549224, 
	DIN9 => N110549225, 
	DIN10 => N110549226, 
	DIN11 => N110549227, 
	DIN12 => N110549228, 
	DIN13 => N110549229, 
	DIN14 => N110549230, 
	DIN15 => N110549231, 
	DOUT0 => N110577316, 
	DOUT1 => N110577317, 
	DOUT2 => N110577318, 
	DOUT3 => N110577319, 
	DOUT4 => N110577320, 
	DOUT5 => N110577321, 
	DOUT6 => N110577322, 
	DOUT7 => N110577323, 
	DOUT8 => N110577324, 
	DOUT9 => N110577325, 
	DOUT10 => N110577326, 
	DOUT11 => N110577327, 
	DOUT12 => N110577328, 
	DOUT13 => N110577329, 
	DOUT14 => N110577330, 
	DOUT15 => N110577331, 
	SIGNEDIN => N110549233, 
	SIGNEDOUT => N110577333
);
U196 : \16adderBalanced\	PORT MAP(
	A0 => N1146684, 
	A1 => N1146644, 
	A2 => N1146680, 
	A3 => N1146652, 
	A4 => N1146636, 
	A5 => N1146664, 
	A6 => N1146692, 
	A7 => N1146688, 
	A8 => N1146672, 
	A9 => N1146660, 
	A10 => N1146676, 
	A11 => N1146668, 
	A12 => N1146648, 
	A13 => N1146656, 
	A14 => N1146628, 
	A15 => N1146632, 
	B0 => TC0, 
	B1 => TC1, 
	B2 => TC2, 
	B3 => TC3, 
	B4 => TC4, 
	B5 => TC5, 
	B6 => TC6, 
	B7 => TC7, 
	B8 => TC8, 
	B9 => TC9, 
	B10 => TC10, 
	B11 => TC11, 
	B12 => TC12, 
	B13 => TC13, 
	B14 => TC14, 
	B15 => TC15, 
	CIN => N1146640, 
	COUT => N1058643, 
	Y0 => N100889, 
	Y1 => N101361, 
	Y2 => N100897, 
	Y3 => N101369, 
	Y4 => N101357, 
	Y5 => N100905, 
	Y6 => N100893, 
	Y7 => N101365, 
	Y8 => N101353, 
	Y9 => N101349, 
	Y10 => N101345, 
	Y11 => N101341, 
	Y12 => N101337, 
	Y13 => N100909, 
	Y14 => N100913, 
	Y15 => N100901
);
U165 : ADDERDELAY	PORT MAP(
	DIN0 => N112178116, 
	DIN1 => N112178117, 
	DIN2 => N112178118, 
	DIN3 => N112178119, 
	DIN4 => N112178120, 
	DIN5 => N112178121, 
	DIN6 => N112178122, 
	DIN7 => N112178123, 
	DIN8 => N112178124, 
	DIN9 => N112178125, 
	DIN10 => N112178126, 
	DIN11 => N112178127, 
	DIN12 => N112178128, 
	DIN13 => N112178129, 
	DIN14 => N112178130, 
	DIN15 => N112178131, 
	DOUT0 => N112202416, 
	DOUT1 => N112202417, 
	DOUT2 => N112202418, 
	DOUT3 => N112202419, 
	DOUT4 => N112202420, 
	DOUT5 => N112202421, 
	DOUT6 => N112202422, 
	DOUT7 => N112202423, 
	DOUT8 => N112202424, 
	DOUT9 => N112202425, 
	DOUT10 => N112202426, 
	DOUT11 => N112202427, 
	DOUT12 => N112202428, 
	DOUT13 => N112202429, 
	DOUT14 => N112202430, 
	DOUT15 => N112202431, 
	SIGNEDIN => N112178133, 
	SIGNEDOUT => N112202433
);
U197 : \16adderBalanced\	PORT MAP(
	A0 => N1145131, 
	A1 => N1145091, 
	A2 => N1145127, 
	A3 => N1145099, 
	A4 => N1145083, 
	A5 => N1145111, 
	A6 => N1145139, 
	A7 => N1145135, 
	A8 => N1145119, 
	A9 => N1145107, 
	A10 => N1145123, 
	A11 => N1145115, 
	A12 => N1145095, 
	A13 => N1145103, 
	A14 => N1145075, 
	A15 => N1145079, 
	B0 => TB0, 
	B1 => TB1, 
	B2 => TB2, 
	B3 => TB3, 
	B4 => TB4, 
	B5 => TB5, 
	B6 => TB6, 
	B7 => TB7, 
	B8 => TB8, 
	B9 => TB9, 
	B10 => TB10, 
	B11 => TB11, 
	B12 => TB12, 
	B13 => TB13, 
	B14 => TB14, 
	B15 => TB15, 
	CIN => N1145087, 
	COUT => N1066581, 
	Y0 => N91218, 
	Y1 => N91220, 
	Y2 => N91190, 
	Y3 => N91192, 
	Y4 => N91194, 
	Y5 => N91196, 
	Y6 => N91198, 
	Y7 => N91200, 
	Y8 => N91202, 
	Y9 => N91204, 
	Y10 => N91206, 
	Y11 => N91208, 
	Y12 => N91210, 
	Y13 => N91212, 
	Y14 => N91214, 
	Y15 => N91216
);
U133 : ADDERDELAY	PORT MAP(
	DIN0 => N110678316, 
	DIN1 => N110678317, 
	DIN2 => N110678318, 
	DIN3 => N110678319, 
	DIN4 => N110678320, 
	DIN5 => N110678321, 
	DIN6 => N110678322, 
	DIN7 => N110678323, 
	DIN8 => N110678324, 
	DIN9 => N110678325, 
	DIN10 => N110678326, 
	DIN11 => N110678327, 
	DIN12 => N110678328, 
	DIN13 => N110678329, 
	DIN14 => N110678330, 
	DIN15 => N110678331, 
	DOUT0 => N111424816, 
	DOUT1 => N111424817, 
	DOUT2 => N111424818, 
	DOUT3 => N111424819, 
	DOUT4 => N111424820, 
	DOUT5 => N111424821, 
	DOUT6 => N111424822, 
	DOUT7 => N111424823, 
	DOUT8 => N111424824, 
	DOUT9 => N111424825, 
	DOUT10 => N111424826, 
	DOUT11 => N111424827, 
	DOUT12 => N111424828, 
	DOUT13 => N111424829, 
	DOUT14 => N111424830, 
	DOUT15 => N111424831, 
	SIGNEDIN => N110678333, 
	SIGNEDOUT => N111424833
);
U101 : ADDERDELAY	PORT MAP(
	DIN0 => N110577316, 
	DIN1 => N110577317, 
	DIN2 => N110577318, 
	DIN3 => N110577319, 
	DIN4 => N110577320, 
	DIN5 => N110577321, 
	DIN6 => N110577322, 
	DIN7 => N110577323, 
	DIN8 => N110577324, 
	DIN9 => N110577325, 
	DIN10 => N110577326, 
	DIN11 => N110577327, 
	DIN12 => N110577328, 
	DIN13 => N110577329, 
	DIN14 => N110577330, 
	DIN15 => N110577331, 
	DOUT0 => N110601616, 
	DOUT1 => N110601617, 
	DOUT2 => N110601618, 
	DOUT3 => N110601619, 
	DOUT4 => N110601620, 
	DOUT5 => N110601621, 
	DOUT6 => N110601622, 
	DOUT7 => N110601623, 
	DOUT8 => N110601624, 
	DOUT9 => N110601625, 
	DOUT10 => N110601626, 
	DOUT11 => N110601627, 
	DOUT12 => N110601628, 
	DOUT13 => N110601629, 
	DOUT14 => N110601630, 
	DOUT15 => N110601631, 
	SIGNEDIN => N110577333, 
	SIGNEDOUT => N110601633
);
U198 : \16adderBalanced\	PORT MAP(
	A0 => N1143146, 
	A1 => N1143067, 
	A2 => N1142988, 
	A3 => N1142909, 
	A4 => N1142830, 
	A5 => N1142751, 
	A6 => N1142672, 
	A7 => N1142593, 
	A8 => N1142514, 
	A9 => N1142435, 
	A10 => N1142356, 
	A11 => N1142277, 
	A12 => N1142198, 
	A13 => N1142119, 
	A14 => N1142040, 
	A15 => N1141961, 
	B0 => TA0, 
	B1 => TA1, 
	B2 => TA2, 
	B3 => TA3, 
	B4 => TA4, 
	B5 => TA5, 
	B6 => TA6, 
	B7 => TA7, 
	B8 => TA8, 
	B9 => TA9, 
	B10 => TA10, 
	B11 => TA11, 
	B12 => TA12, 
	B13 => TA13, 
	B14 => TA14, 
	B15 => TA15, 
	CIN => N1141882, 
	COUT => N1063489, 
	Y0 => N99924, 
	Y1 => N100396, 
	Y2 => N99932, 
	Y3 => N100404, 
	Y4 => N100392, 
	Y5 => N99940, 
	Y6 => N99928, 
	Y7 => N100400, 
	Y8 => N100388, 
	Y9 => N100384, 
	Y10 => N100380, 
	Y11 => N100376, 
	Y12 => N100372, 
	Y13 => N99944, 
	Y14 => N99948, 
	Y15 => N99936
);
U166 : ADDERDELAY	PORT MAP(
	DIN0 => N112202416, 
	DIN1 => N112202417, 
	DIN2 => N112202418, 
	DIN3 => N112202419, 
	DIN4 => N112202420, 
	DIN5 => N112202421, 
	DIN6 => N112202422, 
	DIN7 => N112202423, 
	DIN8 => N112202424, 
	DIN9 => N112202425, 
	DIN10 => N112202426, 
	DIN11 => N112202427, 
	DIN12 => N112202428, 
	DIN13 => N112202429, 
	DIN14 => N112202430, 
	DIN15 => N112202431, 
	DOUT0 => N1147489, 
	DOUT1 => N1147449, 
	DOUT2 => N1147485, 
	DOUT3 => N1147457, 
	DOUT4 => N1147441, 
	DOUT5 => N1147469, 
	DOUT6 => N1147497, 
	DOUT7 => N1147493, 
	DOUT8 => N1147477, 
	DOUT9 => N1147465, 
	DOUT10 => N1268884, 
	DOUT11 => N1257378, 
	DOUT12 => N1147453, 
	DOUT13 => N1147461, 
	DOUT14 => N1147433, 
	DOUT15 => N1147437, 
	SIGNEDIN => N112202433, 
	SIGNEDOUT => N1147445
);
U134 : ADDERDELAY	PORT MAP(
	DIN0 => N111424816, 
	DIN1 => N111424817, 
	DIN2 => N111424818, 
	DIN3 => N111424819, 
	DIN4 => N111424820, 
	DIN5 => N111424821, 
	DIN6 => N111424822, 
	DIN7 => N111424823, 
	DIN8 => N111424824, 
	DIN9 => N111424825, 
	DIN10 => N111424826, 
	DIN11 => N111424827, 
	DIN12 => N111424828, 
	DIN13 => N111424829, 
	DIN14 => N111424830, 
	DIN15 => N111424831, 
	DOUT0 => N111449116, 
	DOUT1 => N111449117, 
	DOUT2 => N111449118, 
	DOUT3 => N111449119, 
	DOUT4 => N111449120, 
	DOUT5 => N111449121, 
	DOUT6 => N111449122, 
	DOUT7 => N111449123, 
	DOUT8 => N111449124, 
	DOUT9 => N111449125, 
	DOUT10 => N111449126, 
	DOUT11 => N111449127, 
	DOUT12 => N111449128, 
	DOUT13 => N111449129, 
	DOUT14 => N111449130, 
	DOUT15 => N111449131, 
	SIGNEDIN => N111424833, 
	SIGNEDOUT => N111449133
);
U102 : ADDERDELAY	PORT MAP(
	DIN0 => N11062590, 
	DIN1 => N11062591, 
	DIN2 => N11062592, 
	DIN3 => N11062593, 
	DIN4 => N11062594, 
	DIN5 => N11062595, 
	DIN6 => N11062596, 
	DIN7 => N11062597, 
	DIN8 => N11062598, 
	DIN9 => N11062599, 
	DIN10 => N110625910, 
	DIN11 => N110625911, 
	DIN12 => N110625912, 
	DIN13 => N110625913, 
	DIN14 => N110625914, 
	DIN15 => N110625915, 
	DOUT0 => N110625916, 
	DOUT1 => N110625917, 
	DOUT2 => N110625918, 
	DOUT3 => N110625919, 
	DOUT4 => N110625920, 
	DOUT5 => N110625921, 
	DOUT6 => N110625922, 
	DOUT7 => N110625923, 
	DOUT8 => N110625924, 
	DOUT9 => N110625925, 
	DOUT10 => N110625926, 
	DOUT11 => N110625927, 
	DOUT12 => N110625928, 
	DOUT13 => N110625929, 
	DOUT14 => N110625930, 
	DOUT15 => N110625931, 
	SIGNEDIN => N110625932, 
	SIGNEDOUT => N110625933
);
U167 : ADDERDELAY	PORT MAP(
	DIN0 => N111765016, 
	DIN1 => N111765017, 
	DIN2 => N111765018, 
	DIN3 => N111765019, 
	DIN4 => N111765020, 
	DIN5 => N111765021, 
	DIN6 => N111765022, 
	DIN7 => N111765023, 
	DIN8 => N111765024, 
	DIN9 => N111765025, 
	DIN10 => N111765026, 
	DIN11 => N111765027, 
	DIN12 => N111765028, 
	DIN13 => N111765029, 
	DIN14 => N111765030, 
	DIN15 => N111765031, 
	DOUT0 => N112251016, 
	DOUT1 => N112251017, 
	DOUT2 => N112251018, 
	DOUT3 => N112251019, 
	DOUT4 => N112251020, 
	DOUT5 => N112251021, 
	DOUT6 => N112251022, 
	DOUT7 => N112251023, 
	DOUT8 => N112251024, 
	DOUT9 => N112251025, 
	DOUT10 => N112251026, 
	DOUT11 => N112251027, 
	DOUT12 => N112251028, 
	DOUT13 => N112251029, 
	DOUT14 => N112251030, 
	DOUT15 => N112251031, 
	SIGNEDIN => N111765033, 
	SIGNEDOUT => N112251033
);
U103 : ADDERDELAY	PORT MAP(
	DIN0 => N110625916, 
	DIN1 => N110625917, 
	DIN2 => N110625918, 
	DIN3 => N110625919, 
	DIN4 => N110625920, 
	DIN5 => N110625921, 
	DIN6 => N110625922, 
	DIN7 => N110625923, 
	DIN8 => N110625924, 
	DIN9 => N110625925, 
	DIN10 => N110625926, 
	DIN11 => N110625927, 
	DIN12 => N110625928, 
	DIN13 => N110625929, 
	DIN14 => N110625930, 
	DIN15 => N110625931, 
	DOUT0 => N110654016, 
	DOUT1 => N110654017, 
	DOUT2 => N110654018, 
	DOUT3 => N110654019, 
	DOUT4 => N110654020, 
	DOUT5 => N110654021, 
	DOUT6 => N110654022, 
	DOUT7 => N110654023, 
	DOUT8 => N110654024, 
	DOUT9 => N110654025, 
	DOUT10 => N110654026, 
	DOUT11 => N110654027, 
	DOUT12 => N110654028, 
	DOUT13 => N110654029, 
	DOUT14 => N110654030, 
	DOUT15 => N110654031, 
	SIGNEDIN => N110625933, 
	SIGNEDOUT => N110654033
);
U135 : ADDERDELAY	PORT MAP(
	DIN0 => N111449116, 
	DIN1 => N111449117, 
	DIN2 => N111449118, 
	DIN3 => N111449119, 
	DIN4 => N111449120, 
	DIN5 => N111449121, 
	DIN6 => N111449122, 
	DIN7 => N111449123, 
	DIN8 => N111449124, 
	DIN9 => N111449125, 
	DIN10 => N111449126, 
	DIN11 => N111449127, 
	DIN12 => N111449128, 
	DIN13 => N111449129, 
	DIN14 => N111449130, 
	DIN15 => N111449131, 
	DOUT0 => N111473416, 
	DOUT1 => N111473417, 
	DOUT2 => N111473418, 
	DOUT3 => N111473419, 
	DOUT4 => N111473420, 
	DOUT5 => N111473421, 
	DOUT6 => N111473422, 
	DOUT7 => N111473423, 
	DOUT8 => N111473424, 
	DOUT9 => N111473425, 
	DOUT10 => N111473426, 
	DOUT11 => N111473427, 
	DOUT12 => N111473428, 
	DOUT13 => N111473429, 
	DOUT14 => N111473430, 
	DOUT15 => N111473431, 
	SIGNEDIN => N111449133, 
	SIGNEDOUT => N111473433
);
U199 : TAPADDER	PORT MAP(
	A0 => N113753616, 
	A1 => N113753617, 
	A2 => N113753618, 
	A3 => N113753619, 
	A4 => N113753620, 
	A5 => N113753621, 
	A6 => N113753622, 
	A7 => N113753623, 
	A8 => N113753624, 
	A9 => N113753625, 
	A10 => N113753626, 
	A11 => N113753627, 
	A12 => N113753628, 
	A13 => N113753629, 
	A14 => N113753630, 
	A15 => N113753631, 
	AND1 => N94145, 
	AND2 => N94147, 
	AND3 => N94157, 
	B0 => N108992, 
	B1 => N109348, 
	B2 => N109000, 
	B3 => N109356, 
	B4 => N109344, 
	B5 => N109008, 
	B6 => N108996, 
	B7 => N109352, 
	B8 => N109340, 
	B9 => N109336, 
	B10 => N109332, 
	B11 => N109328, 
	B12 => N109324, 
	B13 => N109012, 
	B14 => N109016, 
	B15 => N109004, 
	CIN => N113753633, 
	COUT => MONITOR16, 
	O0 => H0, 
	O1 => H1, 
	O2 => H2, 
	O3 => H3, 
	O4 => H4, 
	O5 => H5, 
	O6 => H6, 
	O7 => H7, 
	O8 => H8, 
	O9 => H9, 
	O10 => H10, 
	O11 => H11, 
	O12 => H12, 
	O13 => H13, 
	O14 => H14, 
	O15 => H15, 
	OR1 => N94153, 
	OR2 => N94155, 
	OR3 => N94149, 
	Y0 => MONITOR0, 
	Y1 => MONITOR1, 
	Y2 => MONITOR2, 
	Y3 => MONITOR3, 
	Y4 => MONITOR4, 
	Y5 => MONITOR5, 
	Y6 => MONITOR6, 
	Y7 => MONITOR7, 
	Y8 => MONITOR8, 
	Y9 => MONITOR9, 
	Y10 => MONITOR10, 
	Y11 => MONITOR11, 
	Y12 => MONITOR12, 
	Y13 => MONITOR13, 
	Y14 => MONITOR14, 
	Y15 => MONITOR15
);
U168 : ADDERDELAY	PORT MAP(
	DIN0 => N112251016, 
	DIN1 => N112251017, 
	DIN2 => N112251018, 
	DIN3 => N112251019, 
	DIN4 => N112251020, 
	DIN5 => N112251021, 
	DIN6 => N112251022, 
	DIN7 => N112251023, 
	DIN8 => N112251024, 
	DIN9 => N112251025, 
	DIN10 => N112251026, 
	DIN11 => N112251027, 
	DIN12 => N112251028, 
	DIN13 => N112251029, 
	DIN14 => N112251030, 
	DIN15 => N112251031, 
	DOUT0 => N112275316, 
	DOUT1 => N112275317, 
	DOUT2 => N112275318, 
	DOUT3 => N112275319, 
	DOUT4 => N112275320, 
	DOUT5 => N112275321, 
	DOUT6 => N112275322, 
	DOUT7 => N112275323, 
	DOUT8 => N112275324, 
	DOUT9 => N112275325, 
	DOUT10 => N112275326, 
	DOUT11 => N112275327, 
	DOUT12 => N112275328, 
	DOUT13 => N112275329, 
	DOUT14 => N112275330, 
	DOUT15 => N112275331, 
	SIGNEDIN => N112251033, 
	SIGNEDOUT => N112275333
);
U104 : ADDERDELAY	PORT MAP(
	DIN0 => N110654016, 
	DIN1 => N110654017, 
	DIN2 => N110654018, 
	DIN3 => N110654019, 
	DIN4 => N110654020, 
	DIN5 => N110654021, 
	DIN6 => N110654022, 
	DIN7 => N110654023, 
	DIN8 => N110654024, 
	DIN9 => N110654025, 
	DIN10 => N110654026, 
	DIN11 => N110654027, 
	DIN12 => N110654028, 
	DIN13 => N110654029, 
	DIN14 => N110654030, 
	DIN15 => N110654031, 
	DOUT0 => N110678316, 
	DOUT1 => N110678317, 
	DOUT2 => N110678318, 
	DOUT3 => N110678319, 
	DOUT4 => N110678320, 
	DOUT5 => N110678321, 
	DOUT6 => N110678322, 
	DOUT7 => N110678323, 
	DOUT8 => N110678324, 
	DOUT9 => N110678325, 
	DOUT10 => N110678326, 
	DOUT11 => N110678327, 
	DOUT12 => N110678328, 
	DOUT13 => N110678329, 
	DOUT14 => N110678330, 
	DOUT15 => N110678331, 
	SIGNEDIN => N110654033, 
	SIGNEDOUT => N110678333
);
U136 : ADDERDELAY	PORT MAP(
	DIN0 => N110755016, 
	DIN1 => N110755017, 
	DIN2 => N110755018, 
	DIN3 => N110755019, 
	DIN4 => N110755020, 
	DIN5 => N110755021, 
	DIN6 => N110755022, 
	DIN7 => N110755023, 
	DIN8 => N110755024, 
	DIN9 => N110755025, 
	DIN10 => N110755026, 
	DIN11 => N110755027, 
	DIN12 => N110755028, 
	DIN13 => N110755029, 
	DIN14 => N110755030, 
	DIN15 => N110755031, 
	DOUT0 => N111497716, 
	DOUT1 => N111497717, 
	DOUT2 => N111497718, 
	DOUT3 => N111497719, 
	DOUT4 => N111497720, 
	DOUT5 => N111497721, 
	DOUT6 => N111497722, 
	DOUT7 => N111497723, 
	DOUT8 => N111497724, 
	DOUT9 => N111497725, 
	DOUT10 => N111497726, 
	DOUT11 => N111497727, 
	DOUT12 => N111497728, 
	DOUT13 => N111497729, 
	DOUT14 => N111497730, 
	DOUT15 => N111497731, 
	SIGNEDIN => N110755033, 
	SIGNEDOUT => N111497733
);
U169 : ADDERDELAY	PORT MAP(
	DIN0 => N112275316, 
	DIN1 => N112275317, 
	DIN2 => N112275318, 
	DIN3 => N112275319, 
	DIN4 => N112275320, 
	DIN5 => N112275321, 
	DIN6 => N112275322, 
	DIN7 => N112275323, 
	DIN8 => N112275324, 
	DIN9 => N112275325, 
	DIN10 => N112275326, 
	DIN11 => N112275327, 
	DIN12 => N112275328, 
	DIN13 => N112275329, 
	DIN14 => N112275330, 
	DIN15 => N112275331, 
	DOUT0 => N112299616, 
	DOUT1 => N112299617, 
	DOUT2 => N112299618, 
	DOUT3 => N112299619, 
	DOUT4 => N112299620, 
	DOUT5 => N112299621, 
	DOUT6 => N112299622, 
	DOUT7 => N112299623, 
	DOUT8 => N112299624, 
	DOUT9 => N112299625, 
	DOUT10 => N112299626, 
	DOUT11 => N112299627, 
	DOUT12 => N112299628, 
	DOUT13 => N112299629, 
	DOUT14 => N112299630, 
	DOUT15 => N112299631, 
	SIGNEDIN => N112275333, 
	SIGNEDOUT => N112299633
);
U105 : ADDERDELAY	PORT MAP(
	DIN0 => N11070260, 
	DIN1 => N11070261, 
	DIN2 => N11070262, 
	DIN3 => N11070263, 
	DIN4 => N11070264, 
	DIN5 => N11070265, 
	DIN6 => N11070266, 
	DIN7 => N11070267, 
	DIN8 => N11070268, 
	DIN9 => N11070269, 
	DIN10 => N110702610, 
	DIN11 => N110702611, 
	DIN12 => N110702612, 
	DIN13 => N110702613, 
	DIN14 => N110702614, 
	DIN15 => N110702615, 
	DOUT0 => N110702616, 
	DOUT1 => N110702617, 
	DOUT2 => N110702618, 
	DOUT3 => N110702619, 
	DOUT4 => N110702620, 
	DOUT5 => N110702621, 
	DOUT6 => N110702622, 
	DOUT7 => N110702623, 
	DOUT8 => N110702624, 
	DOUT9 => N110702625, 
	DOUT10 => N110702626, 
	DOUT11 => N110702627, 
	DOUT12 => N110702628, 
	DOUT13 => N110702629, 
	DOUT14 => N110702630, 
	DOUT15 => N110702631, 
	SIGNEDIN => N110702632, 
	SIGNEDOUT => N110702633
);
U137 : ADDERDELAY	PORT MAP(
	DIN0 => N111497716, 
	DIN1 => N111497717, 
	DIN2 => N111497718, 
	DIN3 => N111497719, 
	DIN4 => N111497720, 
	DIN5 => N111497721, 
	DIN6 => N111497722, 
	DIN7 => N111497723, 
	DIN8 => N111497724, 
	DIN9 => N111497725, 
	DIN10 => N111497726, 
	DIN11 => N111497727, 
	DIN12 => N111497728, 
	DIN13 => N111497729, 
	DIN14 => N111497730, 
	DIN15 => N111497731, 
	DOUT0 => N111522016, 
	DOUT1 => N111522017, 
	DOUT2 => N111522018, 
	DOUT3 => N111522019, 
	DOUT4 => N111522020, 
	DOUT5 => N111522021, 
	DOUT6 => N111522022, 
	DOUT7 => N111522023, 
	DOUT8 => N111522024, 
	DOUT9 => N111522025, 
	DOUT10 => N111522026, 
	DOUT11 => N111522027, 
	DOUT12 => N111522028, 
	DOUT13 => N111522029, 
	DOUT14 => N111522030, 
	DOUT15 => N111522031, 
	SIGNEDIN => N111497733, 
	SIGNEDOUT => N111522033
);
U106 : ADDERDELAY	PORT MAP(
	DIN0 => N110702616, 
	DIN1 => N110702617, 
	DIN2 => N110702618, 
	DIN3 => N110702619, 
	DIN4 => N110702620, 
	DIN5 => N110702621, 
	DIN6 => N110702622, 
	DIN7 => N110702623, 
	DIN8 => N110702624, 
	DIN9 => N110702625, 
	DIN10 => N110702626, 
	DIN11 => N110702627, 
	DIN12 => N110702628, 
	DIN13 => N110702629, 
	DIN14 => N110702630, 
	DIN15 => N110702631, 
	DOUT0 => N110730716, 
	DOUT1 => N110730717, 
	DOUT2 => N110730718, 
	DOUT3 => N110730719, 
	DOUT4 => N110730720, 
	DOUT5 => N110730721, 
	DOUT6 => N110730722, 
	DOUT7 => N110730723, 
	DOUT8 => N110730724, 
	DOUT9 => N110730725, 
	DOUT10 => N110730726, 
	DOUT11 => N110730727, 
	DOUT12 => N110730728, 
	DOUT13 => N110730729, 
	DOUT14 => N110730730, 
	DOUT15 => N110730731, 
	SIGNEDIN => N110702633, 
	SIGNEDOUT => N110730733
);
U138 : ADDERDELAY	PORT MAP(
	DIN0 => N111522016, 
	DIN1 => N111522017, 
	DIN2 => N111522018, 
	DIN3 => N111522019, 
	DIN4 => N111522020, 
	DIN5 => N111522021, 
	DIN6 => N111522022, 
	DIN7 => N111522023, 
	DIN8 => N111522024, 
	DIN9 => N111522025, 
	DIN10 => N111522026, 
	DIN11 => N111522027, 
	DIN12 => N111522028, 
	DIN13 => N111522029, 
	DIN14 => N111522030, 
	DIN15 => N111522031, 
	DOUT0 => N111546316, 
	DOUT1 => N111546317, 
	DOUT2 => N111546318, 
	DOUT3 => N111546319, 
	DOUT4 => N111546320, 
	DOUT5 => N111546321, 
	DOUT6 => N111546322, 
	DOUT7 => N111546323, 
	DOUT8 => N111546324, 
	DOUT9 => N111546325, 
	DOUT10 => N111546326, 
	DOUT11 => N111546327, 
	DOUT12 => N111546328, 
	DOUT13 => N111546329, 
	DOUT14 => N111546330, 
	DOUT15 => N111546331, 
	SIGNEDIN => N111522033, 
	SIGNEDOUT => N111546333
);
U107 : ADDERDELAY	PORT MAP(
	DIN0 => N110730716, 
	DIN1 => N110730717, 
	DIN2 => N110730718, 
	DIN3 => N110730719, 
	DIN4 => N110730720, 
	DIN5 => N110730721, 
	DIN6 => N110730722, 
	DIN7 => N110730723, 
	DIN8 => N110730724, 
	DIN9 => N110730725, 
	DIN10 => N110730726, 
	DIN11 => N110730727, 
	DIN12 => N110730728, 
	DIN13 => N110730729, 
	DIN14 => N110730730, 
	DIN15 => N110730731, 
	DOUT0 => N110755016, 
	DOUT1 => N110755017, 
	DOUT2 => N110755018, 
	DOUT3 => N110755019, 
	DOUT4 => N110755020, 
	DOUT5 => N110755021, 
	DOUT6 => N110755022, 
	DOUT7 => N110755023, 
	DOUT8 => N110755024, 
	DOUT9 => N110755025, 
	DOUT10 => N110755026, 
	DOUT11 => N110755027, 
	DOUT12 => N110755028, 
	DOUT13 => N110755029, 
	DOUT14 => N110755030, 
	DOUT15 => N110755031, 
	SIGNEDIN => N110730733, 
	SIGNEDOUT => N110755033
);
U139 : ADDERDELAY	PORT MAP(
	DIN0 => N110831716, 
	DIN1 => N110831717, 
	DIN2 => N110831718, 
	DIN3 => N110831719, 
	DIN4 => N110831720, 
	DIN5 => N110831721, 
	DIN6 => N110831722, 
	DIN7 => N110831723, 
	DIN8 => N110831724, 
	DIN9 => N110831725, 
	DIN10 => N110831726, 
	DIN11 => N110831727, 
	DIN12 => N110831728, 
	DIN13 => N110831729, 
	DIN14 => N110831730, 
	DIN15 => N110831731, 
	DOUT0 => N111570616, 
	DOUT1 => N111570617, 
	DOUT2 => N111570618, 
	DOUT3 => N111570619, 
	DOUT4 => N111570620, 
	DOUT5 => N111570621, 
	DOUT6 => N111570622, 
	DOUT7 => N111570623, 
	DOUT8 => N111570624, 
	DOUT9 => N111570625, 
	DOUT10 => N111570626, 
	DOUT11 => N111570627, 
	DOUT12 => N111570628, 
	DOUT13 => N111570629, 
	DOUT14 => N111570630, 
	DOUT15 => N111570631, 
	SIGNEDIN => N110831733, 
	SIGNEDOUT => N111570633
);
U108 : ADDERDELAY	PORT MAP(
	DIN0 => N11077930, 
	DIN1 => N11077931, 
	DIN2 => N11077932, 
	DIN3 => N11077933, 
	DIN4 => N11077934, 
	DIN5 => N11077935, 
	DIN6 => N11077936, 
	DIN7 => N11077937, 
	DIN8 => N11077938, 
	DIN9 => N11077939, 
	DIN10 => N110779310, 
	DIN11 => N110779311, 
	DIN12 => N110779312, 
	DIN13 => N110779313, 
	DIN14 => N110779314, 
	DIN15 => N110779315, 
	DOUT0 => N110779316, 
	DOUT1 => N110779317, 
	DOUT2 => N110779318, 
	DOUT3 => N110779319, 
	DOUT4 => N110779320, 
	DOUT5 => N110779321, 
	DOUT6 => N110779322, 
	DOUT7 => N110779323, 
	DOUT8 => N110779324, 
	DOUT9 => N110779325, 
	DOUT10 => N110779326, 
	DOUT11 => N110779327, 
	DOUT12 => N110779328, 
	DOUT13 => N110779329, 
	DOUT14 => N110779330, 
	DOUT15 => N110779331, 
	SIGNEDIN => N110779332, 
	SIGNEDOUT => N110779333
);
U109 : ADDERDELAY	PORT MAP(
	DIN0 => N110779316, 
	DIN1 => N110779317, 
	DIN2 => N110779318, 
	DIN3 => N110779319, 
	DIN4 => N110779320, 
	DIN5 => N110779321, 
	DIN6 => N110779322, 
	DIN7 => N110779323, 
	DIN8 => N110779324, 
	DIN9 => N110779325, 
	DIN10 => N110779326, 
	DIN11 => N110779327, 
	DIN12 => N110779328, 
	DIN13 => N110779329, 
	DIN14 => N110779330, 
	DIN15 => N110779331, 
	DOUT0 => N110807416, 
	DOUT1 => N110807417, 
	DOUT2 => N110807418, 
	DOUT3 => N110807419, 
	DOUT4 => N110807420, 
	DOUT5 => N110807421, 
	DOUT6 => N110807422, 
	DOUT7 => N110807423, 
	DOUT8 => N110807424, 
	DOUT9 => N110807425, 
	DOUT10 => N110807426, 
	DOUT11 => N110807427, 
	DOUT12 => N110807428, 
	DOUT13 => N110807429, 
	DOUT14 => N110807430, 
	DOUT15 => N110807431, 
	SIGNEDIN => N110779333, 
	SIGNEDOUT => N110807433
);
U90 : ADDERDELAY	PORT MAP(
	DIN0 => N11031910, 
	DIN1 => N11031911, 
	DIN2 => N11031912, 
	DIN3 => N11031913, 
	DIN4 => N11031914, 
	DIN5 => N11031915, 
	DIN6 => N11031916, 
	DIN7 => N11031917, 
	DIN8 => N11031918, 
	DIN9 => N11031919, 
	DIN10 => N110319110, 
	DIN11 => N110319111, 
	DIN12 => N110319112, 
	DIN13 => N110319113, 
	DIN14 => N110319114, 
	DIN15 => N110319115, 
	DOUT0 => N110319116, 
	DOUT1 => N110319117, 
	DOUT2 => N110319118, 
	DOUT3 => N110319119, 
	DOUT4 => N110319120, 
	DOUT5 => N110319121, 
	DOUT6 => N110319122, 
	DOUT7 => N110319123, 
	DOUT8 => N110319124, 
	DOUT9 => N110319125, 
	DOUT10 => N110319126, 
	DOUT11 => N110319127, 
	DOUT12 => N110319128, 
	DOUT13 => N110319129, 
	DOUT14 => N110319130, 
	DOUT15 => N110319131, 
	SIGNEDIN => N110319132, 
	SIGNEDOUT => N110319133
);
U91 : ADDERDELAY	PORT MAP(
	DIN0 => N110319116, 
	DIN1 => N110319117, 
	DIN2 => N110319118, 
	DIN3 => N110319119, 
	DIN4 => N110319120, 
	DIN5 => N110319121, 
	DIN6 => N110319122, 
	DIN7 => N110319123, 
	DIN8 => N110319124, 
	DIN9 => N110319125, 
	DIN10 => N110319126, 
	DIN11 => N110319127, 
	DIN12 => N110319128, 
	DIN13 => N110319129, 
	DIN14 => N110319130, 
	DIN15 => N110319131, 
	DOUT0 => N110347216, 
	DOUT1 => N110347217, 
	DOUT2 => N110347218, 
	DOUT3 => N110347219, 
	DOUT4 => N110347220, 
	DOUT5 => N110347221, 
	DOUT6 => N110347222, 
	DOUT7 => N110347223, 
	DOUT8 => N110347224, 
	DOUT9 => N110347225, 
	DOUT10 => N110347226, 
	DOUT11 => N110347227, 
	DOUT12 => N110347228, 
	DOUT13 => N110347229, 
	DOUT14 => N110347230, 
	DOUT15 => N110347231, 
	SIGNEDIN => N110319133, 
	SIGNEDOUT => N110347233
);
U92 : ADDERDELAY	PORT MAP(
	DIN0 => N110347216, 
	DIN1 => N110347217, 
	DIN2 => N110347218, 
	DIN3 => N110347219, 
	DIN4 => N110347220, 
	DIN5 => N110347221, 
	DIN6 => N110347222, 
	DIN7 => N110347223, 
	DIN8 => N110347224, 
	DIN9 => N110347225, 
	DIN10 => N110347226, 
	DIN11 => N110347227, 
	DIN12 => N110347228, 
	DIN13 => N110347229, 
	DIN14 => N110347230, 
	DIN15 => N110347231, 
	DOUT0 => N1145131, 
	DOUT1 => N1145091, 
	DOUT2 => N1145127, 
	DOUT3 => N1145099, 
	DOUT4 => N1145083, 
	DOUT5 => N1145111, 
	DOUT6 => N1145139, 
	DOUT7 => N1145135, 
	DOUT8 => N1145119, 
	DOUT9 => N1145107, 
	DOUT10 => N1145123, 
	DOUT11 => N1145115, 
	DOUT12 => N1145095, 
	DOUT13 => N1145103, 
	DOUT14 => N1145075, 
	DOUT15 => N1145079, 
	SIGNEDIN => N110347233, 
	SIGNEDOUT => N1145087
);
U93 : ADDERDELAY	PORT MAP(
	DIN0 => N11039580, 
	DIN1 => N11039581, 
	DIN2 => N11039582, 
	DIN3 => N11039583, 
	DIN4 => N11039584, 
	DIN5 => N11039585, 
	DIN6 => N11039586, 
	DIN7 => N11039587, 
	DIN8 => N11039588, 
	DIN9 => N11039589, 
	DIN10 => N110395810, 
	DIN11 => N110395811, 
	DIN12 => N110395812, 
	DIN13 => N110395813, 
	DIN14 => N110395814, 
	DIN15 => N110395815, 
	DOUT0 => N110395816, 
	DOUT1 => N110395817, 
	DOUT2 => N110395818, 
	DOUT3 => N110395819, 
	DOUT4 => N110395820, 
	DOUT5 => N110395821, 
	DOUT6 => N110395822, 
	DOUT7 => N110395823, 
	DOUT8 => N110395824, 
	DOUT9 => N110395825, 
	DOUT10 => N110395826, 
	DOUT11 => N110395827, 
	DOUT12 => N110395828, 
	DOUT13 => N110395829, 
	DOUT14 => N110395830, 
	DOUT15 => N110395831, 
	SIGNEDIN => N110395832, 
	SIGNEDOUT => N110395833
);
U94 : ADDERDELAY	PORT MAP(
	DIN0 => N110395816, 
	DIN1 => N110395817, 
	DIN2 => N110395818, 
	DIN3 => N110395819, 
	DIN4 => N110395820, 
	DIN5 => N110395821, 
	DIN6 => N110395822, 
	DIN7 => N110395823, 
	DIN8 => N110395824, 
	DIN9 => N110395825, 
	DIN10 => N110395826, 
	DIN11 => N110395827, 
	DIN12 => N110395828, 
	DIN13 => N110395829, 
	DIN14 => N110395830, 
	DIN15 => N110395831, 
	DOUT0 => N110423916, 
	DOUT1 => N110423917, 
	DOUT2 => N110423918, 
	DOUT3 => N110423919, 
	DOUT4 => N110423920, 
	DOUT5 => N110423921, 
	DOUT6 => N110423922, 
	DOUT7 => N110423923, 
	DOUT8 => N110423924, 
	DOUT9 => N110423925, 
	DOUT10 => N110423926, 
	DOUT11 => N110423927, 
	DOUT12 => N110423928, 
	DOUT13 => N110423929, 
	DOUT14 => N110423930, 
	DOUT15 => N110423931, 
	SIGNEDIN => N110395833, 
	SIGNEDOUT => N110423933
);
U95 : ADDERDELAY	PORT MAP(
	DIN0 => N110423916, 
	DIN1 => N110423917, 
	DIN2 => N110423918, 
	DIN3 => N110423919, 
	DIN4 => N110423920, 
	DIN5 => N110423921, 
	DIN6 => N110423922, 
	DIN7 => N110423923, 
	DIN8 => N110423924, 
	DIN9 => N110423925, 
	DIN10 => N110423926, 
	DIN11 => N110423927, 
	DIN12 => N110423928, 
	DIN13 => N110423929, 
	DIN14 => N110423930, 
	DIN15 => N110423931, 
	DOUT0 => N110448216, 
	DOUT1 => N110448217, 
	DOUT2 => N110448218, 
	DOUT3 => N110448219, 
	DOUT4 => N110448220, 
	DOUT5 => N110448221, 
	DOUT6 => N110448222, 
	DOUT7 => N110448223, 
	DOUT8 => N110448224, 
	DOUT9 => N110448225, 
	DOUT10 => N110448226, 
	DOUT11 => N110448227, 
	DOUT12 => N110448228, 
	DOUT13 => N110448229, 
	DOUT14 => N110448230, 
	DOUT15 => N110448231, 
	SIGNEDIN => N110423933, 
	SIGNEDOUT => N110448233
);
U31 : COUNTER	PORT MAP(
	CLK => LOAD, 
	NCLR => NRST, 
	NPRE => VCC, 
	NQ0 => N94143, 
	NQ1 => N94145, 
	NQ2 => N94147, 
	NQ3 => N94149, 
	Q0 => N94151, 
	Q1 => N94153, 
	Q2 => N94155, 
	Q3 => N94157
);
U96 : ADDERDELAY	PORT MAP(
	DIN0 => N11047250, 
	DIN1 => N11047251, 
	DIN2 => N11047252, 
	DIN3 => N11047253, 
	DIN4 => N11047254, 
	DIN5 => N11047255, 
	DIN6 => N11047256, 
	DIN7 => N11047257, 
	DIN8 => N11047258, 
	DIN9 => N11047259, 
	DIN10 => N110472510, 
	DIN11 => N110472511, 
	DIN12 => N110472512, 
	DIN13 => N110472513, 
	DIN14 => N110472514, 
	DIN15 => N110472515, 
	DOUT0 => N110472516, 
	DOUT1 => N110472517, 
	DOUT2 => N110472518, 
	DOUT3 => N110472519, 
	DOUT4 => N110472520, 
	DOUT5 => N110472521, 
	DOUT6 => N110472522, 
	DOUT7 => N110472523, 
	DOUT8 => N110472524, 
	DOUT9 => N110472525, 
	DOUT10 => N110472526, 
	DOUT11 => N110472527, 
	DOUT12 => N110472528, 
	DOUT13 => N110472529, 
	DOUT14 => N110472530, 
	DOUT15 => N110472531, 
	SIGNEDIN => N110472532, 
	SIGNEDOUT => N110472533
);
U32 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => DCO0, 
	DCO1 => DCO1, 
	DCO2 => DCO2, 
	DCO3 => DCO3, 
	DCO4 => DCO4, 
	DCO5 => DCO5, 
	DCO6 => DCO6, 
	DCO7 => DCO7, 
	DSG0 => DSG0, 
	DSG1 => DSG1, 
	DSG2 => DSG2, 
	DSG3 => DSG3, 
	DSG4 => DSG4, 
	DSG5 => DSG5, 
	DSG6 => DSG6, 
	DSG7 => DSG7, 
	ENABLE => ENABLE1, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => COONETEST0, 
	QCO1 => COONETEST1, 
	QCO2 => COONETEST2, 
	QCO3 => COONETEST3, 
	QCO4 => COONETEST4, 
	QCO5 => COONETEST5, 
	QCO6 => COONETEST6, 
	QCO7 => COONETEST7, 
	QSG0 => N06027, 
	QSG1 => N06029, 
	QSG2 => N06031, 
	QSG3 => N06033, 
	QSG4 => N06035, 
	QSG5 => N06037, 
	QSG6 => N06039, 
	QSG7 => N06041, 
	S0 => N1078467, 
	S1 => N1078469, 
	S2 => N1078471, 
	S3 => N1078473, 
	S4 => N1078475, 
	S5 => N1078477, 
	S6 => N1078479, 
	S7 => N1078481, 
	S8 => N1078483, 
	S9 => N1078485, 
	S10 => N1078487, 
	S11 => N1078489, 
	S12 => N1078491, 
	S13 => N1078493, 
	S14 => N1078495, 
	S15 => N1078497, 
	SIGNED => N1078499
);
U1761607403 : ORBLOCK	PORT MAP(
	A0 => A0, 
	A1 => A1, 
	A2 => A2, 
	A3 => A3, 
	A4 => A4, 
	A5 => A5, 
	A6 => A6, 
	A7 => A7, 
	A8 => A8, 
	A9 => A9, 
	A10 => A10, 
	A11 => A11, 
	A12 => A12, 
	A13 => A13, 
	A14 => A14, 
	A15 => A15, 
	B0 => B0, 
	B1 => B1, 
	B2 => B2, 
	B3 => B3, 
	B4 => B4, 
	B5 => B5, 
	B6 => B6, 
	B7 => B7, 
	B8 => B8, 
	B9 => B9, 
	B10 => B10, 
	B11 => B11, 
	B12 => B12, 
	B13 => B13, 
	B14 => B14, 
	B15 => B15, 
	C0 => C0, 
	C1 => C1, 
	C2 => C2, 
	C3 => C3, 
	C4 => C4, 
	C5 => C5, 
	C6 => C6, 
	C7 => C7, 
	C8 => C8, 
	C9 => C9, 
	C10 => C10, 
	C11 => C11, 
	C12 => C12, 
	C13 => C13, 
	C14 => C14, 
	C15 => C15, 
	D0 => D0, 
	D1 => D1, 
	D2 => D2, 
	D3 => D3, 
	D4 => D4, 
	D5 => D5, 
	D6 => D6, 
	D7 => D7, 
	D8 => D8, 
	D9 => D9, 
	D10 => D10, 
	D11 => D11, 
	D12 => D12, 
	D13 => D13, 
	D14 => D14, 
	D15 => D15, 
	E0 => E0, 
	E1 => E1, 
	E2 => E2, 
	E3 => E3, 
	E4 => E4, 
	E5 => E5, 
	E6 => E6, 
	E7 => E7, 
	E8 => E8, 
	E9 => E9, 
	E10 => E10, 
	E11 => E11, 
	E12 => E12, 
	E13 => E13, 
	E14 => E14, 
	E15 => E15, 
	F0 => F0, 
	F1 => F1, 
	F2 => F2, 
	F3 => F3, 
	F4 => F4, 
	F5 => F5, 
	F6 => F6, 
	F7 => F7, 
	F8 => F8, 
	F9 => F9, 
	F10 => F10, 
	F11 => F11, 
	F12 => F12, 
	F13 => F13, 
	F14 => F14, 
	F15 => F15, 
	G0 => G0, 
	G1 => G1, 
	G2 => G2, 
	G3 => G3, 
	G4 => G4, 
	G5 => G5, 
	G6 => G6, 
	G7 => G7, 
	G8 => G8, 
	G9 => G9, 
	G10 => G10, 
	G11 => G11, 
	G12 => G12, 
	G13 => G13, 
	G14 => G14, 
	G15 => G15, 
	H0 => H0, 
	H1 => H1, 
	H2 => H2, 
	H3 => H3, 
	H4 => H4, 
	H5 => H5, 
	H6 => H6, 
	H7 => H7, 
	H8 => H8, 
	H9 => H9, 
	H10 => H10, 
	H11 => H11, 
	H12 => H12, 
	H13 => H13, 
	H14 => H14, 
	H15 => H15, 
	OUTPUT0 => CHECK0, 
	OUTPUT1 => CHECK1, 
	OUTPUT2 => CHECK2, 
	OUTPUT3 => CHECK3, 
	OUTPUT4 => CHECK4, 
	OUTPUT5 => CHECK5, 
	OUTPUT6 => CHECK6, 
	OUTPUT7 => CHECK7, 
	OUTPUT8 => CHECK8, 
	OUTPUT9 => CHECK9, 
	OUTPUT10 => CHECK10, 
	OUTPUT11 => CHECK11, 
	OUTPUT12 => CHECK12, 
	OUTPUT13 => CHECK13, 
	OUTPUT14 => CHECK14, 
	OUTPUT15 => CHECK15
);
U33 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => COONETEST0, 
	DCO1 => COONETEST1, 
	DCO2 => COONETEST2, 
	DCO3 => COONETEST3, 
	DCO4 => COONETEST4, 
	DCO5 => COONETEST5, 
	DCO6 => COONETEST6, 
	DCO7 => COONETEST7, 
	DSG0 => N06027, 
	DSG1 => N06029, 
	DSG2 => N06031, 
	DSG3 => N06033, 
	DSG4 => N06035, 
	DSG5 => N06037, 
	DSG6 => N06039, 
	DSG7 => N06041, 
	ENABLE => ENABLE2, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => COTEST0, 
	QCO1 => COTEST1, 
	QCO2 => COTEST2, 
	QCO3 => COTEST3, 
	QCO4 => COTEST4, 
	QCO5 => COTEST5, 
	QCO6 => COTEST6, 
	QCO7 => COTEST7, 
	QSG0 => N93230, 
	QSG1 => N93232, 
	QSG2 => N93234, 
	QSG3 => N93236, 
	QSG4 => N93238, 
	QSG5 => N93240, 
	QSG6 => N93242, 
	QSG7 => N93244, 
	S0 => N10716200, 
	S1 => N10716201, 
	S2 => N10716202, 
	S3 => N10716203, 
	S4 => N10716204, 
	S5 => N10716205, 
	S6 => N10716206, 
	S7 => N10716207, 
	S8 => N10716208, 
	S9 => N10716209, 
	S10 => N107162010, 
	S11 => N107162011, 
	S12 => N107162012, 
	S13 => N107162013, 
	S14 => N107162014, 
	S15 => N107162015, 
	SIGNED => N107162032
);
U97 : ADDERDELAY	PORT MAP(
	DIN0 => N110472516, 
	DIN1 => N110472517, 
	DIN2 => N110472518, 
	DIN3 => N110472519, 
	DIN4 => N110472520, 
	DIN5 => N110472521, 
	DIN6 => N110472522, 
	DIN7 => N110472523, 
	DIN8 => N110472524, 
	DIN9 => N110472525, 
	DIN10 => N110472526, 
	DIN11 => N110472527, 
	DIN12 => N110472528, 
	DIN13 => N110472529, 
	DIN14 => N110472530, 
	DIN15 => N110472531, 
	DOUT0 => N110500616, 
	DOUT1 => N110500617, 
	DOUT2 => N110500618, 
	DOUT3 => N110500619, 
	DOUT4 => N110500620, 
	DOUT5 => N110500621, 
	DOUT6 => N110500622, 
	DOUT7 => N110500623, 
	DOUT8 => N110500624, 
	DOUT9 => N110500625, 
	DOUT10 => N110500626, 
	DOUT11 => N110500627, 
	DOUT12 => N110500628, 
	DOUT13 => N110500629, 
	DOUT14 => N110500630, 
	DOUT15 => N110500631, 
	SIGNEDIN => N110472533, 
	SIGNEDOUT => N110500633
);
U34 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => COTEST0, 
	DCO1 => COTEST1, 
	DCO2 => COTEST2, 
	DCO3 => COTEST3, 
	DCO4 => COTEST4, 
	DCO5 => COTEST5, 
	DCO6 => COTEST6, 
	DCO7 => COTEST7, 
	DSG0 => N93230, 
	DSG1 => N93232, 
	DSG2 => N93234, 
	DSG3 => N93236, 
	DSG4 => N93238, 
	DSG5 => N93240, 
	DSG6 => N93242, 
	DSG7 => N93244, 
	ENABLE => ENABLE3, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => TEST0, 
	QCO1 => TEST1, 
	QCO2 => TEST2, 
	QCO3 => TEST3, 
	QCO4 => TEST4, 
	QCO5 => TEST5, 
	QCO6 => TEST6, 
	QCO7 => TEST7, 
	QSG0 => SGTEST0, 
	QSG1 => SGTEST1, 
	QSG2 => SGTEST2, 
	QSG3 => SGTEST3, 
	QSG4 => SGTEST4, 
	QSG5 => SGTEST5, 
	QSG6 => SGTEST6, 
	QSG7 => SGTEST7, 
	S0 => N11026670, 
	S1 => N11026671, 
	S2 => N11026672, 
	S3 => N11026673, 
	S4 => N11026674, 
	S5 => N11026675, 
	S6 => N11026676, 
	S7 => N11026677, 
	S8 => N11026678, 
	S9 => N11026679, 
	S10 => N110266710, 
	S11 => N110266711, 
	S12 => N110266712, 
	S13 => N110266713, 
	S14 => N110266714, 
	S15 => N110266715, 
	SIGNED => N110266732
);
U98 : ADDERDELAY	PORT MAP(
	DIN0 => N110500616, 
	DIN1 => N110500617, 
	DIN2 => N110500618, 
	DIN3 => N110500619, 
	DIN4 => N110500620, 
	DIN5 => N110500621, 
	DIN6 => N110500622, 
	DIN7 => N110500623, 
	DIN8 => N110500624, 
	DIN9 => N110500625, 
	DIN10 => N110500626, 
	DIN11 => N110500627, 
	DIN12 => N110500628, 
	DIN13 => N110500629, 
	DIN14 => N110500630, 
	DIN15 => N110500631, 
	DOUT0 => N110524916, 
	DOUT1 => N110524917, 
	DOUT2 => N110524918, 
	DOUT3 => N110524919, 
	DOUT4 => N110524920, 
	DOUT5 => N110524921, 
	DOUT6 => N110524922, 
	DOUT7 => N110524923, 
	DOUT8 => N110524924, 
	DOUT9 => N110524925, 
	DOUT10 => N110524926, 
	DOUT11 => N110524927, 
	DOUT12 => N110524928, 
	DOUT13 => N110524929, 
	DOUT14 => N110524930, 
	DOUT15 => N110524931, 
	SIGNEDIN => N110500633, 
	SIGNEDOUT => N110524933
);
U35 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => TEST0, 
	DCO1 => TEST1, 
	DCO2 => TEST2, 
	DCO3 => TEST3, 
	DCO4 => TEST4, 
	DCO5 => TEST5, 
	DCO6 => TEST6, 
	DCO7 => TEST7, 
	DSG0 => SGTEST0, 
	DSG1 => SGTEST1, 
	DSG2 => SGTEST2, 
	DSG3 => SGTEST3, 
	DSG4 => SGTEST4, 
	DSG5 => SGTEST5, 
	DSG6 => SGTEST6, 
	DSG7 => SGTEST7, 
	ENABLE => ENABLE4, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => N91222, 
	QCO1 => N91224, 
	QCO2 => N91226, 
	QCO3 => N91228, 
	QCO4 => N91230, 
	QCO5 => N91232, 
	QCO6 => N91234, 
	QCO7 => N91236, 
	QSG0 => N91238, 
	QSG1 => N91240, 
	QSG2 => N91242, 
	QSG3 => N91244, 
	QSG4 => N91246, 
	QSG5 => N91248, 
	QSG6 => N91250, 
	QSG7 => N91252, 
	S0 => N11031910, 
	S1 => N11031911, 
	S2 => N11031912, 
	S3 => N11031913, 
	S4 => N11031914, 
	S5 => N11031915, 
	S6 => N11031916, 
	S7 => N11031917, 
	S8 => N11031918, 
	S9 => N11031919, 
	S10 => N110319110, 
	S11 => N110319111, 
	S12 => N110319112, 
	S13 => N110319113, 
	S14 => N110319114, 
	S15 => N110319115, 
	SIGNED => N110319132
);
U99 : ADDERDELAY	PORT MAP(
	DIN0 => N11054920, 
	DIN1 => N11054921, 
	DIN2 => N11054922, 
	DIN3 => N11054923, 
	DIN4 => N11054924, 
	DIN5 => N11054925, 
	DIN6 => N11054926, 
	DIN7 => N11054927, 
	DIN8 => N11054928, 
	DIN9 => N11054929, 
	DIN10 => N110549210, 
	DIN11 => N110549211, 
	DIN12 => N110549212, 
	DIN13 => N110549213, 
	DIN14 => N110549214, 
	DIN15 => N110549215, 
	DOUT0 => N110549216, 
	DOUT1 => N110549217, 
	DOUT2 => N110549218, 
	DOUT3 => N110549219, 
	DOUT4 => N110549220, 
	DOUT5 => N110549221, 
	DOUT6 => N110549222, 
	DOUT7 => N110549223, 
	DOUT8 => N110549224, 
	DOUT9 => N110549225, 
	DOUT10 => N110549226, 
	DOUT11 => N110549227, 
	DOUT12 => N110549228, 
	DOUT13 => N110549229, 
	DOUT14 => N110549230, 
	DOUT15 => N110549231, 
	SIGNEDIN => N110549232, 
	SIGNEDOUT => N110549233
);
U36 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => N91222, 
	DCO1 => N91224, 
	DCO2 => N91226, 
	DCO3 => N91228, 
	DCO4 => N91230, 
	DCO5 => N91232, 
	DCO6 => N91234, 
	DCO7 => N91236, 
	DSG0 => N91238, 
	DSG1 => N91240, 
	DSG2 => N91242, 
	DSG3 => N91244, 
	DSG4 => N91246, 
	DSG5 => N91248, 
	DSG6 => N91250, 
	DSG7 => N91252, 
	ENABLE => ENABLE5, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => N84206, 
	QCO1 => N84208, 
	QCO2 => N84210, 
	QCO3 => N84212, 
	QCO4 => N84214, 
	QCO5 => N84216, 
	QCO6 => N84218, 
	QCO7 => N84220, 
	QSG0 => N84222, 
	QSG1 => N84224, 
	QSG2 => N84226, 
	QSG3 => N84228, 
	QSG4 => N84230, 
	QSG5 => N84232, 
	QSG6 => N84234, 
	QSG7 => N84236, 
	S0 => N11039580, 
	S1 => N11039581, 
	S2 => N11039582, 
	S3 => N11039583, 
	S4 => N11039584, 
	S5 => N11039585, 
	S6 => N11039586, 
	S7 => N11039587, 
	S8 => N11039588, 
	S9 => N11039589, 
	S10 => N110395810, 
	S11 => N110395811, 
	S12 => N110395812, 
	S13 => N110395813, 
	S14 => N110395814, 
	S15 => N110395815, 
	SIGNED => N110395832
);
U69 : \7404\	PORT MAP(
	A_A => N955836, 
	Y_A => N955599, 
	GND => GND, 
	VCC => VCC, 
	A_B => 'Z', 
	Y_B => OPEN, 
	A_C => 'Z', 
	Y_C => OPEN, 
	A_D => 'Z', 
	Y_D => OPEN, 
	A_E => 'Z', 
	Y_E => OPEN, 
	A_F => 'Z', 
	Y_F => OPEN
);
U37 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => N84206, 
	DCO1 => N84208, 
	DCO2 => N84210, 
	DCO3 => N84212, 
	DCO4 => N84214, 
	DCO5 => N84216, 
	DCO6 => N84218, 
	DCO7 => N84220, 
	DSG0 => N84222, 
	DSG1 => N84224, 
	DSG2 => N84226, 
	DSG3 => N84228, 
	DSG4 => N84230, 
	DSG5 => N84232, 
	DSG6 => N84234, 
	DSG7 => N84236, 
	ENABLE => ENABLE6, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => N83393, 
	QCO1 => N83395, 
	QCO2 => N83397, 
	QCO3 => N83399, 
	QCO4 => N83401, 
	QCO5 => N83403, 
	QCO6 => N83405, 
	QCO7 => N83407, 
	QSG0 => N83409, 
	QSG1 => N83411, 
	QSG2 => N83413, 
	QSG3 => N83415, 
	QSG4 => N83417, 
	QSG5 => N83419, 
	QSG6 => N83421, 
	QSG7 => N83423, 
	S0 => N11047250, 
	S1 => N11047251, 
	S2 => N11047252, 
	S3 => N11047253, 
	S4 => N11047254, 
	S5 => N11047255, 
	S6 => N11047256, 
	S7 => N11047257, 
	S8 => N11047258, 
	S9 => N11047259, 
	S10 => N110472510, 
	S11 => N110472511, 
	S12 => N110472512, 
	S13 => N110472513, 
	S14 => N110472514, 
	S15 => N110472515, 
	SIGNED => N110472532
);
U38 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => N83393, 
	DCO1 => N83395, 
	DCO2 => N83397, 
	DCO3 => N83399, 
	DCO4 => N83401, 
	DCO5 => N83403, 
	DCO6 => N83405, 
	DCO7 => N83407, 
	DSG0 => N83409, 
	DSG1 => N83411, 
	DSG2 => N83413, 
	DSG3 => N83415, 
	DSG4 => N83417, 
	DSG5 => N83419, 
	DSG6 => N83421, 
	DSG7 => N83423, 
	ENABLE => ENABLE7, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => N82578, 
	QCO1 => N82580, 
	QCO2 => N82582, 
	QCO3 => N82584, 
	QCO4 => N82586, 
	QCO5 => N82588, 
	QCO6 => N82590, 
	QCO7 => N82592, 
	QSG0 => N82594, 
	QSG1 => N82596, 
	QSG2 => N82598, 
	QSG3 => N82600, 
	QSG4 => N82602, 
	QSG5 => N82604, 
	QSG6 => N82606, 
	QSG7 => N82608, 
	S0 => N11054920, 
	S1 => N11054921, 
	S2 => N11054922, 
	S3 => N11054923, 
	S4 => N11054924, 
	S5 => N11054925, 
	S6 => N11054926, 
	S7 => N11054927, 
	S8 => N11054928, 
	S9 => N11054929, 
	S10 => N110549210, 
	S11 => N110549211, 
	S12 => N110549212, 
	S13 => N110549213, 
	S14 => N110549214, 
	S15 => N110549215, 
	SIGNED => N110549232
);
U39 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => N82578, 
	DCO1 => N82580, 
	DCO2 => N82582, 
	DCO3 => N82584, 
	DCO4 => N82586, 
	DCO5 => N82588, 
	DCO6 => N82590, 
	DCO7 => N82592, 
	DSG0 => N82594, 
	DSG1 => N82596, 
	DSG2 => N82598, 
	DSG3 => N82600, 
	DSG4 => N82602, 
	DSG5 => N82604, 
	DSG6 => N82606, 
	DSG7 => N82608, 
	ENABLE => N94157, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => N81765, 
	QCO1 => N81767, 
	QCO2 => N81769, 
	QCO3 => N81771, 
	QCO4 => N81773, 
	QCO5 => N81775, 
	QCO6 => N81777, 
	QCO7 => N81779, 
	QSG0 => N81781, 
	QSG1 => N81783, 
	QSG2 => N81785, 
	QSG3 => N81787, 
	QSG4 => N81789, 
	QSG5 => N81791, 
	QSG6 => N81793, 
	QSG7 => N81795, 
	S0 => N11062590, 
	S1 => N11062591, 
	S2 => N11062592, 
	S3 => N11062593, 
	S4 => N11062594, 
	S5 => N11062595, 
	S6 => N11062596, 
	S7 => N11062597, 
	S8 => N11062598, 
	S9 => N11062599, 
	S10 => N110625910, 
	S11 => N110625911, 
	S12 => N110625912, 
	S13 => N110625913, 
	S14 => N110625914, 
	S15 => N110625915, 
	SIGNED => N110625932
);
U170 : ADDERDELAY	PORT MAP(
	DIN0 => N112299616, 
	DIN1 => N112299617, 
	DIN2 => N112299618, 
	DIN3 => N112299619, 
	DIN4 => N112299620, 
	DIN5 => N112299621, 
	DIN6 => N112299622, 
	DIN7 => N112299623, 
	DIN8 => N112299624, 
	DIN9 => N112299625, 
	DIN10 => N112299626, 
	DIN11 => N112299627, 
	DIN12 => N112299628, 
	DIN13 => N112299629, 
	DIN14 => N112299630, 
	DIN15 => N112299631, 
	DOUT0 => N112323916, 
	DOUT1 => N112323917, 
	DOUT2 => N112323918, 
	DOUT3 => N112323919, 
	DOUT4 => N112323920, 
	DOUT5 => N112323921, 
	DOUT6 => N112323922, 
	DOUT7 => N112323923, 
	DOUT8 => N112323924, 
	DOUT9 => N112323925, 
	DOUT10 => N112323926, 
	DOUT11 => N112323927, 
	DOUT12 => N112323928, 
	DOUT13 => N112323929, 
	DOUT14 => N112323930, 
	DOUT15 => N112323931, 
	SIGNEDIN => N112299633, 
	SIGNEDOUT => N112323933
);
U171 : ADDERDELAY	PORT MAP(
	DIN0 => N111837916, 
	DIN1 => N111837917, 
	DIN2 => N111837918, 
	DIN3 => N111837919, 
	DIN4 => N111837920, 
	DIN5 => N111837921, 
	DIN6 => N111837922, 
	DIN7 => N111837923, 
	DIN8 => N111837924, 
	DIN9 => N111837925, 
	DIN10 => N111837926, 
	DIN11 => N111837927, 
	DIN12 => N111837928, 
	DIN13 => N111837929, 
	DIN14 => N111837930, 
	DIN15 => N111837931, 
	DOUT0 => N112348216, 
	DOUT1 => N112348217, 
	DOUT2 => N112348218, 
	DOUT3 => N112348219, 
	DOUT4 => N112348220, 
	DOUT5 => N112348221, 
	DOUT6 => N112348222, 
	DOUT7 => N112348223, 
	DOUT8 => N112348224, 
	DOUT9 => N112348225, 
	DOUT10 => N112348226, 
	DOUT11 => N112348227, 
	DOUT12 => N112348228, 
	DOUT13 => N112348229, 
	DOUT14 => N112348230, 
	DOUT15 => N112348231, 
	SIGNEDIN => N111837933, 
	SIGNEDOUT => N112348233
);
U172 : ADDERDELAY	PORT MAP(
	DIN0 => N112348216, 
	DIN1 => N112348217, 
	DIN2 => N112348218, 
	DIN3 => N112348219, 
	DIN4 => N112348220, 
	DIN5 => N112348221, 
	DIN6 => N112348222, 
	DIN7 => N112348223, 
	DIN8 => N112348224, 
	DIN9 => N112348225, 
	DIN10 => N112348226, 
	DIN11 => N112348227, 
	DIN12 => N112348228, 
	DIN13 => N112348229, 
	DIN14 => N112348230, 
	DIN15 => N112348231, 
	DOUT0 => N112372516, 
	DOUT1 => N112372517, 
	DOUT2 => N112372518, 
	DOUT3 => N112372519, 
	DOUT4 => N112372520, 
	DOUT5 => N112372521, 
	DOUT6 => N112372522, 
	DOUT7 => N112372523, 
	DOUT8 => N112372524, 
	DOUT9 => N112372525, 
	DOUT10 => N112372526, 
	DOUT11 => N112372527, 
	DOUT12 => N112372528, 
	DOUT13 => N112372529, 
	DOUT14 => N112372530, 
	DOUT15 => N112372531, 
	SIGNEDIN => N112348233, 
	SIGNEDOUT => N112372533
);
U140 : ADDERDELAY	PORT MAP(
	DIN0 => N111570616, 
	DIN1 => N111570617, 
	DIN2 => N111570618, 
	DIN3 => N111570619, 
	DIN4 => N111570620, 
	DIN5 => N111570621, 
	DIN6 => N111570622, 
	DIN7 => N111570623, 
	DIN8 => N111570624, 
	DIN9 => N111570625, 
	DIN10 => N111570626, 
	DIN11 => N111570627, 
	DIN12 => N111570628, 
	DIN13 => N111570629, 
	DIN14 => N111570630, 
	DIN15 => N111570631, 
	DOUT0 => N111594916, 
	DOUT1 => N111594917, 
	DOUT2 => N111594918, 
	DOUT3 => N111594919, 
	DOUT4 => N111594920, 
	DOUT5 => N111594921, 
	DOUT6 => N111594922, 
	DOUT7 => N111594923, 
	DOUT8 => N111594924, 
	DOUT9 => N111594925, 
	DOUT10 => N111594926, 
	DOUT11 => N111594927, 
	DOUT12 => N111594928, 
	DOUT13 => N111594929, 
	DOUT14 => N111594930, 
	DOUT15 => N111594931, 
	SIGNEDIN => N111570633, 
	SIGNEDOUT => N111594933
);
U173 : ADDERDELAY	PORT MAP(
	DIN0 => N112372516, 
	DIN1 => N112372517, 
	DIN2 => N112372518, 
	DIN3 => N112372519, 
	DIN4 => N112372520, 
	DIN5 => N112372521, 
	DIN6 => N112372522, 
	DIN7 => N112372523, 
	DIN8 => N112372524, 
	DIN9 => N112372525, 
	DIN10 => N112372526, 
	DIN11 => N112372527, 
	DIN12 => N112372528, 
	DIN13 => N112372529, 
	DIN14 => N112372530, 
	DIN15 => N112372531, 
	DOUT0 => N112396816, 
	DOUT1 => N112396817, 
	DOUT2 => N112396818, 
	DOUT3 => N112396819, 
	DOUT4 => N112396820, 
	DOUT5 => N112396821, 
	DOUT6 => N112396822, 
	DOUT7 => N112396823, 
	DOUT8 => N112396824, 
	DOUT9 => N112396825, 
	DOUT10 => N112396826, 
	DOUT11 => N112396827, 
	DOUT12 => N112396828, 
	DOUT13 => N112396829, 
	DOUT14 => N112396830, 
	DOUT15 => N112396831, 
	SIGNEDIN => N112372533, 
	SIGNEDOUT => N112396833
);
U141 : ADDERDELAY	PORT MAP(
	DIN0 => N111594916, 
	DIN1 => N111594917, 
	DIN2 => N111594918, 
	DIN3 => N111594919, 
	DIN4 => N111594920, 
	DIN5 => N111594921, 
	DIN6 => N111594922, 
	DIN7 => N111594923, 
	DIN8 => N111594924, 
	DIN9 => N111594925, 
	DIN10 => N111594926, 
	DIN11 => N111594927, 
	DIN12 => N111594928, 
	DIN13 => N111594929, 
	DIN14 => N111594930, 
	DIN15 => N111594931, 
	DOUT0 => N111619216, 
	DOUT1 => N111619217, 
	DOUT2 => N111619218, 
	DOUT3 => N111619219, 
	DOUT4 => N111619220, 
	DOUT5 => N111619221, 
	DOUT6 => N111619222, 
	DOUT7 => N111619223, 
	DOUT8 => N111619224, 
	DOUT9 => N111619225, 
	DOUT10 => N111619226, 
	DOUT11 => N111619227, 
	DOUT12 => N111619228, 
	DOUT13 => N111619229, 
	DOUT14 => N111619230, 
	DOUT15 => N111619231, 
	SIGNEDIN => N111594933, 
	SIGNEDOUT => N111619233
);
U110 : ADDERDELAY	PORT MAP(
	DIN0 => N110807416, 
	DIN1 => N110807417, 
	DIN2 => N110807418, 
	DIN3 => N110807419, 
	DIN4 => N110807420, 
	DIN5 => N110807421, 
	DIN6 => N110807422, 
	DIN7 => N110807423, 
	DIN8 => N110807424, 
	DIN9 => N110807425, 
	DIN10 => N110807426, 
	DIN11 => N110807427, 
	DIN12 => N110807428, 
	DIN13 => N110807429, 
	DIN14 => N110807430, 
	DIN15 => N110807431, 
	DOUT0 => N110831716, 
	DOUT1 => N110831717, 
	DOUT2 => N110831718, 
	DOUT3 => N110831719, 
	DOUT4 => N110831720, 
	DOUT5 => N110831721, 
	DOUT6 => N110831722, 
	DOUT7 => N110831723, 
	DOUT8 => N110831724, 
	DOUT9 => N110831725, 
	DOUT10 => N110831726, 
	DOUT11 => N110831727, 
	DOUT12 => N110831728, 
	DOUT13 => N110831729, 
	DOUT14 => N110831730, 
	DOUT15 => N110831731, 
	SIGNEDIN => N110807433, 
	SIGNEDOUT => N110831733
);
U174 : ADDERDELAY	PORT MAP(
	DIN0 => N112396816, 
	DIN1 => N112396817, 
	DIN2 => N112396818, 
	DIN3 => N112396819, 
	DIN4 => N112396820, 
	DIN5 => N112396821, 
	DIN6 => N112396822, 
	DIN7 => N112396823, 
	DIN8 => N112396824, 
	DIN9 => N112396825, 
	DIN10 => N112396826, 
	DIN11 => N112396827, 
	DIN12 => N112396828, 
	DIN13 => N112396829, 
	DIN14 => N112396830, 
	DIN15 => N112396831, 
	DOUT0 => N112421116, 
	DOUT1 => N112421117, 
	DOUT2 => N112421118, 
	DOUT3 => N112421119, 
	DOUT4 => N112421120, 
	DOUT5 => N112421121, 
	DOUT6 => N112421122, 
	DOUT7 => N112421123, 
	DOUT8 => N112421124, 
	DOUT9 => N112421125, 
	DOUT10 => N112421126, 
	DOUT11 => N112421127, 
	DOUT12 => N112421128, 
	DOUT13 => N112421129, 
	DOUT14 => N112421130, 
	DOUT15 => N112421131, 
	SIGNEDIN => N112396833, 
	SIGNEDOUT => N112421133
);
U142 : ADDERDELAY	PORT MAP(
	DIN0 => N110908416, 
	DIN1 => N110908417, 
	DIN2 => N110908418, 
	DIN3 => N110908419, 
	DIN4 => N110908420, 
	DIN5 => N110908421, 
	DIN6 => N110908422, 
	DIN7 => N110908423, 
	DIN8 => N110908424, 
	DIN9 => N110908425, 
	DIN10 => N110908426, 
	DIN11 => N110908427, 
	DIN12 => N110908428, 
	DIN13 => N110908429, 
	DIN14 => N110908430, 
	DIN15 => N110908431, 
	DOUT0 => N111643516, 
	DOUT1 => N111643517, 
	DOUT2 => N111643518, 
	DOUT3 => N111643519, 
	DOUT4 => N111643520, 
	DOUT5 => N111643521, 
	DOUT6 => N111643522, 
	DOUT7 => N111643523, 
	DOUT8 => N111643524, 
	DOUT9 => N111643525, 
	DOUT10 => N111643526, 
	DOUT11 => N111643527, 
	DOUT12 => N111643528, 
	DOUT13 => N111643529, 
	DOUT14 => N111643530, 
	DOUT15 => N111643531, 
	SIGNEDIN => N110908433, 
	SIGNEDOUT => N111643533
);
U111 : ADDERDELAY	PORT MAP(
	DIN0 => N11085600, 
	DIN1 => N11085601, 
	DIN2 => N11085602, 
	DIN3 => N11085603, 
	DIN4 => N11085604, 
	DIN5 => N11085605, 
	DIN6 => N11085606, 
	DIN7 => N11085607, 
	DIN8 => N11085608, 
	DIN9 => N11085609, 
	DIN10 => N110856010, 
	DIN11 => N110856011, 
	DIN12 => N110856012, 
	DIN13 => N110856013, 
	DIN14 => N110856014, 
	DIN15 => N110856015, 
	DOUT0 => N110856016, 
	DOUT1 => N110856017, 
	DOUT2 => N110856018, 
	DOUT3 => N110856019, 
	DOUT4 => N110856020, 
	DOUT5 => N110856021, 
	DOUT6 => N110856022, 
	DOUT7 => N110856023, 
	DOUT8 => N110856024, 
	DOUT9 => N110856025, 
	DOUT10 => N110856026, 
	DOUT11 => N110856027, 
	DOUT12 => N110856028, 
	DOUT13 => N110856029, 
	DOUT14 => N110856030, 
	DOUT15 => N110856031, 
	SIGNEDIN => N110856032, 
	SIGNEDOUT => N110856033
);
U175 : ADDERDELAY	PORT MAP(
	DIN0 => N111910816, 
	DIN1 => N111910817, 
	DIN2 => N111910818, 
	DIN3 => N111910819, 
	DIN4 => N111910820, 
	DIN5 => N111910821, 
	DIN6 => N111910822, 
	DIN7 => N111910823, 
	DIN8 => N111910824, 
	DIN9 => N111910825, 
	DIN10 => N111910826, 
	DIN11 => N111910827, 
	DIN12 => N111910828, 
	DIN13 => N111910829, 
	DIN14 => N111910830, 
	DIN15 => N111910831, 
	DOUT0 => N112445416, 
	DOUT1 => N112445417, 
	DOUT2 => N112445418, 
	DOUT3 => N112445419, 
	DOUT4 => N112445420, 
	DOUT5 => N112445421, 
	DOUT6 => N112445422, 
	DOUT7 => N112445423, 
	DOUT8 => N112445424, 
	DOUT9 => N112445425, 
	DOUT10 => N112445426, 
	DOUT11 => N112445427, 
	DOUT12 => N112445428, 
	DOUT13 => N112445429, 
	DOUT14 => N112445430, 
	DOUT15 => N112445431, 
	SIGNEDIN => N111910833, 
	SIGNEDOUT => N112445433
);
U143 : ADDERDELAY	PORT MAP(
	DIN0 => N111643516, 
	DIN1 => N111643517, 
	DIN2 => N111643518, 
	DIN3 => N111643519, 
	DIN4 => N111643520, 
	DIN5 => N111643521, 
	DIN6 => N111643522, 
	DIN7 => N111643523, 
	DIN8 => N111643524, 
	DIN9 => N111643525, 
	DIN10 => N111643526, 
	DIN11 => N111643527, 
	DIN12 => N111643528, 
	DIN13 => N111643529, 
	DIN14 => N111643530, 
	DIN15 => N111643531, 
	DOUT0 => N111667816, 
	DOUT1 => N111667817, 
	DOUT2 => N111667818, 
	DOUT3 => N111667819, 
	DOUT4 => N111667820, 
	DOUT5 => N111667821, 
	DOUT6 => N111667822, 
	DOUT7 => N111667823, 
	DOUT8 => N111667824, 
	DOUT9 => N111667825, 
	DOUT10 => N111667826, 
	DOUT11 => N111667827, 
	DOUT12 => N111667828, 
	DOUT13 => N111667829, 
	DOUT14 => N111667830, 
	DOUT15 => N111667831, 
	SIGNEDIN => N111643533, 
	SIGNEDOUT => N111667833
);
U176 : ADDERDELAY	PORT MAP(
	DIN0 => N112445416, 
	DIN1 => N112445417, 
	DIN2 => N112445418, 
	DIN3 => N112445419, 
	DIN4 => N112445420, 
	DIN5 => N112445421, 
	DIN6 => N112445422, 
	DIN7 => N112445423, 
	DIN8 => N112445424, 
	DIN9 => N112445425, 
	DIN10 => N112445426, 
	DIN11 => N112445427, 
	DIN12 => N112445428, 
	DIN13 => N112445429, 
	DIN14 => N112445430, 
	DIN15 => N112445431, 
	DOUT0 => N112469716, 
	DOUT1 => N112469717, 
	DOUT2 => N112469718, 
	DOUT3 => N112469719, 
	DOUT4 => N112469720, 
	DOUT5 => N112469721, 
	DOUT6 => N112469722, 
	DOUT7 => N112469723, 
	DOUT8 => N112469724, 
	DOUT9 => N112469725, 
	DOUT10 => N112469726, 
	DOUT11 => N112469727, 
	DOUT12 => N112469728, 
	DOUT13 => N112469729, 
	DOUT14 => N112469730, 
	DOUT15 => N112469731, 
	SIGNEDIN => N112445433, 
	SIGNEDOUT => N112469733
);
U144 : ADDERDELAY	PORT MAP(
	DIN0 => N111667816, 
	DIN1 => N111667817, 
	DIN2 => N111667818, 
	DIN3 => N111667819, 
	DIN4 => N111667820, 
	DIN5 => N111667821, 
	DIN6 => N111667822, 
	DIN7 => N111667823, 
	DIN8 => N111667824, 
	DIN9 => N111667825, 
	DIN10 => N111667826, 
	DIN11 => N111667827, 
	DIN12 => N111667828, 
	DIN13 => N111667829, 
	DIN14 => N111667830, 
	DIN15 => N111667831, 
	DOUT0 => N111692116, 
	DOUT1 => N111692117, 
	DOUT2 => N111692118, 
	DOUT3 => N111692119, 
	DOUT4 => N111692120, 
	DOUT5 => N111692121, 
	DOUT6 => N111692122, 
	DOUT7 => N111692123, 
	DOUT8 => N111692124, 
	DOUT9 => N111692125, 
	DOUT10 => N111692126, 
	DOUT11 => N111692127, 
	DOUT12 => N111692128, 
	DOUT13 => N111692129, 
	DOUT14 => N111692130, 
	DOUT15 => N111692131, 
	SIGNEDIN => N111667833, 
	SIGNEDOUT => N111692133
);
U112 : ADDERDELAY	PORT MAP(
	DIN0 => N110856016, 
	DIN1 => N110856017, 
	DIN2 => N110856018, 
	DIN3 => N110856019, 
	DIN4 => N110856020, 
	DIN5 => N110856021, 
	DIN6 => N110856022, 
	DIN7 => N110856023, 
	DIN8 => N110856024, 
	DIN9 => N110856025, 
	DIN10 => N110856026, 
	DIN11 => N110856027, 
	DIN12 => N110856028, 
	DIN13 => N110856029, 
	DIN14 => N110856030, 
	DIN15 => N110856031, 
	DOUT0 => N110884116, 
	DOUT1 => N110884117, 
	DOUT2 => N110884118, 
	DOUT3 => N110884119, 
	DOUT4 => N110884120, 
	DOUT5 => N110884121, 
	DOUT6 => N110884122, 
	DOUT7 => N110884123, 
	DOUT8 => N110884124, 
	DOUT9 => N110884125, 
	DOUT10 => N110884126, 
	DOUT11 => N110884127, 
	DOUT12 => N110884128, 
	DOUT13 => N110884129, 
	DOUT14 => N110884130, 
	DOUT15 => N110884131, 
	SIGNEDIN => N110856033, 
	SIGNEDOUT => N110884133
);
U177 : ADDERDELAY	PORT MAP(
	DIN0 => N112469716, 
	DIN1 => N112469717, 
	DIN2 => N112469718, 
	DIN3 => N112469719, 
	DIN4 => N112469720, 
	DIN5 => N112469721, 
	DIN6 => N112469722, 
	DIN7 => N112469723, 
	DIN8 => N112469724, 
	DIN9 => N112469725, 
	DIN10 => N112469726, 
	DIN11 => N112469727, 
	DIN12 => N112469728, 
	DIN13 => N112469729, 
	DIN14 => N112469730, 
	DIN15 => N112469731, 
	DOUT0 => N112494016, 
	DOUT1 => N112494017, 
	DOUT2 => N112494018, 
	DOUT3 => N112494019, 
	DOUT4 => N112494020, 
	DOUT5 => N112494021, 
	DOUT6 => N112494022, 
	DOUT7 => N112494023, 
	DOUT8 => N112494024, 
	DOUT9 => N112494025, 
	DOUT10 => N112494026, 
	DOUT11 => N112494027, 
	DOUT12 => N112494028, 
	DOUT13 => N112494029, 
	DOUT14 => N112494030, 
	DOUT15 => N112494031, 
	SIGNEDIN => N112469733, 
	SIGNEDOUT => N112494033
);
U145 : ADDERDELAY	PORT MAP(
	DIN0 => N110985116, 
	DIN1 => N110985117, 
	DIN2 => N110985118, 
	DIN3 => N110985119, 
	DIN4 => N110985120, 
	DIN5 => N110985121, 
	DIN6 => N110985122, 
	DIN7 => N110985123, 
	DIN8 => N110985124, 
	DIN9 => N110985125, 
	DIN10 => N110985126, 
	DIN11 => N110985127, 
	DIN12 => N110985128, 
	DIN13 => N110985129, 
	DIN14 => N110985130, 
	DIN15 => N110985131, 
	DOUT0 => N111716416, 
	DOUT1 => N111716417, 
	DOUT2 => N111716418, 
	DOUT3 => N111716419, 
	DOUT4 => N111716420, 
	DOUT5 => N111716421, 
	DOUT6 => N111716422, 
	DOUT7 => N111716423, 
	DOUT8 => N111716424, 
	DOUT9 => N111716425, 
	DOUT10 => N111716426, 
	DOUT11 => N111716427, 
	DOUT12 => N111716428, 
	DOUT13 => N111716429, 
	DOUT14 => N111716430, 
	DOUT15 => N111716431, 
	SIGNEDIN => N110985133, 
	SIGNEDOUT => N111716433
);
U113 : ADDERDELAY	PORT MAP(
	DIN0 => N110884116, 
	DIN1 => N110884117, 
	DIN2 => N110884118, 
	DIN3 => N110884119, 
	DIN4 => N110884120, 
	DIN5 => N110884121, 
	DIN6 => N110884122, 
	DIN7 => N110884123, 
	DIN8 => N110884124, 
	DIN9 => N110884125, 
	DIN10 => N110884126, 
	DIN11 => N110884127, 
	DIN12 => N110884128, 
	DIN13 => N110884129, 
	DIN14 => N110884130, 
	DIN15 => N110884131, 
	DOUT0 => N110908416, 
	DOUT1 => N110908417, 
	DOUT2 => N110908418, 
	DOUT3 => N110908419, 
	DOUT4 => N110908420, 
	DOUT5 => N110908421, 
	DOUT6 => N110908422, 
	DOUT7 => N110908423, 
	DOUT8 => N110908424, 
	DOUT9 => N110908425, 
	DOUT10 => N110908426, 
	DOUT11 => N110908427, 
	DOUT12 => N110908428, 
	DOUT13 => N110908429, 
	DOUT14 => N110908430, 
	DOUT15 => N110908431, 
	SIGNEDIN => N110884133, 
	SIGNEDOUT => N110908433
);
U178 : ADDERDELAY	PORT MAP(
	DIN0 => N112494016, 
	DIN1 => N112494017, 
	DIN2 => N112494018, 
	DIN3 => N112494019, 
	DIN4 => N112494020, 
	DIN5 => N112494021, 
	DIN6 => N112494022, 
	DIN7 => N112494023, 
	DIN8 => N112494024, 
	DIN9 => N112494025, 
	DIN10 => N112494026, 
	DIN11 => N112494027, 
	DIN12 => N112494028, 
	DIN13 => N112494029, 
	DIN14 => N112494030, 
	DIN15 => N112494031, 
	DOUT0 => N112518316, 
	DOUT1 => N112518317, 
	DOUT2 => N112518318, 
	DOUT3 => N112518319, 
	DOUT4 => N112518320, 
	DOUT5 => N112518321, 
	DOUT6 => N112518322, 
	DOUT7 => N112518323, 
	DOUT8 => N112518324, 
	DOUT9 => N112518325, 
	DOUT10 => N112518326, 
	DOUT11 => N112518327, 
	DOUT12 => N112518328, 
	DOUT13 => N112518329, 
	DOUT14 => N112518330, 
	DOUT15 => N112518331, 
	SIGNEDIN => N112494033, 
	SIGNEDOUT => N112518333
);
U146 : ADDERDELAY	PORT MAP(
	DIN0 => N111716416, 
	DIN1 => N111716417, 
	DIN2 => N111716418, 
	DIN3 => N111716419, 
	DIN4 => N111716420, 
	DIN5 => N111716421, 
	DIN6 => N111716422, 
	DIN7 => N111716423, 
	DIN8 => N111716424, 
	DIN9 => N111716425, 
	DIN10 => N111716426, 
	DIN11 => N111716427, 
	DIN12 => N111716428, 
	DIN13 => N111716429, 
	DIN14 => N111716430, 
	DIN15 => N111716431, 
	DOUT0 => N111740716, 
	DOUT1 => N111740717, 
	DOUT2 => N111740718, 
	DOUT3 => N111740719, 
	DOUT4 => N111740720, 
	DOUT5 => N111740721, 
	DOUT6 => N111740722, 
	DOUT7 => N111740723, 
	DOUT8 => N111740724, 
	DOUT9 => N111740725, 
	DOUT10 => N111740726, 
	DOUT11 => N111740727, 
	DOUT12 => N111740728, 
	DOUT13 => N111740729, 
	DOUT14 => N111740730, 
	DOUT15 => N111740731, 
	SIGNEDIN => N111716433, 
	SIGNEDOUT => N111740733
);
U114 : ADDERDELAY	PORT MAP(
	DIN0 => N11093270, 
	DIN1 => N11093271, 
	DIN2 => N11093272, 
	DIN3 => N11093273, 
	DIN4 => N11093274, 
	DIN5 => N11093275, 
	DIN6 => N11093276, 
	DIN7 => N11093277, 
	DIN8 => N11093278, 
	DIN9 => N11093279, 
	DIN10 => N110932710, 
	DIN11 => N110932711, 
	DIN12 => N110932712, 
	DIN13 => N110932713, 
	DIN14 => N110932714, 
	DIN15 => N110932715, 
	DOUT0 => N110932716, 
	DOUT1 => N110932717, 
	DOUT2 => N110932718, 
	DOUT3 => N110932719, 
	DOUT4 => N110932720, 
	DOUT5 => N110932721, 
	DOUT6 => N110932722, 
	DOUT7 => N110932723, 
	DOUT8 => N110932724, 
	DOUT9 => N110932725, 
	DOUT10 => N110932726, 
	DOUT11 => N110932727, 
	DOUT12 => N110932728, 
	DOUT13 => N110932729, 
	DOUT14 => N110932730, 
	DOUT15 => N110932731, 
	SIGNEDIN => N110932732, 
	SIGNEDOUT => N110932733
);
U179 : ADDERDELAY	PORT MAP(
	DIN0 => N111983716, 
	DIN1 => N111983717, 
	DIN2 => N111983718, 
	DIN3 => N111983719, 
	DIN4 => N111983720, 
	DIN5 => N111983721, 
	DIN6 => N111983722, 
	DIN7 => N111983723, 
	DIN8 => N111983724, 
	DIN9 => N111983725, 
	DIN10 => N111983726, 
	DIN11 => N111983727, 
	DIN12 => N111983728, 
	DIN13 => N111983729, 
	DIN14 => N111983730, 
	DIN15 => N111983731, 
	DOUT0 => N112542616, 
	DOUT1 => N112542617, 
	DOUT2 => N112542618, 
	DOUT3 => N112542619, 
	DOUT4 => N112542620, 
	DOUT5 => N112542621, 
	DOUT6 => N112542622, 
	DOUT7 => N112542623, 
	DOUT8 => N112542624, 
	DOUT9 => N112542625, 
	DOUT10 => N112542626, 
	DOUT11 => N112542627, 
	DOUT12 => N112542628, 
	DOUT13 => N112542629, 
	DOUT14 => N112542630, 
	DOUT15 => N112542631, 
	SIGNEDIN => N111983733, 
	SIGNEDOUT => N112542633
);
U147 : ADDERDELAY	PORT MAP(
	DIN0 => N111740716, 
	DIN1 => N111740717, 
	DIN2 => N111740718, 
	DIN3 => N111740719, 
	DIN4 => N111740720, 
	DIN5 => N111740721, 
	DIN6 => N111740722, 
	DIN7 => N111740723, 
	DIN8 => N111740724, 
	DIN9 => N111740725, 
	DIN10 => N111740726, 
	DIN11 => N111740727, 
	DIN12 => N111740728, 
	DIN13 => N111740729, 
	DIN14 => N111740730, 
	DIN15 => N111740731, 
	DOUT0 => N111765016, 
	DOUT1 => N111765017, 
	DOUT2 => N111765018, 
	DOUT3 => N111765019, 
	DOUT4 => N111765020, 
	DOUT5 => N111765021, 
	DOUT6 => N111765022, 
	DOUT7 => N111765023, 
	DOUT8 => N111765024, 
	DOUT9 => N111765025, 
	DOUT10 => N111765026, 
	DOUT11 => N111765027, 
	DOUT12 => N111765028, 
	DOUT13 => N111765029, 
	DOUT14 => N111765030, 
	DOUT15 => N111765031, 
	SIGNEDIN => N111740733, 
	SIGNEDOUT => N111765033
);
U115 : ADDERDELAY	PORT MAP(
	DIN0 => N110932716, 
	DIN1 => N110932717, 
	DIN2 => N110932718, 
	DIN3 => N110932719, 
	DIN4 => N110932720, 
	DIN5 => N110932721, 
	DIN6 => N110932722, 
	DIN7 => N110932723, 
	DIN8 => N110932724, 
	DIN9 => N110932725, 
	DIN10 => N110932726, 
	DIN11 => N110932727, 
	DIN12 => N110932728, 
	DIN13 => N110932729, 
	DIN14 => N110932730, 
	DIN15 => N110932731, 
	DOUT0 => N110960816, 
	DOUT1 => N110960817, 
	DOUT2 => N110960818, 
	DOUT3 => N110960819, 
	DOUT4 => N110960820, 
	DOUT5 => N110960821, 
	DOUT6 => N110960822, 
	DOUT7 => N110960823, 
	DOUT8 => N110960824, 
	DOUT9 => N110960825, 
	DOUT10 => N110960826, 
	DOUT11 => N110960827, 
	DOUT12 => N110960828, 
	DOUT13 => N110960829, 
	DOUT14 => N110960830, 
	DOUT15 => N110960831, 
	SIGNEDIN => N110932733, 
	SIGNEDOUT => N110960833
);
U148 : ADDERDELAY	PORT MAP(
	DIN0 => N111061816, 
	DIN1 => N111061817, 
	DIN2 => N111061818, 
	DIN3 => N111061819, 
	DIN4 => N111061820, 
	DIN5 => N111061821, 
	DIN6 => N111061822, 
	DIN7 => N111061823, 
	DIN8 => N111061824, 
	DIN9 => N111061825, 
	DIN10 => N111061826, 
	DIN11 => N111061827, 
	DIN12 => N111061828, 
	DIN13 => N111061829, 
	DIN14 => N111061830, 
	DIN15 => N111061831, 
	DOUT0 => N111789316, 
	DOUT1 => N111789317, 
	DOUT2 => N111789318, 
	DOUT3 => N111789319, 
	DOUT4 => N111789320, 
	DOUT5 => N111789321, 
	DOUT6 => N111789322, 
	DOUT7 => N111789323, 
	DOUT8 => N111789324, 
	DOUT9 => N111789325, 
	DOUT10 => N111789326, 
	DOUT11 => N111789327, 
	DOUT12 => N111789328, 
	DOUT13 => N111789329, 
	DOUT14 => N111789330, 
	DOUT15 => N111789331, 
	SIGNEDIN => N111061833, 
	SIGNEDOUT => N111789333
);
U116 : ADDERDELAY	PORT MAP(
	DIN0 => N110960816, 
	DIN1 => N110960817, 
	DIN2 => N110960818, 
	DIN3 => N110960819, 
	DIN4 => N110960820, 
	DIN5 => N110960821, 
	DIN6 => N110960822, 
	DIN7 => N110960823, 
	DIN8 => N110960824, 
	DIN9 => N110960825, 
	DIN10 => N110960826, 
	DIN11 => N110960827, 
	DIN12 => N110960828, 
	DIN13 => N110960829, 
	DIN14 => N110960830, 
	DIN15 => N110960831, 
	DOUT0 => N110985116, 
	DOUT1 => N110985117, 
	DOUT2 => N110985118, 
	DOUT3 => N110985119, 
	DOUT4 => N110985120, 
	DOUT5 => N110985121, 
	DOUT6 => N110985122, 
	DOUT7 => N110985123, 
	DOUT8 => N110985124, 
	DOUT9 => N110985125, 
	DOUT10 => N110985126, 
	DOUT11 => N110985127, 
	DOUT12 => N110985128, 
	DOUT13 => N110985129, 
	DOUT14 => N110985130, 
	DOUT15 => N110985131, 
	SIGNEDIN => N110960833, 
	SIGNEDOUT => N110985133
);
U149 : ADDERDELAY	PORT MAP(
	DIN0 => N111789316, 
	DIN1 => N111789317, 
	DIN2 => N111789318, 
	DIN3 => N111789319, 
	DIN4 => N111789320, 
	DIN5 => N111789321, 
	DIN6 => N111789322, 
	DIN7 => N111789323, 
	DIN8 => N111789324, 
	DIN9 => N111789325, 
	DIN10 => N111789326, 
	DIN11 => N111789327, 
	DIN12 => N111789328, 
	DIN13 => N111789329, 
	DIN14 => N111789330, 
	DIN15 => N111789331, 
	DOUT0 => N111813616, 
	DOUT1 => N111813617, 
	DOUT2 => N111813618, 
	DOUT3 => N111813619, 
	DOUT4 => N111813620, 
	DOUT5 => N111813621, 
	DOUT6 => N111813622, 
	DOUT7 => N111813623, 
	DOUT8 => N111813624, 
	DOUT9 => N111813625, 
	DOUT10 => N111813626, 
	DOUT11 => N111813627, 
	DOUT12 => N111813628, 
	DOUT13 => N111813629, 
	DOUT14 => N111813630, 
	DOUT15 => N111813631, 
	SIGNEDIN => N111789333, 
	SIGNEDOUT => N111813633
);
U117 : ADDERDELAY	PORT MAP(
	DIN0 => N11100940, 
	DIN1 => N11100941, 
	DIN2 => N11100942, 
	DIN3 => N11100943, 
	DIN4 => N11100944, 
	DIN5 => N11100945, 
	DIN6 => N11100946, 
	DIN7 => N11100947, 
	DIN8 => N11100948, 
	DIN9 => N11100949, 
	DIN10 => N111009410, 
	DIN11 => N111009411, 
	DIN12 => N111009412, 
	DIN13 => N111009413, 
	DIN14 => N111009414, 
	DIN15 => N111009415, 
	DOUT0 => N111009416, 
	DOUT1 => N111009417, 
	DOUT2 => N111009418, 
	DOUT3 => N111009419, 
	DOUT4 => N111009420, 
	DOUT5 => N111009421, 
	DOUT6 => N111009422, 
	DOUT7 => N111009423, 
	DOUT8 => N111009424, 
	DOUT9 => N111009425, 
	DOUT10 => N111009426, 
	DOUT11 => N111009427, 
	DOUT12 => N111009428, 
	DOUT13 => N111009429, 
	DOUT14 => N111009430, 
	DOUT15 => N111009431, 
	SIGNEDIN => N111009432, 
	SIGNEDOUT => N111009433
);
U118 : ADDERDELAY	PORT MAP(
	DIN0 => N111009416, 
	DIN1 => N111009417, 
	DIN2 => N111009418, 
	DIN3 => N111009419, 
	DIN4 => N111009420, 
	DIN5 => N111009421, 
	DIN6 => N111009422, 
	DIN7 => N111009423, 
	DIN8 => N111009424, 
	DIN9 => N111009425, 
	DIN10 => N111009426, 
	DIN11 => N111009427, 
	DIN12 => N111009428, 
	DIN13 => N111009429, 
	DIN14 => N111009430, 
	DIN15 => N111009431, 
	DOUT0 => N111037516, 
	DOUT1 => N111037517, 
	DOUT2 => N111037518, 
	DOUT3 => N111037519, 
	DOUT4 => N111037520, 
	DOUT5 => N111037521, 
	DOUT6 => N111037522, 
	DOUT7 => N111037523, 
	DOUT8 => N111037524, 
	DOUT9 => N111037525, 
	DOUT10 => N111037526, 
	DOUT11 => N111037527, 
	DOUT12 => N111037528, 
	DOUT13 => N111037529, 
	DOUT14 => N111037530, 
	DOUT15 => N111037531, 
	SIGNEDIN => N111009433, 
	SIGNEDOUT => N111037533
);
U119 : ADDERDELAY	PORT MAP(
	DIN0 => N111037516, 
	DIN1 => N111037517, 
	DIN2 => N111037518, 
	DIN3 => N111037519, 
	DIN4 => N111037520, 
	DIN5 => N111037521, 
	DIN6 => N111037522, 
	DIN7 => N111037523, 
	DIN8 => N111037524, 
	DIN9 => N111037525, 
	DIN10 => N111037526, 
	DIN11 => N111037527, 
	DIN12 => N111037528, 
	DIN13 => N111037529, 
	DIN14 => N111037530, 
	DIN15 => N111037531, 
	DOUT0 => N111061816, 
	DOUT1 => N111061817, 
	DOUT2 => N111061818, 
	DOUT3 => N111061819, 
	DOUT4 => N111061820, 
	DOUT5 => N111061821, 
	DOUT6 => N111061822, 
	DOUT7 => N111061823, 
	DOUT8 => N111061824, 
	DOUT9 => N111061825, 
	DOUT10 => N111061826, 
	DOUT11 => N111061827, 
	DOUT12 => N111061828, 
	DOUT13 => N111061829, 
	DOUT14 => N111061830, 
	DOUT15 => N111061831, 
	SIGNEDIN => N111037533, 
	SIGNEDOUT => N111061833
);
U70 : \7408\	PORT MAP(
	A_A => N94151, 
	B_A => N94145, 
	Y_A => N955836, 
	VCC => VCC, 
	GND => GND, 
	A_B => 'Z', 
	B_B => 'Z', 
	Y_B => OPEN, 
	A_C => 'Z', 
	B_C => 'Z', 
	Y_C => OPEN, 
	A_D => 'Z', 
	B_D => 'Z', 
	Y_D => OPEN
);
U71 : ADDERDELAY	PORT MAP(
	DIN0 => N10716200, 
	DIN1 => N10716201, 
	DIN2 => N10716202, 
	DIN3 => N10716203, 
	DIN4 => N10716204, 
	DIN5 => N10716205, 
	DIN6 => N10716206, 
	DIN7 => N10716207, 
	DIN8 => N10716208, 
	DIN9 => N10716209, 
	DIN10 => N107162010, 
	DIN11 => N107162011, 
	DIN12 => N107162012, 
	DIN13 => N107162013, 
	DIN14 => N107162014, 
	DIN15 => N107162015, 
	DOUT0 => N1143146, 
	DOUT1 => N1143067, 
	DOUT2 => N1142988, 
	DOUT3 => N1142909, 
	DOUT4 => N1142830, 
	DOUT5 => N1142751, 
	DOUT6 => N1142672, 
	DOUT7 => N1142593, 
	DOUT8 => N1142514, 
	DOUT9 => N1142435, 
	DOUT10 => N1142356, 
	DOUT11 => N1142277, 
	DOUT12 => N1142198, 
	DOUT13 => N1142119, 
	DOUT14 => N1142040, 
	DOUT15 => N1141961, 
	SIGNEDIN => N107162032, 
	SIGNEDOUT => N1141882
);
U40 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => N81765, 
	DCO1 => N81767, 
	DCO2 => N81769, 
	DCO3 => N81771, 
	DCO4 => N81773, 
	DCO5 => N81775, 
	DCO6 => N81777, 
	DCO7 => N81779, 
	DSG0 => N81781, 
	DSG1 => N81783, 
	DSG2 => N81785, 
	DSG3 => N81787, 
	DSG4 => N81789, 
	DSG5 => N81791, 
	DSG6 => N81793, 
	DSG7 => N81795, 
	ENABLE => ENABLE9, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => N80950, 
	QCO1 => N80952, 
	QCO2 => N80954, 
	QCO3 => N80956, 
	QCO4 => N80958, 
	QCO5 => N80960, 
	QCO6 => N80962, 
	QCO7 => N80964, 
	QSG0 => N80966, 
	QSG1 => N80968, 
	QSG2 => N80970, 
	QSG3 => N80972, 
	QSG4 => N80974, 
	QSG5 => N80976, 
	QSG6 => N80978, 
	QSG7 => N80980, 
	S0 => N11070260, 
	S1 => N11070261, 
	S2 => N11070262, 
	S3 => N11070263, 
	S4 => N11070264, 
	S5 => N11070265, 
	S6 => N11070266, 
	S7 => N11070267, 
	S8 => N11070268, 
	S9 => N11070269, 
	S10 => N110702610, 
	S11 => N110702611, 
	S12 => N110702612, 
	S13 => N110702613, 
	S14 => N110702614, 
	S15 => N110702615, 
	SIGNED => N110702632
);
U41 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => N80950, 
	DCO1 => N80952, 
	DCO2 => N80954, 
	DCO3 => N80956, 
	DCO4 => N80958, 
	DCO5 => N80960, 
	DCO6 => N80962, 
	DCO7 => N80964, 
	DSG0 => N80966, 
	DSG1 => N80968, 
	DSG2 => N80970, 
	DSG3 => N80972, 
	DSG4 => N80974, 
	DSG5 => N80976, 
	DSG6 => N80978, 
	DSG7 => N80980, 
	ENABLE => ENABLE10, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => N80137, 
	QCO1 => N80139, 
	QCO2 => N80141, 
	QCO3 => N80143, 
	QCO4 => N80145, 
	QCO5 => N80147, 
	QCO6 => N80149, 
	QCO7 => N80151, 
	QSG0 => N80153, 
	QSG1 => N80155, 
	QSG2 => N80157, 
	QSG3 => N80159, 
	QSG4 => N80161, 
	QSG5 => N80163, 
	QSG6 => N80165, 
	QSG7 => N80167, 
	S0 => N11077930, 
	S1 => N11077931, 
	S2 => N11077932, 
	S3 => N11077933, 
	S4 => N11077934, 
	S5 => N11077935, 
	S6 => N11077936, 
	S7 => N11077937, 
	S8 => N11077938, 
	S9 => N11077939, 
	S10 => N110779310, 
	S11 => N110779311, 
	S12 => N110779312, 
	S13 => N110779313, 
	S14 => N110779314, 
	S15 => N110779315, 
	SIGNED => N110779332
);
U74 : ENABLEALL	PORT MAP(
	C0 => N94151, 
	C1 => N94153, 
	C2 => N94155, 
	C3 => N94157, 
	ENABLEELEVEN => ENABLE11, 
	ENABLEFIFTEEN => ENABLE15, 
	ENABLEFIVE => ENABLE5, 
	ENABLEFOUR => ENABLE4, 
	ENABLEFOURTEEN => ENABLE14, 
	ENABLENINE => ENABLE9, 
	ENABLEONE => ENABLE1, 
	ENABLESEVEN => ENABLE7, 
	ENABLESIX => ENABLE6, 
	ENABLETEN => ENABLE10, 
	ENABLETHIRTEEN => ENABLE13, 
	ENABLETHREE => ENABLE3, 
	ENABLETWELVE => ENABLE12, 
	ENABLETWO => ENABLE2, 
	NC0 => N94143, 
	NC1 => N94145, 
	NC2 => N94147
);
U42 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => N80137, 
	DCO1 => N80139, 
	DCO2 => N80141, 
	DCO3 => N80143, 
	DCO4 => N80145, 
	DCO5 => N80147, 
	DCO6 => N80149, 
	DCO7 => N80151, 
	DSG0 => N80153, 
	DSG1 => N80155, 
	DSG2 => N80157, 
	DSG3 => N80159, 
	DSG4 => N80161, 
	DSG5 => N80163, 
	DSG6 => N80165, 
	DSG7 => N80167, 
	ENABLE => ENABLE11, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => N79322, 
	QCO1 => N79324, 
	QCO2 => N79326, 
	QCO3 => N79328, 
	QCO4 => N79330, 
	QCO5 => N79332, 
	QCO6 => N79334, 
	QCO7 => N79336, 
	QSG0 => N79338, 
	QSG1 => N79340, 
	QSG2 => N79342, 
	QSG3 => N79344, 
	QSG4 => N79346, 
	QSG5 => N79348, 
	QSG6 => N79350, 
	QSG7 => N79352, 
	S0 => N11085600, 
	S1 => N11085601, 
	S2 => N11085602, 
	S3 => N11085603, 
	S4 => N11085604, 
	S5 => N11085605, 
	S6 => N11085606, 
	S7 => N11085607, 
	S8 => N11085608, 
	S9 => N11085609, 
	S10 => N110856010, 
	S11 => N110856011, 
	S12 => N110856012, 
	S13 => N110856013, 
	S14 => N110856014, 
	S15 => N110856015, 
	SIGNED => N110856032
);
U43 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => N79322, 
	DCO1 => N79324, 
	DCO2 => N79326, 
	DCO3 => N79328, 
	DCO4 => N79330, 
	DCO5 => N79332, 
	DCO6 => N79334, 
	DCO7 => N79336, 
	DSG0 => N79338, 
	DSG1 => N79340, 
	DSG2 => N79342, 
	DSG3 => N79344, 
	DSG4 => N79346, 
	DSG5 => N79348, 
	DSG6 => N79350, 
	DSG7 => N79352, 
	ENABLE => ENABLE12, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => N78509, 
	QCO1 => N78511, 
	QCO2 => N78513, 
	QCO3 => N78515, 
	QCO4 => N78517, 
	QCO5 => N78519, 
	QCO6 => N78521, 
	QCO7 => N78523, 
	QSG0 => N78525, 
	QSG1 => N78527, 
	QSG2 => N78529, 
	QSG3 => N78531, 
	QSG4 => N78533, 
	QSG5 => N78535, 
	QSG6 => N78537, 
	QSG7 => N78539, 
	S0 => N11093270, 
	S1 => N11093271, 
	S2 => N11093272, 
	S3 => N11093273, 
	S4 => N11093274, 
	S5 => N11093275, 
	S6 => N11093276, 
	S7 => N11093277, 
	S8 => N11093278, 
	S9 => N11093279, 
	S10 => N110932710, 
	S11 => N110932711, 
	S12 => N110932712, 
	S13 => N110932713, 
	S14 => N110932714, 
	S15 => N110932715, 
	SIGNED => N110932732
);
U44 : NEWSLICE	PORT MAP(
	CLK => CLK, 
	DCO0 => N78509, 
	DCO1 => N78511, 
	DCO2 => N78513, 
	DCO3 => N78515, 
	DCO4 => N78517, 
	DCO5 => N78519, 
	DCO6 => N78521, 
	DCO7 => N78523, 
	DSG0 => N78525, 
	DSG1 => N78527, 
	DSG2 => N78529, 
	DSG3 => N78531, 
	DSG4 => N78533, 
	DSG5 => N78535, 
	DSG6 => N78537, 
	DSG7 => N78539, 
	ENABLE => ENABLE13, 
	LOAD => LOAD, 
	NRST => NRST, 
	QCO0 => N77694, 
	QCO1 => N77696, 
	QCO2 => N77698, 
	QCO3 => N77700, 
	QCO4 => N77702, 
	QCO5 => N77704, 
	QCO6 => N77706, 
	QCO7 => N77708, 
	QSG0 => N77710, 
	QSG1 => N77712, 
	QSG2 => N77714, 
	QSG3 => N77716, 
	QSG4 => N77718, 
	QSG5 => N77720, 
	QSG6 => N77722, 
	QSG7 => N77724, 
	S0 => N11100940, 
	S1 => N11100941, 
	S2 => N11100942, 
	S3 => N11100943, 
	S4 => N11100944, 
	S5 => N11100945, 
	S6 => N11100946, 
	S7 => N11100947, 
	S8 => N11100948, 
	S9 => N11100949, 
	S10 => N111009410, 
	S11 => N111009411, 
	S12 => N111009412, 
	S13 => N111009413, 
	S14 => N111009414, 
	S15 => N111009415, 
	SIGNED => N111009432
);
END STRUCTURE;

