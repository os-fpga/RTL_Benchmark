// Copyright (C) 2022, Andes Technology Corp. Confidential Proprietary

module kv_csr_dec #(
    parameter FLEN = 1,
    parameter RVN_SUPPORT_INT = 0,
    parameter RVV_SUPPORT_INT = 0,
    parameter DSP_SUPPORT_INT = 0,
    parameter ACE_SUPPORT_INT = 0,
    parameter NUM_PRIVILEGE_LEVELS = 1,
    parameter PERFORMANCE_MONITOR_INT = 0,
    parameter POWERBRAKE_SUPPORT_INT = 0,
    parameter STACKSAFE_SUPPORT_INT = 0,
    parameter CODENSE_SUPPORT_INT = 0,
    parameter CACHE_SUPPORT_INT = 0,
    parameter ICACHE_ECC_TYPE_INT = 0,
    parameter ECC_SUPPORT_INT = 0,
    parameter MMISC_CTL_EXIST_INT = 0,
    parameter MMSC_CFG2_EXIST_INT = 0,
    parameter ILM_SIZE_KB = 0,
    parameter DLM_SIZE_KB = 0,
    parameter PMA_ENTRIES = 0,
    parameter HAS_VPU_INT = 0,
    parameter XLEN = 64)  (
    existent_csr,
    privileged_csr,
    privileged_csr_ddcause,
    readonly_csr,
    csr_cur_privilege,
    csr_halt_mode,
    cur_privilege_m,
    cur_privilege_s,
    cur_privilege_u,
    csr_mcache_ctl_cctl_suen,
    csr_mstatus_tvm,
    csr_mcounteren,
    csr_mcounterwen,
    csr_scounteren,
    writeonly_csr,
    func_csr,
    csr_ucctlcommand_privileged,
    rd_index,
    csr_addr
);
output existent_csr;
output privileged_csr;
output privileged_csr_ddcause;
output readonly_csr;
input [1:0] csr_cur_privilege;
input csr_halt_mode;
input cur_privilege_m;
input cur_privilege_s;
input cur_privilege_u;
input csr_mcache_ctl_cctl_suen;
input csr_mstatus_tvm;
input [31:0] csr_mcounteren;
input [31:0] csr_mcounterwen;
input [31:0] csr_scounteren;
input writeonly_csr;
input [1:0] func_csr;
input csr_ucctlcommand_privileged;
input [4:0] rd_index;
input [11:0] csr_addr;


localparam PRIVILEGE_USER = 2'b00;
localparam PRIVILEGE_SUPERVISOR = 2'b01;
localparam PRIVILEGE_MACHINE = 2'b11;
wire s0 = (NUM_PRIVILEGE_LEVELS > 2);
wire s1 = (NUM_PRIVILEGE_LEVELS == 2);
wire s2 = (NUM_PRIVILEGE_LEVELS > 1);
wire s3 = cur_privilege_s | cur_privilege_u;
wire s4 = cur_privilege_m | cur_privilege_s;
wire s5;
localparam CSR12_FFLAGS = 12'h001;
localparam CSR12_FRM = 12'h002;
localparam CSR12_FCSR = 12'h003;
localparam CSR12_SSTATUS = 12'h100;
localparam CSR12_SIE = 12'h104;
localparam CSR12_SIP = 12'h144;
localparam CSR12_SIDELEG = 12'h103;
localparam CSR12_SEDELEG = 12'h102;
localparam CSR12_STVEC = 12'h105;
localparam CSR12_SCOUNTEREN = 12'h106;
localparam CSR12_SEPC = 12'h141;
localparam CSR12_SCAUSE = 12'h142;
localparam CSR12_STVAL = 12'h143;
localparam CSR12_SSCRATCH = 12'h140;
localparam CSR12_SATP = 12'h180;
localparam CSR12_SLIE = 12'h9c4;
localparam CSR12_SLIP = 12'h9c5;
localparam CSR12_SDCAUSE = 12'h9c9;
localparam CSR12_MVENDORID = 12'hf11;
localparam CSR12_MARCHID = 12'hf12;
localparam CSR12_MIMPID = 12'hf13;
localparam CSR12_MHARTID = 12'hf14;
localparam CSR12_MSTATUS = 12'h300;
localparam CSR12_MISA = 12'h301;
localparam CSR12_MEDELEG = 12'h302;
localparam CSR12_MIDELEG = 12'h303;
localparam CSR12_MIE = 12'h304;
localparam CSR12_MTVEC = 12'h305;
localparam CSR12_MCOUNTEREN = 12'h306;
localparam CSR12_MCOUNTINHIBIT = 12'h320;
localparam CSR12_MSCRATCH = 12'h340;
localparam CSR12_MEPC = 12'h341;
localparam CSR12_MCAUSE = 12'h342;
localparam CSR12_MTVAL = 12'h343;
localparam CSR12_MIP = 12'h344;
localparam CSR12_MCYCLE = 12'hb00;
localparam CSR12_MINSTRET = 12'hb02;
localparam CSR12_MHPMCOUNTER3 = 12'hb03;
localparam CSR12_MHPMCOUNTER4 = 12'hb04;
localparam CSR12_MHPMCOUNTER5 = 12'hb05;
localparam CSR12_MHPMCOUNTER6 = 12'hb06;
localparam CSR12_MHPMCOUNTER7 = 12'hb07;
localparam CSR12_MHPMCOUNTER8 = 12'hb08;
localparam CSR12_MHPMCOUNTER9 = 12'hb09;
localparam CSR12_MHPMCOUNTER10 = 12'hb0a;
localparam CSR12_MHPMCOUNTER11 = 12'hb0b;
localparam CSR12_MHPMCOUNTER12 = 12'hb0c;
localparam CSR12_MHPMCOUNTER13 = 12'hb0d;
localparam CSR12_MHPMCOUNTER14 = 12'hb0e;
localparam CSR12_MHPMCOUNTER15 = 12'hb0f;
localparam CSR12_MHPMCOUNTER16 = 12'hb10;
localparam CSR12_MHPMCOUNTER17 = 12'hb11;
localparam CSR12_MHPMCOUNTER18 = 12'hb12;
localparam CSR12_MHPMCOUNTER19 = 12'hb13;
localparam CSR12_MHPMCOUNTER20 = 12'hb14;
localparam CSR12_MHPMCOUNTER21 = 12'hb15;
localparam CSR12_MHPMCOUNTER22 = 12'hb16;
localparam CSR12_MHPMCOUNTER23 = 12'hb17;
localparam CSR12_MHPMCOUNTER24 = 12'hb18;
localparam CSR12_MHPMCOUNTER25 = 12'hb19;
localparam CSR12_MHPMCOUNTER26 = 12'hb1a;
localparam CSR12_MHPMCOUNTER27 = 12'hb1b;
localparam CSR12_MHPMCOUNTER28 = 12'hb1c;
localparam CSR12_MHPMCOUNTER29 = 12'hb1d;
localparam CSR12_MHPMCOUNTER30 = 12'hb1e;
localparam CSR12_MHPMCOUNTER31 = 12'hb1f;
localparam CSR12_MCYCLEH = 12'hb80;
localparam CSR12_MINSTRETH = 12'hb82;
localparam CSR12_MHPMCOUNTER3H = 12'hb83;
localparam CSR12_MHPMCOUNTER4H = 12'hb84;
localparam CSR12_MHPMCOUNTER5H = 12'hb85;
localparam CSR12_MHPMCOUNTER6H = 12'hb86;
localparam CSR12_MHPMCOUNTER7H = 12'hb87;
localparam CSR12_MHPMCOUNTER8H = 12'hb88;
localparam CSR12_MHPMCOUNTER9H = 12'hb89;
localparam CSR12_MHPMCOUNTER10H = 12'hb8a;
localparam CSR12_MHPMCOUNTER11H = 12'hb8b;
localparam CSR12_MHPMCOUNTER12H = 12'hb8c;
localparam CSR12_MHPMCOUNTER13H = 12'hb8d;
localparam CSR12_MHPMCOUNTER14H = 12'hb8e;
localparam CSR12_MHPMCOUNTER15H = 12'hb8f;
localparam CSR12_MHPMCOUNTER16H = 12'hb90;
localparam CSR12_MHPMCOUNTER17H = 12'hb91;
localparam CSR12_MHPMCOUNTER18H = 12'hb92;
localparam CSR12_MHPMCOUNTER19H = 12'hb93;
localparam CSR12_MHPMCOUNTER20H = 12'hb94;
localparam CSR12_MHPMCOUNTER21H = 12'hb95;
localparam CSR12_MHPMCOUNTER22H = 12'hb96;
localparam CSR12_MHPMCOUNTER23H = 12'hb97;
localparam CSR12_MHPMCOUNTER24H = 12'hb98;
localparam CSR12_MHPMCOUNTER25H = 12'hb99;
localparam CSR12_MHPMCOUNTER26H = 12'hb9a;
localparam CSR12_MHPMCOUNTER27H = 12'hb9b;
localparam CSR12_MHPMCOUNTER28H = 12'hb9c;
localparam CSR12_MHPMCOUNTER29H = 12'hb9d;
localparam CSR12_MHPMCOUNTER30H = 12'hb9e;
localparam CSR12_MHPMCOUNTER31H = 12'hb9f;
localparam CSR12_HPMEVENT3 = 12'h323;
localparam CSR12_HPMEVENT4 = 12'h324;
localparam CSR12_HPMEVENT5 = 12'h325;
localparam CSR12_HPMEVENT6 = 12'h326;
localparam CSR12_HPMEVENT7 = 12'h327;
localparam CSR12_HPMEVENT8 = 12'h328;
localparam CSR12_HPMEVENT9 = 12'h329;
localparam CSR12_HPMEVENT10 = 12'h32a;
localparam CSR12_HPMEVENT11 = 12'h32b;
localparam CSR12_HPMEVENT12 = 12'h32c;
localparam CSR12_HPMEVENT13 = 12'h32d;
localparam CSR12_HPMEVENT14 = 12'h32e;
localparam CSR12_HPMEVENT15 = 12'h32f;
localparam CSR12_HPMEVENT16 = 12'h330;
localparam CSR12_HPMEVENT17 = 12'h331;
localparam CSR12_HPMEVENT18 = 12'h332;
localparam CSR12_HPMEVENT19 = 12'h333;
localparam CSR12_HPMEVENT20 = 12'h334;
localparam CSR12_HPMEVENT21 = 12'h335;
localparam CSR12_HPMEVENT22 = 12'h336;
localparam CSR12_HPMEVENT23 = 12'h337;
localparam CSR12_HPMEVENT24 = 12'h338;
localparam CSR12_HPMEVENT25 = 12'h339;
localparam CSR12_HPMEVENT26 = 12'h33a;
localparam CSR12_HPMEVENT27 = 12'h33b;
localparam CSR12_HPMEVENT28 = 12'h33c;
localparam CSR12_HPMEVENT29 = 12'h33d;
localparam CSR12_HPMEVENT30 = 12'h33e;
localparam CSR12_HPMEVENT31 = 12'h33f;
localparam CSR12_PMPCFG0 = 12'h3a0;
localparam CSR12_PMPCFG1 = 12'h3a1;
localparam CSR12_PMPCFG2 = 12'h3a2;
localparam CSR12_PMPCFG3 = 12'h3a3;
localparam CSR12_PMPCFG4 = 12'h3a4;
localparam CSR12_PMPCFG5 = 12'h3a5;
localparam CSR12_PMPCFG6 = 12'h3a6;
localparam CSR12_PMPCFG7 = 12'h3a7;
localparam CSR12_PMPCFG8 = 12'h3a8;
localparam CSR12_PMPCFG9 = 12'h3a9;
localparam CSR12_PMPCFG10 = 12'h3aa;
localparam CSR12_PMPCFG11 = 12'h3ab;
localparam CSR12_PMPCFG12 = 12'h3ac;
localparam CSR12_PMPCFG13 = 12'h3ad;
localparam CSR12_PMPCFG14 = 12'h3ae;
localparam CSR12_PMPCFG15 = 12'h3af;
wire s6 = ((csr_addr == CSR12_PMPCFG0)) | (csr_addr == CSR12_PMPCFG1) | (csr_addr == CSR12_PMPCFG2) | (csr_addr == CSR12_PMPCFG3) | (csr_addr == CSR12_PMPCFG4) | (csr_addr == CSR12_PMPCFG5) | (csr_addr == CSR12_PMPCFG6) | (csr_addr == CSR12_PMPCFG7) | (csr_addr == CSR12_PMPCFG8) | (csr_addr == CSR12_PMPCFG9) | (csr_addr == CSR12_PMPCFG10) | (csr_addr == CSR12_PMPCFG11) | (csr_addr == CSR12_PMPCFG12) | (csr_addr == CSR12_PMPCFG13) | (csr_addr == CSR12_PMPCFG14) | (csr_addr == CSR12_PMPCFG15);
localparam CSR12_PMPADDR0 = 12'h3b0;
localparam CSR12_PMPADDR1 = 12'h3b1;
localparam CSR12_PMPADDR2 = 12'h3b2;
localparam CSR12_PMPADDR3 = 12'h3b3;
localparam CSR12_PMPADDR4 = 12'h3b4;
localparam CSR12_PMPADDR5 = 12'h3b5;
localparam CSR12_PMPADDR6 = 12'h3b6;
localparam CSR12_PMPADDR7 = 12'h3b7;
localparam CSR12_PMPADDR8 = 12'h3b8;
localparam CSR12_PMPADDR9 = 12'h3b9;
localparam CSR12_PMPADDR10 = 12'h3ba;
localparam CSR12_PMPADDR11 = 12'h3bb;
localparam CSR12_PMPADDR12 = 12'h3bc;
localparam CSR12_PMPADDR13 = 12'h3bd;
localparam CSR12_PMPADDR14 = 12'h3be;
localparam CSR12_PMPADDR15 = 12'h3bf;
localparam CSR12_PMPADDR16 = 12'h3c0;
localparam CSR12_PMPADDR17 = 12'h3c1;
localparam CSR12_PMPADDR18 = 12'h3c2;
localparam CSR12_PMPADDR19 = 12'h3c3;
localparam CSR12_PMPADDR20 = 12'h3c4;
localparam CSR12_PMPADDR21 = 12'h3c5;
localparam CSR12_PMPADDR22 = 12'h3c6;
localparam CSR12_PMPADDR23 = 12'h3c7;
localparam CSR12_PMPADDR24 = 12'h3c8;
localparam CSR12_PMPADDR25 = 12'h3c9;
localparam CSR12_PMPADDR26 = 12'h3ca;
localparam CSR12_PMPADDR27 = 12'h3cb;
localparam CSR12_PMPADDR28 = 12'h3cc;
localparam CSR12_PMPADDR29 = 12'h3cd;
localparam CSR12_PMPADDR30 = 12'h3ce;
localparam CSR12_PMPADDR31 = 12'h3cf;
localparam CSR12_PMPADDR32 = 12'h3d0;
localparam CSR12_PMPADDR33 = 12'h3d1;
localparam CSR12_PMPADDR34 = 12'h3d2;
localparam CSR12_PMPADDR35 = 12'h3d3;
localparam CSR12_PMPADDR36 = 12'h3d4;
localparam CSR12_PMPADDR37 = 12'h3d5;
localparam CSR12_PMPADDR38 = 12'h3d6;
localparam CSR12_PMPADDR39 = 12'h3d7;
localparam CSR12_PMPADDR40 = 12'h3d8;
localparam CSR12_PMPADDR41 = 12'h3d9;
localparam CSR12_PMPADDR42 = 12'h3da;
localparam CSR12_PMPADDR43 = 12'h3db;
localparam CSR12_PMPADDR44 = 12'h3dc;
localparam CSR12_PMPADDR45 = 12'h3dd;
localparam CSR12_PMPADDR46 = 12'h3de;
localparam CSR12_PMPADDR47 = 12'h3df;
localparam CSR12_PMPADDR48 = 12'h3e0;
localparam CSR12_PMPADDR49 = 12'h3e1;
localparam CSR12_PMPADDR50 = 12'h3e2;
localparam CSR12_PMPADDR51 = 12'h3e3;
localparam CSR12_PMPADDR52 = 12'h3e4;
localparam CSR12_PMPADDR53 = 12'h3e5;
localparam CSR12_PMPADDR54 = 12'h3e6;
localparam CSR12_PMPADDR55 = 12'h3e7;
localparam CSR12_PMPADDR56 = 12'h3e8;
localparam CSR12_PMPADDR57 = 12'h3e9;
localparam CSR12_PMPADDR58 = 12'h3ea;
localparam CSR12_PMPADDR59 = 12'h3eb;
localparam CSR12_PMPADDR60 = 12'h3ec;
localparam CSR12_PMPADDR61 = 12'h3ed;
localparam CSR12_PMPADDR62 = 12'h3ee;
localparam CSR12_PMPADDR63 = 12'h3ef;
wire s7 = ((csr_addr == CSR12_PMPADDR0)) | (csr_addr == CSR12_PMPADDR1) | (csr_addr == CSR12_PMPADDR2) | (csr_addr == CSR12_PMPADDR3) | (csr_addr == CSR12_PMPADDR4) | (csr_addr == CSR12_PMPADDR5) | (csr_addr == CSR12_PMPADDR6) | (csr_addr == CSR12_PMPADDR7) | (csr_addr == CSR12_PMPADDR8) | (csr_addr == CSR12_PMPADDR9) | (csr_addr == CSR12_PMPADDR10) | (csr_addr == CSR12_PMPADDR11) | (csr_addr == CSR12_PMPADDR12) | (csr_addr == CSR12_PMPADDR13) | (csr_addr == CSR12_PMPADDR14) | (csr_addr == CSR12_PMPADDR15) | (csr_addr == CSR12_PMPADDR16) | (csr_addr == CSR12_PMPADDR17) | (csr_addr == CSR12_PMPADDR18) | (csr_addr == CSR12_PMPADDR19) | (csr_addr == CSR12_PMPADDR20) | (csr_addr == CSR12_PMPADDR21) | (csr_addr == CSR12_PMPADDR22) | (csr_addr == CSR12_PMPADDR23) | (csr_addr == CSR12_PMPADDR24) | (csr_addr == CSR12_PMPADDR25) | (csr_addr == CSR12_PMPADDR26) | (csr_addr == CSR12_PMPADDR27) | (csr_addr == CSR12_PMPADDR28) | (csr_addr == CSR12_PMPADDR29) | (csr_addr == CSR12_PMPADDR30) | (csr_addr == CSR12_PMPADDR31) | (csr_addr == CSR12_PMPADDR32) | (csr_addr == CSR12_PMPADDR33) | (csr_addr == CSR12_PMPADDR34) | (csr_addr == CSR12_PMPADDR35) | (csr_addr == CSR12_PMPADDR36) | (csr_addr == CSR12_PMPADDR37) | (csr_addr == CSR12_PMPADDR38) | (csr_addr == CSR12_PMPADDR39) | (csr_addr == CSR12_PMPADDR40) | (csr_addr == CSR12_PMPADDR41) | (csr_addr == CSR12_PMPADDR42) | (csr_addr == CSR12_PMPADDR43) | (csr_addr == CSR12_PMPADDR44) | (csr_addr == CSR12_PMPADDR45) | (csr_addr == CSR12_PMPADDR46) | (csr_addr == CSR12_PMPADDR47) | (csr_addr == CSR12_PMPADDR48) | (csr_addr == CSR12_PMPADDR49) | (csr_addr == CSR12_PMPADDR50) | (csr_addr == CSR12_PMPADDR51) | (csr_addr == CSR12_PMPADDR52) | (csr_addr == CSR12_PMPADDR53) | (csr_addr == CSR12_PMPADDR54) | (csr_addr == CSR12_PMPADDR55) | (csr_addr == CSR12_PMPADDR56) | (csr_addr == CSR12_PMPADDR57) | (csr_addr == CSR12_PMPADDR58) | (csr_addr == CSR12_PMPADDR59) | (csr_addr == CSR12_PMPADDR60) | (csr_addr == CSR12_PMPADDR61) | (csr_addr == CSR12_PMPADDR62) | (csr_addr == CSR12_PMPADDR63);
localparam CSR12_PMACFG0 = 12'hbc0;
localparam CSR12_PMACFG1 = 12'hbc1;
localparam CSR12_PMACFG2 = 12'hbc2;
localparam CSR12_PMACFG3 = 12'hbc3;
localparam CSR12_PMAADDR0 = 12'hbd0;
localparam CSR12_PMAADDR1 = 12'hbd1;
localparam CSR12_PMAADDR2 = 12'hbd2;
localparam CSR12_PMAADDR3 = 12'hbd3;
localparam CSR12_PMAADDR4 = 12'hbd4;
localparam CSR12_PMAADDR5 = 12'hbd5;
localparam CSR12_PMAADDR6 = 12'hbd6;
localparam CSR12_PMAADDR7 = 12'hbd7;
localparam CSR12_PMAADDR8 = 12'hbd8;
localparam CSR12_PMAADDR9 = 12'hbd9;
localparam CSR12_PMAADDR10 = 12'hbda;
localparam CSR12_PMAADDR11 = 12'hbdb;
localparam CSR12_PMAADDR12 = 12'hbdc;
localparam CSR12_PMAADDR13 = 12'hbdd;
localparam CSR12_PMAADDR14 = 12'hbde;
localparam CSR12_PMAADDR15 = 12'hbdf;
localparam CSR12_TSELECT = 12'h7a0;
localparam CSR12_TDATA1 = 12'h7a1;
localparam CSR12_TDATA2 = 12'h7a2;
localparam CSR12_TDATA3 = 12'h7a3;
localparam CSR12_TINFO = 12'h7a4;
localparam CSR12_TCONTROL = 12'h7a5;
localparam CSR12_MCONTEXT = 12'h7a8;
localparam CSR12_SCONTEXT = 12'h7aa;
localparam CSR12_DCSR = 12'h7b0;
localparam CSR12_DPC = 12'h7b1;
localparam CSR12_DSCRATCH0 = 12'h7b2;
localparam CSR12_DSCRATCH1 = 12'h7b3;
localparam CSR12_MICM_CFG = 12'hfc0;
localparam CSR12_MDCM_CFG = 12'hfc1;
localparam CSR12_MMSC_CFG = 12'hfc2;
localparam CSR12_MMSC_CFG2 = 12'hfc3;
localparam CSR12_MMISC_CTL = 12'h7d0;
localparam CSR12_MCLK_CTL = 12'h7df;
localparam CSR12_MILMB = 12'h7c0;
localparam CSR12_MDLMB = 12'h7c1;
localparam CSR12_MECC_CODE = 12'h7c2;
localparam CSR12_MNVEC = 12'h7c3;
localparam CSR12_MXSTATUS = 12'h7c4;
localparam CSR12_MPFT_CTL = 12'h7c5;
localparam CSR12_MHSP_CTL = 12'h7c6;
localparam CSR12_MHSP_BOUND = 12'h7c7;
localparam CSR12_MHSP_BASE = 12'h7c8;
localparam CSR12_MDCAUSE = 12'h7c9;
localparam CSR12_MCACHE_CTL = 12'h7ca;
localparam CSR12_MCCTLBEGINADDR = 12'h7cb;
localparam CSR12_MCCTLCOMMAND = 12'h7cc;
localparam CSR12_MCCTLDATA = 12'h7cd;
localparam CSR12_MCOUNTERWEN = 12'h7ce;
localparam CSR12_MCOUNTERINTEN = 12'h7cf;
localparam CSR12_MCOUNTERMASK_M = 12'h7d1;
localparam CSR12_MCOUNTERMASK_S = 12'h7d2;
localparam CSR12_MCOUNTERMASK_U = 12'h7d3;
localparam CSR12_MCOUNTEROVF = 12'h7d4;
localparam CSR12_MSLIDELEG = 12'h7d5;
localparam CSR12_DEXC2DBG = 12'h7e0;
localparam CSR12_DDCAUSE = 12'h7e1;
localparam CSR12_MRANDSEQ = 12'h7fc;
localparam CSR12_MRANDSEQH = 12'h7fd;
localparam CSR12_MRANDSTATE = 12'h7fe;
localparam CSR12_MRANDSTATEH = 12'h7ff;
localparam CSR12_UITB = 12'h800;
localparam CSR12_UCODE = 12'h801;
localparam CSR12_UDCAUSE = 12'h809;
localparam CSR12_UCCTLBEGINADDR = 12'h80b;
localparam CSR12_UCCTLCOMMAND = 12'h80c;
localparam CSR12_SCOUNTERINTEN = 12'h9cf;
localparam CSR12_SCOUNTERMASK_M = 12'h9d1;
localparam CSR12_SCOUNTERMASK_S = 12'h9d2;
localparam CSR12_SCOUNTERMASK_U = 12'h9d3;
localparam CSR12_SCOUNTEROVF = 12'h9d4;
localparam CSR12_SCCTLDATA = 12'h9cd;
localparam CSR12_SMISC_CTL = 12'h9d0;
localparam CSR12_SCOUNTINHIBIT = 12'h9e0;
localparam CSR12_SHPMEVENT3 = 12'h9e3;
localparam CSR12_SHPMEVENT4 = 12'h9e4;
localparam CSR12_SHPMEVENT5 = 12'h9e5;
localparam CSR12_SHPMEVENT6 = 12'h9e6;
localparam CSR12_USTATUS = 12'h000;
localparam CSR12_UIE = 12'h004;
localparam CSR12_UTVEC = 12'h005;
localparam CSR12_USCRATCH = 12'h040;
localparam CSR12_UEPC = 12'h041;
localparam CSR12_UCAUSE = 12'h042;
localparam CSR12_UTVAL = 12'h043;
localparam CSR12_UIP = 12'h044;
localparam CSR12_CYCLE = 12'hc00;
localparam CSR12_TIME = 12'hc01;
localparam CSR12_INSTRET = 12'hc02;
localparam CSR12_HPMCOUNTER3 = 12'hc03;
localparam CSR12_HPMCOUNTER4 = 12'hc04;
localparam CSR12_HPMCOUNTER5 = 12'hc05;
localparam CSR12_HPMCOUNTER6 = 12'hc06;
localparam CSR12_HPMCOUNTER7 = 12'hc07;
localparam CSR12_HPMCOUNTER8 = 12'hc08;
localparam CSR12_HPMCOUNTER9 = 12'hc09;
localparam CSR12_HPMCOUNTER10 = 12'hc0a;
localparam CSR12_HPMCOUNTER11 = 12'hc0b;
localparam CSR12_HPMCOUNTER12 = 12'hc0c;
localparam CSR12_HPMCOUNTER13 = 12'hc0d;
localparam CSR12_HPMCOUNTER14 = 12'hc0e;
localparam CSR12_HPMCOUNTER15 = 12'hc0f;
localparam CSR12_HPMCOUNTER16 = 12'hc10;
localparam CSR12_HPMCOUNTER17 = 12'hc11;
localparam CSR12_HPMCOUNTER18 = 12'hc12;
localparam CSR12_HPMCOUNTER19 = 12'hc13;
localparam CSR12_HPMCOUNTER20 = 12'hc14;
localparam CSR12_HPMCOUNTER21 = 12'hc15;
localparam CSR12_HPMCOUNTER22 = 12'hc16;
localparam CSR12_HPMCOUNTER23 = 12'hc17;
localparam CSR12_HPMCOUNTER24 = 12'hc18;
localparam CSR12_HPMCOUNTER25 = 12'hc19;
localparam CSR12_HPMCOUNTER26 = 12'hc1a;
localparam CSR12_HPMCOUNTER27 = 12'hc1b;
localparam CSR12_HPMCOUNTER28 = 12'hc1c;
localparam CSR12_HPMCOUNTER29 = 12'hc1d;
localparam CSR12_HPMCOUNTER30 = 12'hc1e;
localparam CSR12_HPMCOUNTER31 = 12'hc1f;
localparam CSR12_CYCLEH = 12'hc80;
localparam CSR12_TIMEH = 12'hc81;
localparam CSR12_INSTRETH = 12'hc82;
localparam CSR12_HPMCOUNTER3H = 12'hc83;
localparam CSR12_HPMCOUNTER4H = 12'hc84;
localparam CSR12_HPMCOUNTER5H = 12'hc85;
localparam CSR12_HPMCOUNTER6H = 12'hc86;
localparam CSR12_HPMCOUNTER7H = 12'hc87;
localparam CSR12_HPMCOUNTER8H = 12'hc88;
localparam CSR12_HPMCOUNTER9H = 12'hc89;
localparam CSR12_HPMCOUNTER10H = 12'hc8a;
localparam CSR12_HPMCOUNTER11H = 12'hc8b;
localparam CSR12_HPMCOUNTER12H = 12'hc8c;
localparam CSR12_HPMCOUNTER13H = 12'hc8d;
localparam CSR12_HPMCOUNTER14H = 12'hc8e;
localparam CSR12_HPMCOUNTER15H = 12'hc8f;
localparam CSR12_HPMCOUNTER16H = 12'hc90;
localparam CSR12_HPMCOUNTER17H = 12'hc91;
localparam CSR12_HPMCOUNTER18H = 12'hc92;
localparam CSR12_HPMCOUNTER19H = 12'hc93;
localparam CSR12_HPMCOUNTER20H = 12'hc94;
localparam CSR12_HPMCOUNTER21H = 12'hc95;
localparam CSR12_HPMCOUNTER22H = 12'hc96;
localparam CSR12_HPMCOUNTER23H = 12'hc97;
localparam CSR12_HPMCOUNTER24H = 12'hc98;
localparam CSR12_HPMCOUNTER25H = 12'hc99;
localparam CSR12_HPMCOUNTER26H = 12'hc9a;
localparam CSR12_HPMCOUNTER27H = 12'hc9b;
localparam CSR12_HPMCOUNTER28H = 12'hc9c;
localparam CSR12_HPMCOUNTER29H = 12'hc9d;
localparam CSR12_HPMCOUNTER30H = 12'hc9e;
localparam CSR12_HPMCOUNTER31H = 12'hc9f;
assign existent_csr = (csr_addr == CSR12_MVENDORID) | (csr_addr == CSR12_MARCHID) | (csr_addr == CSR12_MIMPID) | (csr_addr == CSR12_MHARTID) | (csr_addr == CSR12_MSTATUS) | (csr_addr == CSR12_MISA) | (csr_addr == CSR12_MIE) | ((csr_addr == CSR12_MEDELEG) & (s0 | (s1 & ((RVN_SUPPORT_INT == 1))))) | ((csr_addr == CSR12_MIDELEG) & (s0 | (s1 & ((RVN_SUPPORT_INT == 1))))) | ((csr_addr == CSR12_MSLIDELEG) & s0) | (csr_addr == CSR12_MTVEC) | ((csr_addr == CSR12_MCOUNTEREN) & s2) | (csr_addr == CSR12_MCOUNTINHIBIT) | (csr_addr == CSR12_MSCRATCH) | (csr_addr == CSR12_MEPC) | (csr_addr == CSR12_MCAUSE) | (csr_addr == CSR12_MTVAL) | (csr_addr == CSR12_MIP) | (csr_addr == CSR12_MCYCLE) | (csr_addr == CSR12_MINSTRET) | ((csr_addr == CSR12_MCOUNTERWEN) & (PERFORMANCE_MONITOR_INT == 1) & s2) | ((csr_addr == CSR12_MCOUNTERINTEN) & (PERFORMANCE_MONITOR_INT == 1)) | ((csr_addr == CSR12_MCOUNTERMASK_M) & (PERFORMANCE_MONITOR_INT == 1) & s2) | ((csr_addr == CSR12_MCOUNTERMASK_S) & (PERFORMANCE_MONITOR_INT == 1) & s0) | ((csr_addr == CSR12_MCOUNTERMASK_U) & (PERFORMANCE_MONITOR_INT == 1) & s2) | ((csr_addr == CSR12_MCOUNTEROVF) & (PERFORMANCE_MONITOR_INT == 1)) | (csr_addr == CSR12_MHPMCOUNTER3) | (csr_addr == CSR12_MHPMCOUNTER4) | (csr_addr == CSR12_MHPMCOUNTER5) | (csr_addr == CSR12_MHPMCOUNTER6) | (csr_addr == CSR12_MHPMCOUNTER7) | (csr_addr == CSR12_MHPMCOUNTER8) | (csr_addr == CSR12_MHPMCOUNTER9) | (csr_addr == CSR12_MHPMCOUNTER10) | (csr_addr == CSR12_MHPMCOUNTER11) | (csr_addr == CSR12_MHPMCOUNTER12) | (csr_addr == CSR12_MHPMCOUNTER13) | (csr_addr == CSR12_MHPMCOUNTER14) | (csr_addr == CSR12_MHPMCOUNTER15) | (csr_addr == CSR12_MHPMCOUNTER16) | (csr_addr == CSR12_MHPMCOUNTER17) | (csr_addr == CSR12_MHPMCOUNTER18) | (csr_addr == CSR12_MHPMCOUNTER19) | (csr_addr == CSR12_MHPMCOUNTER20) | (csr_addr == CSR12_MHPMCOUNTER21) | (csr_addr == CSR12_MHPMCOUNTER22) | (csr_addr == CSR12_MHPMCOUNTER23) | (csr_addr == CSR12_MHPMCOUNTER24) | (csr_addr == CSR12_MHPMCOUNTER25) | (csr_addr == CSR12_MHPMCOUNTER26) | (csr_addr == CSR12_MHPMCOUNTER27) | (csr_addr == CSR12_MHPMCOUNTER28) | (csr_addr == CSR12_MHPMCOUNTER29) | (csr_addr == CSR12_MHPMCOUNTER30) | (csr_addr == CSR12_MHPMCOUNTER31) | (csr_addr == CSR12_MCYCLEH) | (csr_addr == CSR12_MINSTRETH) | (csr_addr == CSR12_MHPMCOUNTER3H) | (csr_addr == CSR12_MHPMCOUNTER4H) | (csr_addr == CSR12_MHPMCOUNTER5H) | (csr_addr == CSR12_MHPMCOUNTER6H) | (csr_addr == CSR12_MHPMCOUNTER7H) | (csr_addr == CSR12_MHPMCOUNTER8H) | (csr_addr == CSR12_MHPMCOUNTER9H) | (csr_addr == CSR12_MHPMCOUNTER10H) | (csr_addr == CSR12_MHPMCOUNTER11H) | (csr_addr == CSR12_MHPMCOUNTER12H) | (csr_addr == CSR12_MHPMCOUNTER13H) | (csr_addr == CSR12_MHPMCOUNTER14H) | (csr_addr == CSR12_MHPMCOUNTER15H) | (csr_addr == CSR12_MHPMCOUNTER16H) | (csr_addr == CSR12_MHPMCOUNTER17H) | (csr_addr == CSR12_MHPMCOUNTER18H) | (csr_addr == CSR12_MHPMCOUNTER19H) | (csr_addr == CSR12_MHPMCOUNTER20H) | (csr_addr == CSR12_MHPMCOUNTER21H) | (csr_addr == CSR12_MHPMCOUNTER22H) | (csr_addr == CSR12_MHPMCOUNTER23H) | (csr_addr == CSR12_MHPMCOUNTER24H) | (csr_addr == CSR12_MHPMCOUNTER25H) | (csr_addr == CSR12_MHPMCOUNTER26H) | (csr_addr == CSR12_MHPMCOUNTER27H) | (csr_addr == CSR12_MHPMCOUNTER28H) | (csr_addr == CSR12_MHPMCOUNTER29H) | (csr_addr == CSR12_MHPMCOUNTER30H) | (csr_addr == CSR12_MHPMCOUNTER31H) | (csr_addr == CSR12_HPMEVENT3) | (csr_addr == CSR12_HPMEVENT4) | (csr_addr == CSR12_HPMEVENT5) | (csr_addr == CSR12_HPMEVENT6) | (csr_addr == CSR12_HPMEVENT7) | (csr_addr == CSR12_HPMEVENT8) | (csr_addr == CSR12_HPMEVENT9) | (csr_addr == CSR12_HPMEVENT10) | (csr_addr == CSR12_HPMEVENT11) | (csr_addr == CSR12_HPMEVENT12) | (csr_addr == CSR12_HPMEVENT13) | (csr_addr == CSR12_HPMEVENT14) | (csr_addr == CSR12_HPMEVENT15) | (csr_addr == CSR12_HPMEVENT16) | (csr_addr == CSR12_HPMEVENT17) | (csr_addr == CSR12_HPMEVENT18) | (csr_addr == CSR12_HPMEVENT19) | (csr_addr == CSR12_HPMEVENT20) | (csr_addr == CSR12_HPMEVENT21) | (csr_addr == CSR12_HPMEVENT22) | (csr_addr == CSR12_HPMEVENT23) | (csr_addr == CSR12_HPMEVENT24) | (csr_addr == CSR12_HPMEVENT25) | (csr_addr == CSR12_HPMEVENT26) | (csr_addr == CSR12_HPMEVENT27) | (csr_addr == CSR12_HPMEVENT28) | (csr_addr == CSR12_HPMEVENT29) | (csr_addr == CSR12_HPMEVENT30) | (csr_addr == CSR12_HPMEVENT31) | s6 | s7 | (csr_addr == CSR12_PMACFG0) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMACFG1) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMACFG2) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMACFG3) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR0) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR1) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR2) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR3) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR4) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR5) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR6) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR7) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR8) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR9) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR10) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR11) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR12) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR13) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR14) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_PMAADDR15) & (PMA_ENTRIES != 0) | (csr_addr == CSR12_TSELECT) | (csr_addr == CSR12_TDATA1) | (csr_addr == CSR12_TDATA2) | (csr_addr == CSR12_TDATA3) | (csr_addr == CSR12_TINFO) | (csr_addr == CSR12_TCONTROL) | (csr_addr == CSR12_MCONTEXT) | (csr_addr == CSR12_SCONTEXT) | (csr_addr == CSR12_DCSR) | (csr_addr == CSR12_DPC) | (csr_addr == CSR12_DSCRATCH0) | (csr_addr == CSR12_DSCRATCH1) | (csr_addr == CSR12_MICM_CFG) | (csr_addr == CSR12_MDCM_CFG) | (csr_addr == CSR12_MMSC_CFG) | ((csr_addr == CSR12_MMSC_CFG2) & ((MMSC_CFG2_EXIST_INT == 1))) | ((csr_addr == CSR12_MMISC_CTL) & ((MMISC_CTL_EXIST_INT == 1))) | ((csr_addr == CSR12_MILMB) & (ILM_SIZE_KB != 0)) | ((csr_addr == CSR12_MDLMB) & (DLM_SIZE_KB != 0)) | ((csr_addr == CSR12_MECC_CODE) & ((ECC_SUPPORT_INT == 1) | ((ICACHE_ECC_TYPE_INT != 0)))) | (csr_addr == CSR12_MNVEC) | ((csr_addr == CSR12_MXSTATUS)) | ((csr_addr == CSR12_MPFT_CTL) & ((POWERBRAKE_SUPPORT_INT == 1))) | (csr_addr == CSR12_MDCAUSE) | ((csr_addr == CSR12_MCACHE_CTL) & (CACHE_SUPPORT_INT == 1)) | ((csr_addr == CSR12_MCCTLBEGINADDR) & (CACHE_SUPPORT_INT == 1)) | ((csr_addr == CSR12_MCCTLCOMMAND) & (CACHE_SUPPORT_INT == 1)) | ((csr_addr == CSR12_MCCTLDATA) & (CACHE_SUPPORT_INT == 1)) | (csr_addr == CSR12_DEXC2DBG) | (csr_addr == CSR12_DDCAUSE) | (csr_addr == CSR12_MHSP_CTL) & ((STACKSAFE_SUPPORT_INT == 1)) | (csr_addr == CSR12_MHSP_BOUND) & ((STACKSAFE_SUPPORT_INT == 1)) | (csr_addr == CSR12_MHSP_BASE) & ((STACKSAFE_SUPPORT_INT == 1)) | (csr_addr == CSR12_UITB) | (csr_addr == CSR12_UCODE) & ((DSP_SUPPORT_INT == 1)) | (csr_addr == CSR12_FFLAGS) & (FLEN != 1) | (csr_addr == CSR12_FRM) & (FLEN != 1) | (csr_addr == CSR12_FCSR) & (FLEN != 1) | (csr_addr == CSR12_MCLK_CTL) & ((FLEN != 1)) | ((csr_addr == CSR12_CYCLE) & s2) | ((csr_addr == CSR12_INSTRET) & s2) | ((csr_addr == CSR12_HPMCOUNTER3) & s2) | ((csr_addr == CSR12_HPMCOUNTER4) & s2) | ((csr_addr == CSR12_HPMCOUNTER5) & s2) | ((csr_addr == CSR12_HPMCOUNTER6) & s2) | ((csr_addr == CSR12_HPMCOUNTER7) & s2) | ((csr_addr == CSR12_HPMCOUNTER8) & s2) | ((csr_addr == CSR12_HPMCOUNTER9) & s2) | ((csr_addr == CSR12_HPMCOUNTER10) & s2) | ((csr_addr == CSR12_HPMCOUNTER11) & s2) | ((csr_addr == CSR12_HPMCOUNTER12) & s2) | ((csr_addr == CSR12_HPMCOUNTER13) & s2) | ((csr_addr == CSR12_HPMCOUNTER14) & s2) | ((csr_addr == CSR12_HPMCOUNTER15) & s2) | ((csr_addr == CSR12_HPMCOUNTER16) & s2) | ((csr_addr == CSR12_HPMCOUNTER17) & s2) | ((csr_addr == CSR12_HPMCOUNTER18) & s2) | ((csr_addr == CSR12_HPMCOUNTER19) & s2) | ((csr_addr == CSR12_HPMCOUNTER20) & s2) | ((csr_addr == CSR12_HPMCOUNTER21) & s2) | ((csr_addr == CSR12_HPMCOUNTER22) & s2) | ((csr_addr == CSR12_HPMCOUNTER23) & s2) | ((csr_addr == CSR12_HPMCOUNTER24) & s2) | ((csr_addr == CSR12_HPMCOUNTER25) & s2) | ((csr_addr == CSR12_HPMCOUNTER26) & s2) | ((csr_addr == CSR12_HPMCOUNTER27) & s2) | ((csr_addr == CSR12_HPMCOUNTER28) & s2) | ((csr_addr == CSR12_HPMCOUNTER29) & s2) | ((csr_addr == CSR12_HPMCOUNTER30) & s2) | ((csr_addr == CSR12_HPMCOUNTER31) & s2) | (csr_addr == CSR12_CYCLEH) & s2 | (csr_addr == CSR12_INSTRETH) & s2 | (csr_addr == CSR12_HPMCOUNTER3H) & s2 | (csr_addr == CSR12_HPMCOUNTER4H) & s2 | (csr_addr == CSR12_HPMCOUNTER5H) & s2 | (csr_addr == CSR12_HPMCOUNTER6H) & s2 | (csr_addr == CSR12_HPMCOUNTER7H) & s2 | (csr_addr == CSR12_HPMCOUNTER8H) & s2 | (csr_addr == CSR12_HPMCOUNTER9H) & s2 | (csr_addr == CSR12_HPMCOUNTER10H) & s2 | (csr_addr == CSR12_HPMCOUNTER11H) & s2 | (csr_addr == CSR12_HPMCOUNTER12H) & s2 | (csr_addr == CSR12_HPMCOUNTER13H) & s2 | (csr_addr == CSR12_HPMCOUNTER14H) & s2 | (csr_addr == CSR12_HPMCOUNTER15H) & s2 | (csr_addr == CSR12_HPMCOUNTER16H) & s2 | (csr_addr == CSR12_HPMCOUNTER17H) & s2 | (csr_addr == CSR12_HPMCOUNTER18H) & s2 | (csr_addr == CSR12_HPMCOUNTER19H) & s2 | (csr_addr == CSR12_HPMCOUNTER20H) & s2 | (csr_addr == CSR12_HPMCOUNTER21H) & s2 | (csr_addr == CSR12_HPMCOUNTER22H) & s2 | (csr_addr == CSR12_HPMCOUNTER23H) & s2 | (csr_addr == CSR12_HPMCOUNTER24H) & s2 | (csr_addr == CSR12_HPMCOUNTER25H) & s2 | (csr_addr == CSR12_HPMCOUNTER26H) & s2 | (csr_addr == CSR12_HPMCOUNTER27H) & s2 | (csr_addr == CSR12_HPMCOUNTER28H) & s2 | (csr_addr == CSR12_HPMCOUNTER29H) & s2 | (csr_addr == CSR12_HPMCOUNTER30H) & s2 | (csr_addr == CSR12_HPMCOUNTER31H) & s2 | ((csr_addr == CSR12_SSTATUS) & s0) | ((csr_addr == CSR12_SIE) & s0) | ((csr_addr == CSR12_SLIE) & s0) | ((csr_addr == CSR12_SIP) & s0) | ((csr_addr == CSR12_SLIP) & s0) | ((csr_addr == CSR12_SIDELEG) & s0 & ((RVN_SUPPORT_INT == 1))) | ((csr_addr == CSR12_SEDELEG) & s0 & ((RVN_SUPPORT_INT == 1))) | ((csr_addr == CSR12_STVEC) & s0) | ((csr_addr == CSR12_SEPC) & s0) | ((csr_addr == CSR12_SCAUSE) & s0) | ((csr_addr == CSR12_SDCAUSE) & s0) | ((csr_addr == CSR12_STVAL) & s0) | ((csr_addr == CSR12_SSCRATCH) & s0) | ((csr_addr == CSR12_SATP) & s0) | ((csr_addr == CSR12_SCOUNTEREN) & s0) | ((csr_addr == CSR12_SMISC_CTL) & s0 & ((ACE_SUPPORT_INT == 1))) | ((csr_addr == CSR12_SCOUNTERINTEN) & s0 & (PERFORMANCE_MONITOR_INT == 1)) | ((csr_addr == CSR12_SCOUNTERMASK_M) & s0 & (PERFORMANCE_MONITOR_INT == 1)) | ((csr_addr == CSR12_SCOUNTERMASK_S) & s0 & (PERFORMANCE_MONITOR_INT == 1)) | ((csr_addr == CSR12_SCOUNTERMASK_U) & s0 & (PERFORMANCE_MONITOR_INT == 1)) | ((csr_addr == CSR12_SCOUNTEROVF) & s0 & (PERFORMANCE_MONITOR_INT == 1)) | ((csr_addr == CSR12_SCOUNTINHIBIT) & s0 & (PERFORMANCE_MONITOR_INT == 1)) | ((csr_addr == CSR12_SHPMEVENT3) & s0 & (PERFORMANCE_MONITOR_INT == 1)) | ((csr_addr == CSR12_SHPMEVENT4) & s0 & (PERFORMANCE_MONITOR_INT == 1)) | ((csr_addr == CSR12_SHPMEVENT5) & s0 & (PERFORMANCE_MONITOR_INT == 1)) | ((csr_addr == CSR12_SHPMEVENT6) & s0 & (PERFORMANCE_MONITOR_INT == 1)) | ((csr_addr == CSR12_SCCTLDATA) & s0 & (CACHE_SUPPORT_INT == 1)) | ((csr_addr == CSR12_UCCTLCOMMAND) & s2 & (CACHE_SUPPORT_INT == 1)) | ((csr_addr == CSR12_UCCTLBEGINADDR) & s2 & (CACHE_SUPPORT_INT == 1)) | ((csr_addr == CSR12_USTATUS) & s2 & ((RVN_SUPPORT_INT == 1))) | ((csr_addr == CSR12_UIE) & s2 & ((RVN_SUPPORT_INT == 1))) | ((csr_addr == CSR12_UTVEC) & s2 & ((RVN_SUPPORT_INT == 1))) | ((csr_addr == CSR12_USCRATCH) & s2 & ((RVN_SUPPORT_INT == 1))) | ((csr_addr == CSR12_UEPC) & s2 & ((RVN_SUPPORT_INT == 1))) | ((csr_addr == CSR12_UCAUSE) & s2 & ((RVN_SUPPORT_INT == 1))) | ((csr_addr == CSR12_UTVAL) & s2 & ((RVN_SUPPORT_INT == 1))) | ((csr_addr == CSR12_UIP) & s2 & ((RVN_SUPPORT_INT == 1))) | ((csr_addr == CSR12_UDCAUSE) & s2 & ((RVN_SUPPORT_INT == 1)));
wire s8 = csr_mcounteren[0];
wire s9 = csr_mcounteren[1];
wire s10 = csr_mcounteren[2];
wire s11 = csr_mcounteren[3];
wire s12 = csr_mcounteren[4];
wire s13 = csr_mcounteren[5];
wire s14 = csr_mcounteren[6];
wire s15 = csr_mcounterwen[0];
wire s16 = csr_mcounterwen[1];
wire s17 = csr_mcounterwen[2];
wire s18 = csr_mcounterwen[3];
wire s19 = csr_mcounterwen[4];
wire s20 = csr_mcounterwen[5];
wire s21 = csr_mcounterwen[6];
wire s22 = csr_scounteren[0];
wire s23 = csr_scounteren[1];
wire s24 = csr_scounteren[2];
wire s25 = csr_scounteren[3];
wire s26 = csr_scounteren[4];
wire s27 = csr_scounteren[5];
wire s28 = csr_scounteren[6];
wire s29 = ~(s8 | writeonly_csr);
wire s30 = s1 & cur_privilege_u & s29;
wire s31 = s0 & ((s3 & s29) | (cur_privilege_u & ~s22));
wire s32 = s30 | s31;
wire s33 = ~(s9 | writeonly_csr);
wire s34 = s1 & cur_privilege_u & s33;
wire s35 = s0 & ((s3 & s33) | (cur_privilege_u & ~s23));
wire s36 = s34 | s35;
wire s37 = ~(s10 | writeonly_csr);
wire s38 = s1 & cur_privilege_u & s37;
wire s39 = s0 & ((s3 & s37) | (cur_privilege_u & ~s24));
wire s40 = s38 | s39;
wire s41 = ~(s11 | writeonly_csr);
wire s42 = s1 & cur_privilege_u & s41;
wire s43 = s0 & ((s3 & s41) | (cur_privilege_u & ~s25));
wire s44 = s42 | s43;
wire s45 = ~(s12 | writeonly_csr);
wire s46 = s1 & cur_privilege_u & s45;
wire s47 = s0 & ((s3 & s45) | (cur_privilege_u & ~s26));
wire s48 = s46 | s47;
wire s49 = ~(s13 | writeonly_csr);
wire s50 = s1 & cur_privilege_u & s49;
wire s51 = s0 & ((s3 & s49) | (cur_privilege_u & ~s27));
wire s52 = s50 | s51;
wire s53 = ~(s14 | writeonly_csr);
wire s54 = s1 & cur_privilege_u & s53;
wire s55 = s0 & ((s3 & s53) | (cur_privilege_u & ~s28));
wire s56 = s54 | s55;
assign s5 = ((csr_addr == CSR12_DCSR) & ~csr_halt_mode) | ((csr_addr == CSR12_DPC) & ~csr_halt_mode) | ((csr_addr == CSR12_DSCRATCH0) & ~csr_halt_mode) | ((csr_addr == CSR12_DSCRATCH1) & ~csr_halt_mode) | ((csr_addr == CSR12_DEXC2DBG) & ~csr_halt_mode) | ((csr_addr == CSR12_DDCAUSE) & ~csr_halt_mode) | ((csr_addr == CSR12_SCCTLDATA) & (~cur_privilege_m & ~csr_mcache_ctl_cctl_suen)) | ((csr_addr == CSR12_UCCTLCOMMAND) & ((~cur_privilege_m & ~csr_mcache_ctl_cctl_suen) | csr_ucctlcommand_privileged)) | ((csr_addr == CSR12_UCCTLBEGINADDR) & (~cur_privilege_m & ~csr_mcache_ctl_cctl_suen)) | (~(csr_addr == CSR12_SCONTEXT) & (csr_cur_privilege < csr_addr[9:8]) & s2 & ~csr_halt_mode) | ((csr_addr == CSR12_SCONTEXT) & cur_privilege_u & ~csr_halt_mode) | (((csr_addr == CSR12_HPMCOUNTER7) | (csr_addr == CSR12_HPMCOUNTER7H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER8) | (csr_addr == CSR12_HPMCOUNTER8H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER9) | (csr_addr == CSR12_HPMCOUNTER9H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER10) | (csr_addr == CSR12_HPMCOUNTER10H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER11) | (csr_addr == CSR12_HPMCOUNTER11H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER12) | (csr_addr == CSR12_HPMCOUNTER12H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER13) | (csr_addr == CSR12_HPMCOUNTER13H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER14) | (csr_addr == CSR12_HPMCOUNTER14H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER15) | (csr_addr == CSR12_HPMCOUNTER15H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER16) | (csr_addr == CSR12_HPMCOUNTER16H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER17) | (csr_addr == CSR12_HPMCOUNTER17H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER18) | (csr_addr == CSR12_HPMCOUNTER18H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER19) | (csr_addr == CSR12_HPMCOUNTER19H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER20) | (csr_addr == CSR12_HPMCOUNTER20H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER21) | (csr_addr == CSR12_HPMCOUNTER21H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER22) | (csr_addr == CSR12_HPMCOUNTER22H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER23) | (csr_addr == CSR12_HPMCOUNTER23H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER24) | (csr_addr == CSR12_HPMCOUNTER24H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER25) | (csr_addr == CSR12_HPMCOUNTER25H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER26) | (csr_addr == CSR12_HPMCOUNTER26H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER27) | (csr_addr == CSR12_HPMCOUNTER27H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER28) | (csr_addr == CSR12_HPMCOUNTER28H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER29) | (csr_addr == CSR12_HPMCOUNTER29H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER30) | (csr_addr == CSR12_HPMCOUNTER30H)) & (cur_privilege_s | cur_privilege_u)) | (((csr_addr == CSR12_HPMCOUNTER31) | (csr_addr == CSR12_HPMCOUNTER31H)) & (cur_privilege_s | cur_privilege_u)) | ((csr_addr == CSR12_SATP) & cur_privilege_s & csr_mstatus_tvm);
assign privileged_csr_ddcause = s5 | (((csr_addr == CSR12_CYCLE) | (csr_addr == CSR12_CYCLEH)) & s32 & ~writeonly_csr & ~csr_halt_mode) | (((csr_addr == CSR12_TIME) | (csr_addr == CSR12_TIMEH)) & s36 & ~writeonly_csr & ~csr_halt_mode) | (((csr_addr == CSR12_INSTRET) | (csr_addr == CSR12_INSTRETH)) & s40 & ~writeonly_csr & ~csr_halt_mode) | (((csr_addr == CSR12_HPMCOUNTER3) | (csr_addr == CSR12_HPMCOUNTER3H) | (csr_addr == CSR12_SHPMEVENT3)) & s44 & ~writeonly_csr & ~csr_halt_mode) | (((csr_addr == CSR12_HPMCOUNTER4) | (csr_addr == CSR12_HPMCOUNTER4H) | (csr_addr == CSR12_SHPMEVENT4)) & s48 & ~writeonly_csr & ~csr_halt_mode) | (((csr_addr == CSR12_HPMCOUNTER5) | (csr_addr == CSR12_HPMCOUNTER5H) | (csr_addr == CSR12_SHPMEVENT5)) & s52 & ~writeonly_csr & ~csr_halt_mode) | (((csr_addr == CSR12_HPMCOUNTER6) | (csr_addr == CSR12_HPMCOUNTER6H) | (csr_addr == CSR12_SHPMEVENT6)) & s56 & ~writeonly_csr & ~csr_halt_mode);
assign privileged_csr = s5 | (((csr_addr == CSR12_CYCLE) | (csr_addr == CSR12_CYCLEH)) & s32 & ~csr_halt_mode) | (((csr_addr == CSR12_TIME) | (csr_addr == CSR12_TIMEH)) & s36 & ~csr_halt_mode) | (((csr_addr == CSR12_INSTRET) | (csr_addr == CSR12_INSTRETH)) & s40 & ~csr_halt_mode) | (((csr_addr == CSR12_HPMCOUNTER3) | (csr_addr == CSR12_HPMCOUNTER3H) | (csr_addr == CSR12_SHPMEVENT3)) & s44 & ~csr_halt_mode) | (((csr_addr == CSR12_HPMCOUNTER4) | (csr_addr == CSR12_HPMCOUNTER4H) | (csr_addr == CSR12_SHPMEVENT4)) & s48 & ~csr_halt_mode) | (((csr_addr == CSR12_HPMCOUNTER5) | (csr_addr == CSR12_HPMCOUNTER5H) | (csr_addr == CSR12_SHPMEVENT5)) & s52 & ~csr_halt_mode) | (((csr_addr == CSR12_HPMCOUNTER6) | (csr_addr == CSR12_HPMCOUNTER6H) | (csr_addr == CSR12_SHPMEVENT6)) & s56 & ~csr_halt_mode);
wire s57 = (csr_addr == CSR12_CYCLE) | (csr_addr == CSR12_CYCLEH);
wire s58 = (csr_addr == CSR12_TIME) | (csr_addr == CSR12_TIMEH);
wire s59 = (csr_addr == CSR12_INSTRET) | (csr_addr == CSR12_INSTRETH);
wire s60 = (csr_addr == CSR12_HPMCOUNTER3) | (csr_addr == CSR12_HPMCOUNTER3H) | (csr_addr == CSR12_SHPMEVENT3);
wire s61 = (csr_addr == CSR12_HPMCOUNTER4) | (csr_addr == CSR12_HPMCOUNTER4H) | (csr_addr == CSR12_SHPMEVENT4);
wire s62 = (csr_addr == CSR12_HPMCOUNTER5) | (csr_addr == CSR12_HPMCOUNTER5H) | (csr_addr == CSR12_SHPMEVENT5);
wire s63 = (csr_addr == CSR12_HPMCOUNTER6) | (csr_addr == CSR12_HPMCOUNTER6H) | (csr_addr == CSR12_SHPMEVENT6);
wire s64 = s57 | s58 | s59 | s60 | s61 | s62 | s63;
wire s65 = s15 & (s1 | s4);
wire s66 = s16 & (s1 | s4);
wire s67 = s17 & (s1 | s4);
wire s68 = s18 & (s1 | s4);
wire s69 = s19 & (s1 | s4);
wire s70 = s20 & (s1 | s4);
wire s71 = s21 & (s1 | s4);
assign readonly_csr = (~s64 & (csr_addr[11:10] == 2'b11)) | (s57 & ~s65) | (s58 & ~s66) | (s59 & ~s67) | (s60 & ~s68) | (s61 & ~s69) | (s62 & ~s70) | (s63 & ~s71);
wire [1:0] nds_unused_func_csr = func_csr;
wire [4:0] nds_unused_rd_index = rd_index;
endmodule

