-------------------------------------------------------------------------------
--
-- A testbench model for the
-- GCpad controller core
--
-- Copyright (c) 2004, Arnim Laeuger (arniml@opencores.org)
--
-- $Id: gcpad_mod-c.vhd,v 1.1 2004-10-10 17:26:28 arniml Exp $
--
-------------------------------------------------------------------------------

configuration gcpad_mod_behav_c0 of gcpad_mod is

  for behav
  end for;

end gcpad_mod_behav_c0;
