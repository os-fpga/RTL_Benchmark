library ieee;
use ieee.std_logic_1164.all;

entity top is
	port( a: in std_logic_vector(127 downto 0);
	shift: in std_logic_vector(6 downto 0);
	result: out std_logic_vector(127 downto 0));
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335: std_logic;

begin

w0 <= a(77) and shift(0);
w1 <= shift(1) and w0;
w2 <= a(78) and not shift(0);
w3 <= shift(1) and w2;
w4 <= not w1 and not w3;
w5 <= a(80) and not shift(0);
w6 <= not shift(1) and w5;
w7 <= a(79) and shift(0);
w8 <= not shift(1) and w7;
w9 <= not w6 and not w8;
w10 <= w4 and w9;
w11 <= not shift(2) and not shift(3);
w12 <= not w10 and w11;
w13 <= a(73) and shift(0);
w14 <= shift(1) and w13;
w15 <= a(74) and not shift(0);
w16 <= shift(1) and w15;
w17 <= not w14 and not w16;
w18 <= a(76) and not shift(0);
w19 <= not shift(1) and w18;
w20 <= a(75) and shift(0);
w21 <= not shift(1) and w20;
w22 <= not w19 and not w21;
w23 <= w17 and w22;
w24 <= shift(2) and not shift(3);
w25 <= not w23 and w24;
w26 <= not w12 and not w25;
w27 <= a(65) and shift(0);
w28 <= shift(1) and w27;
w29 <= a(66) and not shift(0);
w30 <= shift(1) and w29;
w31 <= not w28 and not w30;
w32 <= a(68) and not shift(0);
w33 <= not shift(1) and w32;
w34 <= a(67) and shift(0);
w35 <= not shift(1) and w34;
w36 <= not w33 and not w35;
w37 <= w31 and w36;
w38 <= shift(2) and shift(3);
w39 <= not w37 and w38;
w40 <= a(69) and shift(0);
w41 <= shift(1) and w40;
w42 <= a(70) and not shift(0);
w43 <= shift(1) and w42;
w44 <= not w41 and not w43;
w45 <= a(72) and not shift(0);
w46 <= not shift(1) and w45;
w47 <= a(71) and shift(0);
w48 <= not shift(1) and w47;
w49 <= not w46 and not w48;
w50 <= w44 and w49;
w51 <= not shift(2) and shift(3);
w52 <= not w50 and w51;
w53 <= not w39 and not w52;
w54 <= w26 and w53;
w55 <= shift(4) and shift(5);
w56 <= not w54 and w55;
w57 <= a(93) and shift(0);
w58 <= shift(1) and w57;
w59 <= a(94) and not shift(0);
w60 <= shift(1) and w59;
w61 <= not w58 and not w60;
w62 <= a(96) and not shift(0);
w63 <= not shift(1) and w62;
w64 <= a(95) and shift(0);
w65 <= not shift(1) and w64;
w66 <= not w63 and not w65;
w67 <= w61 and w66;
w68 <= w11 and not w67;
w69 <= a(89) and shift(0);
w70 <= shift(1) and w69;
w71 <= a(90) and not shift(0);
w72 <= shift(1) and w71;
w73 <= not w70 and not w72;
w74 <= a(92) and not shift(0);
w75 <= not shift(1) and w74;
w76 <= a(91) and shift(0);
w77 <= not shift(1) and w76;
w78 <= not w75 and not w77;
w79 <= w73 and w78;
w80 <= w24 and not w79;
w81 <= not w68 and not w80;
w82 <= a(81) and shift(0);
w83 <= shift(1) and w82;
w84 <= a(82) and not shift(0);
w85 <= shift(1) and w84;
w86 <= not w83 and not w85;
w87 <= a(84) and not shift(0);
w88 <= not shift(1) and w87;
w89 <= a(83) and shift(0);
w90 <= not shift(1) and w89;
w91 <= not w88 and not w90;
w92 <= w86 and w91;
w93 <= w38 and not w92;
w94 <= a(85) and shift(0);
w95 <= shift(1) and w94;
w96 <= a(86) and not shift(0);
w97 <= shift(1) and w96;
w98 <= not w95 and not w97;
w99 <= a(88) and not shift(0);
w100 <= not shift(1) and w99;
w101 <= a(87) and shift(0);
w102 <= not shift(1) and w101;
w103 <= not w100 and not w102;
w104 <= w98 and w103;
w105 <= w51 and not w104;
w106 <= not w93 and not w105;
w107 <= w81 and w106;
w108 <= not shift(4) and shift(5);
w109 <= not w107 and w108;
w110 <= not w56 and not w109;
w111 <= a(125) and shift(0);
w112 <= shift(1) and w111;
w113 <= a(126) and not shift(0);
w114 <= shift(1) and w113;
w115 <= not w112 and not w114;
w116 <= a(0) and not shift(0);
w117 <= not shift(1) and w116;
w118 <= a(127) and shift(0);
w119 <= not shift(1) and w118;
w120 <= not w117 and not w119;
w121 <= w115 and w120;
w122 <= w11 and not w121;
w123 <= a(121) and shift(0);
w124 <= shift(1) and w123;
w125 <= a(122) and not shift(0);
w126 <= shift(1) and w125;
w127 <= not w124 and not w126;
w128 <= a(124) and not shift(0);
w129 <= not shift(1) and w128;
w130 <= a(123) and shift(0);
w131 <= not shift(1) and w130;
w132 <= not w129 and not w131;
w133 <= w127 and w132;
w134 <= w24 and not w133;
w135 <= not w122 and not w134;
w136 <= a(113) and shift(0);
w137 <= shift(1) and w136;
w138 <= a(114) and not shift(0);
w139 <= shift(1) and w138;
w140 <= not w137 and not w139;
w141 <= a(116) and not shift(0);
w142 <= not shift(1) and w141;
w143 <= a(115) and shift(0);
w144 <= not shift(1) and w143;
w145 <= not w142 and not w144;
w146 <= w140 and w145;
w147 <= w38 and not w146;
w148 <= a(117) and shift(0);
w149 <= shift(1) and w148;
w150 <= a(118) and not shift(0);
w151 <= shift(1) and w150;
w152 <= not w149 and not w151;
w153 <= a(120) and not shift(0);
w154 <= not shift(1) and w153;
w155 <= a(119) and shift(0);
w156 <= not shift(1) and w155;
w157 <= not w154 and not w156;
w158 <= w152 and w157;
w159 <= w51 and not w158;
w160 <= not w147 and not w159;
w161 <= w135 and w160;
w162 <= not shift(4) and not shift(5);
w163 <= not w161 and w162;
w164 <= a(109) and shift(0);
w165 <= shift(1) and w164;
w166 <= a(110) and not shift(0);
w167 <= shift(1) and w166;
w168 <= not w165 and not w167;
w169 <= a(112) and not shift(0);
w170 <= not shift(1) and w169;
w171 <= a(111) and shift(0);
w172 <= not shift(1) and w171;
w173 <= not w170 and not w172;
w174 <= w168 and w173;
w175 <= w11 and not w174;
w176 <= a(105) and shift(0);
w177 <= shift(1) and w176;
w178 <= a(106) and not shift(0);
w179 <= shift(1) and w178;
w180 <= not w177 and not w179;
w181 <= a(108) and not shift(0);
w182 <= not shift(1) and w181;
w183 <= a(107) and shift(0);
w184 <= not shift(1) and w183;
w185 <= not w182 and not w184;
w186 <= w180 and w185;
w187 <= w24 and not w186;
w188 <= not w175 and not w187;
w189 <= a(97) and shift(0);
w190 <= shift(1) and w189;
w191 <= a(98) and not shift(0);
w192 <= shift(1) and w191;
w193 <= not w190 and not w192;
w194 <= a(100) and not shift(0);
w195 <= not shift(1) and w194;
w196 <= a(99) and shift(0);
w197 <= not shift(1) and w196;
w198 <= not w195 and not w197;
w199 <= w193 and w198;
w200 <= w38 and not w199;
w201 <= a(101) and shift(0);
w202 <= shift(1) and w201;
w203 <= a(102) and not shift(0);
w204 <= shift(1) and w203;
w205 <= not w202 and not w204;
w206 <= a(104) and not shift(0);
w207 <= not shift(1) and w206;
w208 <= a(103) and shift(0);
w209 <= not shift(1) and w208;
w210 <= not w207 and not w209;
w211 <= w205 and w210;
w212 <= w51 and not w211;
w213 <= not w200 and not w212;
w214 <= w188 and w213;
w215 <= shift(4) and not shift(5);
w216 <= not w214 and w215;
w217 <= not w163 and not w216;
w218 <= w110 and w217;
w219 <= not shift(6) and not w218;
w220 <= a(13) and shift(0);
w221 <= shift(1) and w220;
w222 <= a(14) and not shift(0);
w223 <= shift(1) and w222;
w224 <= not w221 and not w223;
w225 <= a(16) and not shift(0);
w226 <= not shift(1) and w225;
w227 <= a(15) and shift(0);
w228 <= not shift(1) and w227;
w229 <= not w226 and not w228;
w230 <= w224 and w229;
w231 <= w11 and not w230;
w232 <= a(9) and shift(0);
w233 <= shift(1) and w232;
w234 <= a(10) and not shift(0);
w235 <= shift(1) and w234;
w236 <= not w233 and not w235;
w237 <= a(12) and not shift(0);
w238 <= not shift(1) and w237;
w239 <= a(11) and shift(0);
w240 <= not shift(1) and w239;
w241 <= not w238 and not w240;
w242 <= w236 and w241;
w243 <= w24 and not w242;
w244 <= not w231 and not w243;
w245 <= a(1) and shift(0);
w246 <= shift(1) and w245;
w247 <= a(2) and not shift(0);
w248 <= shift(1) and w247;
w249 <= not w246 and not w248;
w250 <= a(4) and not shift(0);
w251 <= not shift(1) and w250;
w252 <= a(3) and shift(0);
w253 <= not shift(1) and w252;
w254 <= not w251 and not w253;
w255 <= w249 and w254;
w256 <= w38 and not w255;
w257 <= a(5) and shift(0);
w258 <= shift(1) and w257;
w259 <= a(6) and not shift(0);
w260 <= shift(1) and w259;
w261 <= not w258 and not w260;
w262 <= a(8) and not shift(0);
w263 <= not shift(1) and w262;
w264 <= a(7) and shift(0);
w265 <= not shift(1) and w264;
w266 <= not w263 and not w265;
w267 <= w261 and w266;
w268 <= w51 and not w267;
w269 <= not w256 and not w268;
w270 <= w244 and w269;
w271 <= w55 and not w270;
w272 <= a(29) and shift(0);
w273 <= shift(1) and w272;
w274 <= a(30) and not shift(0);
w275 <= shift(1) and w274;
w276 <= not w273 and not w275;
w277 <= a(32) and not shift(0);
w278 <= not shift(1) and w277;
w279 <= a(31) and shift(0);
w280 <= not shift(1) and w279;
w281 <= not w278 and not w280;
w282 <= w276 and w281;
w283 <= w11 and not w282;
w284 <= a(25) and shift(0);
w285 <= shift(1) and w284;
w286 <= a(26) and not shift(0);
w287 <= shift(1) and w286;
w288 <= not w285 and not w287;
w289 <= a(28) and not shift(0);
w290 <= not shift(1) and w289;
w291 <= a(27) and shift(0);
w292 <= not shift(1) and w291;
w293 <= not w290 and not w292;
w294 <= w288 and w293;
w295 <= w24 and not w294;
w296 <= not w283 and not w295;
w297 <= a(17) and shift(0);
w298 <= shift(1) and w297;
w299 <= a(18) and not shift(0);
w300 <= shift(1) and w299;
w301 <= not w298 and not w300;
w302 <= a(20) and not shift(0);
w303 <= not shift(1) and w302;
w304 <= a(19) and shift(0);
w305 <= not shift(1) and w304;
w306 <= not w303 and not w305;
w307 <= w301 and w306;
w308 <= w38 and not w307;
w309 <= a(21) and shift(0);
w310 <= shift(1) and w309;
w311 <= a(22) and not shift(0);
w312 <= shift(1) and w311;
w313 <= not w310 and not w312;
w314 <= a(24) and not shift(0);
w315 <= not shift(1) and w314;
w316 <= a(23) and shift(0);
w317 <= not shift(1) and w316;
w318 <= not w315 and not w317;
w319 <= w313 and w318;
w320 <= w51 and not w319;
w321 <= not w308 and not w320;
w322 <= w296 and w321;
w323 <= w108 and not w322;
w324 <= not w271 and not w323;
w325 <= a(61) and shift(0);
w326 <= shift(1) and w325;
w327 <= a(62) and not shift(0);
w328 <= shift(1) and w327;
w329 <= not w326 and not w328;
w330 <= a(64) and not shift(0);
w331 <= not shift(1) and w330;
w332 <= a(63) and shift(0);
w333 <= not shift(1) and w332;
w334 <= not w331 and not w333;
w335 <= w329 and w334;
w336 <= w11 and not w335;
w337 <= a(57) and shift(0);
w338 <= shift(1) and w337;
w339 <= a(58) and not shift(0);
w340 <= shift(1) and w339;
w341 <= not w338 and not w340;
w342 <= a(60) and not shift(0);
w343 <= not shift(1) and w342;
w344 <= a(59) and shift(0);
w345 <= not shift(1) and w344;
w346 <= not w343 and not w345;
w347 <= w341 and w346;
w348 <= w24 and not w347;
w349 <= not w336 and not w348;
w350 <= a(49) and shift(0);
w351 <= shift(1) and w350;
w352 <= a(50) and not shift(0);
w353 <= shift(1) and w352;
w354 <= not w351 and not w353;
w355 <= a(52) and not shift(0);
w356 <= not shift(1) and w355;
w357 <= a(51) and shift(0);
w358 <= not shift(1) and w357;
w359 <= not w356 and not w358;
w360 <= w354 and w359;
w361 <= w38 and not w360;
w362 <= a(53) and shift(0);
w363 <= shift(1) and w362;
w364 <= a(54) and not shift(0);
w365 <= shift(1) and w364;
w366 <= not w363 and not w365;
w367 <= a(56) and not shift(0);
w368 <= not shift(1) and w367;
w369 <= a(55) and shift(0);
w370 <= not shift(1) and w369;
w371 <= not w368 and not w370;
w372 <= w366 and w371;
w373 <= w51 and not w372;
w374 <= not w361 and not w373;
w375 <= w349 and w374;
w376 <= w162 and not w375;
w377 <= a(45) and shift(0);
w378 <= shift(1) and w377;
w379 <= a(46) and not shift(0);
w380 <= shift(1) and w379;
w381 <= not w378 and not w380;
w382 <= a(48) and not shift(0);
w383 <= not shift(1) and w382;
w384 <= a(47) and shift(0);
w385 <= not shift(1) and w384;
w386 <= not w383 and not w385;
w387 <= w381 and w386;
w388 <= w11 and not w387;
w389 <= a(41) and shift(0);
w390 <= shift(1) and w389;
w391 <= a(42) and not shift(0);
w392 <= shift(1) and w391;
w393 <= not w390 and not w392;
w394 <= a(44) and not shift(0);
w395 <= not shift(1) and w394;
w396 <= a(43) and shift(0);
w397 <= not shift(1) and w396;
w398 <= not w395 and not w397;
w399 <= w393 and w398;
w400 <= w24 and not w399;
w401 <= not w388 and not w400;
w402 <= a(33) and shift(0);
w403 <= shift(1) and w402;
w404 <= a(34) and not shift(0);
w405 <= shift(1) and w404;
w406 <= not w403 and not w405;
w407 <= a(36) and not shift(0);
w408 <= not shift(1) and w407;
w409 <= a(35) and shift(0);
w410 <= not shift(1) and w409;
w411 <= not w408 and not w410;
w412 <= w406 and w411;
w413 <= w38 and not w412;
w414 <= a(40) and not shift(0);
w415 <= not shift(1) and w414;
w416 <= a(37) and shift(0);
w417 <= shift(1) and w416;
w418 <= not w415 and not w417;
w419 <= a(39) and shift(0);
w420 <= not shift(1) and w419;
w421 <= a(38) and not shift(0);
w422 <= shift(1) and w421;
w423 <= not w420 and not w422;
w424 <= w418 and w423;
w425 <= w51 and not w424;
w426 <= not w413 and not w425;
w427 <= w401 and w426;
w428 <= w215 and not w427;
w429 <= not w376 and not w428;
w430 <= w324 and w429;
w431 <= shift(6) and not w430;
w432 <= not w219 and not w431;
w433 <= a(81) and not shift(0);
w434 <= not shift(1) and w433;
w435 <= a(78) and shift(0);
w436 <= shift(1) and w435;
w437 <= not w434 and not w436;
w438 <= a(80) and shift(0);
w439 <= not shift(1) and w438;
w440 <= a(79) and not shift(0);
w441 <= shift(1) and w440;
w442 <= not w439 and not w441;
w443 <= w437 and w442;
w444 <= w11 and not w443;
w445 <= a(77) and not shift(0);
w446 <= not shift(1) and w445;
w447 <= a(74) and shift(0);
w448 <= shift(1) and w447;
w449 <= not w446 and not w448;
w450 <= a(76) and shift(0);
w451 <= not shift(1) and w450;
w452 <= a(75) and not shift(0);
w453 <= shift(1) and w452;
w454 <= not w451 and not w453;
w455 <= w449 and w454;
w456 <= w24 and not w455;
w457 <= not w444 and not w456;
w458 <= a(69) and not shift(0);
w459 <= not shift(1) and w458;
w460 <= a(66) and shift(0);
w461 <= shift(1) and w460;
w462 <= not w459 and not w461;
w463 <= a(68) and shift(0);
w464 <= not shift(1) and w463;
w465 <= a(67) and not shift(0);
w466 <= shift(1) and w465;
w467 <= not w464 and not w466;
w468 <= w462 and w467;
w469 <= w38 and not w468;
w470 <= a(73) and not shift(0);
w471 <= not shift(1) and w470;
w472 <= a(70) and shift(0);
w473 <= shift(1) and w472;
w474 <= not w471 and not w473;
w475 <= a(72) and shift(0);
w476 <= not shift(1) and w475;
w477 <= a(71) and not shift(0);
w478 <= shift(1) and w477;
w479 <= not w476 and not w478;
w480 <= w474 and w479;
w481 <= w51 and not w480;
w482 <= not w469 and not w481;
w483 <= w457 and w482;
w484 <= w55 and not w483;
w485 <= a(97) and not shift(0);
w486 <= not shift(1) and w485;
w487 <= a(94) and shift(0);
w488 <= shift(1) and w487;
w489 <= not w486 and not w488;
w490 <= a(96) and shift(0);
w491 <= not shift(1) and w490;
w492 <= a(95) and not shift(0);
w493 <= shift(1) and w492;
w494 <= not w491 and not w493;
w495 <= w489 and w494;
w496 <= w11 and not w495;
w497 <= a(93) and not shift(0);
w498 <= not shift(1) and w497;
w499 <= a(90) and shift(0);
w500 <= shift(1) and w499;
w501 <= not w498 and not w500;
w502 <= a(92) and shift(0);
w503 <= not shift(1) and w502;
w504 <= a(91) and not shift(0);
w505 <= shift(1) and w504;
w506 <= not w503 and not w505;
w507 <= w501 and w506;
w508 <= w24 and not w507;
w509 <= not w496 and not w508;
w510 <= a(85) and not shift(0);
w511 <= not shift(1) and w510;
w512 <= a(82) and shift(0);
w513 <= shift(1) and w512;
w514 <= not w511 and not w513;
w515 <= a(84) and shift(0);
w516 <= not shift(1) and w515;
w517 <= a(83) and not shift(0);
w518 <= shift(1) and w517;
w519 <= not w516 and not w518;
w520 <= w514 and w519;
w521 <= w38 and not w520;
w522 <= a(89) and not shift(0);
w523 <= not shift(1) and w522;
w524 <= a(86) and shift(0);
w525 <= shift(1) and w524;
w526 <= not w523 and not w525;
w527 <= a(88) and shift(0);
w528 <= not shift(1) and w527;
w529 <= a(87) and not shift(0);
w530 <= shift(1) and w529;
w531 <= not w528 and not w530;
w532 <= w526 and w531;
w533 <= w51 and not w532;
w534 <= not w521 and not w533;
w535 <= w509 and w534;
w536 <= w108 and not w535;
w537 <= not w484 and not w536;
w538 <= a(1) and not shift(0);
w539 <= not shift(1) and w538;
w540 <= a(126) and shift(0);
w541 <= shift(1) and w540;
w542 <= not w539 and not w541;
w543 <= a(0) and shift(0);
w544 <= not shift(1) and w543;
w545 <= a(127) and not shift(0);
w546 <= shift(1) and w545;
w547 <= not w544 and not w546;
w548 <= w542 and w547;
w549 <= w11 and not w548;
w550 <= a(125) and not shift(0);
w551 <= not shift(1) and w550;
w552 <= a(122) and shift(0);
w553 <= shift(1) and w552;
w554 <= not w551 and not w553;
w555 <= a(124) and shift(0);
w556 <= not shift(1) and w555;
w557 <= a(123) and not shift(0);
w558 <= shift(1) and w557;
w559 <= not w556 and not w558;
w560 <= w554 and w559;
w561 <= w24 and not w560;
w562 <= not w549 and not w561;
w563 <= a(117) and not shift(0);
w564 <= not shift(1) and w563;
w565 <= a(114) and shift(0);
w566 <= shift(1) and w565;
w567 <= not w564 and not w566;
w568 <= a(116) and shift(0);
w569 <= not shift(1) and w568;
w570 <= a(115) and not shift(0);
w571 <= shift(1) and w570;
w572 <= not w569 and not w571;
w573 <= w567 and w572;
w574 <= w38 and not w573;
w575 <= a(121) and not shift(0);
w576 <= not shift(1) and w575;
w577 <= a(118) and shift(0);
w578 <= shift(1) and w577;
w579 <= not w576 and not w578;
w580 <= a(120) and shift(0);
w581 <= not shift(1) and w580;
w582 <= a(119) and not shift(0);
w583 <= shift(1) and w582;
w584 <= not w581 and not w583;
w585 <= w579 and w584;
w586 <= w51 and not w585;
w587 <= not w574 and not w586;
w588 <= w562 and w587;
w589 <= w162 and not w588;
w590 <= a(113) and not shift(0);
w591 <= not shift(1) and w590;
w592 <= a(110) and shift(0);
w593 <= shift(1) and w592;
w594 <= not w591 and not w593;
w595 <= a(112) and shift(0);
w596 <= not shift(1) and w595;
w597 <= a(111) and not shift(0);
w598 <= shift(1) and w597;
w599 <= not w596 and not w598;
w600 <= w594 and w599;
w601 <= w11 and not w600;
w602 <= a(109) and not shift(0);
w603 <= not shift(1) and w602;
w604 <= a(106) and shift(0);
w605 <= shift(1) and w604;
w606 <= not w603 and not w605;
w607 <= a(108) and shift(0);
w608 <= not shift(1) and w607;
w609 <= a(107) and not shift(0);
w610 <= shift(1) and w609;
w611 <= not w608 and not w610;
w612 <= w606 and w611;
w613 <= w24 and not w612;
w614 <= not w601 and not w613;
w615 <= a(101) and not shift(0);
w616 <= not shift(1) and w615;
w617 <= a(98) and shift(0);
w618 <= shift(1) and w617;
w619 <= not w616 and not w618;
w620 <= a(100) and shift(0);
w621 <= not shift(1) and w620;
w622 <= a(99) and not shift(0);
w623 <= shift(1) and w622;
w624 <= not w621 and not w623;
w625 <= w619 and w624;
w626 <= w38 and not w625;
w627 <= a(105) and not shift(0);
w628 <= not shift(1) and w627;
w629 <= a(102) and shift(0);
w630 <= shift(1) and w629;
w631 <= not w628 and not w630;
w632 <= a(104) and shift(0);
w633 <= not shift(1) and w632;
w634 <= a(103) and not shift(0);
w635 <= shift(1) and w634;
w636 <= not w633 and not w635;
w637 <= w631 and w636;
w638 <= w51 and not w637;
w639 <= not w626 and not w638;
w640 <= w614 and w639;
w641 <= w215 and not w640;
w642 <= not w589 and not w641;
w643 <= w537 and w642;
w644 <= not shift(6) and not w643;
w645 <= a(65) and not shift(0);
w646 <= not shift(1) and w645;
w647 <= a(62) and shift(0);
w648 <= shift(1) and w647;
w649 <= not w646 and not w648;
w650 <= a(64) and shift(0);
w651 <= not shift(1) and w650;
w652 <= a(63) and not shift(0);
w653 <= shift(1) and w652;
w654 <= not w651 and not w653;
w655 <= w649 and w654;
w656 <= w11 and not w655;
w657 <= a(61) and not shift(0);
w658 <= not shift(1) and w657;
w659 <= a(58) and shift(0);
w660 <= shift(1) and w659;
w661 <= not w658 and not w660;
w662 <= a(60) and shift(0);
w663 <= not shift(1) and w662;
w664 <= a(59) and not shift(0);
w665 <= shift(1) and w664;
w666 <= not w663 and not w665;
w667 <= w661 and w666;
w668 <= w24 and not w667;
w669 <= not w656 and not w668;
w670 <= a(53) and not shift(0);
w671 <= not shift(1) and w670;
w672 <= a(50) and shift(0);
w673 <= shift(1) and w672;
w674 <= not w671 and not w673;
w675 <= a(52) and shift(0);
w676 <= not shift(1) and w675;
w677 <= a(51) and not shift(0);
w678 <= shift(1) and w677;
w679 <= not w676 and not w678;
w680 <= w674 and w679;
w681 <= w38 and not w680;
w682 <= a(57) and not shift(0);
w683 <= not shift(1) and w682;
w684 <= a(54) and shift(0);
w685 <= shift(1) and w684;
w686 <= not w683 and not w685;
w687 <= a(56) and shift(0);
w688 <= not shift(1) and w687;
w689 <= a(55) and not shift(0);
w690 <= shift(1) and w689;
w691 <= not w688 and not w690;
w692 <= w686 and w691;
w693 <= w51 and not w692;
w694 <= not w681 and not w693;
w695 <= w669 and w694;
w696 <= w162 and not w695;
w697 <= a(17) and not shift(0);
w698 <= not shift(1) and w697;
w699 <= a(14) and shift(0);
w700 <= shift(1) and w699;
w701 <= not w698 and not w700;
w702 <= a(16) and shift(0);
w703 <= not shift(1) and w702;
w704 <= a(15) and not shift(0);
w705 <= shift(1) and w704;
w706 <= not w703 and not w705;
w707 <= w701 and w706;
w708 <= w11 and not w707;
w709 <= a(13) and not shift(0);
w710 <= not shift(1) and w709;
w711 <= a(10) and shift(0);
w712 <= shift(1) and w711;
w713 <= not w710 and not w712;
w714 <= a(12) and shift(0);
w715 <= not shift(1) and w714;
w716 <= a(11) and not shift(0);
w717 <= shift(1) and w716;
w718 <= not w715 and not w717;
w719 <= w713 and w718;
w720 <= w24 and not w719;
w721 <= not w708 and not w720;
w722 <= a(5) and not shift(0);
w723 <= not shift(1) and w722;
w724 <= a(2) and shift(0);
w725 <= shift(1) and w724;
w726 <= not w723 and not w725;
w727 <= a(4) and shift(0);
w728 <= not shift(1) and w727;
w729 <= a(3) and not shift(0);
w730 <= shift(1) and w729;
w731 <= not w728 and not w730;
w732 <= w726 and w731;
w733 <= w38 and not w732;
w734 <= a(9) and not shift(0);
w735 <= not shift(1) and w734;
w736 <= a(6) and shift(0);
w737 <= shift(1) and w736;
w738 <= not w735 and not w737;
w739 <= a(8) and shift(0);
w740 <= not shift(1) and w739;
w741 <= a(7) and not shift(0);
w742 <= shift(1) and w741;
w743 <= not w740 and not w742;
w744 <= w738 and w743;
w745 <= w51 and not w744;
w746 <= not w733 and not w745;
w747 <= w721 and w746;
w748 <= w55 and not w747;
w749 <= not w696 and not w748;
w750 <= a(49) and not shift(0);
w751 <= not shift(1) and w750;
w752 <= a(46) and shift(0);
w753 <= shift(1) and w752;
w754 <= not w751 and not w753;
w755 <= a(48) and shift(0);
w756 <= not shift(1) and w755;
w757 <= a(47) and not shift(0);
w758 <= shift(1) and w757;
w759 <= not w756 and not w758;
w760 <= w754 and w759;
w761 <= w11 and not w760;
w762 <= a(42) and shift(0);
w763 <= shift(1) and w762;
w764 <= a(43) and not shift(0);
w765 <= shift(1) and w764;
w766 <= not w763 and not w765;
w767 <= a(45) and not shift(0);
w768 <= not shift(1) and w767;
w769 <= a(44) and shift(0);
w770 <= not shift(1) and w769;
w771 <= not w768 and not w770;
w772 <= w766 and w771;
w773 <= w24 and not w772;
w774 <= not w761 and not w773;
w775 <= a(37) and not shift(0);
w776 <= not shift(1) and w775;
w777 <= a(34) and shift(0);
w778 <= shift(1) and w777;
w779 <= not w776 and not w778;
w780 <= a(36) and shift(0);
w781 <= not shift(1) and w780;
w782 <= a(35) and not shift(0);
w783 <= shift(1) and w782;
w784 <= not w781 and not w783;
w785 <= w779 and w784;
w786 <= w38 and not w785;
w787 <= a(41) and not shift(0);
w788 <= not shift(1) and w787;
w789 <= a(40) and shift(0);
w790 <= not shift(1) and w789;
w791 <= not w788 and not w790;
w792 <= a(39) and not shift(0);
w793 <= shift(1) and w792;
w794 <= a(38) and shift(0);
w795 <= shift(1) and w794;
w796 <= not w793 and not w795;
w797 <= w791 and w796;
w798 <= w51 and not w797;
w799 <= not w786 and not w798;
w800 <= w774 and w799;
w801 <= w215 and not w800;
w802 <= a(33) and not shift(0);
w803 <= not shift(1) and w802;
w804 <= a(30) and shift(0);
w805 <= shift(1) and w804;
w806 <= not w803 and not w805;
w807 <= a(32) and shift(0);
w808 <= not shift(1) and w807;
w809 <= a(31) and not shift(0);
w810 <= shift(1) and w809;
w811 <= not w808 and not w810;
w812 <= w806 and w811;
w813 <= w11 and not w812;
w814 <= a(29) and not shift(0);
w815 <= not shift(1) and w814;
w816 <= a(26) and shift(0);
w817 <= shift(1) and w816;
w818 <= not w815 and not w817;
w819 <= a(28) and shift(0);
w820 <= not shift(1) and w819;
w821 <= a(27) and not shift(0);
w822 <= shift(1) and w821;
w823 <= not w820 and not w822;
w824 <= w818 and w823;
w825 <= w24 and not w824;
w826 <= not w813 and not w825;
w827 <= a(21) and not shift(0);
w828 <= not shift(1) and w827;
w829 <= a(18) and shift(0);
w830 <= shift(1) and w829;
w831 <= not w828 and not w830;
w832 <= a(20) and shift(0);
w833 <= not shift(1) and w832;
w834 <= a(19) and not shift(0);
w835 <= shift(1) and w834;
w836 <= not w833 and not w835;
w837 <= w831 and w836;
w838 <= w38 and not w837;
w839 <= a(25) and not shift(0);
w840 <= not shift(1) and w839;
w841 <= a(22) and shift(0);
w842 <= shift(1) and w841;
w843 <= not w840 and not w842;
w844 <= a(24) and shift(0);
w845 <= not shift(1) and w844;
w846 <= a(23) and not shift(0);
w847 <= shift(1) and w846;
w848 <= not w845 and not w847;
w849 <= w843 and w848;
w850 <= w51 and not w849;
w851 <= not w838 and not w850;
w852 <= w826 and w851;
w853 <= w108 and not w852;
w854 <= not w801 and not w853;
w855 <= w749 and w854;
w856 <= shift(6) and not w855;
w857 <= not w644 and not w856;
w858 <= not shift(1) and w82;
w859 <= not shift(1) and w84;
w860 <= not w858 and not w859;
w861 <= shift(1) and w5;
w862 <= shift(1) and w7;
w863 <= not w861 and not w862;
w864 <= w860 and w863;
w865 <= w11 and not w864;
w866 <= not shift(1) and w0;
w867 <= not shift(1) and w2;
w868 <= not w866 and not w867;
w869 <= shift(1) and w18;
w870 <= shift(1) and w20;
w871 <= not w869 and not w870;
w872 <= w868 and w871;
w873 <= w24 and not w872;
w874 <= not w865 and not w873;
w875 <= not shift(1) and w40;
w876 <= not shift(1) and w42;
w877 <= not w875 and not w876;
w878 <= shift(1) and w32;
w879 <= shift(1) and w34;
w880 <= not w878 and not w879;
w881 <= w877 and w880;
w882 <= w38 and not w881;
w883 <= not shift(1) and w13;
w884 <= not shift(1) and w15;
w885 <= not w883 and not w884;
w886 <= shift(1) and w45;
w887 <= shift(1) and w47;
w888 <= not w886 and not w887;
w889 <= w885 and w888;
w890 <= w51 and not w889;
w891 <= not w882 and not w890;
w892 <= w874 and w891;
w893 <= w55 and not w892;
w894 <= not shift(1) and w189;
w895 <= not shift(1) and w191;
w896 <= not w894 and not w895;
w897 <= shift(1) and w62;
w898 <= shift(1) and w64;
w899 <= not w897 and not w898;
w900 <= w896 and w899;
w901 <= w11 and not w900;
w902 <= not shift(1) and w57;
w903 <= not shift(1) and w59;
w904 <= not w902 and not w903;
w905 <= shift(1) and w74;
w906 <= shift(1) and w76;
w907 <= not w905 and not w906;
w908 <= w904 and w907;
w909 <= w24 and not w908;
w910 <= not w901 and not w909;
w911 <= not shift(1) and w94;
w912 <= not shift(1) and w96;
w913 <= not w911 and not w912;
w914 <= shift(1) and w87;
w915 <= shift(1) and w89;
w916 <= not w914 and not w915;
w917 <= w913 and w916;
w918 <= w38 and not w917;
w919 <= not shift(1) and w69;
w920 <= not shift(1) and w71;
w921 <= not w919 and not w920;
w922 <= shift(1) and w99;
w923 <= shift(1) and w101;
w924 <= not w922 and not w923;
w925 <= w921 and w924;
w926 <= w51 and not w925;
w927 <= not w918 and not w926;
w928 <= w910 and w927;
w929 <= w108 and not w928;
w930 <= not w893 and not w929;
w931 <= not shift(1) and w245;
w932 <= not shift(1) and w247;
w933 <= not w931 and not w932;
w934 <= shift(1) and w116;
w935 <= shift(1) and w118;
w936 <= not w934 and not w935;
w937 <= w933 and w936;
w938 <= w11 and not w937;
w939 <= not shift(1) and w111;
w940 <= not shift(1) and w113;
w941 <= not w939 and not w940;
w942 <= shift(1) and w128;
w943 <= shift(1) and w130;
w944 <= not w942 and not w943;
w945 <= w941 and w944;
w946 <= w24 and not w945;
w947 <= not w938 and not w946;
w948 <= not shift(1) and w148;
w949 <= not shift(1) and w150;
w950 <= not w948 and not w949;
w951 <= shift(1) and w141;
w952 <= shift(1) and w143;
w953 <= not w951 and not w952;
w954 <= w950 and w953;
w955 <= w38 and not w954;
w956 <= not shift(1) and w123;
w957 <= not shift(1) and w125;
w958 <= not w956 and not w957;
w959 <= shift(1) and w153;
w960 <= shift(1) and w155;
w961 <= not w959 and not w960;
w962 <= w958 and w961;
w963 <= w51 and not w962;
w964 <= not w955 and not w963;
w965 <= w947 and w964;
w966 <= w162 and not w965;
w967 <= not shift(1) and w136;
w968 <= not shift(1) and w138;
w969 <= not w967 and not w968;
w970 <= shift(1) and w169;
w971 <= shift(1) and w171;
w972 <= not w970 and not w971;
w973 <= w969 and w972;
w974 <= w11 and not w973;
w975 <= not shift(1) and w164;
w976 <= not shift(1) and w166;
w977 <= not w975 and not w976;
w978 <= shift(1) and w181;
w979 <= shift(1) and w183;
w980 <= not w978 and not w979;
w981 <= w977 and w980;
w982 <= w24 and not w981;
w983 <= not w974 and not w982;
w984 <= not shift(1) and w201;
w985 <= not shift(1) and w203;
w986 <= not w984 and not w985;
w987 <= shift(1) and w194;
w988 <= shift(1) and w196;
w989 <= not w987 and not w988;
w990 <= w986 and w989;
w991 <= w38 and not w990;
w992 <= not shift(1) and w176;
w993 <= not shift(1) and w178;
w994 <= not w992 and not w993;
w995 <= shift(1) and w206;
w996 <= shift(1) and w208;
w997 <= not w995 and not w996;
w998 <= w994 and w997;
w999 <= w51 and not w998;
w1000 <= not w991 and not w999;
w1001 <= w983 and w1000;
w1002 <= w215 and not w1001;
w1003 <= not w966 and not w1002;
w1004 <= w930 and w1003;
w1005 <= not shift(6) and not w1004;
w1006 <= not shift(1) and w27;
w1007 <= not shift(1) and w29;
w1008 <= not w1006 and not w1007;
w1009 <= shift(1) and w330;
w1010 <= shift(1) and w332;
w1011 <= not w1009 and not w1010;
w1012 <= w1008 and w1011;
w1013 <= w11 and not w1012;
w1014 <= not shift(1) and w325;
w1015 <= not shift(1) and w327;
w1016 <= not w1014 and not w1015;
w1017 <= shift(1) and w342;
w1018 <= shift(1) and w344;
w1019 <= not w1017 and not w1018;
w1020 <= w1016 and w1019;
w1021 <= w24 and not w1020;
w1022 <= not w1013 and not w1021;
w1023 <= not shift(1) and w362;
w1024 <= not shift(1) and w364;
w1025 <= not w1023 and not w1024;
w1026 <= shift(1) and w355;
w1027 <= shift(1) and w357;
w1028 <= not w1026 and not w1027;
w1029 <= w1025 and w1028;
w1030 <= w38 and not w1029;
w1031 <= not shift(1) and w337;
w1032 <= not shift(1) and w339;
w1033 <= not w1031 and not w1032;
w1034 <= shift(1) and w367;
w1035 <= shift(1) and w369;
w1036 <= not w1034 and not w1035;
w1037 <= w1033 and w1036;
w1038 <= w51 and not w1037;
w1039 <= not w1030 and not w1038;
w1040 <= w1022 and w1039;
w1041 <= w162 and not w1040;
w1042 <= not shift(1) and w297;
w1043 <= not shift(1) and w299;
w1044 <= not w1042 and not w1043;
w1045 <= shift(1) and w225;
w1046 <= shift(1) and w227;
w1047 <= not w1045 and not w1046;
w1048 <= w1044 and w1047;
w1049 <= w11 and not w1048;
w1050 <= not shift(1) and w220;
w1051 <= not shift(1) and w222;
w1052 <= not w1050 and not w1051;
w1053 <= shift(1) and w237;
w1054 <= shift(1) and w239;
w1055 <= not w1053 and not w1054;
w1056 <= w1052 and w1055;
w1057 <= w24 and not w1056;
w1058 <= not w1049 and not w1057;
w1059 <= not shift(1) and w257;
w1060 <= not shift(1) and w259;
w1061 <= not w1059 and not w1060;
w1062 <= shift(1) and w250;
w1063 <= shift(1) and w252;
w1064 <= not w1062 and not w1063;
w1065 <= w1061 and w1064;
w1066 <= w38 and not w1065;
w1067 <= not shift(1) and w232;
w1068 <= not shift(1) and w234;
w1069 <= not w1067 and not w1068;
w1070 <= shift(1) and w262;
w1071 <= shift(1) and w264;
w1072 <= not w1070 and not w1071;
w1073 <= w1069 and w1072;
w1074 <= w51 and not w1073;
w1075 <= not w1066 and not w1074;
w1076 <= w1058 and w1075;
w1077 <= w55 and not w1076;
w1078 <= not w1041 and not w1077;
w1079 <= not shift(1) and w350;
w1080 <= not shift(1) and w352;
w1081 <= not w1079 and not w1080;
w1082 <= shift(1) and w382;
w1083 <= shift(1) and w384;
w1084 <= not w1082 and not w1083;
w1085 <= w1081 and w1084;
w1086 <= w11 and not w1085;
w1087 <= shift(1) and w396;
w1088 <= shift(1) and w394;
w1089 <= not w1087 and not w1088;
w1090 <= not shift(1) and w379;
w1091 <= not shift(1) and w377;
w1092 <= not w1090 and not w1091;
w1093 <= w1089 and w1092;
w1094 <= w24 and not w1093;
w1095 <= not w1086 and not w1094;
w1096 <= not shift(1) and w416;
w1097 <= not shift(1) and w421;
w1098 <= not w1096 and not w1097;
w1099 <= shift(1) and w407;
w1100 <= shift(1) and w409;
w1101 <= not w1099 and not w1100;
w1102 <= w1098 and w1101;
w1103 <= w38 and not w1102;
w1104 <= not shift(1) and w389;
w1105 <= not shift(1) and w391;
w1106 <= not w1104 and not w1105;
w1107 <= shift(1) and w419;
w1108 <= shift(1) and w414;
w1109 <= not w1107 and not w1108;
w1110 <= w1106 and w1109;
w1111 <= w51 and not w1110;
w1112 <= not w1103 and not w1111;
w1113 <= w1095 and w1112;
w1114 <= w215 and not w1113;
w1115 <= not shift(1) and w402;
w1116 <= not shift(1) and w404;
w1117 <= not w1115 and not w1116;
w1118 <= shift(1) and w277;
w1119 <= shift(1) and w279;
w1120 <= not w1118 and not w1119;
w1121 <= w1117 and w1120;
w1122 <= w11 and not w1121;
w1123 <= not shift(1) and w272;
w1124 <= not shift(1) and w274;
w1125 <= not w1123 and not w1124;
w1126 <= shift(1) and w289;
w1127 <= shift(1) and w291;
w1128 <= not w1126 and not w1127;
w1129 <= w1125 and w1128;
w1130 <= w24 and not w1129;
w1131 <= not w1122 and not w1130;
w1132 <= not shift(1) and w309;
w1133 <= not shift(1) and w311;
w1134 <= not w1132 and not w1133;
w1135 <= shift(1) and w302;
w1136 <= shift(1) and w304;
w1137 <= not w1135 and not w1136;
w1138 <= w1134 and w1137;
w1139 <= w38 and not w1138;
w1140 <= not shift(1) and w284;
w1141 <= not shift(1) and w286;
w1142 <= not w1140 and not w1141;
w1143 <= shift(1) and w314;
w1144 <= shift(1) and w316;
w1145 <= not w1143 and not w1144;
w1146 <= w1142 and w1145;
w1147 <= w51 and not w1146;
w1148 <= not w1139 and not w1147;
w1149 <= w1131 and w1148;
w1150 <= w108 and not w1149;
w1151 <= not w1114 and not w1150;
w1152 <= w1078 and w1151;
w1153 <= shift(6) and not w1152;
w1154 <= not w1005 and not w1153;
w1155 <= shift(1) and w590;
w1156 <= not shift(1) and w565;
w1157 <= not w1155 and not w1156;
w1158 <= shift(1) and w595;
w1159 <= not shift(1) and w570;
w1160 <= not w1158 and not w1159;
w1161 <= w1157 and w1160;
w1162 <= w11 and not w1161;
w1163 <= shift(1) and w602;
w1164 <= not shift(1) and w592;
w1165 <= not w1163 and not w1164;
w1166 <= shift(1) and w607;
w1167 <= not shift(1) and w597;
w1168 <= not w1166 and not w1167;
w1169 <= w1165 and w1168;
w1170 <= w24 and not w1169;
w1171 <= not w1162 and not w1170;
w1172 <= shift(1) and w615;
w1173 <= not shift(1) and w629;
w1174 <= not w1172 and not w1173;
w1175 <= shift(1) and w620;
w1176 <= not shift(1) and w634;
w1177 <= not w1175 and not w1176;
w1178 <= w1174 and w1177;
w1179 <= w38 and not w1178;
w1180 <= shift(1) and w627;
w1181 <= not shift(1) and w604;
w1182 <= not w1180 and not w1181;
w1183 <= shift(1) and w632;
w1184 <= not shift(1) and w609;
w1185 <= not w1183 and not w1184;
w1186 <= w1182 and w1185;
w1187 <= w51 and not w1186;
w1188 <= not w1179 and not w1187;
w1189 <= w1171 and w1188;
w1190 <= w215 and not w1189;
w1191 <= shift(1) and w485;
w1192 <= not shift(1) and w617;
w1193 <= not w1191 and not w1192;
w1194 <= shift(1) and w490;
w1195 <= not shift(1) and w622;
w1196 <= not w1194 and not w1195;
w1197 <= w1193 and w1196;
w1198 <= w11 and not w1197;
w1199 <= shift(1) and w497;
w1200 <= not shift(1) and w487;
w1201 <= not w1199 and not w1200;
w1202 <= shift(1) and w502;
w1203 <= not shift(1) and w492;
w1204 <= not w1202 and not w1203;
w1205 <= w1201 and w1204;
w1206 <= w24 and not w1205;
w1207 <= not w1198 and not w1206;
w1208 <= shift(1) and w510;
w1209 <= not shift(1) and w524;
w1210 <= not w1208 and not w1209;
w1211 <= shift(1) and w515;
w1212 <= not shift(1) and w529;
w1213 <= not w1211 and not w1212;
w1214 <= w1210 and w1213;
w1215 <= w38 and not w1214;
w1216 <= shift(1) and w522;
w1217 <= not shift(1) and w499;
w1218 <= not w1216 and not w1217;
w1219 <= shift(1) and w527;
w1220 <= not shift(1) and w504;
w1221 <= not w1219 and not w1220;
w1222 <= w1218 and w1221;
w1223 <= w51 and not w1222;
w1224 <= not w1215 and not w1223;
w1225 <= w1207 and w1224;
w1226 <= w108 and not w1225;
w1227 <= not w1190 and not w1226;
w1228 <= shift(1) and w538;
w1229 <= not shift(1) and w724;
w1230 <= not w1228 and not w1229;
w1231 <= shift(1) and w543;
w1232 <= not shift(1) and w729;
w1233 <= not w1231 and not w1232;
w1234 <= w1230 and w1233;
w1235 <= w11 and not w1234;
w1236 <= shift(1) and w550;
w1237 <= not shift(1) and w540;
w1238 <= not w1236 and not w1237;
w1239 <= shift(1) and w555;
w1240 <= not shift(1) and w545;
w1241 <= not w1239 and not w1240;
w1242 <= w1238 and w1241;
w1243 <= w24 and not w1242;
w1244 <= not w1235 and not w1243;
w1245 <= shift(1) and w563;
w1246 <= not shift(1) and w577;
w1247 <= not w1245 and not w1246;
w1248 <= shift(1) and w568;
w1249 <= not shift(1) and w582;
w1250 <= not w1248 and not w1249;
w1251 <= w1247 and w1250;
w1252 <= w38 and not w1251;
w1253 <= shift(1) and w575;
w1254 <= not shift(1) and w552;
w1255 <= not w1253 and not w1254;
w1256 <= shift(1) and w580;
w1257 <= not shift(1) and w557;
w1258 <= not w1256 and not w1257;
w1259 <= w1255 and w1258;
w1260 <= w51 and not w1259;
w1261 <= not w1252 and not w1260;
w1262 <= w1244 and w1261;
w1263 <= w162 and not w1262;
w1264 <= shift(1) and w433;
w1265 <= not shift(1) and w512;
w1266 <= not w1264 and not w1265;
w1267 <= shift(1) and w438;
w1268 <= not shift(1) and w517;
w1269 <= not w1267 and not w1268;
w1270 <= w1266 and w1269;
w1271 <= w11 and not w1270;
w1272 <= shift(1) and w445;
w1273 <= not shift(1) and w435;
w1274 <= not w1272 and not w1273;
w1275 <= shift(1) and w450;
w1276 <= not shift(1) and w440;
w1277 <= not w1275 and not w1276;
w1278 <= w1274 and w1277;
w1279 <= w24 and not w1278;
w1280 <= not w1271 and not w1279;
w1281 <= shift(1) and w458;
w1282 <= not shift(1) and w472;
w1283 <= not w1281 and not w1282;
w1284 <= shift(1) and w463;
w1285 <= not shift(1) and w477;
w1286 <= not w1284 and not w1285;
w1287 <= w1283 and w1286;
w1288 <= w38 and not w1287;
w1289 <= shift(1) and w470;
w1290 <= not shift(1) and w447;
w1291 <= not w1289 and not w1290;
w1292 <= shift(1) and w475;
w1293 <= not shift(1) and w452;
w1294 <= not w1292 and not w1293;
w1295 <= w1291 and w1294;
w1296 <= w51 and not w1295;
w1297 <= not w1288 and not w1296;
w1298 <= w1280 and w1297;
w1299 <= w55 and not w1298;
w1300 <= not w1263 and not w1299;
w1301 <= w1227 and w1300;
w1302 <= not shift(6) and not w1301;
w1303 <= shift(1) and w645;
w1304 <= not shift(1) and w460;
w1305 <= not w1303 and not w1304;
w1306 <= shift(1) and w650;
w1307 <= not shift(1) and w465;
w1308 <= not w1306 and not w1307;
w1309 <= w1305 and w1308;
w1310 <= w11 and not w1309;
w1311 <= shift(1) and w657;
w1312 <= not shift(1) and w647;
w1313 <= not w1311 and not w1312;
w1314 <= shift(1) and w662;
w1315 <= not shift(1) and w652;
w1316 <= not w1314 and not w1315;
w1317 <= w1313 and w1316;
w1318 <= w24 and not w1317;
w1319 <= not w1310 and not w1318;
w1320 <= shift(1) and w670;
w1321 <= not shift(1) and w684;
w1322 <= not w1320 and not w1321;
w1323 <= shift(1) and w675;
w1324 <= not shift(1) and w689;
w1325 <= not w1323 and not w1324;
w1326 <= w1322 and w1325;
w1327 <= w38 and not w1326;
w1328 <= shift(1) and w682;
w1329 <= not shift(1) and w659;
w1330 <= not w1328 and not w1329;
w1331 <= shift(1) and w687;
w1332 <= not shift(1) and w664;
w1333 <= not w1331 and not w1332;
w1334 <= w1330 and w1333;
w1335 <= w51 and not w1334;
w1336 <= not w1327 and not w1335;
w1337 <= w1319 and w1336;
w1338 <= w162 and not w1337;
w1339 <= shift(1) and w750;
w1340 <= not shift(1) and w672;
w1341 <= not w1339 and not w1340;
w1342 <= shift(1) and w755;
w1343 <= not shift(1) and w677;
w1344 <= not w1342 and not w1343;
w1345 <= w1341 and w1344;
w1346 <= w11 and not w1345;
w1347 <= shift(1) and w769;
w1348 <= shift(1) and w767;
w1349 <= not w1347 and not w1348;
w1350 <= not shift(1) and w757;
w1351 <= not shift(1) and w752;
w1352 <= not w1350 and not w1351;
w1353 <= w1349 and w1352;
w1354 <= w24 and not w1353;
w1355 <= not w1346 and not w1354;
w1356 <= shift(1) and w775;
w1357 <= not shift(1) and w794;
w1358 <= not w1356 and not w1357;
w1359 <= shift(1) and w780;
w1360 <= not shift(1) and w792;
w1361 <= not w1359 and not w1360;
w1362 <= w1358 and w1361;
w1363 <= w38 and not w1362;
w1364 <= shift(1) and w787;
w1365 <= not shift(1) and w762;
w1366 <= not w1364 and not w1365;
w1367 <= shift(1) and w789;
w1368 <= not shift(1) and w764;
w1369 <= not w1367 and not w1368;
w1370 <= w1366 and w1369;
w1371 <= w51 and not w1370;
w1372 <= not w1363 and not w1371;
w1373 <= w1355 and w1372;
w1374 <= w215 and not w1373;
w1375 <= not w1338 and not w1374;
w1376 <= shift(1) and w697;
w1377 <= not shift(1) and w829;
w1378 <= not w1376 and not w1377;
w1379 <= shift(1) and w702;
w1380 <= not shift(1) and w834;
w1381 <= not w1379 and not w1380;
w1382 <= w1378 and w1381;
w1383 <= w11 and not w1382;
w1384 <= shift(1) and w709;
w1385 <= not shift(1) and w699;
w1386 <= not w1384 and not w1385;
w1387 <= shift(1) and w714;
w1388 <= not shift(1) and w704;
w1389 <= not w1387 and not w1388;
w1390 <= w1386 and w1389;
w1391 <= w24 and not w1390;
w1392 <= not w1383 and not w1391;
w1393 <= shift(1) and w722;
w1394 <= not shift(1) and w736;
w1395 <= not w1393 and not w1394;
w1396 <= shift(1) and w727;
w1397 <= not shift(1) and w741;
w1398 <= not w1396 and not w1397;
w1399 <= w1395 and w1398;
w1400 <= w38 and not w1399;
w1401 <= shift(1) and w734;
w1402 <= not shift(1) and w711;
w1403 <= not w1401 and not w1402;
w1404 <= shift(1) and w739;
w1405 <= not shift(1) and w716;
w1406 <= not w1404 and not w1405;
w1407 <= w1403 and w1406;
w1408 <= w51 and not w1407;
w1409 <= not w1400 and not w1408;
w1410 <= w1392 and w1409;
w1411 <= w55 and not w1410;
w1412 <= shift(1) and w802;
w1413 <= not shift(1) and w777;
w1414 <= not w1412 and not w1413;
w1415 <= shift(1) and w807;
w1416 <= not shift(1) and w782;
w1417 <= not w1415 and not w1416;
w1418 <= w1414 and w1417;
w1419 <= w11 and not w1418;
w1420 <= shift(1) and w814;
w1421 <= not shift(1) and w804;
w1422 <= not w1420 and not w1421;
w1423 <= shift(1) and w819;
w1424 <= not shift(1) and w809;
w1425 <= not w1423 and not w1424;
w1426 <= w1422 and w1425;
w1427 <= w24 and not w1426;
w1428 <= not w1419 and not w1427;
w1429 <= shift(1) and w827;
w1430 <= not shift(1) and w841;
w1431 <= not w1429 and not w1430;
w1432 <= shift(1) and w832;
w1433 <= not shift(1) and w846;
w1434 <= not w1432 and not w1433;
w1435 <= w1431 and w1434;
w1436 <= w38 and not w1435;
w1437 <= shift(1) and w839;
w1438 <= not shift(1) and w816;
w1439 <= not w1437 and not w1438;
w1440 <= shift(1) and w844;
w1441 <= not shift(1) and w821;
w1442 <= not w1440 and not w1441;
w1443 <= w1439 and w1442;
w1444 <= w51 and not w1443;
w1445 <= not w1436 and not w1444;
w1446 <= w1428 and w1445;
w1447 <= w108 and not w1446;
w1448 <= not w1411 and not w1447;
w1449 <= w1375 and w1448;
w1450 <= shift(6) and not w1449;
w1451 <= not w1302 and not w1450;
w1452 <= w11 and not w92;
w1453 <= not w10 and w24;
w1454 <= not w1452 and not w1453;
w1455 <= w38 and not w50;
w1456 <= not w23 and w51;
w1457 <= not w1455 and not w1456;
w1458 <= w1454 and w1457;
w1459 <= w55 and not w1458;
w1460 <= w11 and not w199;
w1461 <= w24 and not w67;
w1462 <= not w1460 and not w1461;
w1463 <= w38 and not w104;
w1464 <= w51 and not w79;
w1465 <= not w1463 and not w1464;
w1466 <= w1462 and w1465;
w1467 <= w108 and not w1466;
w1468 <= not w1459 and not w1467;
w1469 <= w11 and not w255;
w1470 <= w24 and not w121;
w1471 <= not w1469 and not w1470;
w1472 <= w38 and not w158;
w1473 <= w51 and not w133;
w1474 <= not w1472 and not w1473;
w1475 <= w1471 and w1474;
w1476 <= w162 and not w1475;
w1477 <= w11 and not w146;
w1478 <= w24 and not w174;
w1479 <= not w1477 and not w1478;
w1480 <= w38 and not w211;
w1481 <= w51 and not w186;
w1482 <= not w1480 and not w1481;
w1483 <= w1479 and w1482;
w1484 <= w215 and not w1483;
w1485 <= not w1476 and not w1484;
w1486 <= w1468 and w1485;
w1487 <= not shift(6) and not w1486;
w1488 <= w11 and not w360;
w1489 <= w24 and not w387;
w1490 <= not w1488 and not w1489;
w1491 <= w38 and not w424;
w1492 <= w51 and not w399;
w1493 <= not w1491 and not w1492;
w1494 <= w1490 and w1493;
w1495 <= w215 and not w1494;
w1496 <= w11 and not w37;
w1497 <= w24 and not w335;
w1498 <= not w1496 and not w1497;
w1499 <= w38 and not w372;
w1500 <= w51 and not w347;
w1501 <= not w1499 and not w1500;
w1502 <= w1498 and w1501;
w1503 <= w162 and not w1502;
w1504 <= not w1495 and not w1503;
w1505 <= w11 and not w412;
w1506 <= w24 and not w282;
w1507 <= not w1505 and not w1506;
w1508 <= w38 and not w319;
w1509 <= w51 and not w294;
w1510 <= not w1508 and not w1509;
w1511 <= w1507 and w1510;
w1512 <= w108 and not w1511;
w1513 <= w11 and not w307;
w1514 <= w24 and not w230;
w1515 <= not w1513 and not w1514;
w1516 <= w38 and not w267;
w1517 <= w51 and not w242;
w1518 <= not w1516 and not w1517;
w1519 <= w1515 and w1518;
w1520 <= w55 and not w1519;
w1521 <= not w1512 and not w1520;
w1522 <= w1504 and w1521;
w1523 <= shift(6) and not w1522;
w1524 <= not w1487 and not w1523;
w1525 <= w11 and not w520;
w1526 <= w24 and not w443;
w1527 <= not w1525 and not w1526;
w1528 <= w38 and not w480;
w1529 <= w51 and not w455;
w1530 <= not w1528 and not w1529;
w1531 <= w1527 and w1530;
w1532 <= w55 and not w1531;
w1533 <= w11 and not w625;
w1534 <= w24 and not w495;
w1535 <= not w1533 and not w1534;
w1536 <= w38 and not w532;
w1537 <= w51 and not w507;
w1538 <= not w1536 and not w1537;
w1539 <= w1535 and w1538;
w1540 <= w108 and not w1539;
w1541 <= not w1532 and not w1540;
w1542 <= w11 and not w732;
w1543 <= w24 and not w548;
w1544 <= not w1542 and not w1543;
w1545 <= w38 and not w585;
w1546 <= w51 and not w560;
w1547 <= not w1545 and not w1546;
w1548 <= w1544 and w1547;
w1549 <= w162 and not w1548;
w1550 <= w11 and not w573;
w1551 <= w24 and not w600;
w1552 <= not w1550 and not w1551;
w1553 <= w38 and not w637;
w1554 <= w51 and not w612;
w1555 <= not w1553 and not w1554;
w1556 <= w1552 and w1555;
w1557 <= w215 and not w1556;
w1558 <= not w1549 and not w1557;
w1559 <= w1541 and w1558;
w1560 <= not shift(6) and not w1559;
w1561 <= w11 and not w680;
w1562 <= w24 and not w760;
w1563 <= not w1561 and not w1562;
w1564 <= w38 and not w797;
w1565 <= w51 and not w772;
w1566 <= not w1564 and not w1565;
w1567 <= w1563 and w1566;
w1568 <= w215 and not w1567;
w1569 <= w11 and not w468;
w1570 <= w24 and not w655;
w1571 <= not w1569 and not w1570;
w1572 <= w38 and not w692;
w1573 <= w51 and not w667;
w1574 <= not w1572 and not w1573;
w1575 <= w1571 and w1574;
w1576 <= w162 and not w1575;
w1577 <= not w1568 and not w1576;
w1578 <= w11 and not w785;
w1579 <= w24 and not w812;
w1580 <= not w1578 and not w1579;
w1581 <= w38 and not w849;
w1582 <= w51 and not w824;
w1583 <= not w1581 and not w1582;
w1584 <= w1580 and w1583;
w1585 <= w108 and not w1584;
w1586 <= w11 and not w837;
w1587 <= w24 and not w707;
w1588 <= not w1586 and not w1587;
w1589 <= w38 and not w744;
w1590 <= w51 and not w719;
w1591 <= not w1589 and not w1590;
w1592 <= w1588 and w1591;
w1593 <= w55 and not w1592;
w1594 <= not w1585 and not w1593;
w1595 <= w1577 and w1594;
w1596 <= shift(6) and not w1595;
w1597 <= not w1560 and not w1596;
w1598 <= w11 and not w917;
w1599 <= w24 and not w864;
w1600 <= not w1598 and not w1599;
w1601 <= w38 and not w889;
w1602 <= w51 and not w872;
w1603 <= not w1601 and not w1602;
w1604 <= w1600 and w1603;
w1605 <= w55 and not w1604;
w1606 <= w11 and not w990;
w1607 <= w24 and not w900;
w1608 <= not w1606 and not w1607;
w1609 <= w38 and not w925;
w1610 <= w51 and not w908;
w1611 <= not w1609 and not w1610;
w1612 <= w1608 and w1611;
w1613 <= w108 and not w1612;
w1614 <= not w1605 and not w1613;
w1615 <= w11 and not w1065;
w1616 <= w24 and not w937;
w1617 <= not w1615 and not w1616;
w1618 <= w38 and not w962;
w1619 <= w51 and not w945;
w1620 <= not w1618 and not w1619;
w1621 <= w1617 and w1620;
w1622 <= w162 and not w1621;
w1623 <= w11 and not w954;
w1624 <= w24 and not w973;
w1625 <= not w1623 and not w1624;
w1626 <= w38 and not w998;
w1627 <= w51 and not w981;
w1628 <= not w1626 and not w1627;
w1629 <= w1625 and w1628;
w1630 <= w215 and not w1629;
w1631 <= not w1622 and not w1630;
w1632 <= w1614 and w1631;
w1633 <= not shift(6) and not w1632;
w1634 <= w11 and not w1029;
w1635 <= w24 and not w1085;
w1636 <= not w1634 and not w1635;
w1637 <= w38 and not w1110;
w1638 <= w51 and not w1093;
w1639 <= not w1637 and not w1638;
w1640 <= w1636 and w1639;
w1641 <= w215 and not w1640;
w1642 <= w11 and not w881;
w1643 <= w24 and not w1012;
w1644 <= not w1642 and not w1643;
w1645 <= w38 and not w1037;
w1646 <= w51 and not w1020;
w1647 <= not w1645 and not w1646;
w1648 <= w1644 and w1647;
w1649 <= w162 and not w1648;
w1650 <= not w1641 and not w1649;
w1651 <= w11 and not w1102;
w1652 <= w24 and not w1121;
w1653 <= not w1651 and not w1652;
w1654 <= w38 and not w1146;
w1655 <= w51 and not w1129;
w1656 <= not w1654 and not w1655;
w1657 <= w1653 and w1656;
w1658 <= w108 and not w1657;
w1659 <= w11 and not w1138;
w1660 <= w24 and not w1048;
w1661 <= not w1659 and not w1660;
w1662 <= w38 and not w1073;
w1663 <= w51 and not w1056;
w1664 <= not w1662 and not w1663;
w1665 <= w1661 and w1664;
w1666 <= w55 and not w1665;
w1667 <= not w1658 and not w1666;
w1668 <= w1650 and w1667;
w1669 <= shift(6) and not w1668;
w1670 <= not w1633 and not w1669;
w1671 <= w11 and not w1214;
w1672 <= w24 and not w1270;
w1673 <= not w1671 and not w1672;
w1674 <= w38 and not w1295;
w1675 <= w51 and not w1278;
w1676 <= not w1674 and not w1675;
w1677 <= w1673 and w1676;
w1678 <= w55 and not w1677;
w1679 <= w11 and not w1178;
w1680 <= w24 and not w1197;
w1681 <= not w1679 and not w1680;
w1682 <= w38 and not w1222;
w1683 <= w51 and not w1205;
w1684 <= not w1682 and not w1683;
w1685 <= w1681 and w1684;
w1686 <= w108 and not w1685;
w1687 <= not w1678 and not w1686;
w1688 <= w11 and not w1399;
w1689 <= w24 and not w1234;
w1690 <= not w1688 and not w1689;
w1691 <= w38 and not w1259;
w1692 <= w51 and not w1242;
w1693 <= not w1691 and not w1692;
w1694 <= w1690 and w1693;
w1695 <= w162 and not w1694;
w1696 <= w11 and not w1251;
w1697 <= w24 and not w1161;
w1698 <= not w1696 and not w1697;
w1699 <= w38 and not w1186;
w1700 <= w51 and not w1169;
w1701 <= not w1699 and not w1700;
w1702 <= w1698 and w1701;
w1703 <= w215 and not w1702;
w1704 <= not w1695 and not w1703;
w1705 <= w1687 and w1704;
w1706 <= not shift(6) and not w1705;
w1707 <= w24 and not w1345;
w1708 <= w51 and not w1353;
w1709 <= not w1707 and not w1708;
w1710 <= w38 and not w1370;
w1711 <= w11 and not w1326;
w1712 <= not w1710 and not w1711;
w1713 <= w1709 and w1712;
w1714 <= w215 and not w1713;
w1715 <= w11 and not w1287;
w1716 <= w24 and not w1309;
w1717 <= not w1715 and not w1716;
w1718 <= w38 and not w1334;
w1719 <= w51 and not w1317;
w1720 <= not w1718 and not w1719;
w1721 <= w1717 and w1720;
w1722 <= w162 and not w1721;
w1723 <= not w1714 and not w1722;
w1724 <= w11 and not w1362;
w1725 <= w24 and not w1418;
w1726 <= not w1724 and not w1725;
w1727 <= w38 and not w1443;
w1728 <= w51 and not w1426;
w1729 <= not w1727 and not w1728;
w1730 <= w1726 and w1729;
w1731 <= w108 and not w1730;
w1732 <= w11 and not w1435;
w1733 <= w24 and not w1382;
w1734 <= not w1732 and not w1733;
w1735 <= w38 and not w1407;
w1736 <= w51 and not w1390;
w1737 <= not w1735 and not w1736;
w1738 <= w1734 and w1737;
w1739 <= w55 and not w1738;
w1740 <= not w1731 and not w1739;
w1741 <= w1723 and w1740;
w1742 <= shift(6) and not w1741;
w1743 <= not w1706 and not w1742;
w1744 <= w11 and not w104;
w1745 <= w24 and not w92;
w1746 <= not w1744 and not w1745;
w1747 <= not w23 and w38;
w1748 <= not w10 and w51;
w1749 <= not w1747 and not w1748;
w1750 <= w1746 and w1749;
w1751 <= w55 and not w1750;
w1752 <= w11 and not w211;
w1753 <= w24 and not w199;
w1754 <= not w1752 and not w1753;
w1755 <= w38 and not w79;
w1756 <= w51 and not w67;
w1757 <= not w1755 and not w1756;
w1758 <= w1754 and w1757;
w1759 <= w108 and not w1758;
w1760 <= not w1751 and not w1759;
w1761 <= w11 and not w267;
w1762 <= w24 and not w255;
w1763 <= not w1761 and not w1762;
w1764 <= w38 and not w133;
w1765 <= w51 and not w121;
w1766 <= not w1764 and not w1765;
w1767 <= w1763 and w1766;
w1768 <= w162 and not w1767;
w1769 <= w11 and not w158;
w1770 <= w24 and not w146;
w1771 <= not w1769 and not w1770;
w1772 <= w38 and not w186;
w1773 <= w51 and not w174;
w1774 <= not w1772 and not w1773;
w1775 <= w1771 and w1774;
w1776 <= w215 and not w1775;
w1777 <= not w1768 and not w1776;
w1778 <= w1760 and w1777;
w1779 <= not shift(6) and not w1778;
w1780 <= w11 and not w372;
w1781 <= w24 and not w360;
w1782 <= not w1780 and not w1781;
w1783 <= w38 and not w399;
w1784 <= w51 and not w387;
w1785 <= not w1783 and not w1784;
w1786 <= w1782 and w1785;
w1787 <= w215 and not w1786;
w1788 <= w11 and not w50;
w1789 <= w24 and not w37;
w1790 <= not w1788 and not w1789;
w1791 <= w38 and not w347;
w1792 <= w51 and not w335;
w1793 <= not w1791 and not w1792;
w1794 <= w1790 and w1793;
w1795 <= w162 and not w1794;
w1796 <= not w1787 and not w1795;
w1797 <= w11 and not w424;
w1798 <= w24 and not w412;
w1799 <= not w1797 and not w1798;
w1800 <= w38 and not w294;
w1801 <= w51 and not w282;
w1802 <= not w1800 and not w1801;
w1803 <= w1799 and w1802;
w1804 <= w108 and not w1803;
w1805 <= w11 and not w319;
w1806 <= w24 and not w307;
w1807 <= not w1805 and not w1806;
w1808 <= w38 and not w242;
w1809 <= w51 and not w230;
w1810 <= not w1808 and not w1809;
w1811 <= w1807 and w1810;
w1812 <= w55 and not w1811;
w1813 <= not w1804 and not w1812;
w1814 <= w1796 and w1813;
w1815 <= shift(6) and not w1814;
w1816 <= not w1779 and not w1815;
w1817 <= w11 and not w532;
w1818 <= w24 and not w520;
w1819 <= not w1817 and not w1818;
w1820 <= w38 and not w455;
w1821 <= w51 and not w443;
w1822 <= not w1820 and not w1821;
w1823 <= w1819 and w1822;
w1824 <= w55 and not w1823;
w1825 <= w11 and not w637;
w1826 <= w24 and not w625;
w1827 <= not w1825 and not w1826;
w1828 <= w38 and not w507;
w1829 <= w51 and not w495;
w1830 <= not w1828 and not w1829;
w1831 <= w1827 and w1830;
w1832 <= w108 and not w1831;
w1833 <= not w1824 and not w1832;
w1834 <= w11 and not w744;
w1835 <= w24 and not w732;
w1836 <= not w1834 and not w1835;
w1837 <= w38 and not w560;
w1838 <= w51 and not w548;
w1839 <= not w1837 and not w1838;
w1840 <= w1836 and w1839;
w1841 <= w162 and not w1840;
w1842 <= w11 and not w585;
w1843 <= w24 and not w573;
w1844 <= not w1842 and not w1843;
w1845 <= w38 and not w612;
w1846 <= w51 and not w600;
w1847 <= not w1845 and not w1846;
w1848 <= w1844 and w1847;
w1849 <= w215 and not w1848;
w1850 <= not w1841 and not w1849;
w1851 <= w1833 and w1850;
w1852 <= not shift(6) and not w1851;
w1853 <= w11 and not w692;
w1854 <= w24 and not w680;
w1855 <= not w1853 and not w1854;
w1856 <= w38 and not w772;
w1857 <= w51 and not w760;
w1858 <= not w1856 and not w1857;
w1859 <= w1855 and w1858;
w1860 <= w215 and not w1859;
w1861 <= w11 and not w480;
w1862 <= w24 and not w468;
w1863 <= not w1861 and not w1862;
w1864 <= w38 and not w667;
w1865 <= w51 and not w655;
w1866 <= not w1864 and not w1865;
w1867 <= w1863 and w1866;
w1868 <= w162 and not w1867;
w1869 <= not w1860 and not w1868;
w1870 <= w11 and not w797;
w1871 <= w24 and not w785;
w1872 <= not w1870 and not w1871;
w1873 <= w38 and not w824;
w1874 <= w51 and not w812;
w1875 <= not w1873 and not w1874;
w1876 <= w1872 and w1875;
w1877 <= w108 and not w1876;
w1878 <= w11 and not w849;
w1879 <= w24 and not w837;
w1880 <= not w1878 and not w1879;
w1881 <= w38 and not w719;
w1882 <= w51 and not w707;
w1883 <= not w1881 and not w1882;
w1884 <= w1880 and w1883;
w1885 <= w55 and not w1884;
w1886 <= not w1877 and not w1885;
w1887 <= w1869 and w1886;
w1888 <= shift(6) and not w1887;
w1889 <= not w1852 and not w1888;
w1890 <= w11 and not w925;
w1891 <= w24 and not w917;
w1892 <= not w1890 and not w1891;
w1893 <= w38 and not w872;
w1894 <= w51 and not w864;
w1895 <= not w1893 and not w1894;
w1896 <= w1892 and w1895;
w1897 <= w55 and not w1896;
w1898 <= w11 and not w998;
w1899 <= w24 and not w990;
w1900 <= not w1898 and not w1899;
w1901 <= w38 and not w908;
w1902 <= w51 and not w900;
w1903 <= not w1901 and not w1902;
w1904 <= w1900 and w1903;
w1905 <= w108 and not w1904;
w1906 <= not w1897 and not w1905;
w1907 <= w11 and not w1073;
w1908 <= w24 and not w1065;
w1909 <= not w1907 and not w1908;
w1910 <= w38 and not w945;
w1911 <= w51 and not w937;
w1912 <= not w1910 and not w1911;
w1913 <= w1909 and w1912;
w1914 <= w162 and not w1913;
w1915 <= w11 and not w962;
w1916 <= w24 and not w954;
w1917 <= not w1915 and not w1916;
w1918 <= w38 and not w981;
w1919 <= w51 and not w973;
w1920 <= not w1918 and not w1919;
w1921 <= w1917 and w1920;
w1922 <= w215 and not w1921;
w1923 <= not w1914 and not w1922;
w1924 <= w1906 and w1923;
w1925 <= not shift(6) and not w1924;
w1926 <= w11 and not w1037;
w1927 <= w24 and not w1029;
w1928 <= not w1926 and not w1927;
w1929 <= w38 and not w1093;
w1930 <= w51 and not w1085;
w1931 <= not w1929 and not w1930;
w1932 <= w1928 and w1931;
w1933 <= w215 and not w1932;
w1934 <= w11 and not w889;
w1935 <= w24 and not w881;
w1936 <= not w1934 and not w1935;
w1937 <= w38 and not w1020;
w1938 <= w51 and not w1012;
w1939 <= not w1937 and not w1938;
w1940 <= w1936 and w1939;
w1941 <= w162 and not w1940;
w1942 <= not w1933 and not w1941;
w1943 <= w11 and not w1110;
w1944 <= w24 and not w1102;
w1945 <= not w1943 and not w1944;
w1946 <= w38 and not w1129;
w1947 <= w51 and not w1121;
w1948 <= not w1946 and not w1947;
w1949 <= w1945 and w1948;
w1950 <= w108 and not w1949;
w1951 <= w11 and not w1146;
w1952 <= w24 and not w1138;
w1953 <= not w1951 and not w1952;
w1954 <= w38 and not w1056;
w1955 <= w51 and not w1048;
w1956 <= not w1954 and not w1955;
w1957 <= w1953 and w1956;
w1958 <= w55 and not w1957;
w1959 <= not w1950 and not w1958;
w1960 <= w1942 and w1959;
w1961 <= shift(6) and not w1960;
w1962 <= not w1925 and not w1961;
w1963 <= w11 and not w1222;
w1964 <= w24 and not w1214;
w1965 <= not w1963 and not w1964;
w1966 <= w38 and not w1278;
w1967 <= w51 and not w1270;
w1968 <= not w1966 and not w1967;
w1969 <= w1965 and w1968;
w1970 <= w55 and not w1969;
w1971 <= w11 and not w1186;
w1972 <= w24 and not w1178;
w1973 <= not w1971 and not w1972;
w1974 <= w38 and not w1205;
w1975 <= w51 and not w1197;
w1976 <= not w1974 and not w1975;
w1977 <= w1973 and w1976;
w1978 <= w108 and not w1977;
w1979 <= not w1970 and not w1978;
w1980 <= w11 and not w1407;
w1981 <= w24 and not w1399;
w1982 <= not w1980 and not w1981;
w1983 <= w38 and not w1242;
w1984 <= w51 and not w1234;
w1985 <= not w1983 and not w1984;
w1986 <= w1982 and w1985;
w1987 <= w162 and not w1986;
w1988 <= w11 and not w1259;
w1989 <= w24 and not w1251;
w1990 <= not w1988 and not w1989;
w1991 <= w38 and not w1169;
w1992 <= w51 and not w1161;
w1993 <= not w1991 and not w1992;
w1994 <= w1990 and w1993;
w1995 <= w215 and not w1994;
w1996 <= not w1987 and not w1995;
w1997 <= w1979 and w1996;
w1998 <= not shift(6) and not w1997;
w1999 <= w11 and not w1334;
w2000 <= w51 and not w1345;
w2001 <= not w1999 and not w2000;
w2002 <= w38 and not w1353;
w2003 <= w24 and not w1326;
w2004 <= not w2002 and not w2003;
w2005 <= w2001 and w2004;
w2006 <= w215 and not w2005;
w2007 <= w11 and not w1295;
w2008 <= w24 and not w1287;
w2009 <= not w2007 and not w2008;
w2010 <= w38 and not w1317;
w2011 <= w51 and not w1309;
w2012 <= not w2010 and not w2011;
w2013 <= w2009 and w2012;
w2014 <= w162 and not w2013;
w2015 <= not w2006 and not w2014;
w2016 <= w11 and not w1370;
w2017 <= w24 and not w1362;
w2018 <= not w2016 and not w2017;
w2019 <= w38 and not w1426;
w2020 <= w51 and not w1418;
w2021 <= not w2019 and not w2020;
w2022 <= w2018 and w2021;
w2023 <= w108 and not w2022;
w2024 <= w11 and not w1443;
w2025 <= w24 and not w1435;
w2026 <= not w2024 and not w2025;
w2027 <= w38 and not w1390;
w2028 <= w51 and not w1382;
w2029 <= not w2027 and not w2028;
w2030 <= w2026 and w2029;
w2031 <= w55 and not w2030;
w2032 <= not w2023 and not w2031;
w2033 <= w2015 and w2032;
w2034 <= shift(6) and not w2033;
w2035 <= not w1998 and not w2034;
w2036 <= w11 and not w79;
w2037 <= w24 and not w104;
w2038 <= not w2036 and not w2037;
w2039 <= not w10 and w38;
w2040 <= w51 and not w92;
w2041 <= not w2039 and not w2040;
w2042 <= w2038 and w2041;
w2043 <= w55 and not w2042;
w2044 <= w11 and not w186;
w2045 <= w24 and not w211;
w2046 <= not w2044 and not w2045;
w2047 <= w38 and not w67;
w2048 <= w51 and not w199;
w2049 <= not w2047 and not w2048;
w2050 <= w2046 and w2049;
w2051 <= w108 and not w2050;
w2052 <= not w2043 and not w2051;
w2053 <= w11 and not w242;
w2054 <= w24 and not w267;
w2055 <= not w2053 and not w2054;
w2056 <= w38 and not w121;
w2057 <= w51 and not w255;
w2058 <= not w2056 and not w2057;
w2059 <= w2055 and w2058;
w2060 <= w162 and not w2059;
w2061 <= w11 and not w133;
w2062 <= w24 and not w158;
w2063 <= not w2061 and not w2062;
w2064 <= w38 and not w174;
w2065 <= w51 and not w146;
w2066 <= not w2064 and not w2065;
w2067 <= w2063 and w2066;
w2068 <= w215 and not w2067;
w2069 <= not w2060 and not w2068;
w2070 <= w2052 and w2069;
w2071 <= not shift(6) and not w2070;
w2072 <= w11 and not w347;
w2073 <= w24 and not w372;
w2074 <= not w2072 and not w2073;
w2075 <= w38 and not w387;
w2076 <= w51 and not w360;
w2077 <= not w2075 and not w2076;
w2078 <= w2074 and w2077;
w2079 <= w215 and not w2078;
w2080 <= w11 and not w23;
w2081 <= w24 and not w50;
w2082 <= not w2080 and not w2081;
w2083 <= w38 and not w335;
w2084 <= not w37 and w51;
w2085 <= not w2083 and not w2084;
w2086 <= w2082 and w2085;
w2087 <= w162 and not w2086;
w2088 <= not w2079 and not w2087;
w2089 <= w11 and not w399;
w2090 <= w24 and not w424;
w2091 <= not w2089 and not w2090;
w2092 <= w38 and not w282;
w2093 <= w51 and not w412;
w2094 <= not w2092 and not w2093;
w2095 <= w2091 and w2094;
w2096 <= w108 and not w2095;
w2097 <= w11 and not w294;
w2098 <= w24 and not w319;
w2099 <= not w2097 and not w2098;
w2100 <= w38 and not w230;
w2101 <= w51 and not w307;
w2102 <= not w2100 and not w2101;
w2103 <= w2099 and w2102;
w2104 <= w55 and not w2103;
w2105 <= not w2096 and not w2104;
w2106 <= w2088 and w2105;
w2107 <= shift(6) and not w2106;
w2108 <= not w2071 and not w2107;
w2109 <= w11 and not w507;
w2110 <= w24 and not w532;
w2111 <= not w2109 and not w2110;
w2112 <= w38 and not w443;
w2113 <= w51 and not w520;
w2114 <= not w2112 and not w2113;
w2115 <= w2111 and w2114;
w2116 <= w55 and not w2115;
w2117 <= w11 and not w612;
w2118 <= w24 and not w637;
w2119 <= not w2117 and not w2118;
w2120 <= w38 and not w495;
w2121 <= w51 and not w625;
w2122 <= not w2120 and not w2121;
w2123 <= w2119 and w2122;
w2124 <= w108 and not w2123;
w2125 <= not w2116 and not w2124;
w2126 <= w11 and not w719;
w2127 <= w24 and not w744;
w2128 <= not w2126 and not w2127;
w2129 <= w38 and not w548;
w2130 <= w51 and not w732;
w2131 <= not w2129 and not w2130;
w2132 <= w2128 and w2131;
w2133 <= w162 and not w2132;
w2134 <= w11 and not w560;
w2135 <= w24 and not w585;
w2136 <= not w2134 and not w2135;
w2137 <= w38 and not w600;
w2138 <= w51 and not w573;
w2139 <= not w2137 and not w2138;
w2140 <= w2136 and w2139;
w2141 <= w215 and not w2140;
w2142 <= not w2133 and not w2141;
w2143 <= w2125 and w2142;
w2144 <= not shift(6) and not w2143;
w2145 <= w11 and not w667;
w2146 <= w24 and not w692;
w2147 <= not w2145 and not w2146;
w2148 <= w38 and not w760;
w2149 <= w51 and not w680;
w2150 <= not w2148 and not w2149;
w2151 <= w2147 and w2150;
w2152 <= w215 and not w2151;
w2153 <= w11 and not w455;
w2154 <= w24 and not w480;
w2155 <= not w2153 and not w2154;
w2156 <= w38 and not w655;
w2157 <= w51 and not w468;
w2158 <= not w2156 and not w2157;
w2159 <= w2155 and w2158;
w2160 <= w162 and not w2159;
w2161 <= not w2152 and not w2160;
w2162 <= w11 and not w772;
w2163 <= w24 and not w797;
w2164 <= not w2162 and not w2163;
w2165 <= w38 and not w812;
w2166 <= w51 and not w785;
w2167 <= not w2165 and not w2166;
w2168 <= w2164 and w2167;
w2169 <= w108 and not w2168;
w2170 <= w11 and not w824;
w2171 <= w24 and not w849;
w2172 <= not w2170 and not w2171;
w2173 <= w38 and not w707;
w2174 <= w51 and not w837;
w2175 <= not w2173 and not w2174;
w2176 <= w2172 and w2175;
w2177 <= w55 and not w2176;
w2178 <= not w2169 and not w2177;
w2179 <= w2161 and w2178;
w2180 <= shift(6) and not w2179;
w2181 <= not w2144 and not w2180;
w2182 <= w11 and not w908;
w2183 <= w24 and not w925;
w2184 <= not w2182 and not w2183;
w2185 <= w38 and not w864;
w2186 <= w51 and not w917;
w2187 <= not w2185 and not w2186;
w2188 <= w2184 and w2187;
w2189 <= w55 and not w2188;
w2190 <= w11 and not w981;
w2191 <= w24 and not w998;
w2192 <= not w2190 and not w2191;
w2193 <= w38 and not w900;
w2194 <= w51 and not w990;
w2195 <= not w2193 and not w2194;
w2196 <= w2192 and w2195;
w2197 <= w108 and not w2196;
w2198 <= not w2189 and not w2197;
w2199 <= w11 and not w1056;
w2200 <= w24 and not w1073;
w2201 <= not w2199 and not w2200;
w2202 <= w38 and not w937;
w2203 <= w51 and not w1065;
w2204 <= not w2202 and not w2203;
w2205 <= w2201 and w2204;
w2206 <= w162 and not w2205;
w2207 <= w11 and not w945;
w2208 <= w24 and not w962;
w2209 <= not w2207 and not w2208;
w2210 <= w38 and not w973;
w2211 <= w51 and not w954;
w2212 <= not w2210 and not w2211;
w2213 <= w2209 and w2212;
w2214 <= w215 and not w2213;
w2215 <= not w2206 and not w2214;
w2216 <= w2198 and w2215;
w2217 <= not shift(6) and not w2216;
w2218 <= w11 and not w1020;
w2219 <= w24 and not w1037;
w2220 <= not w2218 and not w2219;
w2221 <= w38 and not w1085;
w2222 <= w51 and not w1029;
w2223 <= not w2221 and not w2222;
w2224 <= w2220 and w2223;
w2225 <= w215 and not w2224;
w2226 <= w11 and not w872;
w2227 <= w24 and not w889;
w2228 <= not w2226 and not w2227;
w2229 <= w38 and not w1012;
w2230 <= w51 and not w881;
w2231 <= not w2229 and not w2230;
w2232 <= w2228 and w2231;
w2233 <= w162 and not w2232;
w2234 <= not w2225 and not w2233;
w2235 <= w11 and not w1093;
w2236 <= w24 and not w1110;
w2237 <= not w2235 and not w2236;
w2238 <= w38 and not w1121;
w2239 <= w51 and not w1102;
w2240 <= not w2238 and not w2239;
w2241 <= w2237 and w2240;
w2242 <= w108 and not w2241;
w2243 <= w11 and not w1129;
w2244 <= w24 and not w1146;
w2245 <= not w2243 and not w2244;
w2246 <= w38 and not w1048;
w2247 <= w51 and not w1138;
w2248 <= not w2246 and not w2247;
w2249 <= w2245 and w2248;
w2250 <= w55 and not w2249;
w2251 <= not w2242 and not w2250;
w2252 <= w2234 and w2251;
w2253 <= shift(6) and not w2252;
w2254 <= not w2217 and not w2253;
w2255 <= w11 and not w1205;
w2256 <= w24 and not w1222;
w2257 <= not w2255 and not w2256;
w2258 <= w38 and not w1270;
w2259 <= w51 and not w1214;
w2260 <= not w2258 and not w2259;
w2261 <= w2257 and w2260;
w2262 <= w55 and not w2261;
w2263 <= w11 and not w1169;
w2264 <= w24 and not w1186;
w2265 <= not w2263 and not w2264;
w2266 <= w38 and not w1197;
w2267 <= w51 and not w1178;
w2268 <= not w2266 and not w2267;
w2269 <= w2265 and w2268;
w2270 <= w108 and not w2269;
w2271 <= not w2262 and not w2270;
w2272 <= w11 and not w1390;
w2273 <= w24 and not w1407;
w2274 <= not w2272 and not w2273;
w2275 <= w38 and not w1234;
w2276 <= w51 and not w1399;
w2277 <= not w2275 and not w2276;
w2278 <= w2274 and w2277;
w2279 <= w162 and not w2278;
w2280 <= w11 and not w1242;
w2281 <= w24 and not w1259;
w2282 <= not w2280 and not w2281;
w2283 <= w38 and not w1161;
w2284 <= w51 and not w1251;
w2285 <= not w2283 and not w2284;
w2286 <= w2282 and w2285;
w2287 <= w215 and not w2286;
w2288 <= not w2279 and not w2287;
w2289 <= w2271 and w2288;
w2290 <= not shift(6) and not w2289;
w2291 <= w11 and not w1317;
w2292 <= w24 and not w1334;
w2293 <= not w2291 and not w2292;
w2294 <= w38 and not w1345;
w2295 <= w51 and not w1326;
w2296 <= not w2294 and not w2295;
w2297 <= w2293 and w2296;
w2298 <= w215 and not w2297;
w2299 <= w11 and not w1278;
w2300 <= w24 and not w1295;
w2301 <= not w2299 and not w2300;
w2302 <= w38 and not w1309;
w2303 <= w51 and not w1287;
w2304 <= not w2302 and not w2303;
w2305 <= w2301 and w2304;
w2306 <= w162 and not w2305;
w2307 <= not w2298 and not w2306;
w2308 <= w11 and not w1353;
w2309 <= w24 and not w1370;
w2310 <= not w2308 and not w2309;
w2311 <= w38 and not w1418;
w2312 <= w51 and not w1362;
w2313 <= not w2311 and not w2312;
w2314 <= w2310 and w2313;
w2315 <= w108 and not w2314;
w2316 <= w11 and not w1426;
w2317 <= w24 and not w1443;
w2318 <= not w2316 and not w2317;
w2319 <= w38 and not w1382;
w2320 <= w51 and not w1435;
w2321 <= not w2319 and not w2320;
w2322 <= w2318 and w2321;
w2323 <= w55 and not w2322;
w2324 <= not w2315 and not w2323;
w2325 <= w2307 and w2324;
w2326 <= shift(6) and not w2325;
w2327 <= not w2290 and not w2326;
w2328 <= w55 and not w107;
w2329 <= w108 and not w214;
w2330 <= not w2328 and not w2329;
w2331 <= w162 and not w270;
w2332 <= not w161 and w215;
w2333 <= not w2331 and not w2332;
w2334 <= w2330 and w2333;
w2335 <= not shift(6) and not w2334;
w2336 <= not w54 and w162;
w2337 <= w55 and not w322;
w2338 <= not w2336 and not w2337;
w2339 <= w215 and not w375;
w2340 <= w108 and not w427;
w2341 <= not w2339 and not w2340;
w2342 <= w2338 and w2341;
w2343 <= shift(6) and not w2342;
w2344 <= not w2335 and not w2343;
w2345 <= w55 and not w535;
w2346 <= w108 and not w640;
w2347 <= not w2345 and not w2346;
w2348 <= w162 and not w747;
w2349 <= w215 and not w588;
w2350 <= not w2348 and not w2349;
w2351 <= w2347 and w2350;
w2352 <= not shift(6) and not w2351;
w2353 <= w215 and not w695;
w2354 <= w162 and not w483;
w2355 <= not w2353 and not w2354;
w2356 <= w108 and not w800;
w2357 <= w55 and not w852;
w2358 <= not w2356 and not w2357;
w2359 <= w2355 and w2358;
w2360 <= shift(6) and not w2359;
w2361 <= not w2352 and not w2360;
w2362 <= w55 and not w928;
w2363 <= w108 and not w1001;
w2364 <= not w2362 and not w2363;
w2365 <= w162 and not w1076;
w2366 <= w215 and not w965;
w2367 <= not w2365 and not w2366;
w2368 <= w2364 and w2367;
w2369 <= not shift(6) and not w2368;
w2370 <= w215 and not w1040;
w2371 <= w162 and not w892;
w2372 <= not w2370 and not w2371;
w2373 <= w108 and not w1113;
w2374 <= w55 and not w1149;
w2375 <= not w2373 and not w2374;
w2376 <= w2372 and w2375;
w2377 <= shift(6) and not w2376;
w2378 <= not w2369 and not w2377;
w2379 <= w108 and not w1189;
w2380 <= w55 and not w1225;
w2381 <= not w2379 and not w2380;
w2382 <= w215 and not w1262;
w2383 <= w162 and not w1410;
w2384 <= not w2382 and not w2383;
w2385 <= w2381 and w2384;
w2386 <= not shift(6) and not w2385;
w2387 <= w215 and not w1337;
w2388 <= w162 and not w1298;
w2389 <= not w2387 and not w2388;
w2390 <= w55 and not w1446;
w2391 <= w108 and not w1373;
w2392 <= not w2390 and not w2391;
w2393 <= w2389 and w2392;
w2394 <= shift(6) and not w2393;
w2395 <= not w2386 and not w2394;
w2396 <= w55 and not w1466;
w2397 <= w108 and not w1483;
w2398 <= not w2396 and not w2397;
w2399 <= w162 and not w1519;
w2400 <= w215 and not w1475;
w2401 <= not w2399 and not w2400;
w2402 <= w2398 and w2401;
w2403 <= not shift(6) and not w2402;
w2404 <= w162 and not w1458;
w2405 <= w108 and not w1494;
w2406 <= not w2404 and not w2405;
w2407 <= w55 and not w1511;
w2408 <= w215 and not w1502;
w2409 <= not w2407 and not w2408;
w2410 <= w2406 and w2409;
w2411 <= shift(6) and not w2410;
w2412 <= not w2403 and not w2411;
w2413 <= w55 and not w1539;
w2414 <= w108 and not w1556;
w2415 <= not w2413 and not w2414;
w2416 <= w162 and not w1592;
w2417 <= w215 and not w1548;
w2418 <= not w2416 and not w2417;
w2419 <= w2415 and w2418;
w2420 <= not shift(6) and not w2419;
w2421 <= w162 and not w1531;
w2422 <= w108 and not w1567;
w2423 <= not w2421 and not w2422;
w2424 <= w55 and not w1584;
w2425 <= w215 and not w1575;
w2426 <= not w2424 and not w2425;
w2427 <= w2423 and w2426;
w2428 <= shift(6) and not w2427;
w2429 <= not w2420 and not w2428;
w2430 <= w55 and not w1612;
w2431 <= w108 and not w1629;
w2432 <= not w2430 and not w2431;
w2433 <= w162 and not w1665;
w2434 <= w215 and not w1621;
w2435 <= not w2433 and not w2434;
w2436 <= w2432 and w2435;
w2437 <= not shift(6) and not w2436;
w2438 <= w162 and not w1604;
w2439 <= w108 and not w1640;
w2440 <= not w2438 and not w2439;
w2441 <= w55 and not w1657;
w2442 <= w215 and not w1648;
w2443 <= not w2441 and not w2442;
w2444 <= w2440 and w2443;
w2445 <= shift(6) and not w2444;
w2446 <= not w2437 and not w2445;
w2447 <= w55 and not w1685;
w2448 <= w162 and not w1738;
w2449 <= not w2447 and not w2448;
w2450 <= w215 and not w1694;
w2451 <= w108 and not w1702;
w2452 <= not w2450 and not w2451;
w2453 <= w2449 and w2452;
w2454 <= not shift(6) and not w2453;
w2455 <= w108 and not w1713;
w2456 <= w215 and not w1721;
w2457 <= not w2455 and not w2456;
w2458 <= w55 and not w1730;
w2459 <= w162 and not w1677;
w2460 <= not w2458 and not w2459;
w2461 <= w2457 and w2460;
w2462 <= shift(6) and not w2461;
w2463 <= not w2454 and not w2462;
w2464 <= w55 and not w1758;
w2465 <= w162 and not w1811;
w2466 <= not w2464 and not w2465;
w2467 <= w215 and not w1767;
w2468 <= w108 and not w1775;
w2469 <= not w2467 and not w2468;
w2470 <= w2466 and w2469;
w2471 <= not shift(6) and not w2470;
w2472 <= w108 and not w1786;
w2473 <= w215 and not w1794;
w2474 <= not w2472 and not w2473;
w2475 <= w55 and not w1803;
w2476 <= w162 and not w1750;
w2477 <= not w2475 and not w2476;
w2478 <= w2474 and w2477;
w2479 <= shift(6) and not w2478;
w2480 <= not w2471 and not w2479;
w2481 <= w55 and not w1831;
w2482 <= w162 and not w1884;
w2483 <= not w2481 and not w2482;
w2484 <= w215 and not w1840;
w2485 <= w108 and not w1848;
w2486 <= not w2484 and not w2485;
w2487 <= w2483 and w2486;
w2488 <= not shift(6) and not w2487;
w2489 <= w108 and not w1859;
w2490 <= w215 and not w1867;
w2491 <= not w2489 and not w2490;
w2492 <= w55 and not w1876;
w2493 <= w162 and not w1823;
w2494 <= not w2492 and not w2493;
w2495 <= w2491 and w2494;
w2496 <= shift(6) and not w2495;
w2497 <= not w2488 and not w2496;
w2498 <= w55 and not w1904;
w2499 <= w108 and not w1921;
w2500 <= not w2498 and not w2499;
w2501 <= w162 and not w1957;
w2502 <= w215 and not w1913;
w2503 <= not w2501 and not w2502;
w2504 <= w2500 and w2503;
w2505 <= not shift(6) and not w2504;
w2506 <= w108 and not w1932;
w2507 <= w215 and not w1940;
w2508 <= not w2506 and not w2507;
w2509 <= w55 and not w1949;
w2510 <= w162 and not w1896;
w2511 <= not w2509 and not w2510;
w2512 <= w2508 and w2511;
w2513 <= shift(6) and not w2512;
w2514 <= not w2505 and not w2513;
w2515 <= w55 and not w1977;
w2516 <= w108 and not w1994;
w2517 <= not w2515 and not w2516;
w2518 <= w162 and not w2030;
w2519 <= w215 and not w1986;
w2520 <= not w2518 and not w2519;
w2521 <= w2517 and w2520;
w2522 <= not shift(6) and not w2521;
w2523 <= w108 and not w2005;
w2524 <= w215 and not w2013;
w2525 <= not w2523 and not w2524;
w2526 <= w55 and not w2022;
w2527 <= w162 and not w1969;
w2528 <= not w2526 and not w2527;
w2529 <= w2525 and w2528;
w2530 <= shift(6) and not w2529;
w2531 <= not w2522 and not w2530;
w2532 <= w55 and not w2050;
w2533 <= w108 and not w2067;
w2534 <= not w2532 and not w2533;
w2535 <= w162 and not w2103;
w2536 <= w215 and not w2059;
w2537 <= not w2535 and not w2536;
w2538 <= w2534 and w2537;
w2539 <= not shift(6) and not w2538;
w2540 <= w108 and not w2078;
w2541 <= w215 and not w2086;
w2542 <= not w2540 and not w2541;
w2543 <= w55 and not w2095;
w2544 <= w162 and not w2042;
w2545 <= not w2543 and not w2544;
w2546 <= w2542 and w2545;
w2547 <= shift(6) and not w2546;
w2548 <= not w2539 and not w2547;
w2549 <= w55 and not w2123;
w2550 <= w108 and not w2140;
w2551 <= not w2549 and not w2550;
w2552 <= w162 and not w2176;
w2553 <= w215 and not w2132;
w2554 <= not w2552 and not w2553;
w2555 <= w2551 and w2554;
w2556 <= not shift(6) and not w2555;
w2557 <= w108 and not w2151;
w2558 <= w215 and not w2159;
w2559 <= not w2557 and not w2558;
w2560 <= w55 and not w2168;
w2561 <= w162 and not w2115;
w2562 <= not w2560 and not w2561;
w2563 <= w2559 and w2562;
w2564 <= shift(6) and not w2563;
w2565 <= not w2556 and not w2564;
w2566 <= w55 and not w2196;
w2567 <= w108 and not w2213;
w2568 <= not w2566 and not w2567;
w2569 <= w162 and not w2249;
w2570 <= w215 and not w2205;
w2571 <= not w2569 and not w2570;
w2572 <= w2568 and w2571;
w2573 <= not shift(6) and not w2572;
w2574 <= w108 and not w2224;
w2575 <= w215 and not w2232;
w2576 <= not w2574 and not w2575;
w2577 <= w55 and not w2241;
w2578 <= w162 and not w2188;
w2579 <= not w2577 and not w2578;
w2580 <= w2576 and w2579;
w2581 <= shift(6) and not w2580;
w2582 <= not w2573 and not w2581;
w2583 <= w55 and not w2269;
w2584 <= w108 and not w2286;
w2585 <= not w2583 and not w2584;
w2586 <= w162 and not w2322;
w2587 <= w215 and not w2278;
w2588 <= not w2586 and not w2587;
w2589 <= w2585 and w2588;
w2590 <= not shift(6) and not w2589;
w2591 <= w108 and not w2297;
w2592 <= w215 and not w2305;
w2593 <= not w2591 and not w2592;
w2594 <= w55 and not w2314;
w2595 <= w162 and not w2261;
w2596 <= not w2594 and not w2595;
w2597 <= w2593 and w2596;
w2598 <= shift(6) and not w2597;
w2599 <= not w2590 and not w2598;
w2600 <= w55 and not w214;
w2601 <= w108 and not w161;
w2602 <= not w2600 and not w2601;
w2603 <= w162 and not w322;
w2604 <= w215 and not w270;
w2605 <= not w2603 and not w2604;
w2606 <= w2602 and w2605;
w2607 <= not shift(6) and not w2606;
w2608 <= not w54 and w215;
w2609 <= not w107 and w162;
w2610 <= not w2608 and not w2609;
w2611 <= w108 and not w375;
w2612 <= w55 and not w427;
w2613 <= not w2611 and not w2612;
w2614 <= w2610 and w2613;
w2615 <= shift(6) and not w2614;
w2616 <= not w2607 and not w2615;
w2617 <= w55 and not w640;
w2618 <= w108 and not w588;
w2619 <= not w2617 and not w2618;
w2620 <= w162 and not w852;
w2621 <= w215 and not w747;
w2622 <= not w2620 and not w2621;
w2623 <= w2619 and w2622;
w2624 <= not shift(6) and not w2623;
w2625 <= w108 and not w695;
w2626 <= w215 and not w483;
w2627 <= not w2625 and not w2626;
w2628 <= w55 and not w800;
w2629 <= w162 and not w535;
w2630 <= not w2628 and not w2629;
w2631 <= w2627 and w2630;
w2632 <= shift(6) and not w2631;
w2633 <= not w2624 and not w2632;
w2634 <= w55 and not w1001;
w2635 <= w108 and not w965;
w2636 <= not w2634 and not w2635;
w2637 <= w162 and not w1149;
w2638 <= w215 and not w1076;
w2639 <= not w2637 and not w2638;
w2640 <= w2636 and w2639;
w2641 <= not shift(6) and not w2640;
w2642 <= w108 and not w1040;
w2643 <= w215 and not w892;
w2644 <= not w2642 and not w2643;
w2645 <= w55 and not w1113;
w2646 <= w162 and not w928;
w2647 <= not w2645 and not w2646;
w2648 <= w2644 and w2647;
w2649 <= shift(6) and not w2648;
w2650 <= not w2641 and not w2649;
w2651 <= w55 and not w1189;
w2652 <= w162 and not w1446;
w2653 <= not w2651 and not w2652;
w2654 <= w108 and not w1262;
w2655 <= w215 and not w1410;
w2656 <= not w2654 and not w2655;
w2657 <= w2653 and w2656;
w2658 <= not shift(6) and not w2657;
w2659 <= w108 and not w1337;
w2660 <= w162 and not w1225;
w2661 <= not w2659 and not w2660;
w2662 <= w55 and not w1373;
w2663 <= w215 and not w1298;
w2664 <= not w2662 and not w2663;
w2665 <= w2661 and w2664;
w2666 <= shift(6) and not w2665;
w2667 <= not w2658 and not w2666;
w2668 <= w55 and not w1483;
w2669 <= w108 and not w1475;
w2670 <= not w2668 and not w2669;
w2671 <= w162 and not w1511;
w2672 <= w215 and not w1519;
w2673 <= not w2671 and not w2672;
w2674 <= w2670 and w2673;
w2675 <= not shift(6) and not w2674;
w2676 <= w215 and not w1458;
w2677 <= w162 and not w1466;
w2678 <= not w2676 and not w2677;
w2679 <= w108 and not w1502;
w2680 <= w55 and not w1494;
w2681 <= not w2679 and not w2680;
w2682 <= w2678 and w2681;
w2683 <= shift(6) and not w2682;
w2684 <= not w2675 and not w2683;
w2685 <= w55 and not w1556;
w2686 <= w108 and not w1548;
w2687 <= not w2685 and not w2686;
w2688 <= w162 and not w1584;
w2689 <= w215 and not w1592;
w2690 <= not w2688 and not w2689;
w2691 <= w2687 and w2690;
w2692 <= not shift(6) and not w2691;
w2693 <= w215 and not w1531;
w2694 <= w162 and not w1539;
w2695 <= not w2693 and not w2694;
w2696 <= w108 and not w1575;
w2697 <= w55 and not w1567;
w2698 <= not w2696 and not w2697;
w2699 <= w2695 and w2698;
w2700 <= shift(6) and not w2699;
w2701 <= not w2692 and not w2700;
w2702 <= w55 and not w1629;
w2703 <= w108 and not w1621;
w2704 <= not w2702 and not w2703;
w2705 <= w162 and not w1657;
w2706 <= w215 and not w1665;
w2707 <= not w2705 and not w2706;
w2708 <= w2704 and w2707;
w2709 <= not shift(6) and not w2708;
w2710 <= w215 and not w1604;
w2711 <= w162 and not w1612;
w2712 <= not w2710 and not w2711;
w2713 <= w108 and not w1648;
w2714 <= w55 and not w1640;
w2715 <= not w2713 and not w2714;
w2716 <= w2712 and w2715;
w2717 <= shift(6) and not w2716;
w2718 <= not w2709 and not w2717;
w2719 <= w215 and not w1738;
w2720 <= w162 and not w1730;
w2721 <= not w2719 and not w2720;
w2722 <= w108 and not w1694;
w2723 <= w55 and not w1702;
w2724 <= not w2722 and not w2723;
w2725 <= w2721 and w2724;
w2726 <= not shift(6) and not w2725;
w2727 <= w55 and not w1713;
w2728 <= w108 and not w1721;
w2729 <= not w2727 and not w2728;
w2730 <= w162 and not w1685;
w2731 <= w215 and not w1677;
w2732 <= not w2730 and not w2731;
w2733 <= w2729 and w2732;
w2734 <= shift(6) and not w2733;
w2735 <= not w2726 and not w2734;
w2736 <= w215 and not w1811;
w2737 <= w162 and not w1803;
w2738 <= not w2736 and not w2737;
w2739 <= w108 and not w1767;
w2740 <= w55 and not w1775;
w2741 <= not w2739 and not w2740;
w2742 <= w2738 and w2741;
w2743 <= not shift(6) and not w2742;
w2744 <= w55 and not w1786;
w2745 <= w108 and not w1794;
w2746 <= not w2744 and not w2745;
w2747 <= w162 and not w1758;
w2748 <= w215 and not w1750;
w2749 <= not w2747 and not w2748;
w2750 <= w2746 and w2749;
w2751 <= shift(6) and not w2750;
w2752 <= not w2743 and not w2751;
w2753 <= w215 and not w1884;
w2754 <= w162 and not w1876;
w2755 <= not w2753 and not w2754;
w2756 <= w108 and not w1840;
w2757 <= w55 and not w1848;
w2758 <= not w2756 and not w2757;
w2759 <= w2755 and w2758;
w2760 <= not shift(6) and not w2759;
w2761 <= w55 and not w1859;
w2762 <= w108 and not w1867;
w2763 <= not w2761 and not w2762;
w2764 <= w162 and not w1831;
w2765 <= w215 and not w1823;
w2766 <= not w2764 and not w2765;
w2767 <= w2763 and w2766;
w2768 <= shift(6) and not w2767;
w2769 <= not w2760 and not w2768;
w2770 <= w55 and not w1921;
w2771 <= w108 and not w1913;
w2772 <= not w2770 and not w2771;
w2773 <= w162 and not w1949;
w2774 <= w215 and not w1957;
w2775 <= not w2773 and not w2774;
w2776 <= w2772 and w2775;
w2777 <= not shift(6) and not w2776;
w2778 <= w55 and not w1932;
w2779 <= w108 and not w1940;
w2780 <= not w2778 and not w2779;
w2781 <= w162 and not w1904;
w2782 <= w215 and not w1896;
w2783 <= not w2781 and not w2782;
w2784 <= w2780 and w2783;
w2785 <= shift(6) and not w2784;
w2786 <= not w2777 and not w2785;
w2787 <= w55 and not w1994;
w2788 <= w108 and not w1986;
w2789 <= not w2787 and not w2788;
w2790 <= w162 and not w2022;
w2791 <= w215 and not w2030;
w2792 <= not w2790 and not w2791;
w2793 <= w2789 and w2792;
w2794 <= not shift(6) and not w2793;
w2795 <= w55 and not w2005;
w2796 <= w108 and not w2013;
w2797 <= not w2795 and not w2796;
w2798 <= w162 and not w1977;
w2799 <= w215 and not w1969;
w2800 <= not w2798 and not w2799;
w2801 <= w2797 and w2800;
w2802 <= shift(6) and not w2801;
w2803 <= not w2794 and not w2802;
w2804 <= w55 and not w2067;
w2805 <= w108 and not w2059;
w2806 <= not w2804 and not w2805;
w2807 <= w162 and not w2095;
w2808 <= w215 and not w2103;
w2809 <= not w2807 and not w2808;
w2810 <= w2806 and w2809;
w2811 <= not shift(6) and not w2810;
w2812 <= w55 and not w2078;
w2813 <= w108 and not w2086;
w2814 <= not w2812 and not w2813;
w2815 <= w162 and not w2050;
w2816 <= w215 and not w2042;
w2817 <= not w2815 and not w2816;
w2818 <= w2814 and w2817;
w2819 <= shift(6) and not w2818;
w2820 <= not w2811 and not w2819;
w2821 <= w55 and not w2140;
w2822 <= w108 and not w2132;
w2823 <= not w2821 and not w2822;
w2824 <= w162 and not w2168;
w2825 <= w215 and not w2176;
w2826 <= not w2824 and not w2825;
w2827 <= w2823 and w2826;
w2828 <= not shift(6) and not w2827;
w2829 <= w55 and not w2151;
w2830 <= w108 and not w2159;
w2831 <= not w2829 and not w2830;
w2832 <= w162 and not w2123;
w2833 <= w215 and not w2115;
w2834 <= not w2832 and not w2833;
w2835 <= w2831 and w2834;
w2836 <= shift(6) and not w2835;
w2837 <= not w2828 and not w2836;
w2838 <= w55 and not w2213;
w2839 <= w108 and not w2205;
w2840 <= not w2838 and not w2839;
w2841 <= w162 and not w2241;
w2842 <= w215 and not w2249;
w2843 <= not w2841 and not w2842;
w2844 <= w2840 and w2843;
w2845 <= not shift(6) and not w2844;
w2846 <= w55 and not w2224;
w2847 <= w108 and not w2232;
w2848 <= not w2846 and not w2847;
w2849 <= w162 and not w2196;
w2850 <= w215 and not w2188;
w2851 <= not w2849 and not w2850;
w2852 <= w2848 and w2851;
w2853 <= shift(6) and not w2852;
w2854 <= not w2845 and not w2853;
w2855 <= w55 and not w2286;
w2856 <= w108 and not w2278;
w2857 <= not w2855 and not w2856;
w2858 <= w162 and not w2314;
w2859 <= w215 and not w2322;
w2860 <= not w2858 and not w2859;
w2861 <= w2857 and w2860;
w2862 <= not shift(6) and not w2861;
w2863 <= w55 and not w2297;
w2864 <= w108 and not w2305;
w2865 <= not w2863 and not w2864;
w2866 <= w162 and not w2269;
w2867 <= w215 and not w2261;
w2868 <= not w2866 and not w2867;
w2869 <= w2865 and w2868;
w2870 <= shift(6) and not w2869;
w2871 <= not w2862 and not w2870;
w2872 <= w55 and not w161;
w2873 <= w108 and not w270;
w2874 <= not w2872 and not w2873;
w2875 <= w162 and not w427;
w2876 <= w215 and not w322;
w2877 <= not w2875 and not w2876;
w2878 <= w2874 and w2877;
w2879 <= not shift(6) and not w2878;
w2880 <= not w54 and w108;
w2881 <= not w107 and w215;
w2882 <= not w2880 and not w2881;
w2883 <= w55 and not w375;
w2884 <= w162 and not w214;
w2885 <= not w2883 and not w2884;
w2886 <= w2882 and w2885;
w2887 <= shift(6) and not w2886;
w2888 <= not w2879 and not w2887;
w2889 <= w55 and not w588;
w2890 <= w108 and not w747;
w2891 <= not w2889 and not w2890;
w2892 <= w162 and not w800;
w2893 <= w215 and not w852;
w2894 <= not w2892 and not w2893;
w2895 <= w2891 and w2894;
w2896 <= not shift(6) and not w2895;
w2897 <= w55 and not w695;
w2898 <= w108 and not w483;
w2899 <= not w2897 and not w2898;
w2900 <= w162 and not w640;
w2901 <= w215 and not w535;
w2902 <= not w2900 and not w2901;
w2903 <= w2899 and w2902;
w2904 <= shift(6) and not w2903;
w2905 <= not w2896 and not w2904;
w2906 <= w55 and not w965;
w2907 <= w108 and not w1076;
w2908 <= not w2906 and not w2907;
w2909 <= w162 and not w1113;
w2910 <= w215 and not w1149;
w2911 <= not w2909 and not w2910;
w2912 <= w2908 and w2911;
w2913 <= not shift(6) and not w2912;
w2914 <= w55 and not w1040;
w2915 <= w108 and not w892;
w2916 <= not w2914 and not w2915;
w2917 <= w162 and not w1001;
w2918 <= w215 and not w928;
w2919 <= not w2917 and not w2918;
w2920 <= w2916 and w2919;
w2921 <= shift(6) and not w2920;
w2922 <= not w2913 and not w2921;
w2923 <= w162 and not w1373;
w2924 <= w215 and not w1446;
w2925 <= not w2923 and not w2924;
w2926 <= w55 and not w1262;
w2927 <= w108 and not w1410;
w2928 <= not w2926 and not w2927;
w2929 <= w2925 and w2928;
w2930 <= not shift(6) and not w2929;
w2931 <= w55 and not w1337;
w2932 <= w162 and not w1189;
w2933 <= not w2931 and not w2932;
w2934 <= w108 and not w1298;
w2935 <= w215 and not w1225;
w2936 <= not w2934 and not w2935;
w2937 <= w2933 and w2936;
w2938 <= shift(6) and not w2937;
w2939 <= not w2930 and not w2938;
w2940 <= w162 and not w1494;
w2941 <= w55 and not w1475;
w2942 <= not w2940 and not w2941;
w2943 <= w215 and not w1511;
w2944 <= w108 and not w1519;
w2945 <= not w2943 and not w2944;
w2946 <= w2942 and w2945;
w2947 <= not shift(6) and not w2946;
w2948 <= w108 and not w1458;
w2949 <= w215 and not w1466;
w2950 <= not w2948 and not w2949;
w2951 <= w162 and not w1483;
w2952 <= w55 and not w1502;
w2953 <= not w2951 and not w2952;
w2954 <= w2950 and w2953;
w2955 <= shift(6) and not w2954;
w2956 <= not w2947 and not w2955;
w2957 <= w162 and not w1567;
w2958 <= w55 and not w1548;
w2959 <= not w2957 and not w2958;
w2960 <= w215 and not w1584;
w2961 <= w108 and not w1592;
w2962 <= not w2960 and not w2961;
w2963 <= w2959 and w2962;
w2964 <= not shift(6) and not w2963;
w2965 <= w108 and not w1531;
w2966 <= w215 and not w1539;
w2967 <= not w2965 and not w2966;
w2968 <= w162 and not w1556;
w2969 <= w55 and not w1575;
w2970 <= not w2968 and not w2969;
w2971 <= w2967 and w2970;
w2972 <= shift(6) and not w2971;
w2973 <= not w2964 and not w2972;
w2974 <= w162 and not w1640;
w2975 <= w55 and not w1621;
w2976 <= not w2974 and not w2975;
w2977 <= w215 and not w1657;
w2978 <= w108 and not w1665;
w2979 <= not w2977 and not w2978;
w2980 <= w2976 and w2979;
w2981 <= not shift(6) and not w2980;
w2982 <= w108 and not w1604;
w2983 <= w215 and not w1612;
w2984 <= not w2982 and not w2983;
w2985 <= w162 and not w1629;
w2986 <= w55 and not w1648;
w2987 <= not w2985 and not w2986;
w2988 <= w2984 and w2987;
w2989 <= shift(6) and not w2988;
w2990 <= not w2981 and not w2989;
w2991 <= w162 and not w1713;
w2992 <= w108 and not w1738;
w2993 <= not w2991 and not w2992;
w2994 <= w55 and not w1694;
w2995 <= w215 and not w1730;
w2996 <= not w2994 and not w2995;
w2997 <= w2993 and w2996;
w2998 <= not shift(6) and not w2997;
w2999 <= w55 and not w1721;
w3000 <= w108 and not w1677;
w3001 <= not w2999 and not w3000;
w3002 <= w162 and not w1702;
w3003 <= w215 and not w1685;
w3004 <= not w3002 and not w3003;
w3005 <= w3001 and w3004;
w3006 <= shift(6) and not w3005;
w3007 <= not w2998 and not w3006;
w3008 <= w162 and not w1786;
w3009 <= w108 and not w1811;
w3010 <= not w3008 and not w3009;
w3011 <= w55 and not w1767;
w3012 <= w215 and not w1803;
w3013 <= not w3011 and not w3012;
w3014 <= w3010 and w3013;
w3015 <= not shift(6) and not w3014;
w3016 <= w55 and not w1794;
w3017 <= w108 and not w1750;
w3018 <= not w3016 and not w3017;
w3019 <= w162 and not w1775;
w3020 <= w215 and not w1758;
w3021 <= not w3019 and not w3020;
w3022 <= w3018 and w3021;
w3023 <= shift(6) and not w3022;
w3024 <= not w3015 and not w3023;
w3025 <= w162 and not w1859;
w3026 <= w108 and not w1884;
w3027 <= not w3025 and not w3026;
w3028 <= w55 and not w1840;
w3029 <= w215 and not w1876;
w3030 <= not w3028 and not w3029;
w3031 <= w3027 and w3030;
w3032 <= not shift(6) and not w3031;
w3033 <= w55 and not w1867;
w3034 <= w108 and not w1823;
w3035 <= not w3033 and not w3034;
w3036 <= w162 and not w1848;
w3037 <= w215 and not w1831;
w3038 <= not w3036 and not w3037;
w3039 <= w3035 and w3038;
w3040 <= shift(6) and not w3039;
w3041 <= not w3032 and not w3040;
w3042 <= w162 and not w1932;
w3043 <= w55 and not w1913;
w3044 <= not w3042 and not w3043;
w3045 <= w215 and not w1949;
w3046 <= w108 and not w1957;
w3047 <= not w3045 and not w3046;
w3048 <= w3044 and w3047;
w3049 <= not shift(6) and not w3048;
w3050 <= w55 and not w1940;
w3051 <= w108 and not w1896;
w3052 <= not w3050 and not w3051;
w3053 <= w162 and not w1921;
w3054 <= w215 and not w1904;
w3055 <= not w3053 and not w3054;
w3056 <= w3052 and w3055;
w3057 <= shift(6) and not w3056;
w3058 <= not w3049 and not w3057;
w3059 <= w162 and not w2005;
w3060 <= w55 and not w1986;
w3061 <= not w3059 and not w3060;
w3062 <= w215 and not w2022;
w3063 <= w108 and not w2030;
w3064 <= not w3062 and not w3063;
w3065 <= w3061 and w3064;
w3066 <= not shift(6) and not w3065;
w3067 <= w55 and not w2013;
w3068 <= w108 and not w1969;
w3069 <= not w3067 and not w3068;
w3070 <= w162 and not w1994;
w3071 <= w215 and not w1977;
w3072 <= not w3070 and not w3071;
w3073 <= w3069 and w3072;
w3074 <= shift(6) and not w3073;
w3075 <= not w3066 and not w3074;
w3076 <= w162 and not w2078;
w3077 <= w55 and not w2059;
w3078 <= not w3076 and not w3077;
w3079 <= w215 and not w2095;
w3080 <= w108 and not w2103;
w3081 <= not w3079 and not w3080;
w3082 <= w3078 and w3081;
w3083 <= not shift(6) and not w3082;
w3084 <= w55 and not w2086;
w3085 <= w108 and not w2042;
w3086 <= not w3084 and not w3085;
w3087 <= w162 and not w2067;
w3088 <= w215 and not w2050;
w3089 <= not w3087 and not w3088;
w3090 <= w3086 and w3089;
w3091 <= shift(6) and not w3090;
w3092 <= not w3083 and not w3091;
w3093 <= w162 and not w2151;
w3094 <= w55 and not w2132;
w3095 <= not w3093 and not w3094;
w3096 <= w215 and not w2168;
w3097 <= w108 and not w2176;
w3098 <= not w3096 and not w3097;
w3099 <= w3095 and w3098;
w3100 <= not shift(6) and not w3099;
w3101 <= w55 and not w2159;
w3102 <= w108 and not w2115;
w3103 <= not w3101 and not w3102;
w3104 <= w162 and not w2140;
w3105 <= w215 and not w2123;
w3106 <= not w3104 and not w3105;
w3107 <= w3103 and w3106;
w3108 <= shift(6) and not w3107;
w3109 <= not w3100 and not w3108;
w3110 <= w162 and not w2224;
w3111 <= w55 and not w2205;
w3112 <= not w3110 and not w3111;
w3113 <= w215 and not w2241;
w3114 <= w108 and not w2249;
w3115 <= not w3113 and not w3114;
w3116 <= w3112 and w3115;
w3117 <= not shift(6) and not w3116;
w3118 <= w55 and not w2232;
w3119 <= w108 and not w2188;
w3120 <= not w3118 and not w3119;
w3121 <= w162 and not w2213;
w3122 <= w215 and not w2196;
w3123 <= not w3121 and not w3122;
w3124 <= w3120 and w3123;
w3125 <= shift(6) and not w3124;
w3126 <= not w3117 and not w3125;
w3127 <= w162 and not w2297;
w3128 <= w55 and not w2278;
w3129 <= not w3127 and not w3128;
w3130 <= w215 and not w2314;
w3131 <= w108 and not w2322;
w3132 <= not w3130 and not w3131;
w3133 <= w3129 and w3132;
w3134 <= not shift(6) and not w3133;
w3135 <= w55 and not w2305;
w3136 <= w108 and not w2261;
w3137 <= not w3135 and not w3136;
w3138 <= w162 and not w2286;
w3139 <= w215 and not w2269;
w3140 <= not w3138 and not w3139;
w3141 <= w3137 and w3140;
w3142 <= shift(6) and not w3141;
w3143 <= not w3134 and not w3142;
w3144 <= not shift(6) and not w430;
w3145 <= shift(6) and not w218;
w3146 <= not w3144 and not w3145;
w3147 <= not shift(6) and not w855;
w3148 <= shift(6) and not w643;
w3149 <= not w3147 and not w3148;
w3150 <= not shift(6) and not w1152;
w3151 <= shift(6) and not w1004;
w3152 <= not w3150 and not w3151;
w3153 <= not shift(6) and not w1449;
w3154 <= shift(6) and not w1301;
w3155 <= not w3153 and not w3154;
w3156 <= not shift(6) and not w1522;
w3157 <= shift(6) and not w1486;
w3158 <= not w3156 and not w3157;
w3159 <= not shift(6) and not w1595;
w3160 <= shift(6) and not w1559;
w3161 <= not w3159 and not w3160;
w3162 <= not shift(6) and not w1668;
w3163 <= shift(6) and not w1632;
w3164 <= not w3162 and not w3163;
w3165 <= not shift(6) and not w1741;
w3166 <= shift(6) and not w1705;
w3167 <= not w3165 and not w3166;
w3168 <= not shift(6) and not w1814;
w3169 <= shift(6) and not w1778;
w3170 <= not w3168 and not w3169;
w3171 <= not shift(6) and not w1887;
w3172 <= shift(6) and not w1851;
w3173 <= not w3171 and not w3172;
w3174 <= not shift(6) and not w1960;
w3175 <= shift(6) and not w1924;
w3176 <= not w3174 and not w3175;
w3177 <= not shift(6) and not w2033;
w3178 <= shift(6) and not w1997;
w3179 <= not w3177 and not w3178;
w3180 <= not shift(6) and not w2106;
w3181 <= shift(6) and not w2070;
w3182 <= not w3180 and not w3181;
w3183 <= not shift(6) and not w2179;
w3184 <= shift(6) and not w2143;
w3185 <= not w3183 and not w3184;
w3186 <= not shift(6) and not w2252;
w3187 <= shift(6) and not w2216;
w3188 <= not w3186 and not w3187;
w3189 <= not shift(6) and not w2325;
w3190 <= shift(6) and not w2289;
w3191 <= not w3189 and not w3190;
w3192 <= not shift(6) and not w2342;
w3193 <= shift(6) and not w2334;
w3194 <= not w3192 and not w3193;
w3195 <= not shift(6) and not w2359;
w3196 <= shift(6) and not w2351;
w3197 <= not w3195 and not w3196;
w3198 <= not shift(6) and not w2376;
w3199 <= shift(6) and not w2368;
w3200 <= not w3198 and not w3199;
w3201 <= not shift(6) and not w2393;
w3202 <= shift(6) and not w2385;
w3203 <= not w3201 and not w3202;
w3204 <= not shift(6) and not w2410;
w3205 <= shift(6) and not w2402;
w3206 <= not w3204 and not w3205;
w3207 <= not shift(6) and not w2427;
w3208 <= shift(6) and not w2419;
w3209 <= not w3207 and not w3208;
w3210 <= not shift(6) and not w2444;
w3211 <= shift(6) and not w2436;
w3212 <= not w3210 and not w3211;
w3213 <= not shift(6) and not w2461;
w3214 <= shift(6) and not w2453;
w3215 <= not w3213 and not w3214;
w3216 <= not shift(6) and not w2478;
w3217 <= shift(6) and not w2470;
w3218 <= not w3216 and not w3217;
w3219 <= not shift(6) and not w2495;
w3220 <= shift(6) and not w2487;
w3221 <= not w3219 and not w3220;
w3222 <= not shift(6) and not w2512;
w3223 <= shift(6) and not w2504;
w3224 <= not w3222 and not w3223;
w3225 <= not shift(6) and not w2529;
w3226 <= shift(6) and not w2521;
w3227 <= not w3225 and not w3226;
w3228 <= not shift(6) and not w2546;
w3229 <= shift(6) and not w2538;
w3230 <= not w3228 and not w3229;
w3231 <= not shift(6) and not w2563;
w3232 <= shift(6) and not w2555;
w3233 <= not w3231 and not w3232;
w3234 <= not shift(6) and not w2580;
w3235 <= shift(6) and not w2572;
w3236 <= not w3234 and not w3235;
w3237 <= not shift(6) and not w2597;
w3238 <= shift(6) and not w2589;
w3239 <= not w3237 and not w3238;
w3240 <= not shift(6) and not w2614;
w3241 <= shift(6) and not w2606;
w3242 <= not w3240 and not w3241;
w3243 <= not shift(6) and not w2631;
w3244 <= shift(6) and not w2623;
w3245 <= not w3243 and not w3244;
w3246 <= not shift(6) and not w2648;
w3247 <= shift(6) and not w2640;
w3248 <= not w3246 and not w3247;
w3249 <= not shift(6) and not w2665;
w3250 <= shift(6) and not w2657;
w3251 <= not w3249 and not w3250;
w3252 <= not shift(6) and not w2682;
w3253 <= shift(6) and not w2674;
w3254 <= not w3252 and not w3253;
w3255 <= not shift(6) and not w2699;
w3256 <= shift(6) and not w2691;
w3257 <= not w3255 and not w3256;
w3258 <= not shift(6) and not w2716;
w3259 <= shift(6) and not w2708;
w3260 <= not w3258 and not w3259;
w3261 <= not shift(6) and not w2733;
w3262 <= shift(6) and not w2725;
w3263 <= not w3261 and not w3262;
w3264 <= not shift(6) and not w2750;
w3265 <= shift(6) and not w2742;
w3266 <= not w3264 and not w3265;
w3267 <= not shift(6) and not w2767;
w3268 <= shift(6) and not w2759;
w3269 <= not w3267 and not w3268;
w3270 <= not shift(6) and not w2784;
w3271 <= shift(6) and not w2776;
w3272 <= not w3270 and not w3271;
w3273 <= not shift(6) and not w2801;
w3274 <= shift(6) and not w2793;
w3275 <= not w3273 and not w3274;
w3276 <= not shift(6) and not w2818;
w3277 <= shift(6) and not w2810;
w3278 <= not w3276 and not w3277;
w3279 <= not shift(6) and not w2835;
w3280 <= shift(6) and not w2827;
w3281 <= not w3279 and not w3280;
w3282 <= not shift(6) and not w2852;
w3283 <= shift(6) and not w2844;
w3284 <= not w3282 and not w3283;
w3285 <= not shift(6) and not w2869;
w3286 <= shift(6) and not w2861;
w3287 <= not w3285 and not w3286;
w3288 <= not shift(6) and not w2886;
w3289 <= shift(6) and not w2878;
w3290 <= not w3288 and not w3289;
w3291 <= not shift(6) and not w2903;
w3292 <= shift(6) and not w2895;
w3293 <= not w3291 and not w3292;
w3294 <= not shift(6) and not w2920;
w3295 <= shift(6) and not w2912;
w3296 <= not w3294 and not w3295;
w3297 <= not shift(6) and not w2937;
w3298 <= shift(6) and not w2929;
w3299 <= not w3297 and not w3298;
w3300 <= not shift(6) and not w2954;
w3301 <= shift(6) and not w2946;
w3302 <= not w3300 and not w3301;
w3303 <= not shift(6) and not w2971;
w3304 <= shift(6) and not w2963;
w3305 <= not w3303 and not w3304;
w3306 <= not shift(6) and not w2988;
w3307 <= shift(6) and not w2980;
w3308 <= not w3306 and not w3307;
w3309 <= not shift(6) and not w3005;
w3310 <= shift(6) and not w2997;
w3311 <= not w3309 and not w3310;
w3312 <= not shift(6) and not w3022;
w3313 <= shift(6) and not w3014;
w3314 <= not w3312 and not w3313;
w3315 <= not shift(6) and not w3039;
w3316 <= shift(6) and not w3031;
w3317 <= not w3315 and not w3316;
w3318 <= not shift(6) and not w3056;
w3319 <= shift(6) and not w3048;
w3320 <= not w3318 and not w3319;
w3321 <= not shift(6) and not w3073;
w3322 <= shift(6) and not w3065;
w3323 <= not w3321 and not w3322;
w3324 <= not shift(6) and not w3090;
w3325 <= shift(6) and not w3082;
w3326 <= not w3324 and not w3325;
w3327 <= not shift(6) and not w3107;
w3328 <= shift(6) and not w3099;
w3329 <= not w3327 and not w3328;
w3330 <= not shift(6) and not w3124;
w3331 <= shift(6) and not w3116;
w3332 <= not w3330 and not w3331;
w3333 <= not shift(6) and not w3141;
w3334 <= shift(6) and not w3133;
w3335 <= not w3333 and not w3334;
one <= '1';
result(0) <= not w432;-- level 12
result(1) <= not w857;-- level 12
result(2) <= not w1154;-- level 12
result(3) <= not w1451;-- level 12
result(4) <= not w1524;-- level 12
result(5) <= not w1597;-- level 12
result(6) <= not w1670;-- level 12
result(7) <= not w1743;-- level 12
result(8) <= not w1816;-- level 12
result(9) <= not w1889;-- level 12
result(10) <= not w1962;-- level 12
result(11) <= not w2035;-- level 12
result(12) <= not w2108;-- level 12
result(13) <= not w2181;-- level 12
result(14) <= not w2254;-- level 12
result(15) <= not w2327;-- level 12
result(16) <= not w2344;-- level 12
result(17) <= not w2361;-- level 12
result(18) <= not w2378;-- level 12
result(19) <= not w2395;-- level 12
result(20) <= not w2412;-- level 12
result(21) <= not w2429;-- level 12
result(22) <= not w2446;-- level 12
result(23) <= not w2463;-- level 12
result(24) <= not w2480;-- level 12
result(25) <= not w2497;-- level 12
result(26) <= not w2514;-- level 12
result(27) <= not w2531;-- level 12
result(28) <= not w2548;-- level 12
result(29) <= not w2565;-- level 12
result(30) <= not w2582;-- level 12
result(31) <= not w2599;-- level 12
result(32) <= not w2616;-- level 12
result(33) <= not w2633;-- level 12
result(34) <= not w2650;-- level 12
result(35) <= not w2667;-- level 12
result(36) <= not w2684;-- level 12
result(37) <= not w2701;-- level 12
result(38) <= not w2718;-- level 12
result(39) <= not w2735;-- level 12
result(40) <= not w2752;-- level 12
result(41) <= not w2769;-- level 12
result(42) <= not w2786;-- level 12
result(43) <= not w2803;-- level 12
result(44) <= not w2820;-- level 12
result(45) <= not w2837;-- level 12
result(46) <= not w2854;-- level 12
result(47) <= not w2871;-- level 12
result(48) <= not w2888;-- level 12
result(49) <= not w2905;-- level 12
result(50) <= not w2922;-- level 12
result(51) <= not w2939;-- level 12
result(52) <= not w2956;-- level 12
result(53) <= not w2973;-- level 12
result(54) <= not w2990;-- level 12
result(55) <= not w3007;-- level 12
result(56) <= not w3024;-- level 12
result(57) <= not w3041;-- level 12
result(58) <= not w3058;-- level 12
result(59) <= not w3075;-- level 12
result(60) <= not w3092;-- level 12
result(61) <= not w3109;-- level 12
result(62) <= not w3126;-- level 12
result(63) <= not w3143;-- level 12
result(64) <= not w3146;-- level 12
result(65) <= not w3149;-- level 12
result(66) <= not w3152;-- level 12
result(67) <= not w3155;-- level 12
result(68) <= not w3158;-- level 12
result(69) <= not w3161;-- level 12
result(70) <= not w3164;-- level 12
result(71) <= not w3167;-- level 12
result(72) <= not w3170;-- level 12
result(73) <= not w3173;-- level 12
result(74) <= not w3176;-- level 12
result(75) <= not w3179;-- level 12
result(76) <= not w3182;-- level 12
result(77) <= not w3185;-- level 12
result(78) <= not w3188;-- level 12
result(79) <= not w3191;-- level 12
result(80) <= not w3194;-- level 12
result(81) <= not w3197;-- level 12
result(82) <= not w3200;-- level 12
result(83) <= not w3203;-- level 12
result(84) <= not w3206;-- level 12
result(85) <= not w3209;-- level 12
result(86) <= not w3212;-- level 12
result(87) <= not w3215;-- level 12
result(88) <= not w3218;-- level 12
result(89) <= not w3221;-- level 12
result(90) <= not w3224;-- level 12
result(91) <= not w3227;-- level 12
result(92) <= not w3230;-- level 12
result(93) <= not w3233;-- level 12
result(94) <= not w3236;-- level 12
result(95) <= not w3239;-- level 12
result(96) <= not w3242;-- level 12
result(97) <= not w3245;-- level 12
result(98) <= not w3248;-- level 12
result(99) <= not w3251;-- level 12
result(100) <= not w3254;-- level 12
result(101) <= not w3257;-- level 12
result(102) <= not w3260;-- level 12
result(103) <= not w3263;-- level 12
result(104) <= not w3266;-- level 12
result(105) <= not w3269;-- level 12
result(106) <= not w3272;-- level 12
result(107) <= not w3275;-- level 12
result(108) <= not w3278;-- level 12
result(109) <= not w3281;-- level 12
result(110) <= not w3284;-- level 12
result(111) <= not w3287;-- level 12
result(112) <= not w3290;-- level 12
result(113) <= not w3293;-- level 12
result(114) <= not w3296;-- level 12
result(115) <= not w3299;-- level 12
result(116) <= not w3302;-- level 12
result(117) <= not w3305;-- level 12
result(118) <= not w3308;-- level 12
result(119) <= not w3311;-- level 12
result(120) <= not w3314;-- level 12
result(121) <= not w3317;-- level 12
result(122) <= not w3320;-- level 12
result(123) <= not w3323;-- level 12
result(124) <= not w3326;-- level 12
result(125) <= not w3329;-- level 12
result(126) <= not w3332;-- level 12
result(127) <= not w3335;-- level 12
end Behavioral;