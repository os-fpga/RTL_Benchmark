//-----------------------------------------------------------------------------
//	RapidSilicon
//	Author:	Michael Wood
//	Date:	3/9/2022
//-----------------------------------------------------------------------------
module memss
	#(
	parameter ADDR_WIDTH = 32,
	parameter SRAM_DWIDTH = 32,
	parameter DDR_DWIDTH = 128,
	parameter SRAM_SWIDTH = (SRAM_DWIDTH/8),
	parameter DDR_SWIDTH = (DDR_DWIDTH/8))
	(
	input				ddr_sys_clk,
	input				ddr_phy_clk,
	input				ddr_sys_resetn,
	input				sram_sys_clk,
	input				sram_sys_resetn,
	input 				ddr0_aclk,
	input 				ddr1_aclk,
	input 				ddr2_aclk,
	input 				ddr3_aclk,
	input 				sramb0_aclk,
	input 				sramb1_aclk,
	input 				sramb2_aclk,
	input 				sramb3_aclk,
	input 				cntl_aclk,
	input 				ddr0_aresetn,
	input 				ddr1_aresetn,
	input 				ddr2_aresetn,
	input 				ddr3_aresetn,
	input 				sramb0_aresetn,
	input 				sramb1_aresetn,
	input 				sramb2_aresetn,
	input 				sramb3_aresetn,
	input 				cntl_aresetn,
	input 				ddr0_awvalid,
	output 				ddr0_awready, 
	input 	[ADDR_WIDTH-1:0] 	ddr0_awaddr, 
	input 	[ 2:0] 			ddr0_awsize, 
	input 	[ 1:0]			ddr0_awburst,
	input 	[ 3:0]			ddr0_awcache, 
	input 	[ 2:0]			ddr0_awprot,
	input 				ddr0_awlock,
	input 	[ 3:0]			ddr0_awqos,
 	input 	[ 3:0]			ddr0_awid, 	
	input 	[ 3:0]			ddr0_awlen, 
	input 				ddr0_wvalid, 
	output 				ddr0_wready,
	input 				ddr0_wlast, 	
	input 	[DDR_DWIDTH-1:0]	ddr0_wdata, 
	input 	[DDR_SWIDTH-1:0]	ddr0_wstrb, 
	output 				ddr0_bvalid, 
	input 				ddr0_bready, 
	output 	[ 1:0]			ddr0_bresp, 
	output 	[ 3:0]			ddr0_bid, 	
	input 				ddr0_arvalid, 
	output 				ddr0_arready, 
	input 	[ADDR_WIDTH-1:0]	ddr0_araddr, 
	input 	[ 2:0]			ddr0_arsize, 
	input 	[ 1:0]			ddr0_arburst,
	input 	[ 3:0]			ddr0_arcache, 
	input 	[ 2:0]			ddr0_arprot, 
	input 				ddr0_arlock,
	input 	[ 3:0]			ddr0_arqos,
	input 	[ 3:0]			ddr0_arid, 
	input 	[ 3:0]			ddr0_arlen, 
	output 				ddr0_rvalid, 
	input 				ddr0_rready,
	output 				ddr0_rlast, 
	output 	[DDR_DWIDTH-1:0]	ddr0_rdata, 
	output 	[ 1:0]			ddr0_rresp, 
	output  [ 3:0]			ddr0_rid,
	input 				ddr1_awvalid,
	output 				ddr1_awready, 
	input 	[ADDR_WIDTH-1:0] 	ddr1_awaddr, 
	input 	[ 2:0] 			ddr1_awsize, 
	input 	[ 1:0]			ddr1_awburst,
	input 	[ 3:0]			ddr1_awcache, 
	input 	[ 2:0]			ddr1_awprot,
	input 				ddr1_awlock,
	input 	[ 3:0]			ddr1_awqos,
 	input 	[ 3:0]			ddr1_awid, 	
	input 	[ 3:0]			ddr1_awlen, 
	input 				ddr1_wvalid, 
	output 				ddr1_wready,
	input 				ddr1_wlast, 	
	input 	[DDR_DWIDTH-1:0]	ddr1_wdata, 
	input 	[DDR_SWIDTH-1:0]	ddr1_wstrb, 
	output 				ddr1_bvalid, 
	input 				ddr1_bready, 
	output 	[ 1:0]			ddr1_bresp, 
	output 	[ 3:0]			ddr1_bid, 	
	input 				ddr1_arvalid, 
	output 				ddr1_arready, 
	input 	[ADDR_WIDTH-1:0]	ddr1_araddr, 
	input 	[ 2:0]			ddr1_arsize, 
	input 	[ 1:0]			ddr1_arburst,
	input 	[ 3:0]			ddr1_arcache, 
	input 	[ 2:0]			ddr1_arprot, 
	input 				ddr1_arlock,
	input 	[ 3:0]			ddr1_arqos,
	input 	[ 3:0]			ddr1_arid, 
	input 	[ 3:0]			ddr1_arlen, 
	output 				ddr1_rvalid, 
	input 				ddr1_rready,
	output 				ddr1_rlast, 
	output 	[DDR_DWIDTH-1:0]	ddr1_rdata, 
	output  [ 1:0]			ddr1_rresp, 
	output 	[ 3:0]			ddr1_rid,
	input 				ddr2_awvalid,
	output 				ddr2_awready, 
	input 	[ADDR_WIDTH-1:0] 	ddr2_awaddr, 
	input 	[ 2:0] 			ddr2_awsize, 
	input 	[ 1:0]			ddr2_awburst,
	input 	[ 3:0]			ddr2_awcache, 
	input 	[ 2:0]			ddr2_awprot,
	input 				ddr2_awlock,
	input 	[ 3:0]			ddr2_awqos,
 	input 	[ 3:0]			ddr2_awid, 	
	input 	[ 3:0]			ddr2_awlen, 
	input 				ddr2_wvalid, 
	output 				ddr2_wready,
	input 				ddr2_wlast, 	
	input 	[DDR_DWIDTH-1:0]	ddr2_wdata, 
	input 	[DDR_SWIDTH-1:0]	ddr2_wstrb, 
	output 				ddr2_bvalid, 
	input 				ddr2_bready, 
	output 	[ 1:0]			ddr2_bresp, 
	output 	[ 3:0]			ddr2_bid, 	
	input 				ddr2_arvalid, 
	output 				ddr2_arready, 
	input 	[ADDR_WIDTH-1:0]	ddr2_araddr, 
	input 	[ 2:0]			ddr2_arsize, 
	input 	[ 1:0]			ddr2_arburst,
	input 	[ 3:0]			ddr2_arcache, 
	input 	[ 2:0]			ddr2_arprot, 
	input 				ddr2_arlock,
	input 	[ 3:0]			ddr2_arqos,
	input 	[ 3:0]			ddr2_arid, 
	input 	[ 3:0]			ddr2_arlen, 
	output 				ddr2_rvalid, 
	input 				ddr2_rready,
	output 				ddr2_rlast, 
	output 	[DDR_DWIDTH-1:0]	ddr2_rdata, 
	output 	[ 1:0]			ddr2_rresp, 
	output 	[ 3:0]			ddr2_rid,
	input 				ddr3_awvalid,
	output 				ddr3_awready, 
	input 	[ADDR_WIDTH-1:0] 	ddr3_awaddr, 
	input 	[ 2:0] 			ddr3_awsize, 
	input 	[ 1:0]			ddr3_awburst,
	input 	[ 3:0]			ddr3_awcache, 
	input 	[ 2:0]			ddr3_awprot,
	input 				ddr3_awlock,
	input 	[ 3:0]			ddr3_awqos,
 	input 	[ 3:0]			ddr3_awid, 	
	input 	[ 3:0]			ddr3_awlen, 
	input 				ddr3_wvalid, 
	output 				ddr3_wready,
	input 				ddr3_wlast, 	
	input 	[DDR_DWIDTH-1:0]	ddr3_wdata, 
	input 	[DDR_SWIDTH-1:0]	ddr3_wstrb, 
	output 				ddr3_bvalid, 
	input 				ddr3_bready, 
	output 	[ 1:0]			ddr3_bresp, 
	output 	[ 3:0]			ddr3_bid, 	
	input 				ddr3_arvalid, 
	output 				ddr3_arready, 
	input 	[ADDR_WIDTH-1:0]	ddr3_araddr, 
	input 	[ 2:0]			ddr3_arsize, 
	input 	[ 1:0]			ddr3_arburst,
	input 	[ 3:0]			ddr3_arcache, 
	input 	[ 2:0]			ddr3_arprot, 
	input 				ddr3_arlock,
	input 	[ 3:0]			ddr3_arqos,
	input 	[ 3:0]			ddr3_arid, 
	input 	[ 3:0]			ddr3_arlen, 
	output 				ddr3_rvalid, 
	input 				ddr3_rready,
	output 				ddr3_rlast, 
	output 	[DDR_DWIDTH-1:0]	ddr3_rdata, 
	output 	[ 1:0]			ddr3_rresp, 
	output 	[ 3:0]			ddr3_rid,
	input 				sramb0_awvalid,
	output 				sramb0_awready, 
	input 	[ADDR_WIDTH-1:0] 	sramb0_awaddr, 
	input 	[ 2:0] 			sramb0_awsize, 
	input 	[ 1:0]			sramb0_awburst,
 	input 	[ 3:0]			sramb0_awid, 	
	input 	[ 3:0]			sramb0_awlen, 
	input 				sramb0_wvalid, 
	output 				sramb0_wready,
	input 				sramb0_wlast, 	
	input 	[SRAM_DWIDTH-1:0]	sramb0_wdata, 
	input 	[SRAM_SWIDTH-1:0]	sramb0_wstrb, 
	input 	[ 3:0]			sramb0_wid, 	
	output 				sramb0_bvalid, 
	input 				sramb0_bready, 
	output 	[ 1:0]			sramb0_bresp, 
	output 	[ 3:0]			sramb0_bid, 	
	input 				sramb0_arvalid, 
	output 				sramb0_arready, 
	input 	[ADDR_WIDTH-1:0]	sramb0_araddr, 
	input 	[ 2:0]			sramb0_arsize, 
	input 	[ 1:0]			sramb0_arburst,
	input 	[ 3:0]			sramb0_arid, 
	input 	[ 3:0]			sramb0_arlen, 
	output 				sramb0_rvalid, 
	input 				sramb0_rready,
	output 				sramb0_rlast, 
	output 	[SRAM_DWIDTH-1:0]	sramb0_rdata, 
	output 	[ 1:0]			sramb0_rresp, 
	output 	[ 3:0]			sramb0_rid,
	input 				sramb1_awvalid,
	output 				sramb1_awready, 
	input 	[ADDR_WIDTH-1:0] 	sramb1_awaddr, 
	input 	[ 2:0] 			sramb1_awsize, 
	input 	[ 1:0]			sramb1_awburst,
 	input 	[ 3:0]			sramb1_awid, 	
	input 	[ 3:0]			sramb1_awlen, 
	input 				sramb1_wvalid, 
	output 				sramb1_wready,
	input 				sramb1_wlast, 	
	input 	[SRAM_DWIDTH-1:0]	sramb1_wdata, 
	input 	[SRAM_SWIDTH-1:0]	sramb1_wstrb, 
	input 	[ 3:0]			sramb1_wid, 	
	output 				sramb1_bvalid, 
	input 				sramb1_bready, 
	output 	[ 1:0]			sramb1_bresp, 
	output 	[ 3:0]			sramb1_bid, 	
	input 				sramb1_arvalid, 
	output 				sramb1_arready, 
	input 	[ADDR_WIDTH-1:0]	sramb1_araddr, 
	input 	[ 2:0]			sramb1_arsize, 
	input 	[ 1:0]			sramb1_arburst,
	input 	[ 3:0]			sramb1_arid, 
	input 	[ 3:0]			sramb1_arlen, 
	output 				sramb1_rvalid, 
	input 				sramb1_rready,
	output 				sramb1_rlast, 
	output 	[SRAM_DWIDTH-1:0]	sramb1_rdata, 
	output 	[ 1:0]			sramb1_rresp, 
	output 	[ 3:0]			sramb1_rid,
	input 				sramb2_awvalid,
	output 				sramb2_awready, 
	input 	[ADDR_WIDTH-1:0] 	sramb2_awaddr, 
	input 	[ 2:0] 			sramb2_awsize, 
	input 	[ 1:0]			sramb2_awburst,
 	input 	[ 3:0]			sramb2_awid, 	
	input 	[ 3:0]			sramb2_awlen, 
	input 				sramb2_wvalid, 
	output 				sramb2_wready,
	input 				sramb2_wlast, 	
	input 	[SRAM_DWIDTH-1:0]	sramb2_wdata, 
	input 	[SRAM_SWIDTH-1:0]	sramb2_wstrb, 
	input 	[ 3:0]			sramb2_wid, 	
	output 				sramb2_bvalid, 
	input 				sramb2_bready, 
	output 	[1:0]			sramb2_bresp, 
	output 	[3:0]			sramb2_bid, 	
	input 				sramb2_arvalid, 
	output 				sramb2_arready, 
	input 	[ADDR_WIDTH-1:0]	sramb2_araddr, 
	input 	[ 2:0]			sramb2_arsize, 
	input 	[ 1:0]			sramb2_arburst,
	input 	[ 3:0]			sramb2_arid, 
	input 	[ 3:0]			sramb2_arlen, 
	output 				sramb2_rvalid, 
	input 				sramb2_rready,
	output 				sramb2_rlast, 
	output 	[SRAM_DWIDTH-1:0]	sramb2_rdata, 
	output 	[ 1:0]			sramb2_rresp, 
	output 	[3:0]			sramb2_rid,
	input 				sramb3_awvalid,
	output 				sramb3_awready, 
	input 	[ADDR_WIDTH-1:0] 	sramb3_awaddr, 
	input 	[ 2:0] 			sramb3_awsize, 
	input 	[ 1:0]			sramb3_awburst,
 	input 	[ 3:0]			sramb3_awid, 	
	input 	[ 3:0]			sramb3_awlen, 
	input 				sramb3_wvalid, 
	output 				sramb3_wready,
	input 				sramb3_wlast, 	
	input 	[SRAM_DWIDTH-1:0]	sramb3_wdata, 
	input 	[SRAM_SWIDTH-1:0]	sramb3_wstrb, 
	input 	[ 3:0]			sramb3_wid, 	
	output 				sramb3_bvalid, 
	input 				sramb3_bready, 
	output 	[ 1:0]			sramb3_bresp, 
	output 	[ 3:0]			sramb3_bid, 	
	input 				sramb3_arvalid, 
	output 				sramb3_arready, 
	input 	[ADDR_WIDTH-1:0]	sramb3_araddr, 
	input 	[ 2:0]			sramb3_arsize, 
	input 	[ 1:0]			sramb3_arburst,
	input 	[ 3:0]			sramb3_arid, 
	input 	[ 3:0]			sramb3_arlen, 
	output 				sramb3_rvalid, 
	input 				sramb3_rready,
	output 				sramb3_rlast, 
	output 	[SRAM_DWIDTH-1:0]	sramb3_rdata, 
	output 	[ 1:0]			sramb3_rresp, 
	output 	[ 3:0]			sramb3_rid,
	output				cntl_arready, 
	output				cntl_awready, 
	output	[ 1:0]			cntl_bresp, 
	output				cntl_bvalid, 
	output	[31:0]			cntl_rdata, 
	output	[ 1:0]			cntl_rresp, 
	output				cntl_rvalid, 
	output				cntl_wready, 
	input	[31:0]			cntl_araddr, 
	input				cntl_arvalid, 
	input	[31:0]			cntl_awaddr, 
	input				cntl_awvalid, 
	input				cntl_bready, 
	input				cntl_rready, 
	input	[31:0]			cntl_wdata, 
	input				cntl_wvalid, 	
	output  [ 1:0]			int_gc_fsm,
	input	[ 3:0]			DTI_EXT_VREF,
	output  [29:0]			PAD_MEM_CTL,
	output 	[ 1:0]			PAD_MEM_CLK,
	output  [ 1:0]			PAD_MEM_CLK_N,
	inout  	[ 3:0]			PAD_MEM_DM,
	inout  	[31:0]			PAD_MEM_DQ,
	inout  	[ 3:0]			PAD_MEM_DQS,
	inout	[ 3:0]			PAD_MEM_DQS_N,
	input	[29:0]			CLOCKDR_CTL,
	input 	[ 1:0]			CLOCKDR_CLK,
	input	[ 3:0]			CLOCKDR_DM,
	input   [31:0]			CLOCKDR_DQ,
	input 	[ 3:0]			CLOCKDR_DQS,
	input	[29:0]			JTAG_SI_CTL,
	input 	[ 1:0]			JTAG_SI_CLK,
	input	[ 3:0]			JTAG_SI_DM,
	input   [31:0]			JTAG_SI_DQ,
	input 	[ 3:0]			JTAG_SI_DQS,
	output	[29:0]			JTAG_SO_CTL,
	output 	[ 1:0]			JTAG_SO_CLK,
	output	[ 3:0]			JTAG_SO_DM,
	output  [31:0]			JTAG_SO_DQ,
	output 	[ 3:0]			JTAG_SO_DQS,
	input	[29:0]			MODE_CTL,
	input 	[ 1:0]			MODE_CLK,
	input	[ 3:0]			MODE_DM,
	input   [31:0]			MODE_DQ,
	input 	[ 3:0]			MODE_DQS,
	input	[ 3:0]			MODE_I_DM,
	input   [31:0]			MODE_I_DQ,
	input 	[ 3:0]			MODE_I_DQS,
	input				PAD_REF,
	input				SE,
	input				SE_CK,
	input	[29:0]			SHIFTDR_CTL,
	input 	[ 1:0]			SHIFTDR_CLK,
	input	[ 3:0]			SHIFTDR_DM,
	input   [31:0]			SHIFTDR_DQ,
	input 	[ 3:0]			SHIFTDR_DQS,
	input	[ 1:0]			SI_CLK,
	input	[29:0]			SI_CTL,
	input	[ 3:0]			SI_DM,
	input   [31:0]			SI_DQ,
	input	[ 3:0]			SI_RD,
	input	[ 3:0]			SI_WR,
	output	[ 1:0]			SO_CLK,
	output	[29:0]			SO_CTL,
	output	[ 3:0]			SO_DM,
	output   [31:0]			SO_DQ,
	output	[ 3:0]			SO_RD,
	output	[ 3:0]			SO_WR,
	input				T_CGCTL_CTL,
	input	[ 3:0]			T_CGCTL_DQ,
	input				T_RCTL_CTL,
	input	[ 3:0]			T_RCTL_DQ,
	input				VDD,
	input				VDDO,
	input				VSS,
	input	[29:0]			UPDATEDR_CTL,
	input 	[ 1:0]			UPDATEDR_CLK,
	input	[ 3:0]			UPDATEDR_DM,
	input   [31:0]			UPDATEDR_DQ,
	input 	[ 3:0]			UPDATEDR_DQS,
	inout				PAD_COMP,
	output 	[ 1:0]			YC_CLK,
	output 	[29:0]			YC_CTL,
	output  [ 3:0]			Y_DM, 
	output  [31:0]			Y_DQ, 
	output  [ 3:0]			Y_DQS, 
	inout				PAD_VREF
);


	wire 	[1023:0] 		ddr_rdata;
	wire 	[  39:0]		ddr_bid;
	wire 	[  39:0]		ddr_rid;
	assign ddr0_rdata = ddr_rdata[127:0];
	assign ddr1_rdata = ddr_rdata[383:256];
	assign ddr2_rdata = ddr_rdata[639:512];
	assign ddr3_rdata = ddr_rdata[895:768];

	assign ddr0_bid	  = ddr_bid[3:0];
	assign ddr1_bid	  = ddr_bid[13:10];
	assign ddr2_bid	  = ddr_bid[23:20];
	assign ddr3_bid	  = ddr_bid[33:30];

	assign ddr0_rid	  = ddr_rid[3:0];
	assign ddr1_rid	  = ddr_rid[13:10];
	assign ddr2_rid	  = ddr_rid[23:20];
	assign ddr3_rid	  = ddr_rid[33:30];
	
	

	/*********** SRAM Subsystem  ***********/	
	sram_ss	sram4b(
		.sram_sys_clk		(sram_sys_clk	),
		.sram_sys_resetn	(sram_sys_resetn),
		.sramb0_aclk		(sramb0_aclk	),
		.sramb0_aresetn		(sramb0_aresetn	),
		.sramb1_aclk		(sramb1_aclk	),
		.sramb1_aresetn		(sramb1_aresetn	),
		.sramb2_aclk		(sramb2_aclk	),
		.sramb2_aresetn		(sramb2_aresetn	),
		.sramb3_aclk		(sramb3_aclk	),
		.sramb3_aresetn		(sramb3_aresetn	),
		.sramb0_awvalid		(sramb0_awvalid	),
		.sramb0_awready 	(sramb0_awready	),
		.sramb0_awaddr 		(sramb0_awaddr 	),
		.sramb0_awsize 		(sramb0_awsize 	),
		.sramb0_awburst		(sramb0_awburst	),
 		.sramb0_awid 		(sramb0_awid 	),
		.sramb0_awlen 		(sramb0_awlen 	),
		.sramb0_wvalid 		(sramb0_wvalid 	),
		.sramb0_wready		(sramb0_wready	),
		.sramb0_wlast 		(sramb0_wlast 	),
		.sramb0_wdata 		(sramb0_wdata 	),
		.sramb0_wstrb 		(sramb0_wstrb 	),
		.sramb0_wid 		(sramb0_wid 	),
		.sramb0_bvalid 		(sramb0_bvalid 	),
		.sramb0_bready 		(sramb0_bready 	),
		.sramb0_bresp 		(sramb0_bresp 	),
		.sramb0_bid 		(sramb0_bid 	),
		.sramb0_arvalid 	(sramb0_arvalid	),
		.sramb0_arready 	(sramb0_arready	),
		.sramb0_araddr 		(sramb0_araddr 	),
		.sramb0_arsize 		(sramb0_arsize 	),
		.sramb0_arburst		(sramb0_arburst	),
		.sramb0_arid 		(sramb0_arid 	),
		.sramb0_arlen 		(sramb0_arlen 	),
		.sramb0_rvalid 		(sramb0_rvalid 	),
		.sramb0_rready		(sramb0_rready	),
		.sramb0_rlast 		(sramb0_rlast 	),
		.sramb0_rdata 		(sramb0_rdata 	),
		.sramb0_rresp 		(sramb0_rresp 	),
		.sramb0_rid		(sramb0_rid	),
		.sramb1_awvalid		(sramb1_awvalid	),
		.sramb1_awready 	(sramb1_awready ),
		.sramb1_awaddr 		(sramb1_awaddr 	),
		.sramb1_awsize 		(sramb1_awsize 	),
		.sramb1_awburst		(sramb1_awburst	),
 		.sramb1_awid 		(sramb1_awid 	),
		.sramb1_awlen 		(sramb1_awlen 	),
		.sramb1_wvalid 		(sramb1_wvalid 	),
		.sramb1_wready		(sramb1_wready	),
		.sramb1_wlast 		(sramb1_wlast 	),
		.sramb1_wdata 		(sramb1_wdata 	),
		.sramb1_wstrb 		(sramb1_wstrb 	),
		.sramb1_wid 		(sramb1_wid 	),
		.sramb1_bvalid 		(sramb1_bvalid 	),
		.sramb1_bready 		(sramb1_bready 	),
		.sramb1_bresp 		(sramb1_bresp 	),
		.sramb1_bid 		(sramb1_bid 	),
		.sramb1_arvalid 	(sramb1_arvalid ),
		.sramb1_arready 	(sramb1_arready ),
		.sramb1_araddr 		(sramb1_araddr 	),
		.sramb1_arsize 		(sramb1_arsize 	),
		.sramb1_arburst		(sramb1_arburst	),
		.sramb1_arid 		(sramb1_arid 	),
		.sramb1_arlen 		(sramb1_arlen 	),
		.sramb1_rvalid 		(sramb1_rvalid 	),
		.sramb1_rready		(sramb1_rready	),
		.sramb1_rlast		(sramb1_rlast	),
		.sramb1_rdata 		(sramb1_rdata 	),
		.sramb1_rresp 		(sramb1_rresp 	),
		.sramb1_rid		(sramb1_rid	),
		.sramb2_awvalid		(sramb2_awvalid	),
		.sramb2_awready 	(sramb2_awready ),
		.sramb2_awaddr 		(sramb2_awaddr 	),
		.sramb2_awsize 		(sramb2_awsize 	),
		.sramb2_awburst		(sramb2_awburst	),
 		.sramb2_awid 		(sramb2_awid 	),
		.sramb2_awlen 		(sramb2_awlen 	),
		.sramb2_wvalid 		(sramb2_wvalid 	),
		.sramb2_wready		(sramb2_wready	),
		.sramb2_wlast 		(sramb2_wlast 	),
		.sramb2_wdata 		(sramb2_wdata 	),
		.sramb2_wstrb 		(sramb2_wstrb 	),
		.sramb2_wid 		(sramb2_wid 	),
		.sramb2_bvalid 		(sramb2_bvalid 	),
		.sramb2_bready 		(sramb2_bready 	),
		.sramb2_bresp 		(sramb2_bresp 	),
		.sramb2_bid 		(sramb2_bid 	),
		.sramb2_arvalid 	(sramb2_arvalid ),
		.sramb2_arready 	(sramb2_arready ),
		.sramb2_araddr 		(sramb2_araddr 	),
		.sramb2_arsize 		(sramb2_arsize 	),
		.sramb2_arburst		(sramb2_arburst	),
		.sramb2_arid 		(sramb2_arid 	),
		.sramb2_arlen 		(sramb2_arlen 	),
		.sramb2_rvalid 		(sramb2_rvalid 	),
		.sramb2_rready		(sramb2_rready	),
		.sramb2_rlast 		(sramb2_rlast 	),
		.sramb2_rdata 		(sramb2_rdata 	),
		.sramb2_rresp 		(sramb2_rresp 	),
		.sramb2_rid		(sramb2_rid	),
		.sramb3_awvalid		(sramb3_awvalid	),
		.sramb3_awready 	(sramb3_awready ),
		.sramb3_awaddr 		(sramb3_awaddr 	),
		.sramb3_awsize 		(sramb3_awsize 	),
		.sramb3_awburst		(sramb3_awburst	),
 		.sramb3_awid 		(sramb3_awid 	),
		.sramb3_awlen 		(sramb3_awlen 	),
		.sramb3_wvalid 		(sramb3_wvalid 	),
		.sramb3_wready		(sramb3_wready	),
		.sramb3_wlast 		(sramb3_wlast 	),
		.sramb3_wdata 		(sramb3_wdata 	),
		.sramb3_wstrb 		(sramb3_wstrb 	),
		.sramb3_wid 		(sramb3_wid 	),
		.sramb3_bvalid 		(sramb3_bvalid 	),
		.sramb3_bready 		(sramb3_bready 	),
		.sramb3_bresp 		(sramb3_bresp 	),
		.sramb3_bid 		(sramb3_bid 	),
		.sramb3_arvalid 	(sramb3_arvalid ),
		.sramb3_arready 	(sramb3_arready ),
		.sramb3_araddr 		(sramb3_araddr 	),
		.sramb3_arsize 		(sramb3_arsize 	),
		.sramb3_arburst		(sramb3_arburst	),
		.sramb3_arid 		(sramb3_arid 	),
		.sramb3_arlen 		(sramb3_arlen 	),
		.sramb3_rvalid 		(sramb3_rvalid 	),
		.sramb3_rready		(sramb3_rready	),
		.sramb3_rlast 		(sramb3_rlast 	),
		.sramb3_rdata 		(sramb3_rdata 	),
		.sramb3_rresp 		(sramb3_rresp 	),
		.sramb3_rid		(sramb3_rid	)
	);

	/*********** DDR Subsystem  ***********/	
	dynamo	ddr_wrapper(
		.CLOCKDR_CLK		(CLOCKDR_CLK),
		.CLOCKDR_CTL		(CLOCKDR_CTL),
		.CLOCKDR_DM		(CLOCKDR_DM),
		.CLOCKDR_DQ		(CLOCKDR_DQ),
		.CLOCKDR_DQS		(CLOCKDR_DQS),
		.COMP_CLOCK		(cntl_aclk),
		.COMP_RST_N		(ddr_sys_resetn),
		.DTI_EXT_VREF		(DTI_EXT_VREF),
		.DTI_MC_CLOCK		(ddr_sys_clk),
		.DTI_PHY_CLOCK		(ddr_phy_clk),
		.DTI_SYS_RESET_N	(ddr_sys_resetn),
		.JTAG_SI_CLK		(JTAG_SI_CLK),
		.JTAG_SI_CTL		(JTAG_SI_CTL),
		.JTAG_SI_DM		(JTAG_SI_DM),
		.JTAG_SI_DQ		(JTAG_SI_DQ),
		.JTAG_SI_DQS		(JTAG_SI_DQS),
		.MODE_CLK		(MODE_CLK),
		.MODE_CTL		(MODE_CTL),
		.MODE_DM		(MODE_DM),
		.MODE_DQ		(MODE_DQ),
		.MODE_DQS		(MODE_DQS),
		.MODE_I_DM		(MODE_I_DM),
		.MODE_I_DQ		(MODE_I_DQ),
		.MODE_I_DQS		(MODE_I_DQS),
		.PAD_REF		(PAD_REF),
		.SE			(SE),
		.SE_CK			(SE_CK),
		.SHIFTDR_CLK		(SHIFTDR_CLK),
		.SHIFTDR_CTL		(SHIFTDR_CTL),
		.SHIFTDR_DM		(SHIFTDR_DM),
		.SHIFTDR_DQ		(SHIFTDR_DQ),
		.SHIFTDR_DQS		(SHIFTDR_DQS),
		.SI_CLK			(SI_CLK),
		.SI_CTL			(SI_CTL),
		.SI_DM			(SI_DM),
		.SI_DQ			(SI_DQ),
		.SI_RD			(SI_RD),
		.SI_WR			(SI_WR),
		.T_CGCTL_CTL		(T_CGCTL_CTL),
		.T_CGCTL_DQ		(T_CGCTL_DQ),
		.T_RCTL_CTL		(T_RCTL_CTL),
		.T_RCTL_DQ		(T_RCTL_DQ),
		.UPDATEDR_CLK		(UPDATEDR_CLK),
		.UPDATEDR_CTL		(UPDATEDR_CTL),
		.UPDATEDR_DM		(UPDATEDR_DM),
		.UPDATEDR_DQ		(UPDATEDR_DQ),
		.UPDATEDR_DQS		(UPDATEDR_DQS),
		.VDD			(VDD),
		.VDDO			(VDDO),
		.VSS			(VSS),
		.int_gc_fsm		(int_gc_fsm),
		.aclk_p 		({ddr3_aclk, ddr2_aclk, ddr1_aclk, ddr0_aclk}			),
		.aresetn_p 		({ddr3_aresetn, ddr2_aresetn, ddr1_aresetn, ddr0_aresetn}	),
		.arvalid_p 		({ddr3_arvalid, ddr2_arvalid, ddr1_arvalid, ddr0_arvalid}	),
		.arready_p		({ddr3_arready, ddr2_arready, ddr1_arready, ddr0_arready}	),
		.araddr_p 		({ddr3_araddr[30:0], ddr2_araddr[30:0], ddr1_araddr[30:0], ddr0_araddr[30:0]}),
		.arsize_p 		({ddr3_arsize, ddr2_arsize, ddr1_arsize, ddr0_arsize}		),
		.arburst_p 		({ddr3_arburst, ddr2_arburst, ddr1_arburst, ddr0_arburst}	),
		.arcache_p 		({ddr3_arcache, ddr2_arcache, ddr1_arcache, ddr0_arcache}	),
		.arprot_p 		({ddr3_arprot, ddr2_arprot, ddr1_arprot, ddr0_arprot}		),
		.arlock_p 		({ddr3_arlock, ddr2_arlock, ddr1_arlock, ddr0_arlock}		),
		.arqos_p 		({ddr3_arqos, ddr2_arqos, ddr1_arqos, ddr0_arqos}		),
		.arid_p 		({6'h0, ddr3_arid, 6'h0, ddr2_arid, 6'h0, ddr1_arid, 6'h0, ddr0_arid}			),
		.arlen_p 		({ddr3_arlen, ddr2_arlen, ddr1_arlen, ddr0_arlen}		),
		.rvalid_p		({ddr3_rvalid, ddr2_rvalid, ddr1_rvalid, ddr0_rvalid}		),
		.rready_p 		({ddr3_rready, ddr2_rready, ddr1_rready, ddr0_rready}		),
		.rlast_p		({ddr3_rlast, ddr2_rlast, ddr1_rlast, ddr0_rlast}		),
		.rdata_p 		(ddr_rdata							),
		.rresp_p		({ddr3_rresp, ddr2_rresp, ddr1_rresp, ddr0_rresp}		),
		.rid_p			(ddr_rid							),
		.awvalid_p 		({ddr3_awvalid, ddr2_awvalid, ddr1_awvalid, ddr0_awvalid}	),
		.awready_p		({ddr3_awready, ddr2_awready, ddr1_awready, ddr0_awready}	),
		.awaddr_p 		({ddr3_awaddr[30:0], ddr2_awaddr[30:0], ddr1_awaddr[30:0], ddr0_awaddr[30:0]}		),
		.awsize_p 		({ddr3_awsize, ddr2_awsize, ddr1_awsize, ddr0_awsize}		),
		.awburst_p 		({ddr3_awburst, ddr2_awburst, ddr1_awburst, ddr0_awburst}	),
		.awcache_p 		({ddr3_awcache, ddr2_awcache, ddr1_awcache, ddr0_awcache}	),
		.awprot_p 		({ddr3_awprot, ddr2_awprot, ddr1_awprot, ddr0_awprot}		),
		.awlock_p 		({ddr3_awlock, ddr2_awlock, ddr1_awlock, ddr0_awlock}		),
		.awqos_p 		({ddr3_awqos, ddr2_awqos, ddr1_awqos, ddr0_awqos}		),
		.awid_p 		({6'h0, ddr3_awid, 6'h0, ddr2_awid, 6'h0, ddr1_awid, 6'h0, ddr0_awid}			),
		.awlen_p 		({ddr3_awlen, ddr2_awlen, ddr1_awlen, ddr0_awlen}		),
		.wvalid_p 		({ddr3_wvalid, ddr2_wvalid, ddr1_wvalid, ddr0_wvalid}		),
		.wready_p		({ddr3_wready, ddr2_wready, ddr1_wready, ddr0_wready}		),
		.wlast_p 		({ddr3_wlast, ddr2_wlast, ddr1_wlast, ddr0_wlast}		),
		.wdata_p 		({128'b0, ddr3_wdata, 128'b0, ddr2_wdata, 128'b0, ddr1_wdata, 128'b0, ddr0_wdata}	),
		.wstrb_p 		({16'h0, ddr3_wstrb, 16'h0, ddr2_wstrb, 16'h0, ddr1_wstrb, 16'h0, ddr0_wstrb}		),
		.bvalid_p		({ddr3_bvalid, ddr2_bvalid, ddr1_bvalid, ddr0_bvalid}		),
		.bready_p 		({ddr3_bready, ddr2_bready, ddr1_bready, ddr0_bready}		),
		.bresp_p		({ddr3_bresp, ddr2_bresp, ddr1_bresp, ddr0_bresp}		),
		.bid_p			(ddr_bid							),
		.axi4lite_clk 		(cntl_aclk							),
		.axi4lite_reset_n 	(cntl_aresetn							),
		.axi4lite_arready	(cntl_arready							),	
		.axi4lite_awready	(cntl_awready							),
		.axi4lite_bresp		(cntl_bresp							),
		.axi4lite_bvalid	(cntl_bvalid							),
		.axi4lite_rdata		(cntl_rdata							),
		.axi4lite_rresp		(cntl_rresp							),
		.axi4lite_rvalid	(cntl_rvalid							),
		.axi4lite_wready	(cntl_wready							),
		.axi4lite_araddr 	(cntl_araddr[11:0]						),
		.axi4lite_arvalid 	(cntl_arvalid							),
		.axi4lite_awaddr 	(cntl_awaddr[11:0]						),
		.axi4lite_awvalid 	(cntl_awvalid							),
		.axi4lite_bready 	(cntl_bready							),
		.axi4lite_rready 	(cntl_rready							),
		.axi4lite_wdata 	(cntl_wdata							),
		.axi4lite_wvalid 	(cntl_wvalid							),
		.JTAG_SO_CLK		(JTAG_SO_CLK),
		.JTAG_SO_CTL		(JTAG_SO_CTL),
		.JTAG_SO_DM		(JTAG_SO_DM),
		.JTAG_SO_DQ		(JTAG_SO_DQ),
		.JTAG_SO_DQS		(JTAG_SO_DQS),
		.PAD_MEM_CLK		(PAD_MEM_CLK),
		.PAD_MEM_CLK_N		(PAD_MEM_CLK_N),
		.PAD_MEM_CTL		(PAD_MEM_CTL),
		.SO_CLK			(SO_CLK),
		.SO_CTL			(SO_CTL),
		.SO_DM			(SO_DM),
		.SO_DQ			(SO_DQ),
		.SO_RD			(SO_RD),
		.SO_WR			(SO_WR),
		.YC_CLK			(YC_CLK),
		.YC_CTL			(YC_CTL),
		.Y_DM			(Y_DM),
		.Y_DQ			(Y_DQ),
		.Y_DQS			(Y_DQS),
		.PAD_COMP		(PAD_COMP),
		.PAD_MEM_DM		(PAD_MEM_DM),
		.PAD_MEM_DQ		(PAD_MEM_DQ),
		.PAD_MEM_DQS		(PAD_MEM_DQS),
		.PAD_MEM_DQS_N		(PAD_MEM_DQS_N),
		.PAD_VREF		(PAD_VREF)
	);
endmodule
