-------------------------------------------------------------------------------
-- $Id: ram_loader-c.vhd,v 1.1 2005-04-10 18:02:32 arniml Exp $
-------------------------------------------------------------------------------

configuration ram_loader_rtl_c0 of ram_loader is

  for rtl
  end for;

end ram_loader_rtl_c0;
