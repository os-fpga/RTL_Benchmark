library ieee;
use ieee.std_logic_1164.all;

entity top is
 port( a, b: in std_logic_vector(127 downto 0);
      f: out std_logic_vector(127 downto 0);
      cOut: out std_logic);
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019: std_logic;

begin

w0 <= a(0) and not b(0);
w1 <= not a(0) and b(0);
w2 <= not w0 and not w1;
w3 <= a(0) and b(0);
w4 <= not a(1) and not b(1);
w5 <= a(1) and b(1);
w6 <= not w4 and not w5;
w7 <= w3 and not w6;
w8 <= not w3 and w6;
w9 <= not w7 and not w8;
w10 <= w3 and not w4;
w11 <= not w5 and not w10;
w12 <= not a(2) and not b(2);
w13 <= a(2) and b(2);
w14 <= not w12 and not w13;
w15 <= w11 and not w14;
w16 <= not w11 and w14;
w17 <= not w15 and not w16;
w18 <= not w11 and not w12;
w19 <= not w13 and not w18;
w20 <= not a(3) and not b(3);
w21 <= a(3) and b(3);
w22 <= not w20 and not w21;
w23 <= w19 and not w22;
w24 <= not w19 and w22;
w25 <= not w23 and not w24;
w26 <= not w19 and not w20;
w27 <= not w21 and not w26;
w28 <= not a(4) and not b(4);
w29 <= a(4) and b(4);
w30 <= not w28 and not w29;
w31 <= w27 and not w30;
w32 <= not w27 and w30;
w33 <= not w31 and not w32;
w34 <= not w27 and not w28;
w35 <= not w29 and not w34;
w36 <= not a(5) and not b(5);
w37 <= a(5) and b(5);
w38 <= not w36 and not w37;
w39 <= w35 and not w38;
w40 <= not w35 and w38;
w41 <= not w39 and not w40;
w42 <= not w35 and not w36;
w43 <= not w37 and not w42;
w44 <= not a(6) and not b(6);
w45 <= a(6) and b(6);
w46 <= not w44 and not w45;
w47 <= w43 and not w46;
w48 <= not w43 and w46;
w49 <= not w47 and not w48;
w50 <= not w43 and not w44;
w51 <= not w45 and not w50;
w52 <= not a(7) and not b(7);
w53 <= a(7) and b(7);
w54 <= not w52 and not w53;
w55 <= w51 and not w54;
w56 <= not w51 and w54;
w57 <= not w55 and not w56;
w58 <= not w51 and not w52;
w59 <= not w53 and not w58;
w60 <= not a(8) and not b(8);
w61 <= a(8) and b(8);
w62 <= not w60 and not w61;
w63 <= w59 and not w62;
w64 <= not w59 and w62;
w65 <= not w63 and not w64;
w66 <= not w59 and not w60;
w67 <= not w61 and not w66;
w68 <= not a(9) and not b(9);
w69 <= a(9) and b(9);
w70 <= not w68 and not w69;
w71 <= w67 and not w70;
w72 <= not w67 and w70;
w73 <= not w71 and not w72;
w74 <= not w67 and not w68;
w75 <= not w69 and not w74;
w76 <= not a(10) and not b(10);
w77 <= a(10) and b(10);
w78 <= not w76 and not w77;
w79 <= w75 and not w78;
w80 <= not w75 and w78;
w81 <= not w79 and not w80;
w82 <= not w75 and not w76;
w83 <= not w77 and not w82;
w84 <= not a(11) and not b(11);
w85 <= a(11) and b(11);
w86 <= not w84 and not w85;
w87 <= w83 and not w86;
w88 <= not w83 and w86;
w89 <= not w87 and not w88;
w90 <= not w83 and not w84;
w91 <= not w85 and not w90;
w92 <= not a(12) and not b(12);
w93 <= a(12) and b(12);
w94 <= not w92 and not w93;
w95 <= w91 and not w94;
w96 <= not w91 and w94;
w97 <= not w95 and not w96;
w98 <= not w91 and not w92;
w99 <= not w93 and not w98;
w100 <= not a(13) and not b(13);
w101 <= a(13) and b(13);
w102 <= not w100 and not w101;
w103 <= w99 and not w102;
w104 <= not w99 and w102;
w105 <= not w103 and not w104;
w106 <= not w99 and not w100;
w107 <= not w101 and not w106;
w108 <= not a(14) and not b(14);
w109 <= a(14) and b(14);
w110 <= not w108 and not w109;
w111 <= w107 and not w110;
w112 <= not w107 and w110;
w113 <= not w111 and not w112;
w114 <= not w107 and not w108;
w115 <= not w109 and not w114;
w116 <= not a(15) and not b(15);
w117 <= a(15) and b(15);
w118 <= not w116 and not w117;
w119 <= w115 and not w118;
w120 <= not w115 and w118;
w121 <= not w119 and not w120;
w122 <= not w115 and not w116;
w123 <= not w117 and not w122;
w124 <= not a(16) and not b(16);
w125 <= a(16) and b(16);
w126 <= not w124 and not w125;
w127 <= w123 and not w126;
w128 <= not w123 and w126;
w129 <= not w127 and not w128;
w130 <= not w123 and not w124;
w131 <= not w125 and not w130;
w132 <= not a(17) and not b(17);
w133 <= a(17) and b(17);
w134 <= not w132 and not w133;
w135 <= w131 and not w134;
w136 <= not w131 and w134;
w137 <= not w135 and not w136;
w138 <= not w131 and not w132;
w139 <= not w133 and not w138;
w140 <= not a(18) and not b(18);
w141 <= a(18) and b(18);
w142 <= not w140 and not w141;
w143 <= w139 and not w142;
w144 <= not w139 and w142;
w145 <= not w143 and not w144;
w146 <= not w139 and not w140;
w147 <= not w141 and not w146;
w148 <= not a(19) and not b(19);
w149 <= a(19) and b(19);
w150 <= not w148 and not w149;
w151 <= w147 and not w150;
w152 <= not w147 and w150;
w153 <= not w151 and not w152;
w154 <= not w147 and not w148;
w155 <= not w149 and not w154;
w156 <= not a(20) and not b(20);
w157 <= a(20) and b(20);
w158 <= not w156 and not w157;
w159 <= w155 and not w158;
w160 <= not w155 and w158;
w161 <= not w159 and not w160;
w162 <= not w155 and not w156;
w163 <= not w157 and not w162;
w164 <= not a(21) and not b(21);
w165 <= a(21) and b(21);
w166 <= not w164 and not w165;
w167 <= w163 and not w166;
w168 <= not w163 and w166;
w169 <= not w167 and not w168;
w170 <= not w163 and not w164;
w171 <= not w165 and not w170;
w172 <= not a(22) and not b(22);
w173 <= a(22) and b(22);
w174 <= not w172 and not w173;
w175 <= w171 and not w174;
w176 <= not w171 and w174;
w177 <= not w175 and not w176;
w178 <= not w171 and not w172;
w179 <= not w173 and not w178;
w180 <= not a(23) and not b(23);
w181 <= a(23) and b(23);
w182 <= not w180 and not w181;
w183 <= w179 and not w182;
w184 <= not w179 and w182;
w185 <= not w183 and not w184;
w186 <= not w179 and not w180;
w187 <= not w181 and not w186;
w188 <= not a(24) and not b(24);
w189 <= a(24) and b(24);
w190 <= not w188 and not w189;
w191 <= w187 and not w190;
w192 <= not w187 and w190;
w193 <= not w191 and not w192;
w194 <= not w187 and not w188;
w195 <= not w189 and not w194;
w196 <= not a(25) and not b(25);
w197 <= a(25) and b(25);
w198 <= not w196 and not w197;
w199 <= w195 and not w198;
w200 <= not w195 and w198;
w201 <= not w199 and not w200;
w202 <= not w195 and not w196;
w203 <= not w197 and not w202;
w204 <= not a(26) and not b(26);
w205 <= a(26) and b(26);
w206 <= not w204 and not w205;
w207 <= w203 and not w206;
w208 <= not w203 and w206;
w209 <= not w207 and not w208;
w210 <= not w203 and not w204;
w211 <= not w205 and not w210;
w212 <= not a(27) and not b(27);
w213 <= a(27) and b(27);
w214 <= not w212 and not w213;
w215 <= w211 and not w214;
w216 <= not w211 and w214;
w217 <= not w215 and not w216;
w218 <= not w211 and not w212;
w219 <= not w213 and not w218;
w220 <= not a(28) and not b(28);
w221 <= a(28) and b(28);
w222 <= not w220 and not w221;
w223 <= w219 and not w222;
w224 <= not w219 and w222;
w225 <= not w223 and not w224;
w226 <= not w219 and not w220;
w227 <= not w221 and not w226;
w228 <= not a(29) and not b(29);
w229 <= a(29) and b(29);
w230 <= not w228 and not w229;
w231 <= w227 and not w230;
w232 <= not w227 and w230;
w233 <= not w231 and not w232;
w234 <= not w227 and not w228;
w235 <= not w229 and not w234;
w236 <= not a(30) and not b(30);
w237 <= a(30) and b(30);
w238 <= not w236 and not w237;
w239 <= w235 and not w238;
w240 <= not w235 and w238;
w241 <= not w239 and not w240;
w242 <= not w235 and not w236;
w243 <= not w237 and not w242;
w244 <= not a(31) and not b(31);
w245 <= a(31) and b(31);
w246 <= not w244 and not w245;
w247 <= w243 and not w246;
w248 <= not w243 and w246;
w249 <= not w247 and not w248;
w250 <= not w243 and not w244;
w251 <= not w245 and not w250;
w252 <= not a(32) and not b(32);
w253 <= a(32) and b(32);
w254 <= not w252 and not w253;
w255 <= w251 and not w254;
w256 <= not w251 and w254;
w257 <= not w255 and not w256;
w258 <= not w251 and not w252;
w259 <= not w253 and not w258;
w260 <= not a(33) and not b(33);
w261 <= a(33) and b(33);
w262 <= not w260 and not w261;
w263 <= w259 and not w262;
w264 <= not w259 and w262;
w265 <= not w263 and not w264;
w266 <= not w259 and not w260;
w267 <= not w261 and not w266;
w268 <= not a(34) and not b(34);
w269 <= a(34) and b(34);
w270 <= not w268 and not w269;
w271 <= w267 and not w270;
w272 <= not w267 and w270;
w273 <= not w271 and not w272;
w274 <= not w267 and not w268;
w275 <= not w269 and not w274;
w276 <= not a(35) and not b(35);
w277 <= a(35) and b(35);
w278 <= not w276 and not w277;
w279 <= w275 and not w278;
w280 <= not w275 and w278;
w281 <= not w279 and not w280;
w282 <= not w275 and not w276;
w283 <= not w277 and not w282;
w284 <= not a(36) and not b(36);
w285 <= a(36) and b(36);
w286 <= not w284 and not w285;
w287 <= w283 and not w286;
w288 <= not w283 and w286;
w289 <= not w287 and not w288;
w290 <= not w283 and not w284;
w291 <= not w285 and not w290;
w292 <= not a(37) and not b(37);
w293 <= a(37) and b(37);
w294 <= not w292 and not w293;
w295 <= w291 and not w294;
w296 <= not w291 and w294;
w297 <= not w295 and not w296;
w298 <= not w291 and not w292;
w299 <= not w293 and not w298;
w300 <= not a(38) and not b(38);
w301 <= a(38) and b(38);
w302 <= not w300 and not w301;
w303 <= w299 and not w302;
w304 <= not w299 and w302;
w305 <= not w303 and not w304;
w306 <= not w299 and not w300;
w307 <= not w301 and not w306;
w308 <= not a(39) and not b(39);
w309 <= a(39) and b(39);
w310 <= not w308 and not w309;
w311 <= w307 and not w310;
w312 <= not w307 and w310;
w313 <= not w311 and not w312;
w314 <= not w307 and not w308;
w315 <= not w309 and not w314;
w316 <= not a(40) and not b(40);
w317 <= a(40) and b(40);
w318 <= not w316 and not w317;
w319 <= w315 and not w318;
w320 <= not w315 and w318;
w321 <= not w319 and not w320;
w322 <= not w315 and not w316;
w323 <= not w317 and not w322;
w324 <= not a(41) and not b(41);
w325 <= a(41) and b(41);
w326 <= not w324 and not w325;
w327 <= w323 and not w326;
w328 <= not w323 and w326;
w329 <= not w327 and not w328;
w330 <= not w323 and not w324;
w331 <= not w325 and not w330;
w332 <= not a(42) and not b(42);
w333 <= a(42) and b(42);
w334 <= not w332 and not w333;
w335 <= w331 and not w334;
w336 <= not w331 and w334;
w337 <= not w335 and not w336;
w338 <= not w331 and not w332;
w339 <= not w333 and not w338;
w340 <= not a(43) and not b(43);
w341 <= a(43) and b(43);
w342 <= not w340 and not w341;
w343 <= w339 and not w342;
w344 <= not w339 and w342;
w345 <= not w343 and not w344;
w346 <= not w339 and not w340;
w347 <= not w341 and not w346;
w348 <= not a(44) and not b(44);
w349 <= a(44) and b(44);
w350 <= not w348 and not w349;
w351 <= w347 and not w350;
w352 <= not w347 and w350;
w353 <= not w351 and not w352;
w354 <= not w347 and not w348;
w355 <= not w349 and not w354;
w356 <= not a(45) and not b(45);
w357 <= a(45) and b(45);
w358 <= not w356 and not w357;
w359 <= w355 and not w358;
w360 <= not w355 and w358;
w361 <= not w359 and not w360;
w362 <= not w355 and not w356;
w363 <= not w357 and not w362;
w364 <= not a(46) and not b(46);
w365 <= a(46) and b(46);
w366 <= not w364 and not w365;
w367 <= w363 and not w366;
w368 <= not w363 and w366;
w369 <= not w367 and not w368;
w370 <= not w363 and not w364;
w371 <= not w365 and not w370;
w372 <= not a(47) and not b(47);
w373 <= a(47) and b(47);
w374 <= not w372 and not w373;
w375 <= w371 and not w374;
w376 <= not w371 and w374;
w377 <= not w375 and not w376;
w378 <= not w371 and not w372;
w379 <= not w373 and not w378;
w380 <= not a(48) and not b(48);
w381 <= a(48) and b(48);
w382 <= not w380 and not w381;
w383 <= w379 and not w382;
w384 <= not w379 and w382;
w385 <= not w383 and not w384;
w386 <= not w379 and not w380;
w387 <= not w381 and not w386;
w388 <= not a(49) and not b(49);
w389 <= a(49) and b(49);
w390 <= not w388 and not w389;
w391 <= w387 and not w390;
w392 <= not w387 and w390;
w393 <= not w391 and not w392;
w394 <= not w387 and not w388;
w395 <= not w389 and not w394;
w396 <= not a(50) and not b(50);
w397 <= a(50) and b(50);
w398 <= not w396 and not w397;
w399 <= w395 and not w398;
w400 <= not w395 and w398;
w401 <= not w399 and not w400;
w402 <= not w395 and not w396;
w403 <= not w397 and not w402;
w404 <= not a(51) and not b(51);
w405 <= a(51) and b(51);
w406 <= not w404 and not w405;
w407 <= w403 and not w406;
w408 <= not w403 and w406;
w409 <= not w407 and not w408;
w410 <= not w403 and not w404;
w411 <= not w405 and not w410;
w412 <= not a(52) and not b(52);
w413 <= a(52) and b(52);
w414 <= not w412 and not w413;
w415 <= w411 and not w414;
w416 <= not w411 and w414;
w417 <= not w415 and not w416;
w418 <= not w411 and not w412;
w419 <= not w413 and not w418;
w420 <= not a(53) and not b(53);
w421 <= a(53) and b(53);
w422 <= not w420 and not w421;
w423 <= w419 and not w422;
w424 <= not w419 and w422;
w425 <= not w423 and not w424;
w426 <= not w419 and not w420;
w427 <= not w421 and not w426;
w428 <= not a(54) and not b(54);
w429 <= a(54) and b(54);
w430 <= not w428 and not w429;
w431 <= w427 and not w430;
w432 <= not w427 and w430;
w433 <= not w431 and not w432;
w434 <= not w427 and not w428;
w435 <= not w429 and not w434;
w436 <= not a(55) and not b(55);
w437 <= a(55) and b(55);
w438 <= not w436 and not w437;
w439 <= w435 and not w438;
w440 <= not w435 and w438;
w441 <= not w439 and not w440;
w442 <= not w435 and not w436;
w443 <= not w437 and not w442;
w444 <= not a(56) and not b(56);
w445 <= a(56) and b(56);
w446 <= not w444 and not w445;
w447 <= w443 and not w446;
w448 <= not w443 and w446;
w449 <= not w447 and not w448;
w450 <= not w443 and not w444;
w451 <= not w445 and not w450;
w452 <= not a(57) and not b(57);
w453 <= a(57) and b(57);
w454 <= not w452 and not w453;
w455 <= w451 and not w454;
w456 <= not w451 and w454;
w457 <= not w455 and not w456;
w458 <= not w451 and not w452;
w459 <= not w453 and not w458;
w460 <= not a(58) and not b(58);
w461 <= a(58) and b(58);
w462 <= not w460 and not w461;
w463 <= w459 and not w462;
w464 <= not w459 and w462;
w465 <= not w463 and not w464;
w466 <= not w459 and not w460;
w467 <= not w461 and not w466;
w468 <= not a(59) and not b(59);
w469 <= a(59) and b(59);
w470 <= not w468 and not w469;
w471 <= w467 and not w470;
w472 <= not w467 and w470;
w473 <= not w471 and not w472;
w474 <= not w467 and not w468;
w475 <= not w469 and not w474;
w476 <= not a(60) and not b(60);
w477 <= a(60) and b(60);
w478 <= not w476 and not w477;
w479 <= w475 and not w478;
w480 <= not w475 and w478;
w481 <= not w479 and not w480;
w482 <= not w475 and not w476;
w483 <= not w477 and not w482;
w484 <= not a(61) and not b(61);
w485 <= a(61) and b(61);
w486 <= not w484 and not w485;
w487 <= w483 and not w486;
w488 <= not w483 and w486;
w489 <= not w487 and not w488;
w490 <= not w483 and not w484;
w491 <= not w485 and not w490;
w492 <= not a(62) and not b(62);
w493 <= a(62) and b(62);
w494 <= not w492 and not w493;
w495 <= w491 and not w494;
w496 <= not w491 and w494;
w497 <= not w495 and not w496;
w498 <= not w491 and not w492;
w499 <= not w493 and not w498;
w500 <= not a(63) and not b(63);
w501 <= a(63) and b(63);
w502 <= not w500 and not w501;
w503 <= w499 and not w502;
w504 <= not w499 and w502;
w505 <= not w503 and not w504;
w506 <= not w499 and not w500;
w507 <= not w501 and not w506;
w508 <= not a(64) and not b(64);
w509 <= a(64) and b(64);
w510 <= not w508 and not w509;
w511 <= w507 and not w510;
w512 <= not w507 and w510;
w513 <= not w511 and not w512;
w514 <= not w507 and not w508;
w515 <= not w509 and not w514;
w516 <= not a(65) and not b(65);
w517 <= a(65) and b(65);
w518 <= not w516 and not w517;
w519 <= w515 and not w518;
w520 <= not w515 and w518;
w521 <= not w519 and not w520;
w522 <= not w515 and not w516;
w523 <= not w517 and not w522;
w524 <= not a(66) and not b(66);
w525 <= a(66) and b(66);
w526 <= not w524 and not w525;
w527 <= w523 and not w526;
w528 <= not w523 and w526;
w529 <= not w527 and not w528;
w530 <= not w523 and not w524;
w531 <= not w525 and not w530;
w532 <= not a(67) and not b(67);
w533 <= a(67) and b(67);
w534 <= not w532 and not w533;
w535 <= w531 and not w534;
w536 <= not w531 and w534;
w537 <= not w535 and not w536;
w538 <= not w531 and not w532;
w539 <= not w533 and not w538;
w540 <= not a(68) and not b(68);
w541 <= a(68) and b(68);
w542 <= not w540 and not w541;
w543 <= w539 and not w542;
w544 <= not w539 and w542;
w545 <= not w543 and not w544;
w546 <= not w539 and not w540;
w547 <= not w541 and not w546;
w548 <= not a(69) and not b(69);
w549 <= a(69) and b(69);
w550 <= not w548 and not w549;
w551 <= w547 and not w550;
w552 <= not w547 and w550;
w553 <= not w551 and not w552;
w554 <= not w547 and not w548;
w555 <= not w549 and not w554;
w556 <= not a(70) and not b(70);
w557 <= a(70) and b(70);
w558 <= not w556 and not w557;
w559 <= w555 and not w558;
w560 <= not w555 and w558;
w561 <= not w559 and not w560;
w562 <= not w555 and not w556;
w563 <= not w557 and not w562;
w564 <= not a(71) and not b(71);
w565 <= a(71) and b(71);
w566 <= not w564 and not w565;
w567 <= w563 and not w566;
w568 <= not w563 and w566;
w569 <= not w567 and not w568;
w570 <= not w563 and not w564;
w571 <= not w565 and not w570;
w572 <= not a(72) and not b(72);
w573 <= a(72) and b(72);
w574 <= not w572 and not w573;
w575 <= w571 and not w574;
w576 <= not w571 and w574;
w577 <= not w575 and not w576;
w578 <= not w571 and not w572;
w579 <= not w573 and not w578;
w580 <= not a(73) and not b(73);
w581 <= a(73) and b(73);
w582 <= not w580 and not w581;
w583 <= w579 and not w582;
w584 <= not w579 and w582;
w585 <= not w583 and not w584;
w586 <= not w579 and not w580;
w587 <= not w581 and not w586;
w588 <= not a(74) and not b(74);
w589 <= a(74) and b(74);
w590 <= not w588 and not w589;
w591 <= w587 and not w590;
w592 <= not w587 and w590;
w593 <= not w591 and not w592;
w594 <= not w587 and not w588;
w595 <= not w589 and not w594;
w596 <= not a(75) and not b(75);
w597 <= a(75) and b(75);
w598 <= not w596 and not w597;
w599 <= w595 and not w598;
w600 <= not w595 and w598;
w601 <= not w599 and not w600;
w602 <= not w595 and not w596;
w603 <= not w597 and not w602;
w604 <= not a(76) and not b(76);
w605 <= a(76) and b(76);
w606 <= not w604 and not w605;
w607 <= w603 and not w606;
w608 <= not w603 and w606;
w609 <= not w607 and not w608;
w610 <= not w603 and not w604;
w611 <= not w605 and not w610;
w612 <= not a(77) and not b(77);
w613 <= a(77) and b(77);
w614 <= not w612 and not w613;
w615 <= w611 and not w614;
w616 <= not w611 and w614;
w617 <= not w615 and not w616;
w618 <= not w611 and not w612;
w619 <= not w613 and not w618;
w620 <= not a(78) and not b(78);
w621 <= a(78) and b(78);
w622 <= not w620 and not w621;
w623 <= w619 and not w622;
w624 <= not w619 and w622;
w625 <= not w623 and not w624;
w626 <= not w619 and not w620;
w627 <= not w621 and not w626;
w628 <= not a(79) and not b(79);
w629 <= a(79) and b(79);
w630 <= not w628 and not w629;
w631 <= w627 and not w630;
w632 <= not w627 and w630;
w633 <= not w631 and not w632;
w634 <= not w627 and not w628;
w635 <= not w629 and not w634;
w636 <= not a(80) and not b(80);
w637 <= a(80) and b(80);
w638 <= not w636 and not w637;
w639 <= w635 and not w638;
w640 <= not w635 and w638;
w641 <= not w639 and not w640;
w642 <= not w635 and not w636;
w643 <= not w637 and not w642;
w644 <= not a(81) and not b(81);
w645 <= a(81) and b(81);
w646 <= not w644 and not w645;
w647 <= w643 and not w646;
w648 <= not w643 and w646;
w649 <= not w647 and not w648;
w650 <= not w643 and not w644;
w651 <= not w645 and not w650;
w652 <= not a(82) and not b(82);
w653 <= a(82) and b(82);
w654 <= not w652 and not w653;
w655 <= w651 and not w654;
w656 <= not w651 and w654;
w657 <= not w655 and not w656;
w658 <= not w651 and not w652;
w659 <= not w653 and not w658;
w660 <= not a(83) and not b(83);
w661 <= a(83) and b(83);
w662 <= not w660 and not w661;
w663 <= w659 and not w662;
w664 <= not w659 and w662;
w665 <= not w663 and not w664;
w666 <= not w659 and not w660;
w667 <= not w661 and not w666;
w668 <= not a(84) and not b(84);
w669 <= a(84) and b(84);
w670 <= not w668 and not w669;
w671 <= w667 and not w670;
w672 <= not w667 and w670;
w673 <= not w671 and not w672;
w674 <= not w667 and not w668;
w675 <= not w669 and not w674;
w676 <= not a(85) and not b(85);
w677 <= a(85) and b(85);
w678 <= not w676 and not w677;
w679 <= w675 and not w678;
w680 <= not w675 and w678;
w681 <= not w679 and not w680;
w682 <= not w675 and not w676;
w683 <= not w677 and not w682;
w684 <= not a(86) and not b(86);
w685 <= a(86) and b(86);
w686 <= not w684 and not w685;
w687 <= w683 and not w686;
w688 <= not w683 and w686;
w689 <= not w687 and not w688;
w690 <= not w683 and not w684;
w691 <= not w685 and not w690;
w692 <= not a(87) and not b(87);
w693 <= a(87) and b(87);
w694 <= not w692 and not w693;
w695 <= w691 and not w694;
w696 <= not w691 and w694;
w697 <= not w695 and not w696;
w698 <= not w691 and not w692;
w699 <= not w693 and not w698;
w700 <= not a(88) and not b(88);
w701 <= a(88) and b(88);
w702 <= not w700 and not w701;
w703 <= w699 and not w702;
w704 <= not w699 and w702;
w705 <= not w703 and not w704;
w706 <= not w699 and not w700;
w707 <= not w701 and not w706;
w708 <= not a(89) and not b(89);
w709 <= a(89) and b(89);
w710 <= not w708 and not w709;
w711 <= w707 and not w710;
w712 <= not w707 and w710;
w713 <= not w711 and not w712;
w714 <= not w707 and not w708;
w715 <= not w709 and not w714;
w716 <= not a(90) and not b(90);
w717 <= a(90) and b(90);
w718 <= not w716 and not w717;
w719 <= w715 and not w718;
w720 <= not w715 and w718;
w721 <= not w719 and not w720;
w722 <= not w715 and not w716;
w723 <= not w717 and not w722;
w724 <= not a(91) and not b(91);
w725 <= a(91) and b(91);
w726 <= not w724 and not w725;
w727 <= w723 and not w726;
w728 <= not w723 and w726;
w729 <= not w727 and not w728;
w730 <= not w723 and not w724;
w731 <= not w725 and not w730;
w732 <= not a(92) and not b(92);
w733 <= a(92) and b(92);
w734 <= not w732 and not w733;
w735 <= w731 and not w734;
w736 <= not w731 and w734;
w737 <= not w735 and not w736;
w738 <= not w731 and not w732;
w739 <= not w733 and not w738;
w740 <= not a(93) and not b(93);
w741 <= a(93) and b(93);
w742 <= not w740 and not w741;
w743 <= w739 and not w742;
w744 <= not w739 and w742;
w745 <= not w743 and not w744;
w746 <= not w739 and not w740;
w747 <= not w741 and not w746;
w748 <= not a(94) and not b(94);
w749 <= a(94) and b(94);
w750 <= not w748 and not w749;
w751 <= w747 and not w750;
w752 <= not w747 and w750;
w753 <= not w751 and not w752;
w754 <= not w747 and not w748;
w755 <= not w749 and not w754;
w756 <= not a(95) and not b(95);
w757 <= a(95) and b(95);
w758 <= not w756 and not w757;
w759 <= w755 and not w758;
w760 <= not w755 and w758;
w761 <= not w759 and not w760;
w762 <= not w755 and not w756;
w763 <= not w757 and not w762;
w764 <= not a(96) and not b(96);
w765 <= a(96) and b(96);
w766 <= not w764 and not w765;
w767 <= w763 and not w766;
w768 <= not w763 and w766;
w769 <= not w767 and not w768;
w770 <= not w763 and not w764;
w771 <= not w765 and not w770;
w772 <= not a(97) and not b(97);
w773 <= a(97) and b(97);
w774 <= not w772 and not w773;
w775 <= w771 and not w774;
w776 <= not w771 and w774;
w777 <= not w775 and not w776;
w778 <= not w771 and not w772;
w779 <= not w773 and not w778;
w780 <= not a(98) and not b(98);
w781 <= a(98) and b(98);
w782 <= not w780 and not w781;
w783 <= w779 and not w782;
w784 <= not w779 and w782;
w785 <= not w783 and not w784;
w786 <= not w779 and not w780;
w787 <= not w781 and not w786;
w788 <= not a(99) and not b(99);
w789 <= a(99) and b(99);
w790 <= not w788 and not w789;
w791 <= w787 and not w790;
w792 <= not w787 and w790;
w793 <= not w791 and not w792;
w794 <= not w787 and not w788;
w795 <= not w789 and not w794;
w796 <= not a(100) and not b(100);
w797 <= a(100) and b(100);
w798 <= not w796 and not w797;
w799 <= w795 and not w798;
w800 <= not w795 and w798;
w801 <= not w799 and not w800;
w802 <= not w795 and not w796;
w803 <= not w797 and not w802;
w804 <= not a(101) and not b(101);
w805 <= a(101) and b(101);
w806 <= not w804 and not w805;
w807 <= w803 and not w806;
w808 <= not w803 and w806;
w809 <= not w807 and not w808;
w810 <= not w803 and not w804;
w811 <= not w805 and not w810;
w812 <= not a(102) and not b(102);
w813 <= a(102) and b(102);
w814 <= not w812 and not w813;
w815 <= w811 and not w814;
w816 <= not w811 and w814;
w817 <= not w815 and not w816;
w818 <= not w811 and not w812;
w819 <= not w813 and not w818;
w820 <= not a(103) and not b(103);
w821 <= a(103) and b(103);
w822 <= not w820 and not w821;
w823 <= w819 and not w822;
w824 <= not w819 and w822;
w825 <= not w823 and not w824;
w826 <= not w819 and not w820;
w827 <= not w821 and not w826;
w828 <= not a(104) and not b(104);
w829 <= a(104) and b(104);
w830 <= not w828 and not w829;
w831 <= w827 and not w830;
w832 <= not w827 and w830;
w833 <= not w831 and not w832;
w834 <= not w827 and not w828;
w835 <= not w829 and not w834;
w836 <= not a(105) and not b(105);
w837 <= a(105) and b(105);
w838 <= not w836 and not w837;
w839 <= w835 and not w838;
w840 <= not w835 and w838;
w841 <= not w839 and not w840;
w842 <= not w835 and not w836;
w843 <= not w837 and not w842;
w844 <= not a(106) and not b(106);
w845 <= a(106) and b(106);
w846 <= not w844 and not w845;
w847 <= w843 and not w846;
w848 <= not w843 and w846;
w849 <= not w847 and not w848;
w850 <= not w843 and not w844;
w851 <= not w845 and not w850;
w852 <= not a(107) and not b(107);
w853 <= a(107) and b(107);
w854 <= not w852 and not w853;
w855 <= w851 and not w854;
w856 <= not w851 and w854;
w857 <= not w855 and not w856;
w858 <= not w851 and not w852;
w859 <= not w853 and not w858;
w860 <= not a(108) and not b(108);
w861 <= a(108) and b(108);
w862 <= not w860 and not w861;
w863 <= w859 and not w862;
w864 <= not w859 and w862;
w865 <= not w863 and not w864;
w866 <= not w859 and not w860;
w867 <= not w861 and not w866;
w868 <= not a(109) and not b(109);
w869 <= a(109) and b(109);
w870 <= not w868 and not w869;
w871 <= w867 and not w870;
w872 <= not w867 and w870;
w873 <= not w871 and not w872;
w874 <= not w867 and not w868;
w875 <= not w869 and not w874;
w876 <= not a(110) and not b(110);
w877 <= a(110) and b(110);
w878 <= not w876 and not w877;
w879 <= w875 and not w878;
w880 <= not w875 and w878;
w881 <= not w879 and not w880;
w882 <= not w875 and not w876;
w883 <= not w877 and not w882;
w884 <= not a(111) and not b(111);
w885 <= a(111) and b(111);
w886 <= not w884 and not w885;
w887 <= w883 and not w886;
w888 <= not w883 and w886;
w889 <= not w887 and not w888;
w890 <= not w883 and not w884;
w891 <= not w885 and not w890;
w892 <= not a(112) and not b(112);
w893 <= a(112) and b(112);
w894 <= not w892 and not w893;
w895 <= w891 and not w894;
w896 <= not w891 and w894;
w897 <= not w895 and not w896;
w898 <= not w891 and not w892;
w899 <= not w893 and not w898;
w900 <= not a(113) and not b(113);
w901 <= a(113) and b(113);
w902 <= not w900 and not w901;
w903 <= w899 and not w902;
w904 <= not w899 and w902;
w905 <= not w903 and not w904;
w906 <= not w899 and not w900;
w907 <= not w901 and not w906;
w908 <= not a(114) and not b(114);
w909 <= a(114) and b(114);
w910 <= not w908 and not w909;
w911 <= w907 and not w910;
w912 <= not w907 and w910;
w913 <= not w911 and not w912;
w914 <= not w907 and not w908;
w915 <= not w909 and not w914;
w916 <= not a(115) and not b(115);
w917 <= a(115) and b(115);
w918 <= not w916 and not w917;
w919 <= w915 and not w918;
w920 <= not w915 and w918;
w921 <= not w919 and not w920;
w922 <= not w915 and not w916;
w923 <= not w917 and not w922;
w924 <= not a(116) and not b(116);
w925 <= a(116) and b(116);
w926 <= not w924 and not w925;
w927 <= w923 and not w926;
w928 <= not w923 and w926;
w929 <= not w927 and not w928;
w930 <= not w923 and not w924;
w931 <= not w925 and not w930;
w932 <= not a(117) and not b(117);
w933 <= a(117) and b(117);
w934 <= not w932 and not w933;
w935 <= w931 and not w934;
w936 <= not w931 and w934;
w937 <= not w935 and not w936;
w938 <= not w931 and not w932;
w939 <= not w933 and not w938;
w940 <= not a(118) and not b(118);
w941 <= a(118) and b(118);
w942 <= not w940 and not w941;
w943 <= w939 and not w942;
w944 <= not w939 and w942;
w945 <= not w943 and not w944;
w946 <= not w939 and not w940;
w947 <= not w941 and not w946;
w948 <= not a(119) and not b(119);
w949 <= a(119) and b(119);
w950 <= not w948 and not w949;
w951 <= w947 and not w950;
w952 <= not w947 and w950;
w953 <= not w951 and not w952;
w954 <= not w947 and not w948;
w955 <= not w949 and not w954;
w956 <= not a(120) and not b(120);
w957 <= a(120) and b(120);
w958 <= not w956 and not w957;
w959 <= w955 and not w958;
w960 <= not w955 and w958;
w961 <= not w959 and not w960;
w962 <= not w955 and not w956;
w963 <= not w957 and not w962;
w964 <= not a(121) and not b(121);
w965 <= a(121) and b(121);
w966 <= not w964 and not w965;
w967 <= w963 and not w966;
w968 <= not w963 and w966;
w969 <= not w967 and not w968;
w970 <= not w963 and not w964;
w971 <= not w965 and not w970;
w972 <= not a(122) and not b(122);
w973 <= a(122) and b(122);
w974 <= not w972 and not w973;
w975 <= w971 and not w974;
w976 <= not w971 and w974;
w977 <= not w975 and not w976;
w978 <= not w971 and not w972;
w979 <= not w973 and not w978;
w980 <= not a(123) and not b(123);
w981 <= a(123) and b(123);
w982 <= not w980 and not w981;
w983 <= w979 and not w982;
w984 <= not w979 and w982;
w985 <= not w983 and not w984;
w986 <= not w979 and not w980;
w987 <= not w981 and not w986;
w988 <= not a(124) and not b(124);
w989 <= a(124) and b(124);
w990 <= not w988 and not w989;
w991 <= w987 and not w990;
w992 <= not w987 and w990;
w993 <= not w991 and not w992;
w994 <= not w987 and not w988;
w995 <= not w989 and not w994;
w996 <= not a(125) and not b(125);
w997 <= a(125) and b(125);
w998 <= not w996 and not w997;
w999 <= w995 and not w998;
w1000 <= not w995 and w998;
w1001 <= not w999 and not w1000;
w1002 <= not w995 and not w996;
w1003 <= not w997 and not w1002;
w1004 <= not a(126) and not b(126);
w1005 <= a(126) and b(126);
w1006 <= not w1004 and not w1005;
w1007 <= w1003 and not w1006;
w1008 <= not w1003 and w1006;
w1009 <= not w1007 and not w1008;
w1010 <= not w1003 and not w1004;
w1011 <= not w1005 and not w1010;
w1012 <= not a(127) and not b(127);
w1013 <= a(127) and b(127);
w1014 <= not w1012 and not w1013;
w1015 <= w1011 and not w1014;
w1016 <= not w1011 and w1014;
w1017 <= not w1015 and not w1016;
w1018 <= not w1011 and not w1012;
w1019 <= not w1013 and not w1018;
one <= '1';
f(0) <= not w2;-- level 2
f(1) <= not w9;-- level 4
f(2) <= w17;-- level 5
f(3) <= w25;-- level 7
f(4) <= w33;-- level 9
f(5) <= w41;-- level 11
f(6) <= w49;-- level 13
f(7) <= w57;-- level 15
f(8) <= w65;-- level 17
f(9) <= w73;-- level 19
f(10) <= w81;-- level 21
f(11) <= w89;-- level 23
f(12) <= w97;-- level 25
f(13) <= w105;-- level 27
f(14) <= w113;-- level 29
f(15) <= w121;-- level 31
f(16) <= w129;-- level 33
f(17) <= w137;-- level 35
f(18) <= w145;-- level 37
f(19) <= w153;-- level 39
f(20) <= w161;-- level 41
f(21) <= w169;-- level 43
f(22) <= w177;-- level 45
f(23) <= w185;-- level 47
f(24) <= w193;-- level 49
f(25) <= w201;-- level 51
f(26) <= w209;-- level 53
f(27) <= w217;-- level 55
f(28) <= w225;-- level 57
f(29) <= w233;-- level 59
f(30) <= w241;-- level 61
f(31) <= w249;-- level 63
f(32) <= w257;-- level 65
f(33) <= w265;-- level 67
f(34) <= w273;-- level 69
f(35) <= w281;-- level 71
f(36) <= w289;-- level 73
f(37) <= w297;-- level 75
f(38) <= w305;-- level 77
f(39) <= w313;-- level 79
f(40) <= w321;-- level 81
f(41) <= w329;-- level 83
f(42) <= w337;-- level 85
f(43) <= w345;-- level 87
f(44) <= w353;-- level 89
f(45) <= w361;-- level 91
f(46) <= w369;-- level 93
f(47) <= w377;-- level 95
f(48) <= w385;-- level 97
f(49) <= w393;-- level 99
f(50) <= w401;-- level 101
f(51) <= w409;-- level 103
f(52) <= w417;-- level 105
f(53) <= w425;-- level 107
f(54) <= w433;-- level 109
f(55) <= w441;-- level 111
f(56) <= w449;-- level 113
f(57) <= w457;-- level 115
f(58) <= w465;-- level 117
f(59) <= w473;-- level 119
f(60) <= w481;-- level 121
f(61) <= w489;-- level 123
f(62) <= w497;-- level 125
f(63) <= w505;-- level 127
f(64) <= w513;-- level 129
f(65) <= w521;-- level 131
f(66) <= w529;-- level 133
f(67) <= w537;-- level 135
f(68) <= w545;-- level 137
f(69) <= w553;-- level 139
f(70) <= w561;-- level 141
f(71) <= w569;-- level 143
f(72) <= w577;-- level 145
f(73) <= w585;-- level 147
f(74) <= w593;-- level 149
f(75) <= w601;-- level 151
f(76) <= w609;-- level 153
f(77) <= w617;-- level 155
f(78) <= w625;-- level 157
f(79) <= w633;-- level 159
f(80) <= w641;-- level 161
f(81) <= w649;-- level 163
f(82) <= w657;-- level 165
f(83) <= w665;-- level 167
f(84) <= w673;-- level 169
f(85) <= w681;-- level 171
f(86) <= w689;-- level 173
f(87) <= w697;-- level 175
f(88) <= w705;-- level 177
f(89) <= w713;-- level 179
f(90) <= w721;-- level 181
f(91) <= w729;-- level 183
f(92) <= w737;-- level 185
f(93) <= w745;-- level 187
f(94) <= w753;-- level 189
f(95) <= w761;-- level 191
f(96) <= w769;-- level 193
f(97) <= w777;-- level 195
f(98) <= w785;-- level 197
f(99) <= w793;-- level 199
f(100) <= w801;-- level 201
f(101) <= w809;-- level 203
f(102) <= w817;-- level 205
f(103) <= w825;-- level 207
f(104) <= w833;-- level 209
f(105) <= w841;-- level 211
f(106) <= w849;-- level 213
f(107) <= w857;-- level 215
f(108) <= w865;-- level 217
f(109) <= w873;-- level 219
f(110) <= w881;-- level 221
f(111) <= w889;-- level 223
f(112) <= w897;-- level 225
f(113) <= w905;-- level 227
f(114) <= w913;-- level 229
f(115) <= w921;-- level 231
f(116) <= w929;-- level 233
f(117) <= w937;-- level 235
f(118) <= w945;-- level 237
f(119) <= w953;-- level 239
f(120) <= w961;-- level 241
f(121) <= w969;-- level 243
f(122) <= w977;-- level 245
f(123) <= w985;-- level 247
f(124) <= w993;-- level 249
f(125) <= w1001;-- level 251
f(126) <= w1009;-- level 253
f(127) <= w1017;-- level 255
cOut <= not w1019;-- level 255
end Behavioral;