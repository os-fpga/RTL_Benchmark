// Copyright (C) 2022, Andes Technology Corp. Confidential Proprietary

module kv_dsp_predec (
    instr,
    csr_mmisc_ctl_rvcompm,
    instr_dsp,
    instr_legal_dsp,
    rs1_ren,
    rs2_ren,
    rs3_ren,
    rs4_ren,
    rs1_addr,
    rs2_addr,
    rs3_addr,
    rs4_addr,
    rd1_wen,
    rd2_wen,
    rd1_addr,
    rd2_addr,
    ready_stage
);
parameter OP_DSP = 7'b1111111;
input [31:0] instr;
input csr_mmisc_ctl_rvcompm;
output instr_dsp;
output instr_legal_dsp;
output rs1_ren;
output rs2_ren;
output rs3_ren;
output rs4_ren;
output [4:0] rs1_addr;
output [4:0] rs2_addr;
output [4:0] rs3_addr;
output [4:0] rs4_addr;
output rd1_wen;
output rd2_wen;
output [4:0] rd1_addr;
output [4:0] rd2_addr;
output [2:0] ready_stage;


wire s0;
wire s1;
wire s2;
wire s3;
wire s4;
wire s5;
wire s6;
wire s7;
wire s8;
wire s9;
wire s10;
wire s11;
wire s12;
wire s13;
wire s14;
wire s15;
wire s16;
wire s17;
wire s18;
wire s19;
wire s20;
wire s21;
wire s22;
wire s23;
wire s24;
wire s25;
wire s26;
wire s27;
wire s28;
wire s29;
wire s30;
wire s31;
wire s32;
wire s33;
wire s34;
wire s35;
wire s36;
wire s37;
wire s38;
wire s39;
wire s40;
wire s41;
wire s42;
wire s43;
wire s44;
wire s45;
wire s46;
wire s47;
wire s48;
wire s49;
wire s50;
wire s51;
wire s52;
wire s53;
wire s54;
wire s55;
wire s56;
wire s57;
wire s58;
wire s59;
wire s60;
wire s61;
wire s62;
wire s63;
wire s64;
wire s65;
wire s66;
wire s67;
wire s68;
wire s69;
wire s70;
wire s71;
wire s72;
wire s73;
wire s74;
wire s75;
wire s76;
wire s77;
wire s78;
wire s79;
wire s80;
wire s81;
wire s82;
wire s83;
wire s84;
wire s85;
wire s86;
wire s87;
wire s88;
wire s89;
wire s90;
wire s91;
wire s92;
wire s93;
wire s94;
wire s95;
wire s96;
wire s97;
wire s98;
wire s99;
wire s100;
wire s101;
wire s102;
wire s103;
wire s104;
wire s105;
wire s106;
wire s107;
wire s108;
wire s109;
wire s110;
wire s111;
wire s112;
wire s113;
wire s114;
wire s115;
wire s116;
wire s117;
wire s118;
wire s119;
wire s120;
wire s121;
wire s122;
wire s123;
wire s124;
wire s125;
wire s126;
wire s127;
wire s128;
wire s129;
wire s130;
wire s131;
wire s132;
wire s133;
wire s134;
wire s135;
wire s136;
wire s137;
wire s138;
wire s139;
wire s140;
wire s141;
wire s142;
wire s143;
wire s144;
wire s145;
wire s146;
wire s147;
wire s148;
wire s149;
wire s150;
wire s151;
wire s152;
wire s153;
wire s154;
wire s155;
wire s156;
wire s157;
wire s158;
wire s159;
wire s160;
wire s161;
wire s162;
wire s163;
wire s164;
wire s165;
wire s166;
wire s167;
wire s168;
wire s169;
wire s170;
wire s171;
wire s172;
wire s173;
wire s174;
wire s175;
wire s176;
wire s177;
wire s178;
wire s179;
wire s180;
wire s181;
wire s182;
wire s183;
wire s184;
wire s185;
wire s186;
wire s187;
wire s188;
wire s189;
wire s190;
wire s191;
wire s192;
wire s193;
wire s194;
wire s195;
wire s196;
wire s197;
wire s198;
wire s199;
wire s200;
wire s201;
wire s202;
wire s203;
wire s204;
wire s205;
wire s206;
wire s207;
wire s208;
wire s209;
wire s210;
wire s211;
wire s212;
wire s213;
wire s214;
wire s215;
wire s216;
wire s217;
wire s218;
wire s219;
wire s220;
wire s221;
wire s222;
wire s223;
wire s224;
wire s225;
wire s226;
wire s227;
wire s228;
wire s229;
wire s230;
wire s231;
wire s232;
wire s233;
wire s234;
wire s235;
wire s236;
wire s237;
wire s238;
wire s239;
wire s240;
wire s241;
wire s242;
wire s243;
wire s244;
wire s245;
wire s246;
wire s247;
wire s248;
wire s249;
wire s250;
wire s251;
wire s252;
wire s253;
wire s254;
wire s255;
wire s256;
wire s257;
wire s258;
wire s259;
wire s260;
wire s261;
wire s262;
wire s263;
wire s264;
wire s265;
wire s266;
wire s267;
wire s268;
wire s269;
wire s270;
wire s271;
wire s272;
wire s273;
wire s274;
wire s275;
wire s276;
wire s277;
wire s278;
wire s279;
wire s280;
wire s281;
wire s282;
wire s283;
wire s284;
wire s285;
wire s286;
wire s287;
wire s288;
wire s289;
wire s290;
wire s291;
wire s292;
wire s293;
wire s294;
wire s295;
wire s296;
wire s297;
wire s298;
wire s299;
wire s300;
wire s301;
wire s302;
wire s303;
wire s304;
wire s305;
wire s306;
wire s307;
wire s308;
wire s309;
wire s310;
wire s311;
wire s312;
wire s313;
wire s314;
wire s315;
wire s316;
wire s317;
wire s318;
wire s319;
wire s320;
wire s321;
wire s322;
wire s323;
wire s324;
wire s325;
wire s326;
wire s327;
wire s328;
wire s329;
wire s330;
wire s331;
wire s332;
wire s333;
wire s334;
wire s335;
wire s336;
wire s337;
wire s338;
wire s339;
wire s340;
wire s341;
wire s342;
wire s343;
wire s344;
wire s345;
wire [4:0] s346;
wire [4:0] s347;
wire [4:0] s348;
wire [4:0] s349;
wire [4:0] s350;
wire [4:0] s351;
wire [4:0] s352;
wire [4:0] s353;
wire [4:0] s354;
wire [4:0] s355;
wire [4:0] s356;
wire [4:0] s357;
wire [4:0] s358;
wire [4:0] s359;
assign instr_dsp = (instr[6:0] == OP_DSP);
assign s0 = (instr[31:25] == 7'b0100100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s1 = (instr[31:25] == 7'b0100000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s2 = (instr[31:25] == 7'b1100000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s3 = (instr[31:25] == 7'b1110000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s4 = (instr[31:25] == 7'b1110011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s5 = (instr[31:26] == 6'b111010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s6 = (instr[31:30] == 2'b11) & (instr[14:12] == 3'b010) & (instr[6:0] == OP_DSP);
assign s7 = (instr[31:20] == 12'b101011100000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s8 = (instr[31:20] == 12'b101011101000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s9 = (instr[31:20] == 12'b101011111000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s10 = (instr[31:20] == 12'b101011100011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s11 = (instr[31:20] == 12'b101011101011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s12 = (instr[31:20] == 12'b101011111011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s13 = (instr[31:20] == 12'b101011100001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s14 = (instr[31:20] == 12'b101011101001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s15 = (instr[31:20] == 12'b101011111001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s16 = (instr[31:25] == 7'b0100111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s17 = (instr[31:25] == 7'b0100110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s18 = (instr[31:25] == 7'b0100010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s19 = (instr[31:25] == 7'b0100011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s20 = (instr[31:23] == 9'b101011000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s21 = (instr[31:20] == 12'b101011010000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s22 = (instr[31:20] == 12'b101011010001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s23 = (instr[31:20] == 12'b101011010100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s24 = (instr[31:25] == 7'b0001100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s25 = (instr[31:25] == 7'b0001000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s26 = (instr[31:25] == 7'b1001000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s27 = (instr[31:25] == 7'b0000010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s28 = (instr[31:25] == 7'b0000000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s29 = (instr[31:25] == 7'b0001010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s30 = (instr[31:25] == 7'b0001011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s31 = (instr[31:25] == 7'b0000101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s32 = (instr[31:25] == 7'b0001101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s33 = (instr[31:25] == 7'b0010101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s34 = (instr[31:25] == 7'b1101001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s35 = (instr[31:25] == 7'b1110001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s36 = (instr[31:25] == 7'b1111001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s37 = (instr[31:25] == 7'b1000111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s38 = (instr[31:25] == 7'b1001111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s39 = (instr[31:25] == 7'b1000011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s40 = (instr[31:25] == 7'b1001011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s41 = (instr[31:25] == 7'b0000110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s42 = (instr[31:25] == 7'b0001110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s43 = (instr[31:25] == 7'b0010110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s44 = (instr[31:25] == 7'b0101101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s45 = (instr[31:25] == 7'b0110101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s46 = (instr[31:25] == 7'b0111101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s47 = (instr[31:25] == 7'b0100100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s48 = (instr[31:25] == 7'b0100101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s49 = (instr[31:25] == 7'b0101110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s50 = (instr[31:25] == 7'b0110110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s51 = (instr[31:25] == 7'b0111110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s52 = (instr[31:25] == 7'b1001010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s53 = (instr[31:25] == 7'b0011100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s54 = (instr[31:25] == 7'b0011101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s55 = (instr[31:25] == 7'b0110000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s56 = (instr[31:25] == 7'b0111000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s57 = (instr[31:25] == 7'b0100011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s58 = (instr[31:25] == 7'b0101011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s59 = (instr[31:25] == 7'b1100111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s60 = (instr[31:25] == 7'b1101111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s61 = (instr[31:25] == 7'b0110011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s62 = (instr[31:25] == 7'b0111011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s63 = (instr[31:25] == 7'b1110111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s64 = (instr[31:25] == 7'b1111111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s65 = (instr[31:25] == 7'b0100001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s66 = (instr[31:25] == 7'b0101001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s67 = (instr[31:25] == 7'b1000111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s68 = (instr[31:25] == 7'b1001111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s69 = (instr[31:25] == 7'b1010111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s70 = (instr[31:25] == 7'b1011111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s71 = (instr[31:25] == 7'b0100110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s72 = (instr[31:25] == 7'b0100111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s73 = (instr[31:25] == 7'b1001011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s74 = (instr[31:25] == 7'b0010011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s75 = (instr[31:25] == 7'b0011011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s76 = (instr[31:25] == 7'b0110110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s77 = (instr[31:23] == 9'b011111001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s78 = (instr[31:25] == 7'b0110010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s79 = (instr[31:24] == 8'b01110101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s80 = (instr[31:25] == 7'b0101111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s81 = (instr[31:25] == 7'b0110111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s82 = (instr[31:25] == 7'b0101011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s83 = (instr[31:25] == 7'b0110011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s84 = (instr[31:25] == 7'b0110111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s85 = (instr[31:25] == 7'b0111111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s86 = (instr[31:25] == 7'b0001010) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s87 = (instr[31:25] == 7'b0001011) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s88 = (instr[31:25] == 7'b0001101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s89 = (instr[31:25] == 7'b0001001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s90 = (instr[31:25] == 7'b1001001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s91 = (instr[31:25] == 7'b0000011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s92 = (instr[31:25] == 7'b0000001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s93 = (instr[31:25] == 7'b0110001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s94 = (instr[31:25] == 7'b0111001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s95 = (instr[31:25] == 7'b1100010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s96 = (instr[31:25] == 7'b1111001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s97 = (instr[31:25] == 7'b1111000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s98 = (instr[31:25] == 7'b1100011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s99 = (instr[31:25] == 7'b1111000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s100 = (instr[31:25] == 7'b1110000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s101 = (instr[31:25] == 7'b1111110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s102 = (instr[31:25] == 7'b1111111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s103 = (instr[31:25] == 7'b0000111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s104 = (instr[31:25] == 7'b0001111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s105 = (instr[31:25] == 7'b0010111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s106 = (instr[31:25] == 7'b0011111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s107 = (instr[31:25] == 7'b0000100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s108 = (instr[31:25] == 7'b0000000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s109 = (instr[31:25] == 7'b1000000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s110 = (instr[31:25] == 7'b0010000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s111 = (instr[31:25] == 7'b0000010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s112 = (instr[31:25] == 7'b0000011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s113 = (instr[31:25] == 7'b0000010) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s114 = (instr[31:25] == 7'b0000011) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s115 = (instr[31:25] == 7'b0000101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s116 = (instr[31:25] == 7'b0000001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s117 = (instr[31:25] == 7'b1000001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s118 = (instr[31:25] == 7'b0010001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s119 = (instr[31:23] == 9'b100011000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s120 = (instr[31:24] == 8'b10000100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s121 = (instr[31:25] == 7'b1110010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s122 = (instr[31:25] == 7'b0001111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s123 = (instr[31:25] == 7'b0001110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s124 = (instr[31:25] == 7'b0000111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s125 = (instr[31:25] == 7'b0000110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s126 = (instr[31:25] == 7'b0101110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s127 = (instr[31:23] == 9'b011111000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s128 = (instr[31:25] == 7'b0101010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s129 = (instr[31:24] == 8'b01110100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s130 = (instr[31:25] == 7'b0101111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s131 = (instr[31:25] == 7'b1000100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s132 = (instr[31:25] == 7'b1001100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s133 = (instr[31:25] == 7'b1010100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s134 = (instr[31:25] == 7'b1000110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s135 = (instr[31:25] == 7'b1001110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s136 = (instr[31:25] == 7'b1000101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s137 = (instr[31:25] == 7'b1001101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s138 = (instr[31:25] == 7'b1010101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s139 = (instr[31:25] == 7'b1000010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s140 = (instr[31:25] == 7'b1100100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s141 = (instr[31:25] == 7'b1100101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s142 = (instr[31:25] == 7'b1000101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s143 = (instr[31:25] == 7'b1000001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s144 = (instr[31:25] == 7'b0000100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s145 = (instr[31:25] == 7'b0001100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s146 = (instr[31:25] == 7'b0010100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s147 = (instr[31:25] == 7'b0101100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s148 = (instr[31:25] == 7'b0110100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s149 = (instr[31:25] == 7'b0111100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s150 = (instr[31:25] == 7'b1000100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s151 = (instr[31:25] == 7'b1000000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s152 = (instr[31:25] == 7'b0100000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s153 = (instr[31:25] == 7'b0101000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s154 = (instr[31:25] == 7'b0100010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s155 = (instr[31:25] == 7'b0101010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s156 = (instr[31:25] == 7'b0110010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s157 = (instr[31:25] == 7'b0111010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s158 = (instr[31:25] == 7'b1010110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s159 = (instr[31:25] == 7'b1011110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s160 = (instr[31:25] == 7'b1000011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s161 = (instr[31:25] == 7'b1010100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s162 = (instr[31:25] == 7'b1010101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s163 = (instr[31:25] == 7'b1010000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s164 = (instr[31:25] == 7'b1010001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s165 = (instr[31:25] == 7'b0010010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s166 = (instr[31:26] == 6'b110101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s167 = (instr[31:25] == 7'b0101100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s168 = (instr[31:25] == 7'b0110100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s169 = (instr[31:23] == 9'b011110000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s170 = (instr[31:23] == 9'b011110001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s171 = (instr[31:25] == 7'b0101000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s172 = (instr[31:25] == 7'b0110000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s173 = (instr[31:24] == 8'b01110000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s174 = (instr[31:24] == 8'b01110001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s175 = (instr[31:25] == 7'b0101101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s176 = (instr[31:25] == 7'b0110101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s177 = (instr[31:23] == 9'b011110100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s178 = (instr[31:23] == 9'b011110101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s179 = (instr[31:25] == 7'b0101001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s180 = (instr[31:25] == 7'b0110001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s181 = (instr[31:24] == 8'b01110010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s182 = (instr[31:24] == 8'b01110011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s183 = (instr[31:25] == 7'b0100010) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s184 = (instr[31:25] == 7'b0100011) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s185 = (instr[31:25] == 7'b0100101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s186 = (instr[31:25] == 7'b0100001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s187 = (instr[31:25] == 7'b1100001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s188 = (instr[31:20] == 12'b101011001000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s189 = (instr[31:20] == 12'b101011001001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s190 = (instr[31:20] == 12'b101011001010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s191 = (instr[31:20] == 12'b101011001011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s192 = (instr[31:20] == 12'b101011010011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s193 = (instr[31:20] == 12'b101011011000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s194 = (instr[31:20] == 12'b101011011001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s195 = (instr[31:23] == 9'b100011010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s196 = (instr[31:24] == 8'b10000101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s197 = (instr[31:25] == 7'b1111010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s198 = (instr[31:25] == 7'b0011111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s199 = (instr[31:25] == 7'b0011110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s200 = (instr[31:25] == 7'b0010111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s201 = (instr[31:25] == 7'b0010110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s202 = (instr[31:25] == 7'b0011100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s203 = (instr[31:25] == 7'b0011000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s204 = (instr[31:25] == 7'b1011000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s205 = (instr[31:25] == 7'b0001010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s206 = (instr[31:25] == 7'b0001000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s207 = (instr[31:25] == 7'b0011010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s208 = (instr[31:25] == 7'b0011011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s209 = (instr[31:25] == 7'b1011010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s210 = (instr[31:25] == 7'b1011011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s211 = (instr[31:25] == 7'b0011010) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s212 = (instr[31:25] == 7'b0011011) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s213 = (instr[31:25] == 7'b0011101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s214 = (instr[31:25] == 7'b0011001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s215 = (instr[31:25] == 7'b1011001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s216 = (instr[31:25] == 7'b0001011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s217 = (instr[31:25] == 7'b0001001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s218 = (instr[31:25] == 7'b1010010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s219 = (instr[31:25] == 7'b1100110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s220 = (instr[31:25] == 7'b1001101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s221 = (instr[31:25] == 7'b1001001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s222 = (instr[31:25] == 7'b1001100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s223 = (instr[31:25] == 7'b1001000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s224 = (instr[31:25] == 7'b1010011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s225 = (instr[31:25] == 7'b1011100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s226 = (instr[31:25] == 7'b1011101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s227 = (instr[31:25] == 7'b1011000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s228 = (instr[31:25] == 7'b1011001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s229 = (instr[31:25] == 7'b0010100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s230 = (instr[31:25] == 7'b0010000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s231 = (instr[31:25] == 7'b1010000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s232 = (instr[31:25] == 7'b0011000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s233 = (instr[31:25] == 7'b0010010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s234 = (instr[31:25] == 7'b0010011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s235 = (instr[31:25] == 7'b0010010) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s236 = (instr[31:25] == 7'b0010011) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s237 = (instr[31:25] == 7'b0010101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s238 = (instr[31:25] == 7'b0010001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s239 = (instr[31:25] == 7'b1010001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s240 = (instr[31:25] == 7'b0011001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s241 = (instr[31:25] == 7'b1101111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s242 = (instr[31:25] == 7'b1100111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s243 = (instr[31:20] == 12'b101011001100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s244 = (instr[31:20] == 12'b101011001101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s245 = (instr[31:20] == 12'b101011001110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s246 = (instr[31:20] == 12'b101011001111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s247 = (instr[31:20] == 12'b101011010111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s248 = 1'b0;
assign s249 = 1'b0;
assign s250 = 1'b0;
assign s251 = 1'b0;
assign s252 = 1'b0;
assign s253 = 1'b0;
assign s254 = 1'b0;
assign s255 = 1'b0;
assign s256 = 1'b0;
assign s257 = 1'b0;
assign s258 = 1'b0;
assign s259 = 1'b0;
assign s260 = 1'b0;
assign s261 = 1'b0;
assign s262 = 1'b0;
assign s263 = 1'b0;
assign s264 = 1'b0;
assign s265 = 1'b0;
assign s266 = 1'b0;
assign s267 = 1'b0;
assign s268 = 1'b0;
assign s269 = 1'b0;
assign s270 = 1'b0;
assign s271 = 1'b0;
assign s272 = 1'b0;
assign s273 = 1'b0;
assign s274 = 1'b0;
assign s275 = 1'b0;
assign s276 = 1'b0;
assign s277 = 1'b0;
assign s278 = 1'b0;
assign s279 = 1'b0;
assign s280 = 1'b0;
assign s281 = 1'b0;
assign s282 = 1'b0;
assign s283 = 1'b0;
assign s284 = 1'b0;
assign s285 = 1'b0;
assign s286 = 1'b0;
assign s287 = 1'b0;
assign s288 = 1'b0;
assign s289 = 1'b0;
assign s290 = 1'b0;
assign s291 = 1'b0;
assign s292 = 1'b0;
assign s293 = 1'b0;
assign s294 = 1'b0;
assign s295 = 1'b0;
assign s296 = 1'b0;
assign s297 = 1'b0;
assign s298 = 1'b0;
assign s299 = 1'b0;
assign s300 = 1'b0;
assign s301 = 1'b0;
assign s302 = 1'b0;
assign s303 = 1'b0;
assign s304 = 1'b0;
assign s305 = 1'b0;
assign s306 = 1'b0;
assign s307 = 1'b0;
assign s308 = 1'b0;
assign s309 = 1'b0;
assign s310 = 1'b0;
assign s311 = 1'b0;
assign s312 = 1'b0;
assign s313 = 1'b0;
assign s314 = 1'b0;
assign s315 = 1'b0;
assign s316 = 1'b0;
assign s317 = 1'b0;
assign s318 = 1'b0;
assign s319 = 1'b0;
assign s320 = 1'b0;
assign s321 = 1'b0;
assign s322 = 1'b0;
assign s323 = 1'b0;
assign s324 = 1'b0;
assign s325 = 1'b0;
assign s326 = 1'b0;
assign s327 = 1'b0;
assign s328 = 1'b0;
assign instr_legal_dsp = ~csr_mmisc_ctl_rvcompm & (s0 | s1 | s2 | s3 | s4 | s5 | s6 | s7 | s8 | s9 | s10 | s11 | s12 | s13 | s14 | s15 | s16 | s17 | s18 | s19 | s20 | s21 | s22 | s23 | s24 | s25 | s26 | s27 | s28 | s29 | s30 | s31 | s32 | s33 | s34 | s35 | s36 | s37 | s38 | s39 | s40 | s41 | s42 | s43 | s44 | s45 | s46 | s47 | s48 | s49 | s50 | s51 | s52 | s53 | s54 | s55 | s56 | s57 | s58 | s59 | s60 | s61 | s62 | s63 | s64 | s65 | s66 | s67 | s68 | s69 | s70 | s71 | s72 | s73 | s74 | s75 | s76 | s77 | s78 | s79 | s80 | s81 | s82 | s83 | s84 | s85 | s86 | s87 | s88 | s89 | s90 | s91 | s92 | s93 | s94 | s95 | s96 | s97 | s98 | s99 | s100 | s101 | s102 | s103 | s104 | s105 | s106 | s107 | s108 | s109 | s110 | s111 | s112 | s113 | s114 | s115 | s117 | s116 | s118 | s119 | s120 | s121 | s122 | s123 | s124 | s125 | s126 | s127 | s128 | s129 | s130 | s131 | s132 | s133 | s134 | s135 | s136 | s137 | s138 | s139 | s140 | s141 | s142 | s143 | s144 | s145 | s146 | s147 | s148 | s149 | s150 | s151 | s152 | s153 | s154 | s155 | s156 | s157 | s158 | s159 | s160 | s161 | s162 | s163 | s164 | s165 | s166 | s167 | s168 | s169 | s170 | s171 | s172 | s173 | s174 | s175 | s176 | s177 | s178 | s179 | s180 | s181 | s182 | s183 | s184 | s185 | s186 | s187 | s188 | s189 | s190 | s191 | s192 | s193 | s194 | s195 | s196 | s197 | s198 | s199 | s200 | s201 | s202 | s203 | s204 | s205 | s206 | s207 | s208 | s209 | s210 | s211 | s212 | s213 | s214 | s215 | s216 | s217 | s218 | s219 | s220 | s221 | s222 | s223 | s224 | s225 | s226 | s227 | s228 | s229 | s230 | s231 | s232 | s233 | s234 | s235 | s236 | s237 | s238 | s239 | s240 | s241 | s242 | s243 | s244 | s245 | s246 | s247 | s248 | s249 | s250 | s251 | s252 | s253 | s254 | s255 | s256 | s257 | s258 | s259 | s260 | s261 | s262 | s263 | s264 | s265 | s266 | s267 | s268 | s269 | s270 | s271 | s272 | s273 | s274 | s275 | s276 | s277 | s278 | s279 | s280 | s281 | s282 | s283 | s284 | s285 | s286 | s287 | s288 | s289 | s290 | s291 | s292 | s293 | s294 | s295 | s296 | s297 | s298 | s299 | s300 | s301 | s302 | s303 | s304 | s305 | s306 | s307 | s308 | s309 | s310 | s311 | s312 | s313 | s314 | s315 | s316 | s317 | s318 | s319 | s320 | s321 | s322 | s323 | s324 | s325 | s326 | s327 | s328);
assign rs1_ren = instr_dsp;
assign rs2_ren = instr_dsp & !(s303 | s277 | s290 | s307 | s306 | s302 | s301 | s20 | s241 | s5 | s197 | s121 | s75 | s166 | s247 | s246 | s245 | s244 | s243 | s192 | s191 | s190 | s189 | s188 | s7 | s10 | s13 | s193 | s195 | s119 | s77 | s127 | s178 | s177 | s170 | s169 | s8 | s11 | s14 | s194 | s196 | s120 | s79 | s129 | s182 | s181 | s174 | s173 | s9 | s12 | s15);
assign rs3_ren = s260 | s259 | s258 | s275 | s274 | s272 | s273 | s271 | s268 | s267 | s266 | s265 | s264 | s36 | s35 | s34 | s159 | s158 | s137 | s138 | s136 | s135 | s134 | s133 | s132 | s131 | s210 | s73 | s224 | s160 | s209 | s52 | s218 | s139 | s102 | s141 | s219 | s140 | s72 | s71 | s50 | s51 | s49 | s48 | s47 | s46 | s45 | s44 | s64 | s63 | s60 | s59 | s62 | s61 | s58 | s57 | s98 | s95 | s66 | s65 | s56 | s55 | s20 | s6 | s215 | s90 | s239 | s117 | s187 | s204 | s26 | s231 | s109 | s2 | s130 | s241 | s242;
assign rs4_ren = s159 | s158 | s137 | s138 | s136 | s135 | s134 | s133 | s132 | s131 | s210 | s73 | s224 | s160 | s209 | s52 | s218 | s139 | s215 | s90 | s239 | s117 | s187 | s204 | s26 | s231 | s109 | s2;
assign rs1_addr = ({5{s333}} & s346) | ({5{s332}} & s354);
assign rs2_addr = ({5{s336}} & s352) | ({5{s335}} & s348) | ({5{s334}} & s355);
assign rs3_addr = ({5{s340}} & s353) | ({5{s339}} & s350) | ({5{s338}} & s347) | ({5{s337}} & s357);
assign rs4_addr = ({5{s342}} & s349) | ({5{s341}} & s358);
assign rd1_wen = instr_dsp;
assign rd2_wen = s159 | s158 | s137 | s138 | s136 | s135 | s134 | s133 | s132 | s131 | s210 | s73 | s224 | s160 | s209 | s52 | s218 | s139 | s215 | s90 | s239 | s117 | s187 | s204 | s26 | s231 | s109 | s2 | s100 | s99 | s226 | s225 | s162 | s161 | s228 | s227 | s164 | s163 | s130;
assign rd1_addr = ({5{s344}} & s350) | ({5{s343}} & s356);
assign rd2_addr = ({5{s345}} & s359);
assign s329 = instr_dsp & !(s330 | s331);
assign s330 = s152 | s153 | s55 | s56 | s65 | s66 | s93 | s94 | s95 | s98 | s154 | s155 | s156 | s157 | s57 | s58 | s61 | s62 | s67 | s68 | s69 | s70 | s59 | s60 | s63 | s64 | s53 | s54 | s147 | s149 | s148 | s44 | s45 | s46 | s47 | s48 | s49 | s51 | s50 | s71 | s72 | s140 | s219 | s141 | s101 | s102 | s99 | s100 | s34 | s35 | s36 | s292 | s293 | s294 | s258 | s259 | s260 | s39 | s40 | s144 | s145 | s146 | s163 | s164 | s227 | s228 | s41 | s42 | s43 | s31 | s32 | s33 | s261 | s262 | s263 | s255 | s256 | s257;
assign s331 = s130 | s139 | s218 | s52 | s209 | s160 | s224 | s73 | s210 | s131 | s132 | s133 | s134 | s135 | s136 | s138 | s137 | s158 | s159 | s269 | s270 | s295 | s297 | s296 | s264 | s265 | s266 | s267 | s268 | s271 | s273 | s272 | s274 | s275;
assign ready_stage = {s331,s330,s329};
assign s332 = instr_dsp & !s333;
assign s333 = s215 | s90 | s239 | s117 | s187 | s204 | s26 | s231 | s109 | s2 | s130 | s241 | s242;
assign s334 = instr_dsp & !(s335 | s336);
assign s335 = s215 | s90 | s239 | s117 | s187 | s204 | s26 | s231 | s109 | s2;
assign s336 = s251 | s23 | s21 | s22;
assign s337 = instr_dsp & !(s338 | s339 | s340);
assign s338 = s215 | s90 | s239 | s117 | s187 | s204 | s26 | s231 | s109 | s2 | s130 | s241 | s242;
assign s339 = s159 | s158 | s137 | s138 | s136 | s135 | s134 | s133 | s132 | s131 | s210 | s73 | s224 | s160 | s209 | s52 | s218 | s139;
assign s340 = s6;
assign s341 = instr_dsp & !s342;
assign s342 = s215 | s90 | s239 | s117 | s187 | s204 | s26 | s231 | s109 | s2;
assign s343 = instr_dsp & !s344;
assign s344 = s159 | s158 | s137 | s138 | s136 | s135 | s134 | s133 | s132 | s131 | s210 | s73 | s224 | s160 | s209 | s52 | s218 | s139 | s215 | s90 | s239 | s117 | s187 | s204 | s26 | s231 | s109 | s2 | s100 | s99 | s226 | s225 | s162 | s161 | s228 | s227 | s164 | s163 | s130;
assign s345 = instr_dsp;
assign s346 = {instr[19:16],1'b0};
assign s347 = {instr[19:16],1'b1};
assign s348 = {instr[24:21],1'b0};
assign s349 = {instr[24:21],1'b1};
assign s350 = {instr[11:8],1'b0};
assign s351 = {instr[11:8],1'b1};
assign s352 = 5'd0;
assign s353 = instr[29:25];
assign s354 = instr[19:15];
assign s355 = instr[24:20];
assign s356 = instr[11:7];
assign s357 = s356;
assign s358 = s351;
assign s359 = s351;
endmodule

