// Copyright (C) 2022, Andes Technology Corp. Confidential Proprietary

module kv_mini_dec (
    pp16_support,
    instr_retire,
    instr,
    instr_exec_it,
    instr_pp,
    reso_info,
    pp_ecnt,
    instr_event,
    trace_itype
);
input pp16_support;
input instr_retire;
input [31:0] instr;
input instr_exec_it;
input instr_pp;
input [12:0] reso_info;
input [7:0] pp_ecnt;
output [40:0] instr_event;
output [15:0] trace_itype;
localparam OP_LOAD = 7'b0000011;
localparam OP_IMM = 7'b0010011;
localparam OP_AUIPC = 7'b0010111;
localparam OP_IMM32 = 7'b0011011;
localparam OP_STORE = 7'b0100011;
localparam OP_ATOMIC = 7'b0101111;
localparam OP_OP = 7'b0110011;
localparam OP_LUI = 7'b0110111;
localparam OP_OP32 = 7'b0111011;
localparam OP_BRANCH = 7'b1100011;
localparam OP_JALR = 7'b1100111;
localparam OP_JAL = 7'b1101111;
localparam OP_SYSTEM = 7'b1110011;
localparam OP_DSP = 7'b1111111;
localparam OP_FP_LOAD = 7'b0000111;
localparam OP_FP_STORE = 7'b0100111;
localparam OP_FP = 7'b1010011;
localparam OP_FP_MADD = 7'b1000011;
localparam OP_FP_MSUB = 7'b1000111;
localparam OP_FP_NMADD = 7'b1001111;
localparam OP_FP_NMSUB = 7'b1001011;
localparam FPU_ADD = 5'b00000;
localparam FPU_SUB = 5'b00001;
localparam FPU_MUL = 5'b00010;
localparam FPU_DIV = 5'b00011;
localparam FPU_SQRT = 5'b01011;
localparam ATOMIC_LR = 5'b00010;
localparam ATOMIC_SC = 5'b00011;
localparam OP_C0 = 2'b00;
localparam OP_C1 = 2'b01;
localparam OP_C2 = 2'b10;
localparam OP_CUSTOM0 = 7'b0001011;
localparam OP_CUSTOM1 = 7'b0101011;
localparam OP_CUSTOM2 = 7'b1011011;


wire s0 = reso_info[0];
wire [4:0] s1 = instr[11:7];
wire [4:0] s2 = instr[19:15];
wire s3 = (s1 == 5'd1) | (s1 == 5'd5);
wire s4 = (s2 == 5'd1) | (s2 == 5'd5);
wire [4:0] s5 = instr[11:7];
wire [4:0] s6 = instr[11:7];
wire [4:0] s7 = instr[6:2];
wire s8 = (s5 == 5'd1) | (s5 == 5'd5);
wire s9 = (instr[6:0] == OP_LOAD);
wire s10 = (instr[6:0] == OP_STORE);
wire s11 = (instr[6:0] == OP_ATOMIC);
wire s12 = (instr[6:0] == OP_ATOMIC) & (instr[31:27] == ATOMIC_LR);
wire s13 = (instr[6:0] == OP_ATOMIC) & (instr[31:27] == ATOMIC_SC);
wire s14 = (instr[6:0] == OP_JAL);
wire s15 = (instr[6:0] == OP_JALR);
wire s16 = (instr[6:0] == OP_FP_LOAD);
wire s17 = (instr[6:0] == OP_FP_STORE);
wire s18 = (instr[6:0] == OP_FP_MADD);
wire s19 = (instr[6:0] == OP_FP_MSUB);
wire s20 = (instr[6:0] == OP_FP_NMADD);
wire s21 = (instr[6:0] == OP_FP_NMSUB);
wire s22 = (instr[6:0] == OP_FP) & (instr[31:27] == FPU_ADD);
wire s23 = (instr[6:0] == OP_FP) & (instr[31:27] == FPU_SUB);
wire s24 = (instr[6:0] == OP_FP) & (instr[31:27] == FPU_MUL);
wire s25 = (instr[6:0] == OP_FP) & (instr[31:27] == FPU_DIV);
wire s26 = (instr[6:0] == OP_FP) & (instr[31:27] == FPU_SQRT);
wire s27 = (instr[6:0] == OP_CUSTOM2) & (instr[31:25] == 7'b0000000) & (instr[19:12] == 8'b00010100);
wire s28 = (instr[6:0] == OP_CUSTOM2) & (instr[31:25] == 7'b0000000) & (instr[19:12] == 8'b00011100);
wire s29 = ((instr[6:0] == OP_FP) & ~s22 & ~s23 & ~s24 & ~s25 & ~s26) | s27 | s28;
wire s30 = (instr[6:0] == OP_BRANCH);
wire s31 = (instr[6:0] == OP_OP) & (instr[14] == 1'b0) & (instr[31:25] == 7'b0000001);
wire s32 = (instr[6:0] == OP_OP) & (instr[14] == 1'b1) & (instr[31:25] == 7'b0000001);
wire s33 = 1'b0;
wire s34 = 1'b0;
wire s35 = s31 | s33;
wire s36 = s32 | s34;
wire s37 = (instr[6:0] == OP_DSP);
wire s38 = (instr[31:25] == 7'b0000101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s39 = (instr[31:25] == 7'b0001101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s40 = (instr[31:25] == 7'b0010101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s41 = (instr[31:25] == 7'b1101001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s42 = (instr[31:25] == 7'b1110001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s43 = (instr[31:25] == 7'b1111001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s44 = (instr[31:25] == 7'b1000111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s45 = (instr[31:25] == 7'b1001111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s46 = (instr[31:25] == 7'b1000011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s47 = (instr[31:25] == 7'b1001011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s48 = (instr[31:25] == 7'b0000110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s49 = (instr[31:25] == 7'b0001110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s50 = (instr[31:25] == 7'b0010110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s51 = (instr[31:25] == 7'b0101101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s52 = (instr[31:25] == 7'b0110101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s53 = (instr[31:25] == 7'b0111101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s54 = (instr[31:25] == 7'b0100100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s55 = (instr[31:25] == 7'b0100101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s56 = (instr[31:25] == 7'b0101110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s57 = (instr[31:25] == 7'b0110110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s58 = (instr[31:25] == 7'b0111110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s59 = (instr[31:25] == 7'b1001010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s60 = (instr[31:25] == 7'b0011100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s61 = (instr[31:25] == 7'b0011101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s62 = (instr[31:25] == 7'b0110000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s63 = (instr[31:25] == 7'b0111000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s64 = (instr[31:25] == 7'b0100011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s65 = (instr[31:25] == 7'b0101011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s66 = (instr[31:25] == 7'b1100111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s67 = (instr[31:25] == 7'b1101111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s68 = (instr[31:25] == 7'b0110011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s69 = (instr[31:25] == 7'b0111011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s70 = (instr[31:25] == 7'b1110111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s71 = (instr[31:25] == 7'b1111111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s72 = (instr[31:25] == 7'b0100001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s73 = (instr[31:25] == 7'b0101001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s74 = (instr[31:25] == 7'b1000111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s75 = (instr[31:25] == 7'b1001111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s76 = (instr[31:25] == 7'b1010111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s77 = (instr[31:25] == 7'b1011111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s78 = (instr[31:25] == 7'b0100110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s79 = (instr[31:25] == 7'b0100111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s80 = (instr[31:25] == 7'b1001011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s81 = (instr[31:25] == 7'b0110001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s82 = (instr[31:25] == 7'b0111001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s83 = (instr[31:25] == 7'b1100010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s84 = (instr[31:25] == 7'b1100011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s85 = (instr[31:25] == 7'b1111000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s86 = (instr[31:25] == 7'b1110000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s87 = (instr[31:25] == 7'b0101111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s88 = (instr[31:25] == 7'b1000100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s89 = (instr[31:25] == 7'b1001100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s90 = (instr[31:25] == 7'b1010100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s91 = (instr[31:25] == 7'b1000110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s92 = (instr[31:25] == 7'b1001110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s93 = (instr[31:25] == 7'b1000101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s94 = (instr[31:25] == 7'b1001101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s95 = (instr[31:25] == 7'b1010101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s96 = (instr[31:25] == 7'b1000010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s97 = (instr[31:25] == 7'b1100100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s98 = (instr[31:25] == 7'b1100101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s99 = (instr[31:25] == 7'b0000100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s100 = (instr[31:25] == 7'b0001100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s101 = (instr[31:25] == 7'b0010100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s102 = (instr[31:25] == 7'b0101100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s103 = (instr[31:25] == 7'b0110100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s104 = (instr[31:25] == 7'b0111100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s105 = (instr[31:25] == 7'b0100000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s106 = (instr[31:25] == 7'b0101000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s107 = (instr[31:25] == 7'b0100010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s108 = (instr[31:25] == 7'b0101010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s109 = (instr[31:25] == 7'b0110010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s110 = (instr[31:25] == 7'b0111010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s111 = (instr[31:25] == 7'b1010110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s112 = (instr[31:25] == 7'b1011110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s113 = (instr[31:25] == 7'b1000011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s114 = (instr[31:25] == 7'b1010100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s115 = (instr[31:25] == 7'b1010101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s116 = (instr[31:25] == 7'b1010000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s117 = (instr[31:25] == 7'b1010001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s118 = (instr[31:25] == 7'b1011010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s119 = (instr[31:25] == 7'b1011011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s120 = (instr[31:25] == 7'b1010010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s121 = (instr[31:25] == 7'b1100110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s122 = (instr[31:25] == 7'b1010011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
wire s123 = (instr[31:25] == 7'b1011100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s124 = (instr[31:25] == 7'b1011101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s125 = (instr[31:25] == 7'b1011000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s126 = (instr[31:25] == 7'b1011001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
wire s127 = 1'b0;
wire s128 = 1'b0;
wire s129 = 1'b0;
wire s130 = 1'b0;
wire s131 = 1'b0;
wire s132 = 1'b0;
wire s133 = 1'b0;
wire s134 = 1'b0;
wire s135 = 1'b0;
wire s136 = 1'b0;
wire s137 = 1'b0;
wire s138 = 1'b0;
wire s139 = 1'b0;
wire s140 = 1'b0;
wire s141 = 1'b0;
wire s142 = 1'b0;
wire s143 = 1'b0;
wire s144 = 1'b0;
wire s145 = 1'b0;
wire s146 = 1'b0;
wire s147 = 1'b0;
wire s148 = 1'b0;
wire s149 = 1'b0;
wire s150 = 1'b0;
wire s151 = 1'b0;
wire s152 = 1'b0;
wire s153 = 1'b0;
wire s154 = s46 | s47 | s44 | s45 | s105 | s106 | s81 | s82 | s107 | s108 | s109 | s110 | s74 | s75 | s76 | s77 | s99 | s100 | s101 | s116 | s117 | s125 | s126 | s114 | s115 | s123 | s124 | s85 | s86 | s48 | s49 | s50 | s38 | s39 | s40 | s148 | s149 | s150 | s133 | s134 | s135 | s127 | s128 | s129;
wire s155 = s62 | s63 | s72 | s73 | s83 | s84 | s64 | s65 | s68 | s69 | s66 | s67 | s70 | s71 | s60 | s61 | s102 | s104 | s103 | s51 | s52 | s53 | s54 | s55 | s56 | s58 | s57 | s78 | s79 | s87 | s97 | s121 | s98 | s96 | s120 | s59 | s118 | s113 | s122 | s80 | s119 | s88 | s89 | s90 | s91 | s92 | s93 | s95 | s94 | s111 | s112 | s41 | s42 | s43 | s141 | s142 | s151 | s153 | s152 | s136 | s137 | s138 | s139 | s140 | s143 | s145 | s144 | s146 | s147 | s130 | s131 | s132;
wire s156 = s37 & !(s154 | s155);
wire s157 = (instr[1:0] == OP_C2) & (instr[15:13] == 3'b010);
wire s158 = (instr[1:0] == OP_C2) & (instr[15:13] == 3'b110);
wire s159 = (instr[1:0] == OP_C0) & (instr[15:13] == 3'b010);
wire s160 = (instr[1:0] == OP_C0) & (instr[15:13] == 3'b110);
wire s161 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b101);
wire s162 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b001);
wire s163 = (instr[1:0] == OP_C2) & (instr[12] == 1'b0) & (instr[15:13] == 3'b100) & (s7 == 5'b0);
wire s164 = (instr[1:0] == OP_C2) & (instr[12] == 1'b1) & (instr[15:13] == 3'b100) & (s7 == 5'b0) & (s5 != 5'b0);
wire s165 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b110);
wire s166 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b111);
wire s167 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b010);
wire s168 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b011) & (s6 != 5'b00010);
wire s169 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b000);
wire s170 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b011) & (s6 == 5'b00010);
wire s171 = (instr[1:0] == OP_C0) & (instr[15:13] == 3'b000);
wire s172 = (instr[1:0] == OP_C2) & (instr[15:13] == 3'b000);
wire s173 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b100) & (instr[11:10] == 2'b00);
wire s174 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b100) & (instr[11:10] == 2'b01);
wire s175 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b100) & (instr[11:10] == 2'b10);
wire s176 = (instr[1:0] == OP_C2) & (instr[15:13] == 3'b100) & (instr[12] == 1'b0) & (s7 != 5'b0);
wire s177 = (instr[1:0] == OP_C2) & (instr[15:13] == 3'b100) & (instr[12] == 1'b1) & (s7 != 5'b0);
wire s178 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b100) & (instr[12:10] == 3'b011) & (instr[6:5] == 2'b11);
wire s179 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b100) & (instr[12:10] == 3'b011) & (instr[6:5] == 2'b10);
wire s180 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b100) & (instr[12:10] == 3'b011) & (instr[6:5] == 2'b01);
wire s181 = (instr[1:0] == OP_C1) & (instr[15:13] == 3'b100) & (instr[12:10] == 3'b011) & (instr[6:5] == 2'b00);
wire s182 = (instr[1:0] == OP_C2) & (instr[15:2] == 14'h2400);
wire s183 = instr_exec_it;
wire s184 = 1'b0;
wire s185 = 1'b0;
wire s186 = 1'b0;
wire s187 = 1'b0;
wire s188 = 1'b0;
wire s189 = 1'b0;
wire s190 = 1'b0;
wire s191 = (instr[1:0] == OP_C2) & (instr[15:13] == 3'b011);
wire s192 = (instr[1:0] == OP_C2) & (instr[15:13] == 3'b001) & ~pp16_support;
wire s193 = (instr[1:0] == OP_C0) & (instr[15:13] == 3'b011);
wire s194 = (instr[1:0] == OP_C0) & (instr[15:13] == 3'b001) & ~pp16_support;
wire s195 = (instr[1:0] == OP_C2) & (instr[15:13] == 3'b111);
wire s196 = (instr[1:0] == OP_C2) & (instr[15:13] == 3'b101) & ~pp16_support;
wire s197 = (instr[1:0] == OP_C0) & (instr[15:13] == 3'b111);
wire s198 = (instr[1:0] == OP_C0) & (instr[15:13] == 3'b101) & ~pp16_support;
wire s199 = pp16_support & instr_pp & (instr[6:5] == 2'b10);
wire s200 = pp16_support & instr_pp & (instr[6:5] == 2'b00);
wire s201 = pp16_support & instr_pp & (instr[6:5] == 2'b01);
wire s202 = pp16_support & (instr[1:0] == OP_C2) & (instr[15:13] == 3'b001);
wire s203 = pp16_support & (instr[1:0] == OP_C0) & (instr[15:13] == 3'b001);
wire s204 = pp16_support & (instr[1:0] == OP_C2) & (instr[15:13] == 3'b101);
wire s205 = pp16_support & (instr[1:0] == OP_C0) & (instr[15:13] == 3'b101);
wire s206 = s157 | s184 | s159 | s186 | s202 | s203;
wire s207 = s158 | s185 | s160 | s187 | s204 | s205;
wire s208 = s191 | s192 | s193 | s194;
wire s209 = s195 | s196 | s197 | s198;
wire s210 = s161 | s162 | s163 | s164;
wire s211 = s165 | s166;
wire s212 = s167 | s168 | s169 | s188 | s170 | s171 | s172 | s173 | s174 | s175 | s176 | s177 | s178 | s179 | s180 | s181 | s189 | s190;
wire s213 = (instr[6:0] == OP_CUSTOM0) & (instr[13:12] == 2'b00);
wire s214 = (instr[6:0] == OP_CUSTOM0) & (instr[13:12] == 2'b10);
wire s215 = (instr[6:0] == OP_CUSTOM1) & (instr[14:12] == 3'b001);
wire s216 = (instr[6:0] == OP_CUSTOM1) & (instr[14:12] == 3'b101);
wire s217 = (instr[6:0] == OP_CUSTOM1) & (instr[14:12] == 3'b010);
wire s218 = 1'b0;
wire s219 = 1'b0;
wire s220 = (instr[6:0] == OP_CUSTOM0) & (instr[13:12] == 2'b11);
wire s221 = (instr[6:0] == OP_CUSTOM1) & (instr[14:12] == 3'b000);
wire s222 = (instr[6:0] == OP_CUSTOM1) & (instr[14:12] == 3'b100);
wire s223 = 1'b0;
wire s224 = s214 | s213 | s215 | s216 | s217 | s218 | s219;
wire s225 = s220 | s221 | s222 | s223;
wire s226 = (instr[6:0] == OP_CUSTOM0) & (instr[13:12] == 2'b01);
wire s227 = (instr[6:0] == OP_CUSTOM2) & (instr[14:12] == 3'b000) & (instr[31:25] == 7'b0000101);
wire s228 = (instr[6:0] == OP_CUSTOM2) & (instr[14:12] == 3'b000) & (instr[31:25] == 7'b0000110);
wire s229 = (instr[6:0] == OP_CUSTOM2) & (instr[14:12] == 3'b000) & (instr[31:25] == 7'b0000111);
wire s230 = 1'b0;
wire s231 = s227 | s228 | s229 | s230;
wire s232 = (instr[6:0] == OP_CUSTOM2) & (instr[14:12] == 3'b000) & (instr[31:27] == 5'b00100);
wire s233 = (instr[6:0] == OP_CUSTOM2) & (instr[14:12] == 3'b111) & ((instr[7] == 1'b0));
wire s234 = (instr[6:0] == OP_CUSTOM2) & (instr[14:12] == 3'b101);
wire s235 = (instr[6:0] == OP_CUSTOM2) & (instr[14:12] == 3'b110);
wire s236 = (instr[6:0] == OP_CUSTOM2) & (instr[14:12] == 3'b011) & ((instr[25] == 1'b0)) & ((instr[31] == 1'b0));
wire s237 = (instr[6:0] == OP_CUSTOM2) & (instr[14:12] == 3'b010) & ((instr[25] == 1'b0)) & ((instr[31] == 1'b0));
wire s238 = s236 | s237;
wire s239 = s233 | s234 | s235;
wire s240 = (instr[6:0] == OP_SYSTEM) | s182;
wire s241 = (((instr[6:0] == OP_IMM) | ((instr[6:0] == OP_OP) & (~s31 & ~s32)) | (instr[6:0] == OP_LUI) | (instr[6:0] == OP_AUIPC))) | s226 | s231 | s232 | s238;
wire s242 = (s15 & s4 & (~s3 | (s2 != s1)) & (instr[31:20] == 12'd0)) | (s164 & s8 & (s5 != 5'd1)) | (s163 & s8);
wire s243 = (s30 | s211 | s239);
assign instr_event[21] = instr_retire & (s9 | s12 | s206 | s224 | s200 | s201);
assign instr_event[39] = instr_retire & (s10 | s13 | s207 | s225 | s199);
assign instr_event[1] = instr_retire & (s11 & ~s12 & ~s13);
assign instr_event[40] = instr_retire & (s240);
assign instr_event[0] = instr_retire & (s241 | s212 | s156 | instr_pp);
assign instr_event[19] = instr_retire & (s14 | s162 | s161);
assign instr_event[20] = instr_retire & (s15 | s164 | s163 | s201);
assign instr_event[6] = instr_retire & (s243 | s14 | s15 | s210 | s201);
assign instr_event[24] = instr_retire & (s35 | s154);
assign instr_event[23] = instr_retire & (s155);
assign instr_event[8] = instr_retire & (s36);
assign instr_event[13] = instr_retire & (s16 | s208);
assign instr_event[16] = instr_retire & (s17 | s209);
assign instr_event[10] = instr_retire & (s22 | s23);
assign instr_event[14] = instr_retire & (s24);
assign instr_event[12] = instr_retire & (s18 | s19 | s20 | s21);
assign instr_event[11] = instr_retire & (s25 | s26);
assign instr_event[15] = instr_retire & (s29);
assign instr_event[2] = instr_retire & (s243);
assign instr_event[3] = instr_retire & (s243) & reso_info[11];
assign instr_event[4] = instr_retire & (s243) & reso_info[0];
assign instr_event[5] = instr_retire & (s243) & reso_info[0] & reso_info[11];
assign instr_event[37] = instr_retire & (s242 | s201);
assign instr_event[38] = instr_retire & (s242 | s201) & reso_info[11];
assign instr_event[9] = instr_retire & (s183);
assign instr_event[22] = 1'b0;
assign instr_event[7] = 1'b0;
assign instr_event[17] = 1'b0;
assign instr_event[18] = 1'b0;
assign instr_event[27] = instr_retire & (instr_pp);
assign instr_event[36] = instr_retire & (s199);
assign instr_event[25] = instr_retire & (s200);
assign instr_event[26] = instr_retire & (s201);
assign instr_event[28 +:4] = {4{instr_pp}} & pp_ecnt[0 +:4];
assign instr_event[32 +:4] = {4{instr_pp}} & pp_ecnt[4 +:4];
wire s244 = s243 & ~s0;
wire s245 = s243 & s0;
wire s246 = (s14 & ((s1 == 5'd1) | (s1 == 5'd5))) | s162;
wire s247 = (s14 & (s1 == 5'd0)) | s161;
wire s248 = (s15 & (s1 == 5'd1) & (s2 != 5'd5)) | (s15 & (s1 == 5'd5) & (s2 != 5'd1)) | (s164 & (s5 != 5'd5));
wire s249 = (s15 & (s1 == 5'd0) & (s2 != 5'd1) & (s2 != 5'd5)) | (s163 & (s5 != 5'd1) & (s5 != 5'd5));
wire s250 = (s15 & (s1 != 5'd1) & (s1 != 5'd5) & ((s2 == 5'd1) | (s2 == 5'd5))) | (s163 & ((s5 == 5'd1) | (s5 == 5'd5)));
wire s251 = (s15 & (s1 == 5'd1) & (s2 == 5'd5)) | (s15 & (s1 == 5'd5) & (s2 == 5'd1)) | (s164 & (s5 == 5'd5));
wire s252 = (s14 & (s1 != 5'd0) & (s1 != 5'd1) & (s1 != 5'd5));
wire s253 = (s15 & (s1 != 5'd0) & (s1 != 5'd1) & (s1 != 5'd5) & (s2 != 5'd1) & (s2 != 5'd5));
assign trace_itype[0] = 1'b0;
assign trace_itype[1] = 1'b0;
assign trace_itype[2] = 1'b0;
assign trace_itype[3] = 1'b0;
assign trace_itype[4] = s244;
assign trace_itype[5] = s245;
assign trace_itype[6] = 1'b0;
assign trace_itype[7] = 1'b0;
assign trace_itype[8] = s248;
assign trace_itype[9] = s246;
assign trace_itype[10] = s249;
assign trace_itype[11] = s247;
assign trace_itype[12] = s251;
assign trace_itype[13] = s250;
assign trace_itype[14] = s253;
assign trace_itype[15] = s252;
endmodule

