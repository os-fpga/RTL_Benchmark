--*************************************************************************
-- Project    : 16 Quadrature Amplitude Demodulator    	                  *
--                                                                        *
-- File Name  : QADM_16.vhd                                               *
--                                                                        *
-- Author     : Kaustubh Chaudhari                                        *
--                                                                        *
-- Email      : kaustubhcha305@gmail.com                                  *
--                                                                        *
-- Description: 16 QADM, requires 10 bit QAM i/p and gives 4 bit Demod o/p*
--                                                                        *
--*************************************************************************
--                                                                        *
-- Copyright (C) 2016 Author                                              *
--                                                                        *
-- This program is free software: you can redistribute it and/or modify   *
-- it under the terms of the GNU General Public License as published by   *
-- the Free Software Foundation, either version 3 of the License, or      *
-- (at your option) any later version.                                    *
--                                                                        *
-- This program is distributed in the hope that it will be useful,        *
-- but WITHOUT ANY WARRANTY; without even the implied warranty of         *
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the          *
-- GNU General Public License for more details.                           *
--                                                                        *
-- You should have received a copy of the GNU General Public License      *
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.  *
--*************************************************************************
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity QADM_16 is
PORT(output:  OUT  std_logic_vector(3 downto 0);  --4 bit output depending on i/p QAM wave
     clk:  IN  std_logic; --clock
	 inp: IN  std_logic_vector(9 downto 0) --input in 10bit resolution
    );
end QADM_16;

architecture Behavioral of QADM_16 is
type sine_array is array (0 to 2047) of integer range 0 to 1023;
signal sine1 : sine_array:=(512, 513, 514, 515, 515, 516, 517, 518, 519, 519, 520, 521, 522, 522, 523, 524, 
525, 526, 526, 527, 528, 529, 529, 530, 531, 532, 533, 533, 534, 535, 536, 536, 
537, 538, 539, 539, 540, 541, 542, 542, 543, 544, 545, 546, 546, 547, 548, 549, 
549, 550, 551, 551, 552, 553, 554, 554, 555, 556, 557, 557, 558, 559, 560, 560, 
561, 562, 562, 563, 564, 565, 565, 566, 567, 567, 568, 569, 570, 570, 571, 572, 
572, 573, 574, 574, 575, 576, 576, 577, 578, 578, 579, 580, 580, 581, 582, 582, 
583, 584, 584, 585, 586, 586, 587, 587, 588, 589, 589, 590, 591, 591, 592, 592, 
593, 594, 594, 595, 595, 596, 597, 597, 598, 598, 599, 599, 600, 601, 601, 602, 
602, 603, 603, 604, 604, 605, 605, 606, 606, 607, 608, 608, 609, 609, 610, 610, 
611, 611, 612, 612, 612, 613, 613, 614, 614, 615, 615, 616, 616, 617, 617, 618, 
618, 618, 619, 619, 620, 620, 620, 621, 621, 622, 622, 622, 623, 623, 624, 624, 
624, 625, 625, 625, 626, 626, 626, 627, 627, 627, 628, 628, 628, 629, 629, 629, 
630, 630, 630, 630, 631, 631, 631, 632, 632, 632, 632, 633, 633, 633, 633, 634, 
634, 634, 634, 634, 635, 635, 635, 635, 635, 636, 636, 636, 636, 636, 636, 637, 
637, 637, 637, 637, 637, 637, 638, 638, 638, 638, 638, 638, 638, 638, 638, 638, 
638, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 
639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 638, 638, 
638, 638, 638, 638, 638, 638, 638, 638, 638, 637, 637, 637, 637, 637, 637, 637, 
636, 636, 636, 636, 636, 636, 635, 635, 635, 635, 635, 634, 634, 634, 634, 634, 
633, 633, 633, 633, 632, 632, 632, 632, 631, 631, 631, 630, 630, 630, 630, 629, 
629, 629, 628, 628, 628, 627, 627, 627, 626, 626, 626, 625, 625, 625, 624, 624, 
624, 623, 623, 622, 622, 622, 621, 621, 620, 620, 620, 619, 619, 618, 618, 618, 
617, 617, 616, 616, 615, 615, 614, 614, 613, 613, 612, 612, 612, 611, 611, 610, 
610, 609, 609, 608, 608, 607, 606, 606, 605, 605, 604, 604, 603, 603, 602, 602, 
601, 601, 600, 599, 599, 598, 598, 597, 597, 596, 595, 595, 594, 594, 593, 592, 
592, 591, 591, 590, 589, 589, 588, 587, 587, 586, 586, 585, 584, 584, 583, 582, 
582, 581, 580, 580, 579, 578, 578, 577, 576, 576, 575, 574, 574, 573, 572, 572, 
571, 570, 570, 569, 568, 567, 567, 566, 565, 565, 564, 563, 562, 562, 561, 560, 
560, 559, 558, 557, 557, 556, 555, 554, 554, 553, 552, 551, 551, 550, 549, 549, 
548, 547, 546, 546, 545, 544, 543, 542, 542, 541, 540, 539, 539, 538, 537, 536, 
536, 535, 534, 533, 533, 532, 531, 530, 529, 529, 528, 527, 526, 526, 525, 524, 
523, 522, 522, 521, 520, 519, 519, 518, 517, 516, 515, 515, 514, 513, 512, 512, 
511, 510, 509, 508, 508, 507, 506, 505, 504, 504, 503, 502, 501, 501, 500, 499, 
498, 497, 497, 496, 495, 494, 494, 493, 492, 491, 490, 490, 489, 488, 487, 487, 
486, 485, 484, 484, 483, 482, 481, 481, 480, 479, 478, 477, 477, 476, 475, 474, 
474, 473, 472, 472, 471, 470, 469, 469, 468, 467, 466, 466, 465, 464, 463, 463, 
462, 461, 461, 460, 459, 458, 458, 457, 456, 456, 455, 454, 453, 453, 452, 451, 
451, 450, 449, 449, 448, 447, 447, 446, 445, 445, 444, 443, 443, 442, 441, 441, 
440, 439, 439, 438, 437, 437, 436, 436, 435, 434, 434, 433, 432, 432, 431, 431, 
430, 429, 429, 428, 428, 427, 426, 426, 425, 425, 424, 424, 423, 422, 422, 421, 
421, 420, 420, 419, 419, 418, 418, 417, 417, 416, 415, 415, 414, 414, 413, 413, 
412, 412, 411, 411, 411, 410, 410, 409, 409, 408, 408, 407, 407, 406, 406, 405, 
405, 405, 404, 404, 403, 403, 403, 402, 402, 401, 401, 401, 400, 400, 399, 399, 
399, 398, 398, 398, 397, 397, 397, 396, 396, 396, 395, 395, 395, 394, 394, 394, 
393, 393, 393, 393, 392, 392, 392, 391, 391, 391, 391, 390, 390, 390, 390, 389, 
389, 389, 389, 389, 388, 388, 388, 388, 388, 387, 387, 387, 387, 387, 387, 386, 
386, 386, 386, 386, 386, 386, 385, 385, 385, 385, 385, 385, 385, 385, 385, 385, 
385, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 
384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 385, 385, 
385, 385, 385, 385, 385, 385, 385, 385, 385, 386, 386, 386, 386, 386, 386, 386, 
387, 387, 387, 387, 387, 387, 388, 388, 388, 388, 388, 389, 389, 389, 389, 389, 
390, 390, 390, 390, 391, 391, 391, 391, 392, 392, 392, 393, 393, 393, 393, 394, 
394, 394, 395, 395, 395, 396, 396, 396, 397, 397, 397, 398, 398, 398, 399, 399, 
399, 400, 400, 401, 401, 401, 402, 402, 403, 403, 403, 404, 404, 405, 405, 405, 
406, 406, 407, 407, 408, 408, 409, 409, 410, 410, 411, 411, 411, 412, 412, 413, 
413, 414, 414, 415, 415, 416, 417, 417, 418, 418, 419, 419, 420, 420, 421, 421, 
422, 422, 423, 424, 424, 425, 425, 426, 426, 427, 428, 428, 429, 429, 430, 431, 
431, 432, 432, 433, 434, 434, 435, 436, 436, 437, 437, 438, 439, 439, 440, 441, 
441, 442, 443, 443, 444, 445, 445, 446, 447, 447, 448, 449, 449, 450, 451, 451, 
452, 453, 453, 454, 455, 456, 456, 457, 458, 458, 459, 460, 461, 461, 462, 463, 
463, 464, 465, 466, 466, 467, 468, 469, 469, 470, 471, 472, 472, 473, 474, 474, 
475, 476, 477, 477, 478, 479, 480, 481, 481, 482, 483, 484, 484, 485, 486, 487, 
487, 488, 489, 490, 490, 491, 492, 493, 494, 494, 495, 496, 497, 497, 498, 499, 
500, 501, 501, 502, 503, 504, 504, 505, 506, 507, 508, 508, 509, 510, 511, 512,
512, 513, 514, 515, 515, 516, 517, 518, 519, 519, 520, 521, 522, 522, 523, 524, 
525, 526, 526, 527, 528, 529, 529, 530, 531, 532, 533, 533, 534, 535, 536, 536, 
537, 538, 539, 539, 540, 541, 542, 542, 543, 544, 545, 546, 546, 547, 548, 549, 
549, 550, 551, 551, 552, 553, 554, 554, 555, 556, 557, 557, 558, 559, 560, 560, 
561, 562, 562, 563, 564, 565, 565, 566, 567, 567, 568, 569, 570, 570, 571, 572, 
572, 573, 574, 574, 575, 576, 576, 577, 578, 578, 579, 580, 580, 581, 582, 582, 
583, 584, 584, 585, 586, 586, 587, 587, 588, 589, 589, 590, 591, 591, 592, 592, 
593, 594, 594, 595, 595, 596, 597, 597, 598, 598, 599, 599, 600, 601, 601, 602, 
602, 603, 603, 604, 604, 605, 605, 606, 606, 607, 608, 608, 609, 609, 610, 610, 
611, 611, 612, 612, 612, 613, 613, 614, 614, 615, 615, 616, 616, 617, 617, 618, 
618, 618, 619, 619, 620, 620, 620, 621, 621, 622, 622, 622, 623, 623, 624, 624, 
624, 625, 625, 625, 626, 626, 626, 627, 627, 627, 628, 628, 628, 629, 629, 629, 
630, 630, 630, 630, 631, 631, 631, 632, 632, 632, 632, 633, 633, 633, 633, 634, 
634, 634, 634, 634, 635, 635, 635, 635, 635, 636, 636, 636, 636, 636, 636, 637, 
637, 637, 637, 637, 637, 637, 638, 638, 638, 638, 638, 638, 638, 638, 638, 638, 
638, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 
639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 639, 638, 638, 
638, 638, 638, 638, 638, 638, 638, 638, 638, 637, 637, 637, 637, 637, 637, 637, 
636, 636, 636, 636, 636, 636, 635, 635, 635, 635, 635, 634, 634, 634, 634, 634, 
633, 633, 633, 633, 632, 632, 632, 632, 631, 631, 631, 630, 630, 630, 630, 629, 
629, 629, 628, 628, 628, 627, 627, 627, 626, 626, 626, 625, 625, 625, 624, 624, 
624, 623, 623, 622, 622, 622, 621, 621, 620, 620, 620, 619, 619, 618, 618, 618, 
617, 617, 616, 616, 615, 615, 614, 614, 613, 613, 612, 612, 612, 611, 611, 610, 
610, 609, 609, 608, 608, 607, 606, 606, 605, 605, 604, 604, 603, 603, 602, 602, 
601, 601, 600, 599, 599, 598, 598, 597, 597, 596, 595, 595, 594, 594, 593, 592, 
592, 591, 591, 590, 589, 589, 588, 587, 587, 586, 586, 585, 584, 584, 583, 582, 
582, 581, 580, 580, 579, 578, 578, 577, 576, 576, 575, 574, 574, 573, 572, 572, 
571, 570, 570, 569, 568, 567, 567, 566, 565, 565, 564, 563, 562, 562, 561, 560, 
560, 559, 558, 557, 557, 556, 555, 554, 554, 553, 552, 551, 551, 550, 549, 549, 
548, 547, 546, 546, 545, 544, 543, 542, 542, 541, 540, 539, 539, 538, 537, 536, 
536, 535, 534, 533, 533, 532, 531, 530, 529, 529, 528, 527, 526, 526, 525, 524, 
523, 522, 522, 521, 520, 519, 519, 518, 517, 516, 515, 515, 514, 513, 512, 512, 
511, 510, 509, 508, 508, 507, 506, 505, 504, 504, 503, 502, 501, 501, 500, 499, 
498, 497, 497, 496, 495, 494, 494, 493, 492, 491, 490, 490, 489, 488, 487, 487, 
486, 485, 484, 484, 483, 482, 481, 481, 480, 479, 478, 477, 477, 476, 475, 474, 
474, 473, 472, 472, 471, 470, 469, 469, 468, 467, 466, 466, 465, 464, 463, 463, 
462, 461, 461, 460, 459, 458, 458, 457, 456, 456, 455, 454, 453, 453, 452, 451, 
451, 450, 449, 449, 448, 447, 447, 446, 445, 445, 444, 443, 443, 442, 441, 441, 
440, 439, 439, 438, 437, 437, 436, 436, 435, 434, 434, 433, 432, 432, 431, 431, 
430, 429, 429, 428, 428, 427, 426, 426, 425, 425, 424, 424, 423, 422, 422, 421, 
421, 420, 420, 419, 419, 418, 418, 417, 417, 416, 415, 415, 414, 414, 413, 413, 
412, 412, 411, 411, 411, 410, 410, 409, 409, 408, 408, 407, 407, 406, 406, 405, 
405, 405, 404, 404, 403, 403, 403, 402, 402, 401, 401, 401, 400, 400, 399, 399, 
399, 398, 398, 398, 397, 397, 397, 396, 396, 396, 395, 395, 395, 394, 394, 394, 
393, 393, 393, 393, 392, 392, 392, 391, 391, 391, 391, 390, 390, 390, 390, 389, 
389, 389, 389, 389, 388, 388, 388, 388, 388, 387, 387, 387, 387, 387, 387, 386, 
386, 386, 386, 386, 386, 386, 385, 385, 385, 385, 385, 385, 385, 385, 385, 385, 
385, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 
384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 384, 385, 385, 
385, 385, 385, 385, 385, 385, 385, 385, 385, 386, 386, 386, 386, 386, 386, 386, 
387, 387, 387, 387, 387, 387, 388, 388, 388, 388, 388, 389, 389, 389, 389, 389, 
390, 390, 390, 390, 391, 391, 391, 391, 392, 392, 392, 393, 393, 393, 393, 394, 
394, 394, 395, 395, 395, 396, 396, 396, 397, 397, 397, 398, 398, 398, 399, 399, 
399, 400, 400, 401, 401, 401, 402, 402, 403, 403, 403, 404, 404, 405, 405, 405, 
406, 406, 407, 407, 408, 408, 409, 409, 410, 410, 411, 411, 411, 412, 412, 413, 
413, 414, 414, 415, 415, 416, 417, 417, 418, 418, 419, 419, 420, 420, 421, 421, 
422, 422, 423, 424, 424, 425, 425, 426, 426, 427, 428, 428, 429, 429, 430, 431, 
431, 432, 432, 433, 434, 434, 435, 436, 436, 437, 437, 438, 439, 439, 440, 441, 
441, 442, 443, 443, 444, 445, 445, 446, 447, 447, 448, 449, 449, 450, 451, 451, 
452, 453, 453, 454, 455, 456, 456, 457, 458, 458, 459, 460, 461, 461, 462, 463, 
463, 464, 465, 466, 466, 467, 468, 469, 469, 470, 471, 472, 472, 473, 474, 474, 
475, 476, 477, 477, 478, 479, 480, 481, 481, 482, 483, 484, 484, 485, 486, 487, 
487, 488, 489, 490, 490, 491, 492, 493, 494, 494, 495, 496, 497, 497, 498, 499, 
500, 501, 501, 502, 503, 504, 504, 505, 506, 507, 508, 508, 509, 510, 511, 512);
signal sine2 : sine_array:=(512, 515, 516, 518, 519, 521, 522, 524, 526, 527, 529, 530, 532, 533, 535, 537, 
538, 540, 541, 543, 544, 546, 547, 549, 551, 552, 554, 555, 557, 558, 560, 561, 
563, 564, 566, 567, 569, 571, 572, 574, 575, 577, 578, 580, 581, 583, 584, 586, 
587, 589, 590, 592, 593, 595, 596, 598, 599, 601, 602, 603, 605, 606, 608, 609, 
611, 612, 614, 615, 616, 618, 619, 621, 622, 624, 625, 626, 628, 629, 631, 632, 
633, 635, 636, 637, 639, 640, 642, 643, 644, 646, 647, 648, 650, 651, 652, 653, 
655, 656, 657, 659, 660, 661, 662, 664, 665, 666, 667, 669, 670, 671, 672, 674, 
675, 676, 677, 678, 680, 681, 682, 683, 684, 685, 687, 688, 689, 690, 691, 692, 
693, 694, 695, 697, 698, 699, 700, 701, 702, 703, 704, 705, 706, 707, 708, 709, 
710, 711, 712, 713, 714, 715, 716, 717, 718, 719, 719, 720, 721, 722, 723, 724, 
725, 726, 727, 727, 728, 729, 730, 731, 731, 732, 733, 734, 735, 735, 736, 737, 
738, 738, 739, 740, 740, 741, 742, 742, 743, 744, 744, 745, 746, 746, 747, 748, 
748, 749, 749, 750, 750, 751, 752, 752, 753, 753, 754, 754, 755, 755, 756, 756, 
756, 757, 757, 758, 758, 759, 759, 759, 760, 760, 760, 761, 761, 761, 762, 762, 
762, 763, 763, 763, 764, 764, 764, 764, 764, 765, 765, 765, 765, 765, 766, 766, 
766, 766, 766, 766, 766, 767, 767, 767, 767, 767, 767, 767, 767, 767, 767, 767, 
767, 767, 767, 767, 767, 767, 767, 767, 767, 767, 766, 766, 766, 766, 766, 766, 
766, 765, 765, 765, 765, 765, 764, 764, 764, 764, 764, 763, 763, 763, 762, 762, 
762, 761, 761, 761, 760, 760, 760, 759, 759, 759, 758, 758, 757, 757, 756, 756, 
756, 755, 755, 754, 754, 753, 753, 752, 752, 751, 750, 750, 749, 749, 748, 748, 
747, 746, 746, 745, 744, 744, 743, 742, 742, 741, 740, 740, 739, 738, 738, 737, 
736, 735, 735, 734, 733, 732, 731, 731, 730, 729, 728, 727, 727, 726, 725, 724, 
723, 722, 721, 720, 719, 719, 718, 717, 716, 715, 714, 713, 712, 711, 710, 709, 
708, 707, 706, 705, 704, 703, 702, 701, 700, 699, 698, 697, 695, 694, 693, 692, 
691, 690, 689, 688, 687, 685, 684, 683, 682, 681, 680, 678, 677, 676, 675, 674, 
672, 671, 670, 669, 667, 666, 665, 664, 662, 661, 660, 659, 657, 656, 655, 653, 
652, 651, 650, 648, 647, 646, 644, 643, 642, 640, 639, 637, 636, 635, 633, 632, 
631, 629, 628, 626, 625, 624, 622, 621, 619, 618, 616, 615, 614, 612, 611, 609, 
608, 606, 605, 603, 602, 601, 599, 598, 596, 595, 593, 592, 590, 589, 587, 586, 
584, 583, 581, 580, 578, 577, 575, 574, 572, 571, 569, 567, 566, 564, 563, 561, 
560, 558, 557, 555, 554, 552, 551, 549, 547, 546, 544, 543, 541, 540, 538, 537, 
535, 533, 532, 530, 529, 527, 526, 524, 522, 521, 519, 518, 516, 515, 513, 512, 
510, 508, 507, 505, 504, 502, 501, 499, 497, 496, 494, 493, 491, 490, 488, 486, 
485, 483, 482, 480, 479, 477, 476, 474, 472, 471, 469, 468, 466, 465, 463, 462, 
460, 459, 457, 456, 454, 452, 451, 449, 448, 446, 445, 443, 442, 440, 439, 437, 
436, 434, 433, 431, 430, 428, 427, 425, 424, 422, 421, 420, 418, 417, 415, 414, 
412, 411, 409, 408, 407, 405, 404, 402, 401, 399, 398, 397, 395, 394, 392, 391, 
390, 388, 387, 386, 384, 383, 381, 380, 379, 377, 376, 375, 373, 372, 371, 370, 
368, 367, 366, 364, 363, 362, 361, 359, 358, 357, 356, 354, 353, 352, 351, 349, 
348, 347, 346, 345, 343, 342, 341, 340, 339, 338, 336, 335, 334, 333, 332, 331, 
330, 329, 328, 326, 325, 324, 323, 322, 321, 320, 319, 318, 317, 316, 315, 314, 
313, 312, 311, 310, 309, 308, 307, 306, 305, 304, 304, 303, 302, 301, 300, 299, 
298, 297, 296, 296, 295, 294, 293, 292, 292, 291, 290, 289, 288, 288, 287, 286, 
285, 285, 284, 283, 283, 282, 281, 281, 280, 279, 279, 278, 277, 277, 276, 275, 
275, 274, 274, 273, 273, 272, 271, 271, 270, 270, 269, 269, 268, 268, 267, 267, 
267, 266, 266, 265, 265, 264, 264, 264, 263, 263, 263, 262, 262, 262, 261, 261, 
261, 260, 260, 260, 259, 259, 259, 259, 259, 258, 258, 258, 258, 258, 257, 257, 
257, 257, 257, 257, 257, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 
256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 257, 257, 257, 257, 257, 257, 
257, 258, 258, 258, 258, 258, 259, 259, 259, 259, 259, 260, 260, 260, 261, 261, 
261, 262, 262, 262, 263, 263, 263, 264, 264, 264, 265, 265, 266, 266, 267, 267, 
267, 268, 268, 269, 269, 270, 270, 271, 271, 272, 273, 273, 274, 274, 275, 275, 
276, 277, 277, 278, 279, 279, 280, 281, 281, 282, 283, 283, 284, 285, 285, 286, 
287, 288, 288, 289, 290, 291, 292, 292, 293, 294, 295, 296, 296, 297, 298, 299, 
300, 301, 302, 303, 304, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 
315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 328, 329, 330, 331, 
332, 333, 334, 335, 336, 338, 339, 340, 341, 342, 343, 345, 346, 347, 348, 349, 
351, 352, 353, 354, 356, 357, 358, 359, 361, 362, 363, 364, 366, 367, 368, 370, 
371, 372, 373, 375, 376, 377, 379, 380, 381, 383, 384, 386, 387, 388, 390, 391, 
392, 394, 395, 397, 398, 399, 401, 402, 404, 405, 407, 408, 409, 411, 412, 414, 
415, 417, 418, 420, 421, 422, 424, 425, 427, 428, 430, 431, 433, 434, 436, 437, 
439, 440, 442, 443, 445, 446, 448, 449, 451, 452, 454, 456, 457, 459, 460, 462, 
463, 465, 466, 468, 469, 471, 472, 474, 476, 477, 479, 480, 482, 483, 485, 486, 
488, 490, 491, 493, 494, 496, 497, 499, 501, 502, 504, 505, 507, 508, 510, 512, 
512, 515, 516, 518, 519, 521, 522, 524, 526, 527, 529, 530, 532, 533, 535, 537, 
538, 540, 541, 543, 544, 546, 547, 549, 551, 552, 554, 555, 557, 558, 560, 561, 
563, 564, 566, 567, 569, 571, 572, 574, 575, 577, 578, 580, 581, 583, 584, 586, 
587, 589, 590, 592, 593, 595, 596, 598, 599, 601, 602, 603, 605, 606, 608, 609, 
611, 612, 614, 615, 616, 618, 619, 621, 622, 624, 625, 626, 628, 629, 631, 632, 
633, 635, 636, 637, 639, 640, 642, 643, 644, 646, 647, 648, 650, 651, 652, 653, 
655, 656, 657, 659, 660, 661, 662, 664, 665, 666, 667, 669, 670, 671, 672, 674, 
675, 676, 677, 678, 680, 681, 682, 683, 684, 685, 687, 688, 689, 690, 691, 692, 
693, 694, 695, 697, 698, 699, 700, 701, 702, 703, 704, 705, 706, 707, 708, 709, 
710, 711, 712, 713, 714, 715, 716, 717, 718, 719, 719, 720, 721, 722, 723, 724, 
725, 726, 727, 727, 728, 729, 730, 731, 731, 732, 733, 734, 735, 735, 736, 737, 
738, 738, 739, 740, 740, 741, 742, 742, 743, 744, 744, 745, 746, 746, 747, 748, 
748, 749, 749, 750, 750, 751, 752, 752, 753, 753, 754, 754, 755, 755, 756, 756, 
756, 757, 757, 758, 758, 759, 759, 759, 760, 760, 760, 761, 761, 761, 762, 762, 
762, 763, 763, 763, 764, 764, 764, 764, 764, 765, 765, 765, 765, 765, 766, 766, 
766, 766, 766, 766, 766, 767, 767, 767, 767, 767, 767, 767, 767, 767, 767, 767, 
767, 767, 767, 767, 767, 767, 767, 767, 767, 767, 766, 766, 766, 766, 766, 766, 
766, 765, 765, 765, 765, 765, 764, 764, 764, 764, 764, 763, 763, 763, 762, 762, 
762, 761, 761, 761, 760, 760, 760, 759, 759, 759, 758, 758, 757, 757, 756, 756, 
756, 755, 755, 754, 754, 753, 753, 752, 752, 751, 750, 750, 749, 749, 748, 748, 
747, 746, 746, 745, 744, 744, 743, 742, 742, 741, 740, 740, 739, 738, 738, 737, 
736, 735, 735, 734, 733, 732, 731, 731, 730, 729, 728, 727, 727, 726, 725, 724, 
723, 722, 721, 720, 719, 719, 718, 717, 716, 715, 714, 713, 712, 711, 710, 709, 
708, 707, 706, 705, 704, 703, 702, 701, 700, 699, 698, 697, 695, 694, 693, 692, 
691, 690, 689, 688, 687, 685, 684, 683, 682, 681, 680, 678, 677, 676, 675, 674, 
672, 671, 670, 669, 667, 666, 665, 664, 662, 661, 660, 659, 657, 656, 655, 653, 
652, 651, 650, 648, 647, 646, 644, 643, 642, 640, 639, 637, 636, 635, 633, 632, 
631, 629, 628, 626, 625, 624, 622, 621, 619, 618, 616, 615, 614, 612, 611, 609, 
608, 606, 605, 603, 602, 601, 599, 598, 596, 595, 593, 592, 590, 589, 587, 586, 
584, 583, 581, 580, 578, 577, 575, 574, 572, 571, 569, 567, 566, 564, 563, 561, 
560, 558, 557, 555, 554, 552, 551, 549, 547, 546, 544, 543, 541, 540, 538, 537, 
535, 533, 532, 530, 529, 527, 526, 524, 522, 521, 519, 518, 516, 515, 513, 512, 
510, 508, 507, 505, 504, 502, 501, 499, 497, 496, 494, 493, 491, 490, 488, 486, 
485, 483, 482, 480, 479, 477, 476, 474, 472, 471, 469, 468, 466, 465, 463, 462, 
460, 459, 457, 456, 454, 452, 451, 449, 448, 446, 445, 443, 442, 440, 439, 437, 
436, 434, 433, 431, 430, 428, 427, 425, 424, 422, 421, 420, 418, 417, 415, 414, 
412, 411, 409, 408, 407, 405, 404, 402, 401, 399, 398, 397, 395, 394, 392, 391, 
390, 388, 387, 386, 384, 383, 381, 380, 379, 377, 376, 375, 373, 372, 371, 370, 
368, 367, 366, 364, 363, 362, 361, 359, 358, 357, 356, 354, 353, 352, 351, 349, 
348, 347, 346, 345, 343, 342, 341, 340, 339, 338, 336, 335, 334, 333, 332, 331, 
330, 329, 328, 326, 325, 324, 323, 322, 321, 320, 319, 318, 317, 316, 315, 314, 
313, 312, 311, 310, 309, 308, 307, 306, 305, 304, 304, 303, 302, 301, 300, 299, 
298, 297, 296, 296, 295, 294, 293, 292, 292, 291, 290, 289, 288, 288, 287, 286, 
285, 285, 284, 283, 283, 282, 281, 281, 280, 279, 279, 278, 277, 277, 276, 275, 
275, 274, 274, 273, 273, 272, 271, 271, 270, 270, 269, 269, 268, 268, 267, 267, 
267, 266, 266, 265, 265, 264, 264, 264, 263, 263, 263, 262, 262, 262, 261, 261, 
261, 260, 260, 260, 259, 259, 259, 259, 259, 258, 258, 258, 258, 258, 257, 257, 
257, 257, 257, 257, 257, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 
256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 257, 257, 257, 257, 257, 257, 
257, 258, 258, 258, 258, 258, 259, 259, 259, 259, 259, 260, 260, 260, 261, 261, 
261, 262, 262, 262, 263, 263, 263, 264, 264, 264, 265, 265, 266, 266, 267, 267, 
267, 268, 268, 269, 269, 270, 270, 271, 271, 272, 273, 273, 274, 274, 275, 275, 
276, 277, 277, 278, 279, 279, 280, 281, 281, 282, 283, 283, 284, 285, 285, 286, 
287, 288, 288, 289, 290, 291, 292, 292, 293, 294, 295, 296, 296, 297, 298, 299, 
300, 301, 302, 303, 304, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 
315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 328, 329, 330, 331, 
332, 333, 334, 335, 336, 338, 339, 340, 341, 342, 343, 345, 346, 347, 348, 349, 
351, 352, 353, 354, 356, 357, 358, 359, 361, 362, 363, 364, 366, 367, 368, 370, 
371, 372, 373, 375, 376, 377, 379, 380, 381, 383, 384, 386, 387, 388, 390, 391, 
392, 394, 395, 397, 398, 399, 401, 402, 404, 405, 407, 408, 409, 411, 412, 414, 
415, 417, 418, 420, 421, 422, 424, 425, 427, 428, 430, 431, 433, 434, 436, 437, 
439, 440, 442, 443, 445, 446, 448, 449, 451, 452, 454, 456, 457, 459, 460, 462, 
463, 465, 466, 468, 469, 471, 472, 474, 476, 477, 479, 480, 482, 483, 485, 486, 
488, 490, 491, 493, 494, 496, 497, 499, 501, 502, 504, 505, 507, 508, 510, 512); 
signal buf1,buf2,buf3,buf4,buf5,buf6,buf7,buf8,buf9,buf10,buf11,buf12,buf13,buf14,buf15,buf16 : std_logic_vector(9 downto 0);
signal ctr : integer range 0 to 2047;
BEGIN
process(clk)
begin		
 if rising_edge(clk) then
  if (ctr<1023) then
	buf1 <= std_logic_vector(to_unsigned((sine1(ctr)+sine1(ctr+256)-512),10));
	buf2 <= std_logic_vector(to_unsigned((sine1(ctr)+sine2(ctr+256)-512),10));
	buf3 <= std_logic_vector(to_unsigned((sine1(ctr)+sine1(ctr+512+256)-512),10));
	buf4 <= std_logic_vector(to_unsigned((sine1(ctr)+sine2(ctr+512+256)-512),10));
	buf5 <= std_logic_vector(to_unsigned((sine2(ctr)+sine1(ctr+256)-512),10));
	buf6 <= std_logic_vector(to_unsigned((sine2(ctr)+sine2(ctr+256)-512),10));
	buf7 <= std_logic_vector(to_unsigned((sine2(ctr)+sine1(ctr+512+256)-512),10));
	buf8 <= std_logic_vector(to_unsigned((sine2(ctr)+sine2(ctr+512+256)-512),10));
	buf9 <= std_logic_vector(to_unsigned((sine1(ctr+512)+sine1(ctr+256)-512),10));
	buf10 <= std_logic_vector(to_unsigned((sine1(ctr+512)+sine2(ctr+256)-512),10));
	buf11 <= std_logic_vector(to_unsigned((sine1(ctr+512)+sine1(ctr+512+256)-512),10));
	buf12 <= std_logic_vector(to_unsigned((sine1(ctr+512)+sine2(ctr+512+256)-512),10));
	buf13 <= std_logic_vector(to_unsigned((sine2(ctr+512)+sine1(ctr+256)-512),10));
	buf14 <= std_logic_vector(to_unsigned((sine2(ctr+512)+sine2(ctr+256)-512),10));
	buf15 <= std_logic_vector(to_unsigned((sine2(ctr+512)+sine1(ctr+512+256)-512),10));
	buf16 <= std_logic_vector(to_unsigned((sine2(ctr+512)+sine2(ctr+512+256)-512),10));
	ctr<=ctr+1;
  else
	buf1 <= std_logic_vector(to_unsigned((sine1(ctr)+sine1(ctr+256)-512),10));
	buf2 <= std_logic_vector(to_unsigned((sine1(ctr)+sine2(ctr+256)-512),10));
	buf3 <= std_logic_vector(to_unsigned((sine1(ctr)+sine1(ctr+512+256)-512),10));
	buf4 <= std_logic_vector(to_unsigned((sine1(ctr)+sine2(ctr+512+256)-512),10));
	buf5 <= std_logic_vector(to_unsigned((sine2(ctr)+sine1(ctr+256)-512),10));
	buf6 <= std_logic_vector(to_unsigned((sine2(ctr)+sine2(ctr+256)-512),10));
	buf7 <= std_logic_vector(to_unsigned((sine2(ctr)+sine1(ctr+512+256)-512),10));
	buf8 <= std_logic_vector(to_unsigned((sine2(ctr)+sine2(ctr+512+256)-512),10));
	buf9 <= std_logic_vector(to_unsigned((sine1(ctr+512)+sine1(ctr+256)-512),10));
	buf10 <= std_logic_vector(to_unsigned((sine1(ctr+512)+sine2(ctr+256)-512),10));
	buf11 <= std_logic_vector(to_unsigned((sine1(ctr+512)+sine1(ctr+512+256)-512),10));
	buf12 <= std_logic_vector(to_unsigned((sine1(ctr+512)+sine2(ctr+512+256)-512),10));
	buf13 <= std_logic_vector(to_unsigned((sine2(ctr+512)+sine1(ctr+256)-512),10));
	buf14 <= std_logic_vector(to_unsigned((sine2(ctr+512)+sine2(ctr+256)-512),10));
	buf15 <= std_logic_vector(to_unsigned((sine2(ctr+512)+sine1(ctr+512+256)-512),10));
	buf16 <= std_logic_vector(to_unsigned((sine2(ctr+512)+sine2(ctr+512+256)-512),10));
	ctr<=0;
  end if;
 end if;
 if inp=buf1 then output<="0000";
  elsif inp=buf2 then output<="0001";
  elsif inp=buf3 then output<="0010";
  elsif inp=buf4 then output<="0011";
  elsif inp=buf5 then output<="0100";
  elsif inp=buf6 then output<="0101";
  elsif inp=buf7 then output<="0110";
  elsif inp=buf8 then output<="0111";
  elsif inp=buf9 then output<="1000";
  elsif inp=buf10 then output<="1001";
  elsif inp=buf11 then output<="1010";
  elsif inp=buf12 then output<="1011";
  elsif inp=buf13 then output<="1100";
  elsif inp=buf14 then output<="1101";
  elsif inp=buf15 then output<="1110";
  elsif inp=buf16 then output<="1111";
  else output<="ZZZZ";
 end if;
end process;
END;