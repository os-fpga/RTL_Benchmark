library ieee;
use ieee.std_logic_1164.all;

entity top is
	port( a: in std_logic_vector(23 downto 0);
	sin: out std_logic_vector(24 downto 0));
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415: std_logic;

begin

w0 <= a(21) and a(22);
w1 <= not a(1) and not a(2);
w2 <= not a(0) and w1;
w3 <= not a(3) and w2;
w4 <= not a(4) and w3;
w5 <= not a(5) and w4;
w6 <= not a(6) and w5;
w7 <= not a(7) and w6;
w8 <= not a(8) and w7;
w9 <= not a(9) and w8;
w10 <= not a(10) and w9;
w11 <= not a(11) and w10;
w12 <= not a(12) and w11;
w13 <= not a(13) and w12;
w14 <= not a(14) and w13;
w15 <= not a(15) and w14;
w16 <= not a(16) and w15;
w17 <= not a(17) and w16;
w18 <= not a(18) and w17;
w19 <= not a(19) and w18;
w20 <= not a(20) and w19;
w21 <= not a(21) and w20;
w22 <= a(21) and not w20;
w23 <= not w21 and not w22;
w24 <= not a(22) and w23;
w25 <= not w0 and not w24;
w26 <= a(20) and a(22);
w27 <= a(20) and not w19;
w28 <= not w20 and not w27;
w29 <= not a(22) and w28;
w30 <= not w26 and not w29;
w31 <= w25 and w30;
w32 <= a(15) and a(22);
w33 <= not a(22) and not w15;
w34 <= a(15) and not w14;
w35 <= w33 and not w34;
w36 <= not w32 and not w35;
w37 <= w31 and w36;
w38 <= not a(22) and not w18;
w39 <= a(19) and not w38;
w40 <= not a(19) and w38;
w41 <= not w39 and not w40;
w42 <= a(18) and a(22);
w43 <= a(18) and not w17;
w44 <= w38 and not w43;
w45 <= not w42 and not w44;
w46 <= not w41 and not w45;
w47 <= not a(22) and not w16;
w48 <= a(17) and not w47;
w49 <= not a(17) and w47;
w50 <= not w48 and not w49;
w51 <= a(16) and not w33;
w52 <= not a(16) and w33;
w53 <= not w51 and not w52;
w54 <= not w50 and w53;
w55 <= w46 and w54;
w56 <= w37 and w55;
w57 <= w50 and w53;
w58 <= w46 and w57;
w59 <= w25 and not w30;
w60 <= w36 and w59;
w61 <= w58 and w60;
w62 <= not w41 and w45;
w63 <= w57 and w62;
w64 <= w60 and w63;
w65 <= not w36 and w59;
w66 <= w41 and not w45;
w67 <= w57 and w66;
w68 <= w65 and w67;
w69 <= not w25 and w30;
w70 <= not w36 and w69;
w71 <= w50 and not w53;
w72 <= w62 and w71;
w73 <= w70 and w72;
w74 <= not w25 and not w30;
w75 <= not w36 and w74;
w76 <= w54 and w62;
w77 <= w75 and w76;
w78 <= w36 and w74;
w79 <= w55 and w78;
w80 <= w31 and not w36;
w81 <= w54 and w66;
w82 <= w80 and w81;
w83 <= w55 and w70;
w84 <= w72 and w75;
w85 <= not w50 and not w53;
w86 <= w66 and w85;
w87 <= w75 and w86;
w88 <= w78 and w86;
w89 <= w72 and w78;
w90 <= w78 and w81;
w91 <= not w89 and not w90;
w92 <= w55 and w60;
w93 <= w46 and w71;
w94 <= w78 and w93;
w95 <= not w92 and not w94;
w96 <= w55 and w65;
w97 <= w66 and w71;
w98 <= w60 and w97;
w99 <= not w96 and not w98;
w100 <= w76 and w78;
w101 <= w62 and w85;
w102 <= w78 and w101;
w103 <= not w100 and not w102;
w104 <= w80 and w86;
w105 <= w55 and w75;
w106 <= not w104 and not w105;
w107 <= w103 and w106;
w108 <= w99 and w107;
w109 <= w95 and w108;
w110 <= w91 and w109;
w111 <= not w88 and w110;
w112 <= not w87 and w111;
w113 <= not w84 and w112;
w114 <= not w83 and w113;
w115 <= not w82 and w114;
w116 <= w60 and w93;
w117 <= w70 and w101;
w118 <= w37 and w101;
w119 <= w65 and w72;
w120 <= w41 and w45;
w121 <= w57 and w120;
w122 <= w65 and w121;
w123 <= w36 and w69;
w124 <= w101 and w123;
w125 <= w58 and w75;
w126 <= w75 and w93;
w127 <= w67 and w123;
w128 <= w58 and w78;
w129 <= not w127 and not w128;
w130 <= not w126 and w129;
w131 <= not w125 and w130;
w132 <= not w124 and w131;
w133 <= not w122 and w132;
w134 <= not w119 and w133;
w135 <= not w118 and w134;
w136 <= w58 and w70;
w137 <= w85 and w120;
w138 <= w78 and w137;
w139 <= not w136 and not w138;
w140 <= w60 and w101;
w141 <= w67 and w70;
w142 <= w70 and w76;
w143 <= w71 and w120;
w144 <= w75 and w143;
w145 <= w46 and w85;
w146 <= w78 and w145;
w147 <= not w144 and not w146;
w148 <= not w142 and w147;
w149 <= not w141 and w148;
w150 <= not w140 and w149;
w151 <= w139 and w150;
w152 <= w135 and w151;
w153 <= not w117 and w152;
w154 <= not w116 and w153;
w155 <= w54 and w120;
w156 <= w65 and w155;
w157 <= w70 and w81;
w158 <= w78 and w97;
w159 <= not w157 and not w158;
w160 <= not w156 and w159;
w161 <= w80 and w97;
w162 <= w65 and w145;
w163 <= w121 and w123;
w164 <= w75 and w121;
w165 <= w67 and w80;
w166 <= w60 and w76;
w167 <= w70 and w97;
w168 <= w58 and w123;
w169 <= w75 and w137;
w170 <= w75 and w81;
w171 <= w75 and w97;
w172 <= w78 and w143;
w173 <= w72 and w80;
w174 <= w65 and w76;
w175 <= w70 and w93;
w176 <= w55 and w123;
w177 <= w75 and w101;
w178 <= w63 and w75;
w179 <= not w177 and not w178;
w180 <= not w176 and w179;
w181 <= not w175 and w180;
w182 <= not w174 and w181;
w183 <= not w173 and w182;
w184 <= w65 and w137;
w185 <= w55 and w80;
w186 <= not w184 and not w185;
w187 <= w80 and w137;
w188 <= w80 and w155;
w189 <= not w187 and not w188;
w190 <= w186 and w189;
w191 <= w183 and w190;
w192 <= not w172 and w191;
w193 <= not w171 and w192;
w194 <= not w170 and w193;
w195 <= not w169 and w194;
w196 <= not w168 and w195;
w197 <= not w167 and w196;
w198 <= not w166 and w197;
w199 <= not w165 and w198;
w200 <= not w164 and w199;
w201 <= not w163 and w200;
w202 <= not w162 and w201;
w203 <= not w161 and w202;
w204 <= w123 and w143;
w205 <= w70 and w145;
w206 <= not w204 and not w205;
w207 <= w63 and w123;
w208 <= w37 and w143;
w209 <= not w207 and not w208;
w210 <= w206 and w209;
w211 <= w203 and w210;
w212 <= w160 and w211;
w213 <= w154 and w212;
w214 <= w115 and w213;
w215 <= not w79 and w214;
w216 <= not w77 and w215;
w217 <= not w73 and w216;
w218 <= not w68 and w217;
w219 <= not w64 and w218;
w220 <= not w61 and w219;
w221 <= not w56 and w220;
w222 <= not a(22) and not w4;
w223 <= a(5) and not w222;
w224 <= not a(5) and w222;
w225 <= not w223 and not w224;
w226 <= a(4) and a(22);
w227 <= a(4) and not w3;
w228 <= w222 and not w227;
w229 <= not w226 and not w228;
w230 <= w225 and not w229;
w231 <= not w225 and w229;
w232 <= not w230 and not w231;
w233 <= not a(22) and not w2;
w234 <= a(3) and not w233;
w235 <= not a(3) and w233;
w236 <= not w234 and not w235;
w237 <= a(2) and a(22);
w238 <= not a(0) and not a(1);
w239 <= a(2) and not w238;
w240 <= w233 and not w239;
w241 <= not w237 and not w240;
w242 <= w236 and not w241;
w243 <= not w236 and w241;
w244 <= not w242 and not w243;
w245 <= w232 and not w244;
w246 <= w80 and w101;
w247 <= w58 and w65;
w248 <= w63 and w65;
w249 <= w72 and w123;
w250 <= w70 and w155;
w251 <= not w161 and not w250;
w252 <= w65 and w81;
w253 <= not w61 and not w252;
w254 <= w129 and w253;
w255 <= w251 and w254;
w256 <= not w87 and w255;
w257 <= not w249 and w256;
w258 <= not w141 and w257;
w259 <= not w248 and w258;
w260 <= not w247 and w259;
w261 <= not w246 and w260;
w262 <= w123 and w145;
w263 <= w70 and w86;
w264 <= not w171 and not w263;
w265 <= w60 and w137;
w266 <= not w64 and not w265;
w267 <= w75 and w155;
w268 <= not w79 and not w267;
w269 <= not w157 and w268;
w270 <= w266 and w269;
w271 <= w264 and w270;
w272 <= not w262 and w271;
w273 <= not w162 and w272;
w274 <= w37 and w121;
w275 <= not w73 and not w274;
w276 <= w37 and w97;
w277 <= w86 and w123;
w278 <= w78 and w155;
w279 <= w97 and w123;
w280 <= not w278 and not w279;
w281 <= not w205 and w280;
w282 <= not w277 and w281;
w283 <= not w118 and w282;
w284 <= not w276 and w283;
w285 <= w60 and w143;
w286 <= w63 and w70;
w287 <= w63 and w78;
w288 <= not w138 and not w287;
w289 <= not w125 and w288;
w290 <= not w286 and w289;
w291 <= not w285 and w290;
w292 <= w58 and w80;
w293 <= w123 and w137;
w294 <= not w292 and not w293;
w295 <= w80 and w121;
w296 <= not w100 and not w295;
w297 <= w60 and w145;
w298 <= w81 and w123;
w299 <= not w297 and not w298;
w300 <= w76 and w123;
w301 <= w37 and w63;
w302 <= not w142 and not w176;
w303 <= not w301 and w302;
w304 <= not w167 and w303;
w305 <= not w166 and w304;
w306 <= w60 and w121;
w307 <= w60 and w86;
w308 <= w60 and w155;
w309 <= w60 and w67;
w310 <= w70 and w137;
w311 <= w65 and w97;
w312 <= not w310 and not w311;
w313 <= not w309 and w312;
w314 <= not w308 and w313;
w315 <= not w307 and w314;
w316 <= not w306 and w315;
w317 <= w37 and w145;
w318 <= w37 and w76;
w319 <= not w77 and not w318;
w320 <= w123 and w155;
w321 <= w319 and not w320;
w322 <= not w317 and w321;
w323 <= not w56 and not w165;
w324 <= w322 and w323;
w325 <= w316 and w324;
w326 <= w305 and w325;
w327 <= not w124 and w326;
w328 <= not w83 and w327;
w329 <= not w96 and w328;
w330 <= not w173 and w329;
w331 <= w106 and w330;
w332 <= not w300 and w331;
w333 <= w299 and w332;
w334 <= w296 and w333;
w335 <= w209 and w334;
w336 <= w294 and w335;
w337 <= w291 and w336;
w338 <= w284 and w337;
w339 <= w275 and w338;
w340 <= w273 and w339;
w341 <= w261 and w340;
w342 <= not w158 and w341;
w343 <= not w84 and w342;
w344 <= w75 and w145;
w345 <= not w142 and not w300;
w346 <= not w124 and not w287;
w347 <= not w157 and not w277;
w348 <= w346 and w347;
w349 <= w264 and w348;
w350 <= w91 and w349;
w351 <= not w158 and w350;
w352 <= not w178 and w351;
w353 <= w345 and w352;
w354 <= not w117 and w353;
w355 <= w67 and w75;
w356 <= not w87 and not w207;
w357 <= not w286 and w356;
w358 <= w67 and w78;
w359 <= not w88 and not w358;
w360 <= not w170 and w359;
w361 <= not w249 and w360;
w362 <= w357 and w361;
w363 <= not w355 and w362;
w364 <= not w73 and w363;
w365 <= w78 and w121;
w366 <= not w205 and not w365;
w367 <= w93 and w123;
w368 <= w103 and w139;
w369 <= not w77 and w368;
w370 <= not w169 and w369;
w371 <= not w175 and w370;
w372 <= not w367 and w371;
w373 <= not w168 and w372;
w374 <= w366 and w373;
w375 <= w364 and w374;
w376 <= not w172 and w375;
w377 <= not w94 and w376;
w378 <= not w79 and w377;
w379 <= not w126 and w378;
w380 <= not w164 and w379;
w381 <= not w84 and w380;
w382 <= not w105 and not w144;
w383 <= not w128 and not w177;
w384 <= not w125 and w383;
w385 <= not w262 and w384;
w386 <= not w176 and w385;
w387 <= not w83 and w386;
w388 <= w382 and w387;
w389 <= w381 and w388;
w390 <= w354 and w389;
w391 <= not w278 and w390;
w392 <= not w146 and w391;
w393 <= not w267 and w392;
w394 <= not w344 and w393;
w395 <= w37 and w72;
w396 <= w70 and w121;
w397 <= w65 and w101;
w398 <= not w140 and not w397;
w399 <= w65 and w93;
w400 <= not w247 and not w399;
w401 <= not w116 and w400;
w402 <= w398 and w401;
w403 <= not w96 and w402;
w404 <= not w204 and not w293;
w405 <= not w174 and w404;
w406 <= not w162 and w405;
w407 <= not w92 and w406;
w408 <= w70 and w143;
w409 <= not w250 and not w408;
w410 <= not w310 and not w320;
w411 <= w299 and w410;
w412 <= w409 and w411;
w413 <= w407 and w412;
w414 <= w403 and w413;
w415 <= not w163 and w414;
w416 <= not w396 and w415;
w417 <= not w61 and w416;
w418 <= w63 and w80;
w419 <= w76 and w80;
w420 <= w37 and w58;
w421 <= w80 and w145;
w422 <= w37 and w93;
w423 <= not w127 and not w279;
w424 <= not w185 and not w306;
w425 <= not w141 and not w167;
w426 <= not w122 and w425;
w427 <= w80 and w93;
w428 <= not w292 and not w427;
w429 <= w426 and w428;
w430 <= w424 and w429;
w431 <= w423 and w430;
w432 <= not w56 and w431;
w433 <= not w317 and w432;
w434 <= not w422 and w433;
w435 <= not w421 and w434;
w436 <= not w420 and w435;
w437 <= not w118 and w436;
w438 <= not w246 and w437;
w439 <= not w419 and w438;
w440 <= not w418 and w439;
w441 <= w417 and w440;
w442 <= not w318 and w441;
w443 <= not w395 and w442;
w444 <= not w173 and w443;
w445 <= w65 and w143;
w446 <= not w68 and not w285;
w447 <= not w445 and w446;
w448 <= not w308 and w447;
w449 <= not w265 and w448;
w450 <= not w184 and w449;
w451 <= not w156 and w450;
w452 <= not w309 and w451;
w453 <= w60 and w72;
w454 <= w65 and w86;
w455 <= not w166 and not w454;
w456 <= w60 and w81;
w457 <= not w307 and not w311;
w458 <= not w456 and w457;
w459 <= w455 and w458;
w460 <= not w252 and w459;
w461 <= not w248 and w460;
w462 <= not w119 and w461;
w463 <= not w64 and w462;
w464 <= not w453 and w463;
w465 <= w417 and w464;
w466 <= w425 and w465;
w467 <= w423 and w466;
w468 <= w452 and w467;
w469 <= not w98 and w468;
w470 <= not w444 and not w469;
w471 <= a(14) and a(22);
w472 <= a(14) and not w13;
w473 <= not w14 and not w472;
w474 <= not a(22) and w473;
w475 <= not w471 and not w474;
w476 <= not a(22) and not w12;
w477 <= a(13) and not w476;
w478 <= not a(13) and w476;
w479 <= not w477 and not w478;
w480 <= not w475 and w479;
w481 <= w475 and not w479;
w482 <= not w480 and not w481;
w483 <= w470 and w482;
w484 <= not w470 and not w482;
w485 <= not w483 and not w484;
w486 <= not w394 and w485;
w487 <= w444 and not w469;
w488 <= not w444 and w469;
w489 <= not w487 and not w488;
w490 <= w444 and w469;
w491 <= w394 and not w490;
w492 <= w489 and not w491;
w493 <= not w475 and w492;
w494 <= not w394 and not w470;
w495 <= not w489 and not w494;
w496 <= w475 and not w494;
w497 <= not w495 and not w496;
w498 <= not w493 and w497;
w499 <= not w394 and not w479;
w500 <= w498 and not w499;
w501 <= not w498 and w499;
w502 <= w37 and w86;
w503 <= w37 and w155;
w504 <= w37 and w81;
w505 <= not w188 and not w504;
w506 <= not w158 and w505;
w507 <= not w171 and w506;
w508 <= not w317 and w507;
w509 <= not w175 and not w367;
w510 <= not w246 and w509;
w511 <= not w184 and not w421;
w512 <= not w187 and w511;
w513 <= not w177 and not w344;
w514 <= not w77 and w513;
w515 <= w512 and w514;
w516 <= w510 and w515;
w517 <= w508 and w516;
w518 <= w135 and w517;
w519 <= not w79 and w518;
w520 <= not w298 and w519;
w521 <= not w503 and w520;
w522 <= not w117 and not w170;
w523 <= not w141 and w522;
w524 <= not w287 and w523;
w525 <= not w310 and w524;
w526 <= not w162 and w525;
w527 <= not w420 and w526;
w528 <= not w68 and not w146;
w529 <= not w64 and w528;
w530 <= not w453 and w529;
w531 <= not w419 and w530;
w532 <= not w168 and not w293;
w533 <= not w279 and w532;
w534 <= not w399 and w533;
w535 <= not w248 and not w297;
w536 <= not w306 and w535;
w537 <= w115 and not w178;
w538 <= not w309 and w537;
w539 <= w37 and w137;
w540 <= not w136 and not w539;
w541 <= w538 and w540;
w542 <= w536 and w541;
w543 <= w534 and w542;
w544 <= w531 and w543;
w545 <= w527 and w544;
w546 <= w521 and w545;
w547 <= w305 and w546;
w548 <= not w502 and w547;
w549 <= w37 and w67;
w550 <= w91 and w323;
w551 <= not w170 and w550;
w552 <= not w84 and w551;
w553 <= not w122 and w552;
w554 <= not w248 and w553;
w555 <= not w456 and w554;
w556 <= not w504 and w555;
w557 <= not w172 and not w287;
w558 <= not w64 and w557;
w559 <= not w267 and not w355;
w560 <= w424 and w559;
w561 <= not w177 and w560;
w562 <= not w298 and w561;
w563 <= not w279 and w562;
w564 <= not w104 and w563;
w565 <= w103 and w382;
w566 <= w455 and w565;
w567 <= w564 and w566;
w568 <= not w358 and w567;
w569 <= not w138 and w568;
w570 <= not w79 and w569;
w571 <= not w167 and w570;
w572 <= not w307 and w571;
w573 <= not w276 and w572;
w574 <= not w344 and w573;
w575 <= not w301 and w574;
w576 <= not w158 and not w164;
w577 <= not w87 and w576;
w578 <= not w119 and w577;
w579 <= w575 and w578;
w580 <= w294 and w579;
w581 <= w558 and w580;
w582 <= w556 and w581;
w583 <= not w141 and w582;
w584 <= not w396 and w583;
w585 <= not w549 and w584;
w586 <= not w161 and w585;
w587 <= not w262 and not w365;
w588 <= not w126 and not w453;
w589 <= w587 and w588;
w590 <= not w146 and w589;
w591 <= not w125 and w590;
w592 <= not w250 and w591;
w593 <= not w252 and w592;
w594 <= not w163 and not w422;
w595 <= not w88 and not w178;
w596 <= not w427 and w595;
w597 <= not w77 and not w278;
w598 <= not w320 and w597;
w599 <= w206 and w598;
w600 <= not w94 and w599;
w601 <= not w171 and w600;
w602 <= not w421 and w601;
w603 <= not w82 and w602;
w604 <= not w169 and w603;
w605 <= not w408 and w604;
w606 <= w129 and w605;
w607 <= w596 and w606;
w608 <= w594 and w607;
w609 <= w593 and w608;
w610 <= w586 and w609;
w611 <= w312 and w610;
w612 <= not w502 and w611;
w613 <= not w317 and w612;
w614 <= not w548 and not w613;
w615 <= not w444 and not w614;
w616 <= not a(22) and not w10;
w617 <= a(11) and not w616;
w618 <= not a(11) and w616;
w619 <= not w617 and not w618;
w620 <= not w394 and not w619;
w621 <= not w615 and w620;
w622 <= w615 and not w620;
w623 <= not w621 and not w622;
w624 <= a(12) and a(22);
w625 <= a(12) and not w11;
w626 <= w476 and not w625;
w627 <= not w624 and not w626;
w628 <= not w394 and not w627;
w629 <= w623 and w628;
w630 <= not w621 and not w629;
w631 <= not w500 and not w630;
w632 <= not w501 and w631;
w633 <= not w500 and not w632;
w634 <= not w489 and not w491;
w635 <= not w475 and w634;
w636 <= w475 and w495;
w637 <= w489 and not w494;
w638 <= w479 and w637;
w639 <= not w479 and w492;
w640 <= not w638 and not w639;
w641 <= not w636 and w640;
w642 <= not w635 and w641;
w643 <= w548 and not w613;
w644 <= not w548 and w613;
w645 <= not w643 and not w644;
w646 <= w548 and w613;
w647 <= w444 and not w646;
w648 <= w645 and not w647;
w649 <= not w475 and w648;
w650 <= not w615 and not w645;
w651 <= w475 and not w615;
w652 <= not w650 and not w651;
w653 <= not w649 and w652;
w654 <= not w620 and w653;
w655 <= not w479 and w634;
w656 <= w479 and w495;
w657 <= w627 and w637;
w658 <= w492 and not w627;
w659 <= not w657 and not w658;
w660 <= not w656 and w659;
w661 <= not w655 and w660;
w662 <= w620 and not w653;
w663 <= not w654 and not w662;
w664 <= w661 and w663;
w665 <= not w654 and not w664;
w666 <= w642 and not w665;
w667 <= not w642 and w665;
w668 <= not w666 and not w667;
w669 <= not w623 and not w628;
w670 <= not w629 and not w669;
w671 <= w668 and w670;
w672 <= not w666 and not w671;
w673 <= not w630 and not w632;
w674 <= not w501 and w633;
w675 <= not w673 and not w674;
w676 <= not w672 and w675;
w677 <= w672 and not w675;
w678 <= not w676 and not w677;
w679 <= not w172 and not w365;
w680 <= not w169 and w679;
w681 <= not w309 and w680;
w682 <= not w116 and w681;
w683 <= not w420 and w682;
w684 <= not w318 and w683;
w685 <= not w295 and w684;
w686 <= w80 and w143;
w687 <= not w73 and not w117;
w688 <= not w166 and w687;
w689 <= not w686 and w688;
w690 <= not w287 and not w445;
w691 <= not w453 and w690;
w692 <= not w456 and w691;
w693 <= not w301 and w692;
w694 <= not w185 and w693;
w695 <= w426 and w694;
w696 <= w689 and w695;
w697 <= not w89 and w696;
w698 <= not w454 and w697;
w699 <= not w247 and w698;
w700 <= not w156 and w699;
w701 <= not w56 and w700;
w702 <= not w188 and w701;
w703 <= not w82 and not w248;
w704 <= not w298 and w595;
w705 <= not w300 and w704;
w706 <= not w168 and w705;
w707 <= not w98 and w706;
w708 <= not w127 and not w161;
w709 <= not w165 and w708;
w710 <= not w162 and not w422;
w711 <= w709 and w710;
w712 <= w707 and w711;
w713 <= w703 and w712;
w714 <= not w138 and w713;
w715 <= not w207 and w714;
w716 <= not w92 and w715;
w717 <= not w502 and w716;
w718 <= not w395 and w717;
w719 <= not w87 and not w263;
w720 <= not w397 and w719;
w721 <= not w265 and w720;
w722 <= not w118 and w721;
w723 <= not w421 and w722;
w724 <= not w164 and not w355;
w725 <= not w252 and w724;
w726 <= not w204 and not w250;
w727 <= not w175 and w726;
w728 <= w725 and w727;
w729 <= w723 and w728;
w730 <= w718 and w729;
w731 <= w702 and w730;
w732 <= w685 and w731;
w733 <= not w358 and w732;
w734 <= not w176 and w733;
w735 <= not w83 and w734;
w736 <= not w187 and w735;
w737 <= not w116 and not w176;
w738 <= not w187 and w737;
w739 <= not w427 and w738;
w740 <= not w119 and not w136;
w741 <= not w297 and w740;
w742 <= not w173 and w741;
w743 <= not w61 and not w126;
w744 <= not w420 and w743;
w745 <= not w84 and not w128;
w746 <= not w162 and w745;
w747 <= w744 and w746;
w748 <= w598 and w747;
w749 <= w742 and w748;
w750 <= not w169 and w749;
w751 <= not w300 and w750;
w752 <= not w367 and w751;
w753 <= not w83 and w752;
w754 <= not w265 and w753;
w755 <= not w56 and w754;
w756 <= not w175 and not w249;
w757 <= not w73 and not w125;
w758 <= not w94 and not w286;
w759 <= not w408 and not w539;
w760 <= w251 and w759;
w761 <= w99 and w760;
w762 <= not w208 and w761;
w763 <= not w318 and w762;
w764 <= not w247 and w763;
w765 <= not w156 and w764;
w766 <= w575 and w765;
w767 <= w758 and w766;
w768 <= w757 and w767;
w769 <= w756 and w768;
w770 <= w755 and w769;
w771 <= w739 and w770;
w772 <= not w122 and w771;
w773 <= w528 and w772;
w774 <= not w308 and w773;
w775 <= not w686 and w774;
w776 <= not w246 and w775;
w777 <= not w736 and not w776;
w778 <= not w548 and not w777;
w779 <= not a(22) and not w8;
w780 <= a(9) and not w779;
w781 <= not a(9) and w779;
w782 <= not w780 and not w781;
w783 <= not w394 and not w782;
w784 <= not w778 and w783;
w785 <= w778 and not w783;
w786 <= not w784 and not w785;
w787 <= a(10) and a(22);
w788 <= a(10) and not w9;
w789 <= w616 and not w788;
w790 <= not w787 and not w789;
w791 <= not w394 and not w790;
w792 <= w786 and w791;
w793 <= not w784 and not w792;
w794 <= not w645 and not w647;
w795 <= not w475 and w794;
w796 <= w475 and w650;
w797 <= not w615 and w645;
w798 <= w479 and w797;
w799 <= not w479 and w648;
w800 <= not w798 and not w799;
w801 <= not w796 and w800;
w802 <= not w795 and w801;
w803 <= not w627 and w634;
w804 <= w495 and w627;
w805 <= w619 and w637;
w806 <= w492 and not w619;
w807 <= not w805 and not w806;
w808 <= not w804 and w807;
w809 <= not w803 and w808;
w810 <= w802 and w809;
w811 <= w736 and not w776;
w812 <= not w736 and w776;
w813 <= not w811 and not w812;
w814 <= w736 and w776;
w815 <= w548 and not w814;
w816 <= w813 and not w815;
w817 <= not w475 and w816;
w818 <= not w778 and not w813;
w819 <= w475 and not w778;
w820 <= not w818 and not w819;
w821 <= not w817 and w820;
w822 <= not w783 and w821;
w823 <= not w479 and w794;
w824 <= w479 and w650;
w825 <= w627 and w797;
w826 <= not w627 and w648;
w827 <= not w825 and not w826;
w828 <= not w824 and w827;
w829 <= not w823 and w828;
w830 <= w783 and not w821;
w831 <= not w822 and not w830;
w832 <= w829 and w831;
w833 <= not w822 and not w832;
w834 <= not w802 and not w809;
w835 <= not w810 and not w834;
w836 <= not w833 and w835;
w837 <= not w810 and not w836;
w838 <= not w793 and not w837;
w839 <= not w793 and not w838;
w840 <= not w837 and not w838;
w841 <= not w839 and not w840;
w842 <= not w661 and not w663;
w843 <= not w664 and not w842;
w844 <= not w841 and w843;
w845 <= not w838 and not w844;
w846 <= not w668 and not w670;
w847 <= not w671 and not w846;
w848 <= not w845 and w847;
w849 <= not w619 and w634;
w850 <= w495 and w619;
w851 <= w637 and w790;
w852 <= w492 and not w790;
w853 <= not w851 and not w852;
w854 <= not w850 and w853;
w855 <= not w849 and w854;
w856 <= not w116 and not w396;
w857 <= w95 and w856;
w858 <= not w502 and w857;
w859 <= not w188 and w858;
w860 <= not w246 and w859;
w861 <= not w124 and not w420;
w862 <= not w172 and w861;
w863 <= not w300 and w862;
w864 <= not w295 and w863;
w865 <= w253 and w864;
w866 <= w273 and w865;
w867 <= w860 and w866;
w868 <= not w102 and w867;
w869 <= not w146 and w868;
w870 <= not w136 and w869;
w871 <= not w454 and w870;
w872 <= not w445 and w871;
w873 <= not w104 and w872;
w874 <= not w320 and not w418;
w875 <= not w297 and w874;
w876 <= not w395 and w875;
w877 <= not w77 and w357;
w878 <= not w166 and w877;
w879 <= not w539 and w878;
w880 <= not w317 and w879;
w881 <= not w89 and not w277;
w882 <= w512 and w588;
w883 <= w881 and w882;
w884 <= w880 and w883;
w885 <= w876 and w884;
w886 <= not w169 and w885;
w887 <= not w249 and w886;
w888 <= not w98 and w887;
w889 <= not w127 and not w164;
w890 <= not w168 and w889;
w891 <= not w142 and w890;
w892 <= not w83 and w891;
w893 <= not w686 and w892;
w894 <= not w292 and w893;
w895 <= not w140 and not w344;
w896 <= not w185 and w895;
w897 <= not w105 and not w355;
w898 <= not w301 and w897;
w899 <= w446 and w523;
w900 <= w898 and w899;
w901 <= w896 and w900;
w902 <= w275 and w901;
w903 <= w894 and w902;
w904 <= w888 and w903;
w905 <= w873 and w904;
w906 <= not w250 and w905;
w907 <= not w205 and w906;
w908 <= not w208 and w907;
w909 <= not w503 and w908;
w910 <= not w119 and not w310;
w911 <= not w397 and w910;
w912 <= not w105 and w911;
w913 <= not w300 and w912;
w914 <= not w168 and w913;
w915 <= not w184 and w914;
w916 <= not w309 and w915;
w917 <= not w307 and w916;
w918 <= not w83 and not w207;
w919 <= not w318 and w918;
w920 <= not w419 and not w421;
w921 <= w919 and w920;
w922 <= not w94 and w921;
w923 <= not w277 and w922;
w924 <= not w396 and w923;
w925 <= not w265 and w924;
w926 <= not w140 and not w252;
w927 <= not w124 and w926;
w928 <= not w141 and w927;
w929 <= not w118 and w928;
w930 <= not w172 and not w358;
w931 <= not w344 and w930;
w932 <= not w178 and w931;
w933 <= not w367 and w932;
w934 <= not w79 and not w128;
w935 <= not w146 and w934;
w936 <= not w399 and w935;
w937 <= w206 and w936;
w938 <= w933 and w937;
w939 <= w876 and w938;
w940 <= not w278 and w939;
w941 <= not w126 and w940;
w942 <= not w170 and w941;
w943 <= not w122 and w942;
w944 <= w737 and w943;
w945 <= not w173 and w944;
w946 <= not w287 and w945;
w947 <= not w125 and w946;
w948 <= not w502 and w947;
w949 <= not w301 and w948;
w950 <= w929 and w949;
w951 <= w91 and w950;
w952 <= w925 and w951;
w953 <= w917 and w952;
w954 <= w564 and w953;
w955 <= not w249 and w954;
w956 <= not w453 and w955;
w957 <= not w317 and w956;
w958 <= not w909 and not w957;
w959 <= not w736 and not w958;
w960 <= not a(22) and not w6;
w961 <= a(7) and not w960;
w962 <= not a(7) and w960;
w963 <= not w961 and not w962;
w964 <= not w394 and not w963;
w965 <= not w959 and w964;
w966 <= w959 and not w964;
w967 <= not w965 and not w966;
w968 <= a(8) and a(22);
w969 <= a(8) and not w7;
w970 <= w779 and not w969;
w971 <= not w968 and not w970;
w972 <= w967 and not w971;
w973 <= not w394 and w972;
w974 <= not w965 and not w973;
w975 <= w855 and not w974;
w976 <= w634 and not w790;
w977 <= w495 and w790;
w978 <= w637 and w782;
w979 <= w492 and not w782;
w980 <= not w978 and not w979;
w981 <= not w977 and w980;
w982 <= not w976 and w981;
w983 <= not w813 and not w815;
w984 <= not w475 and w983;
w985 <= w475 and w818;
w986 <= not w778 and w813;
w987 <= w479 and w986;
w988 <= not w479 and w816;
w989 <= not w987 and not w988;
w990 <= not w985 and w989;
w991 <= not w984 and w990;
w992 <= not w627 and w794;
w993 <= w627 and w650;
w994 <= w619 and w797;
w995 <= not w619 and w648;
w996 <= not w994 and not w995;
w997 <= not w993 and w996;
w998 <= not w992 and w997;
w999 <= w991 and not w998;
w1000 <= not w991 and w998;
w1001 <= not w999 and not w1000;
w1002 <= w982 and not w1001;
w1003 <= w991 and w998;
w1004 <= not w1002 and not w1003;
w1005 <= w855 and not w975;
w1006 <= not w974 and not w975;
w1007 <= not w1005 and not w1006;
w1008 <= not w1004 and not w1007;
w1009 <= not w975 and not w1008;
w1010 <= not w786 and not w791;
w1011 <= not w792 and not w1010;
w1012 <= not w1009 and w1011;
w1013 <= w1009 and not w1011;
w1014 <= not w1012 and not w1013;
w1015 <= w833 and not w835;
w1016 <= not w836 and not w1015;
w1017 <= w1014 and w1016;
w1018 <= not w1012 and not w1017;
w1019 <= not w841 and not w844;
w1020 <= w843 and not w844;
w1021 <= not w1019 and not w1020;
w1022 <= not w1018 and w1021;
w1023 <= w1018 and not w1021;
w1024 <= not w1022 and not w1023;
w1025 <= not w619 and w794;
w1026 <= w619 and w650;
w1027 <= w790 and w797;
w1028 <= w648 and not w790;
w1029 <= not w1027 and not w1028;
w1030 <= not w1026 and w1029;
w1031 <= not w1025 and w1030;
w1032 <= w634 and not w782;
w1033 <= w495 and w782;
w1034 <= w637 and w971;
w1035 <= w492 and not w971;
w1036 <= not w1034 and not w1035;
w1037 <= not w1033 and w1036;
w1038 <= not w1032 and w1037;
w1039 <= w1031 and w1038;
w1040 <= not w298 and not w445;
w1041 <= not w285 and w1040;
w1042 <= not w176 and not w396;
w1043 <= not w503 and w1042;
w1044 <= not w125 and not w293;
w1045 <= not w453 and w1044;
w1046 <= not w422 and w1045;
w1047 <= w1043 and w1046;
w1048 <= w1041 and w1047;
w1049 <= w933 and w1048;
w1050 <= w99 and w1049;
w1051 <= not w146 and w1050;
w1052 <= not w277 and w1051;
w1053 <= not w162 and w1052;
w1054 <= not w419 and w1053;
w1055 <= not w68 and w345;
w1056 <= not w185 and w1055;
w1057 <= w398 and w1056;
w1058 <= not w174 and w1057;
w1059 <= w410 and not w418;
w1060 <= not w126 and w1059;
w1061 <= not w164 and w1060;
w1062 <= not w168 and w1061;
w1063 <= not w454 and w1062;
w1064 <= not w308 and w1063;
w1065 <= not w295 and w1064;
w1066 <= not w173 and not w549;
w1067 <= not w90 and not w286;
w1068 <= w1066 and w1067;
w1069 <= w559 and w1068;
w1070 <= w508 and w1069;
w1071 <= w275 and w1070;
w1072 <= w1065 and w1071;
w1073 <= w1058 and w1072;
w1074 <= w261 and w1073;
w1075 <= w1054 and w1074;
w1076 <= not w138 and w1075;
w1077 <= not w83 and w1076;
w1078 <= not w156 and w1077;
w1079 <= not w116 and w1078;
w1080 <= not w502 and w1079;
w1081 <= w409 and w1066;
w1082 <= w757 and w1081;
w1083 <= not w170 and w1082;
w1084 <= not w344 and w1083;
w1085 <= w596 and w898;
w1086 <= w264 and w1085;
w1087 <= w1058 and w1086;
w1088 <= w1084 and w1087;
w1089 <= not w79 and w1088;
w1090 <= not w146 and w1089;
w1091 <= not w100 and w1090;
w1092 <= not w163 and w1091;
w1093 <= not w119 and w1092;
w1094 <= not w265 and w1093;
w1095 <= not w276 and w1094;
w1096 <= w587 and w861;
w1097 <= not w144 and w1096;
w1098 <= not w164 and w1097;
w1099 <= not w298 and w1098;
w1100 <= not w249 and w1099;
w1101 <= not w502 and w1100;
w1102 <= not w686 and w1101;
w1103 <= w510 and w919;
w1104 <= not w274 and w1103;
w1105 <= w1102 and w1104;
w1106 <= w425 and w1105;
w1107 <= not w117 and w1106;
w1108 <= not w286 and w1107;
w1109 <= not w208 and w1108;
w1110 <= not w295 and w1109;
w1111 <= not w104 and w1110;
w1112 <= not w165 and w1111;
w1113 <= not w158 and not w358;
w1114 <= not w92 and w1113;
w1115 <= not w61 and w1114;
w1116 <= w710 and w1115;
w1117 <= w401 and w1116;
w1118 <= w455 and w1117;
w1119 <= w316 and w1118;
w1120 <= w91 and w1119;
w1121 <= w1112 and w1120;
w1122 <= w1095 and w1121;
w1123 <= not w102 and w1122;
w1124 <= not w169 and w1123;
w1125 <= not w285 and w1124;
w1126 <= not w1080 and not w1125;
w1127 <= not w909 and not w1126;
w1128 <= w1080 and not w1127;
w1129 <= not w1080 and w1127;
w1130 <= a(6) and a(22);
w1131 <= a(6) and not w5;
w1132 <= w960 and not w1131;
w1133 <= not w1130 and not w1132;
w1134 <= not w394 and not w1133;
w1135 <= not w1128 and w1134;
w1136 <= not w1129 and w1135;
w1137 <= not w1128 and not w1136;
w1138 <= not w1031 and not w1038;
w1139 <= not w1039 and not w1138;
w1140 <= not w1137 and w1139;
w1141 <= not w1039 and not w1140;
w1142 <= w909 and not w957;
w1143 <= not w909 and w957;
w1144 <= not w1142 and not w1143;
w1145 <= w909 and w957;
w1146 <= w736 and not w1145;
w1147 <= w1144 and not w1146;
w1148 <= not w475 and w1147;
w1149 <= not w959 and not w1144;
w1150 <= w475 and not w959;
w1151 <= not w1149 and not w1150;
w1152 <= not w1148 and w1151;
w1153 <= not w964 and w1152;
w1154 <= not w479 and w983;
w1155 <= w479 and w818;
w1156 <= w627 and w986;
w1157 <= not w627 and w816;
w1158 <= not w1156 and not w1157;
w1159 <= not w1155 and w1158;
w1160 <= not w1154 and w1159;
w1161 <= w964 and not w1152;
w1162 <= not w1153 and not w1161;
w1163 <= w1160 and w1162;
w1164 <= not w1153 and not w1163;
w1165 <= not w1141 and not w1164;
w1166 <= not w1141 and not w1165;
w1167 <= not w1164 and not w1165;
w1168 <= not w1166 and not w1167;
w1169 <= not w394 and not w973;
w1170 <= not w971 and w1169;
w1171 <= w967 and not w973;
w1172 <= not w1170 and not w1171;
w1173 <= not w1168 and not w1172;
w1174 <= not w1165 and not w1173;
w1175 <= not w829 and not w831;
w1176 <= not w832 and not w1175;
w1177 <= not w1174 and w1176;
w1178 <= not w1004 and not w1008;
w1179 <= not w1007 and not w1008;
w1180 <= not w1178 and not w1179;
w1181 <= w1174 and not w1176;
w1182 <= not w1177 and not w1181;
w1183 <= not w1180 and w1182;
w1184 <= not w1177 and not w1183;
w1185 <= not w1014 and not w1016;
w1186 <= not w1017 and not w1185;
w1187 <= not w1184 and w1186;
w1188 <= w1182 and not w1183;
w1189 <= not w1180 and not w1183;
w1190 <= not w1188 and not w1189;
w1191 <= not w1144 and not w1146;
w1192 <= not w475 and w1191;
w1193 <= w475 and w1149;
w1194 <= not w959 and w1144;
w1195 <= w479 and w1194;
w1196 <= not w479 and w1147;
w1197 <= not w1195 and not w1196;
w1198 <= not w1193 and w1197;
w1199 <= not w1192 and w1198;
w1200 <= not w790 and w794;
w1201 <= w650 and w790;
w1202 <= w782 and w797;
w1203 <= w648 and not w782;
w1204 <= not w1202 and not w1203;
w1205 <= not w1201 and w1204;
w1206 <= not w1200 and w1205;
w1207 <= w634 and not w971;
w1208 <= w495 and w971;
w1209 <= w637 and w963;
w1210 <= w492 and not w963;
w1211 <= not w1209 and not w1210;
w1212 <= not w1208 and w1211;
w1213 <= not w1207 and w1212;
w1214 <= w1206 and not w1213;
w1215 <= not w1206 and w1213;
w1216 <= not w1214 and not w1215;
w1217 <= w1199 and not w1216;
w1218 <= w1206 and w1213;
w1219 <= not w1217 and not w1218;
w1220 <= not w1160 and not w1162;
w1221 <= not w1163 and not w1220;
w1222 <= not w1219 and w1221;
w1223 <= not w1219 and not w1222;
w1224 <= w1221 and not w1222;
w1225 <= not w1223 and not w1224;
w1226 <= w1137 and not w1139;
w1227 <= not w1140 and not w1226;
w1228 <= not w1225 and w1227;
w1229 <= not w1222 and not w1228;
w1230 <= w982 and not w1002;
w1231 <= not w1001 and not w1002;
w1232 <= not w1230 and not w1231;
w1233 <= not w1229 and not w1232;
w1234 <= not w1229 and not w1233;
w1235 <= not w1232 and not w1233;
w1236 <= not w1234 and not w1235;
w1237 <= not w1168 and not w1173;
w1238 <= not w1172 and not w1173;
w1239 <= not w1237 and not w1238;
w1240 <= not w1236 and not w1239;
w1241 <= not w1233 and not w1240;
w1242 <= not w1190 and not w1241;
w1243 <= not w1190 and not w1242;
w1244 <= not w1241 and not w1242;
w1245 <= not w1243 and not w1244;
w1246 <= not w627 and w983;
w1247 <= w627 and w818;
w1248 <= w619 and w986;
w1249 <= not w619 and w816;
w1250 <= not w1248 and not w1249;
w1251 <= not w1247 and w1250;
w1252 <= not w1246 and w1251;
w1253 <= not w1129 and w1137;
w1254 <= w1134 and not w1136;
w1255 <= not w1253 and not w1254;
w1256 <= w1252 and not w1255;
w1257 <= not w225 and not w394;
w1258 <= not w1080 and w1257;
w1259 <= w1080 and not w1257;
w1260 <= w1080 and not w1125;
w1261 <= not w1080 and w1125;
w1262 <= not w1260 and not w1261;
w1263 <= w1080 and w1125;
w1264 <= w909 and not w1263;
w1265 <= w1262 and not w1264;
w1266 <= not w475 and w1265;
w1267 <= not w1127 and not w1262;
w1268 <= w475 and not w1127;
w1269 <= not w1267 and not w1268;
w1270 <= not w1266 and w1269;
w1271 <= not w1258 and w1270;
w1272 <= not w1259 and w1271;
w1273 <= not w1258 and not w1272;
w1274 <= not w1252 and w1255;
w1275 <= not w1256 and not w1274;
w1276 <= not w1273 and w1275;
w1277 <= not w1256 and not w1276;
w1278 <= not w479 and w1191;
w1279 <= w479 and w1149;
w1280 <= w627 and w1194;
w1281 <= not w627 and w1147;
w1282 <= not w1280 and not w1281;
w1283 <= not w1279 and w1282;
w1284 <= not w1278 and w1283;
w1285 <= not w619 and w983;
w1286 <= w619 and w818;
w1287 <= w790 and w986;
w1288 <= not w790 and w816;
w1289 <= not w1287 and not w1288;
w1290 <= not w1286 and w1289;
w1291 <= not w1285 and w1290;
w1292 <= w1284 and w1291;
w1293 <= not w782 and w794;
w1294 <= w650 and w782;
w1295 <= w797 and w971;
w1296 <= w648 and not w971;
w1297 <= not w1295 and not w1296;
w1298 <= not w1294 and w1297;
w1299 <= not w1293 and w1298;
w1300 <= w1284 and not w1291;
w1301 <= not w1284 and w1291;
w1302 <= not w1300 and not w1301;
w1303 <= w1299 and not w1302;
w1304 <= not w1292 and not w1303;
w1305 <= not w1199 and w1216;
w1306 <= not w1217 and not w1305;
w1307 <= not w1304 and w1306;
w1308 <= w634 and not w963;
w1309 <= w495 and w963;
w1310 <= w637 and w1133;
w1311 <= w492 and not w1133;
w1312 <= not w1310 and not w1311;
w1313 <= not w1309 and w1312;
w1314 <= not w1308 and w1313;
w1315 <= not w229 and not w394;
w1316 <= not w1080 and w1315;
w1317 <= w1080 and not w1315;
w1318 <= not w1262 and not w1264;
w1319 <= not w475 and w1318;
w1320 <= w475 and w1267;
w1321 <= not w1127 and w1262;
w1322 <= w479 and w1321;
w1323 <= not w479 and w1265;
w1324 <= not w1322 and not w1323;
w1325 <= not w1320 and w1324;
w1326 <= not w1319 and w1325;
w1327 <= not w1316 and w1326;
w1328 <= not w1317 and w1327;
w1329 <= not w1316 and not w1328;
w1330 <= w1314 and not w1329;
w1331 <= not w1314 and w1329;
w1332 <= not w1330 and not w1331;
w1333 <= not w790 and w983;
w1334 <= w790 and w818;
w1335 <= w782 and w986;
w1336 <= not w782 and w816;
w1337 <= not w1335 and not w1336;
w1338 <= not w1334 and w1337;
w1339 <= not w1333 and w1338;
w1340 <= not w627 and w1191;
w1341 <= w627 and w1149;
w1342 <= w619 and w1194;
w1343 <= not w619 and w1147;
w1344 <= not w1342 and not w1343;
w1345 <= not w1341 and w1344;
w1346 <= not w1340 and w1345;
w1347 <= w1339 and w1346;
w1348 <= w794 and not w971;
w1349 <= w650 and w971;
w1350 <= w797 and w963;
w1351 <= w648 and not w963;
w1352 <= not w1350 and not w1351;
w1353 <= not w1349 and w1352;
w1354 <= not w1348 and w1353;
w1355 <= not w1339 and w1346;
w1356 <= w1339 and not w1346;
w1357 <= not w1355 and not w1356;
w1358 <= w1354 and not w1357;
w1359 <= not w1347 and not w1358;
w1360 <= w1332 and not w1359;
w1361 <= not w1330 and not w1360;
w1362 <= w1304 and not w1306;
w1363 <= not w1307 and not w1362;
w1364 <= not w1361 and w1363;
w1365 <= not w1307 and not w1364;
w1366 <= not w1277 and not w1365;
w1367 <= not w1277 and not w1366;
w1368 <= not w1365 and not w1366;
w1369 <= not w1367 and not w1368;
w1370 <= w1227 and not w1228;
w1371 <= not w1225 and not w1228;
w1372 <= not w1370 and not w1371;
w1373 <= not w1369 and not w1372;
w1374 <= not w1366 and not w1373;
w1375 <= not w1236 and w1239;
w1376 <= w1236 and not w1239;
w1377 <= not w1375 and not w1376;
w1378 <= not w1374 and not w1377;
w1379 <= not w1369 and not w1373;
w1380 <= not w1372 and not w1373;
w1381 <= not w1379 and not w1380;
w1382 <= not w1259 and w1273;
w1383 <= w1270 and not w1272;
w1384 <= not w1382 and not w1383;
w1385 <= w1299 and not w1303;
w1386 <= not w1302 and not w1303;
w1387 <= not w1385 and not w1386;
w1388 <= not w1384 and not w1387;
w1389 <= not w1384 and not w1388;
w1390 <= not w1387 and not w1388;
w1391 <= not w1389 and not w1390;
w1392 <= w634 and not w1133;
w1393 <= w495 and w1133;
w1394 <= w225 and w637;
w1395 <= not w225 and w492;
w1396 <= not w1394 and not w1395;
w1397 <= not w1393 and w1396;
w1398 <= not w1392 and w1397;
w1399 <= not w236 and not w394;
w1400 <= not w171 and w759;
w1401 <= not w124 and w1400;
w1402 <= not w250 and w1401;
w1403 <= not w73 and w1402;
w1404 <= not w162 and w1403;
w1405 <= not w297 and w1404;
w1406 <= not w502 and w1405;
w1407 <= not w503 and w1406;
w1408 <= not w170 and not w300;
w1409 <= not w265 and w1408;
w1410 <= w382 and w534;
w1411 <= w1409 and w1410;
w1412 <= w918 and w1411;
w1413 <= w594 and w1412;
w1414 <= not w287 and w1413;
w1415 <= not w164 and w1414;
w1416 <= not w367 and w1415;
w1417 <= not w184 and w1416;
w1418 <= not w317 and w1417;
w1419 <= not w274 and not w310;
w1420 <= not w396 and w1419;
w1421 <= not w122 and w1420;
w1422 <= not w453 and w1421;
w1423 <= not w306 and w1422;
w1424 <= not w166 and w1423;
w1425 <= not w292 and w1424;
w1426 <= not w104 and w1425;
w1427 <= w323 and w1426;
w1428 <= w1418 and w1427;
w1429 <= w371 and w1428;
w1430 <= w1407 and w1429;
w1431 <= not w128 and w1430;
w1432 <= not w158 and w1431;
w1433 <= not w68 and w1432;
w1434 <= not w311 and w1433;
w1435 <= not w208 and w1434;
w1436 <= not w549 and w1435;
w1437 <= not w161 and w1436;
w1438 <= not w475 and w1437;
w1439 <= not w1080 and not w1438;
w1440 <= w1399 and w1439;
w1441 <= not w479 and w1318;
w1442 <= w479 and w1267;
w1443 <= w627 and w1321;
w1444 <= not w627 and w1265;
w1445 <= not w1443 and not w1444;
w1446 <= not w1442 and w1445;
w1447 <= not w1441 and w1446;
w1448 <= not w1399 and not w1439;
w1449 <= not w1440 and not w1448;
w1450 <= w1447 and w1449;
w1451 <= not w1440 and not w1450;
w1452 <= w1398 and not w1451;
w1453 <= not w1398 and w1451;
w1454 <= not w1452 and not w1453;
w1455 <= not w782 and w983;
w1456 <= w782 and w818;
w1457 <= w971 and w986;
w1458 <= w816 and not w971;
w1459 <= not w1457 and not w1458;
w1460 <= not w1456 and w1459;
w1461 <= not w1455 and w1460;
w1462 <= not w619 and w1191;
w1463 <= w619 and w1149;
w1464 <= w790 and w1194;
w1465 <= not w790 and w1147;
w1466 <= not w1464 and not w1465;
w1467 <= not w1463 and w1466;
w1468 <= not w1462 and w1467;
w1469 <= w1461 and w1468;
w1470 <= w794 and not w963;
w1471 <= w650 and w963;
w1472 <= w797 and w1133;
w1473 <= w648 and not w1133;
w1474 <= not w1472 and not w1473;
w1475 <= not w1471 and w1474;
w1476 <= not w1470 and w1475;
w1477 <= not w1461 and w1468;
w1478 <= w1461 and not w1468;
w1479 <= not w1477 and not w1478;
w1480 <= w1476 and not w1479;
w1481 <= not w1469 and not w1480;
w1482 <= w1454 and not w1481;
w1483 <= not w1452 and not w1482;
w1484 <= not w1391 and not w1483;
w1485 <= not w1388 and not w1484;
w1486 <= w1273 and not w1275;
w1487 <= not w1276 and not w1486;
w1488 <= not w1485 and w1487;
w1489 <= w1485 and not w1487;
w1490 <= not w1488 and not w1489;
w1491 <= w1361 and not w1363;
w1492 <= not w1364 and not w1491;
w1493 <= w1490 and w1492;
w1494 <= not w1488 and not w1493;
w1495 <= not w1381 and not w1494;
w1496 <= w1381 and not w1494;
w1497 <= not w1381 and w1494;
w1498 <= not w1496 and not w1497;
w1499 <= w1080 and not w1437;
w1500 <= not w1437 and not w1499;
w1501 <= not w475 and w1500;
w1502 <= w475 and w1499;
w1503 <= w479 and not w1080;
w1504 <= w1437 and not w1503;
w1505 <= not w1502 and not w1504;
w1506 <= not w1501 and w1505;
w1507 <= not w236 and w634;
w1508 <= w236 and not w494;
w1509 <= not w637 and not w1508;
w1510 <= not w1507 and w1509;
w1511 <= w494 and w1510;
w1512 <= w1506 and w1511;
w1513 <= not w225 and w634;
w1514 <= w225 and w495;
w1515 <= w229 and w637;
w1516 <= not w229 and w492;
w1517 <= not w1515 and not w1516;
w1518 <= not w1514 and w1517;
w1519 <= not w1513 and w1518;
w1520 <= w1512 and w1519;
w1521 <= not w790 and w1191;
w1522 <= w790 and w1149;
w1523 <= w782 and w1194;
w1524 <= not w782 and w1147;
w1525 <= not w1523 and not w1524;
w1526 <= not w1522 and w1525;
w1527 <= not w1521 and w1526;
w1528 <= not w971 and w983;
w1529 <= w818 and w971;
w1530 <= w963 and w986;
w1531 <= w816 and not w963;
w1532 <= not w1530 and not w1531;
w1533 <= not w1529 and w1532;
w1534 <= not w1528 and w1533;
w1535 <= w794 and not w1133;
w1536 <= w650 and w1133;
w1537 <= w225 and w797;
w1538 <= not w225 and w648;
w1539 <= not w1537 and not w1538;
w1540 <= not w1536 and w1539;
w1541 <= not w1535 and w1540;
w1542 <= w1534 and not w1541;
w1543 <= not w1534 and w1541;
w1544 <= not w1542 and not w1543;
w1545 <= w1527 and not w1544;
w1546 <= w1534 and w1541;
w1547 <= not w1545 and not w1546;
w1548 <= not w1512 and not w1519;
w1549 <= not w1520 and not w1548;
w1550 <= not w1547 and w1549;
w1551 <= not w1520 and not w1550;
w1552 <= not w1317 and w1329;
w1553 <= w1326 and not w1328;
w1554 <= not w1552 and not w1553;
w1555 <= w1551 and not w1554;
w1556 <= not w1551 and w1554;
w1557 <= not w1555 and not w1556;
w1558 <= w1354 and not w1358;
w1559 <= not w1357 and not w1358;
w1560 <= not w1558 and not w1559;
w1561 <= not w1557 and not w1560;
w1562 <= not w1551 and not w1554;
w1563 <= not w1561 and not w1562;
w1564 <= not w1332 and w1359;
w1565 <= not w1360 and not w1564;
w1566 <= not w1563 and w1565;
w1567 <= w1391 and not w1483;
w1568 <= not w1391 and w1483;
w1569 <= not w1567 and not w1568;
w1570 <= w1563 and not w1565;
w1571 <= not w1566 and not w1570;
w1572 <= not w1569 and w1571;
w1573 <= not w1566 and not w1572;
w1574 <= not w1490 and not w1492;
w1575 <= not w1493 and not w1574;
w1576 <= not w1573 and w1575;
w1577 <= not w627 and w1318;
w1578 <= w627 and w1267;
w1579 <= w619 and w1321;
w1580 <= not w619 and w1265;
w1581 <= not w1579 and not w1580;
w1582 <= not w1578 and w1581;
w1583 <= not w1577 and w1582;
w1584 <= not w229 and w634;
w1585 <= w229 and w495;
w1586 <= w236 and w637;
w1587 <= not w236 and w492;
w1588 <= not w1586 and not w1587;
w1589 <= not w1585 and w1588;
w1590 <= not w1584 and w1589;
w1591 <= w1583 and w1590;
w1592 <= not w1506 and not w1511;
w1593 <= not w1512 and not w1592;
w1594 <= not w1583 and not w1590;
w1595 <= not w1591 and not w1594;
w1596 <= w1593 and w1595;
w1597 <= not w1591 and not w1596;
w1598 <= not w1447 and not w1449;
w1599 <= not w1450 and not w1598;
w1600 <= not w1597 and w1599;
w1601 <= w1597 and not w1599;
w1602 <= not w1600 and not w1601;
w1603 <= w1476 and not w1480;
w1604 <= not w1479 and not w1480;
w1605 <= not w1603 and not w1604;
w1606 <= w1602 and not w1605;
w1607 <= not w1600 and not w1606;
w1608 <= not w1454 and w1481;
w1609 <= not w1482 and not w1608;
w1610 <= not w1607 and w1609;
w1611 <= w1607 and not w1609;
w1612 <= not w1610 and not w1611;
w1613 <= w1557 and w1560;
w1614 <= not w1561 and not w1613;
w1615 <= w1612 and w1614;
w1616 <= not w1610 and not w1615;
w1617 <= w1569 and not w1571;
w1618 <= not w1572 and not w1617;
w1619 <= not w1616 and w1618;
w1620 <= not w627 and w1500;
w1621 <= w627 and w1499;
w1622 <= w619 and not w1080;
w1623 <= w1437 and not w1622;
w1624 <= not w1621 and not w1623;
w1625 <= not w1620 and w1624;
w1626 <= not w236 and w794;
w1627 <= w236 and not w615;
w1628 <= not w797 and not w1627;
w1629 <= not w1626 and w1628;
w1630 <= w615 and w1629;
w1631 <= w1625 and w1630;
w1632 <= not w782 and w1191;
w1633 <= w782 and w1149;
w1634 <= w971 and w1194;
w1635 <= not w971 and w1147;
w1636 <= not w1634 and not w1635;
w1637 <= not w1633 and w1636;
w1638 <= not w1632 and w1637;
w1639 <= not w963 and w983;
w1640 <= w818 and w963;
w1641 <= w986 and w1133;
w1642 <= w816 and not w1133;
w1643 <= not w1641 and not w1642;
w1644 <= not w1640 and w1643;
w1645 <= not w1639 and w1644;
w1646 <= w1638 and not w1645;
w1647 <= not w1638 and w1645;
w1648 <= not w1646 and not w1647;
w1649 <= w1631 and not w1648;
w1650 <= w1638 and w1645;
w1651 <= not w1649 and not w1650;
w1652 <= not w225 and w794;
w1653 <= w225 and w650;
w1654 <= w229 and w797;
w1655 <= not w229 and w648;
w1656 <= not w1654 and not w1655;
w1657 <= not w1653 and w1656;
w1658 <= not w1652 and w1657;
w1659 <= not w479 and w1500;
w1660 <= w479 and w1499;
w1661 <= w627 and not w1080;
w1662 <= w1437 and not w1661;
w1663 <= not w1660 and not w1662;
w1664 <= not w1659 and w1663;
w1665 <= not w619 and w1318;
w1666 <= w619 and w1267;
w1667 <= w790 and w1321;
w1668 <= not w790 and w1265;
w1669 <= not w1667 and not w1668;
w1670 <= not w1666 and w1669;
w1671 <= not w1665 and w1670;
w1672 <= w1664 and not w1671;
w1673 <= not w1664 and w1671;
w1674 <= not w1672 and not w1673;
w1675 <= w1658 and not w1674;
w1676 <= w1664 and w1671;
w1677 <= not w1675 and not w1676;
w1678 <= not w1651 and not w1677;
w1679 <= not w1651 and not w1678;
w1680 <= not w1677 and not w1678;
w1681 <= not w1679 and not w1680;
w1682 <= w1527 and not w1545;
w1683 <= not w1544 and not w1545;
w1684 <= not w1682 and not w1683;
w1685 <= not w1681 and not w1684;
w1686 <= not w1678 and not w1685;
w1687 <= w1547 and not w1549;
w1688 <= not w1550 and not w1687;
w1689 <= not w1686 and w1688;
w1690 <= w1602 and not w1606;
w1691 <= not w1605 and not w1606;
w1692 <= not w1690 and not w1691;
w1693 <= w1686 and not w1688;
w1694 <= not w1689 and not w1693;
w1695 <= not w1692 and w1694;
w1696 <= not w1689 and not w1695;
w1697 <= not w1612 and not w1614;
w1698 <= not w1615 and not w1697;
w1699 <= not w1696 and w1698;
w1700 <= not w494 and not w1510;
w1701 <= not w971 and w1191;
w1702 <= w971 and w1149;
w1703 <= w963 and w1194;
w1704 <= not w963 and w1147;
w1705 <= not w1703 and not w1704;
w1706 <= not w1702 and w1705;
w1707 <= not w1701 and w1706;
w1708 <= not w790 and w1318;
w1709 <= w790 and w1267;
w1710 <= w782 and w1321;
w1711 <= not w782 and w1265;
w1712 <= not w1710 and not w1711;
w1713 <= not w1709 and w1712;
w1714 <= not w1708 and w1713;
w1715 <= w983 and not w1133;
w1716 <= w818 and w1133;
w1717 <= w225 and w986;
w1718 <= not w225 and w816;
w1719 <= not w1717 and not w1718;
w1720 <= not w1716 and w1719;
w1721 <= not w1715 and w1720;
w1722 <= w1714 and not w1721;
w1723 <= not w1714 and w1721;
w1724 <= not w1722 and not w1723;
w1725 <= w1707 and not w1724;
w1726 <= w1714 and w1721;
w1727 <= not w1725 and not w1726;
w1728 <= not w1511 and not w1727;
w1729 <= not w1700 and w1728;
w1730 <= not w1511 and not w1729;
w1731 <= not w1700 and w1730;
w1732 <= not w1727 and not w1729;
w1733 <= not w1731 and not w1732;
w1734 <= not w1631 and w1648;
w1735 <= not w1649 and not w1734;
w1736 <= not w1733 and w1735;
w1737 <= not w1729 and not w1736;
w1738 <= w1593 and not w1596;
w1739 <= not w1594 and w1597;
w1740 <= not w1738 and not w1739;
w1741 <= not w1737 and w1740;
w1742 <= w1737 and not w1740;
w1743 <= not w1741 and not w1742;
w1744 <= not w1681 and not w1685;
w1745 <= not w1684 and not w1685;
w1746 <= not w1744 and not w1745;
w1747 <= not w1743 and not w1746;
w1748 <= not w1737 and not w1740;
w1749 <= not w1747 and not w1748;
w1750 <= w1692 and not w1694;
w1751 <= not w1695 and not w1750;
w1752 <= not w1749 and w1751;
w1753 <= not w619 and w1500;
w1754 <= w619 and w1499;
w1755 <= w790 and not w1080;
w1756 <= w1437 and not w1755;
w1757 <= not w1754 and not w1756;
w1758 <= not w1753 and w1757;
w1759 <= not w782 and w1318;
w1760 <= w782 and w1267;
w1761 <= w971 and w1321;
w1762 <= not w971 and w1265;
w1763 <= not w1761 and not w1762;
w1764 <= not w1760 and w1763;
w1765 <= not w1759 and w1764;
w1766 <= w1758 and w1765;
w1767 <= not w963 and w1191;
w1768 <= w963 and w1149;
w1769 <= w1133 and w1194;
w1770 <= not w1133 and w1147;
w1771 <= not w1769 and not w1770;
w1772 <= not w1768 and w1771;
w1773 <= not w1767 and w1772;
w1774 <= w1758 and not w1765;
w1775 <= not w1758 and w1765;
w1776 <= not w1774 and not w1775;
w1777 <= w1773 and not w1776;
w1778 <= not w1766 and not w1777;
w1779 <= not w229 and w794;
w1780 <= w229 and w650;
w1781 <= w236 and w797;
w1782 <= not w236 and w648;
w1783 <= not w1781 and not w1782;
w1784 <= not w1780 and w1783;
w1785 <= not w1779 and w1784;
w1786 <= not w1625 and not w1630;
w1787 <= not w1631 and not w1786;
w1788 <= w1785 and not w1787;
w1789 <= not w1785 and w1787;
w1790 <= not w1788 and not w1789;
w1791 <= not w1778 and not w1790;
w1792 <= w1785 and w1787;
w1793 <= not w1791 and not w1792;
w1794 <= w1658 and not w1675;
w1795 <= not w1674 and not w1675;
w1796 <= not w1794 and not w1795;
w1797 <= not w1793 and not w1796;
w1798 <= not w1733 and not w1736;
w1799 <= w1735 and not w1736;
w1800 <= not w1798 and not w1799;
w1801 <= not w1793 and not w1797;
w1802 <= not w1796 and not w1797;
w1803 <= not w1801 and not w1802;
w1804 <= not w1800 and not w1803;
w1805 <= not w1797 and not w1804;
w1806 <= not w225 and w983;
w1807 <= w225 and w818;
w1808 <= w229 and w986;
w1809 <= not w229 and w816;
w1810 <= not w1808 and not w1809;
w1811 <= not w1807 and w1810;
w1812 <= not w1806 and w1811;
w1813 <= not w790 and w1500;
w1814 <= w790 and w1499;
w1815 <= w782 and not w1080;
w1816 <= w1437 and not w1815;
w1817 <= not w1814 and not w1816;
w1818 <= not w1813 and w1817;
w1819 <= not w236 and w983;
w1820 <= w236 and not w778;
w1821 <= not w986 and not w1820;
w1822 <= not w1819 and w1821;
w1823 <= w778 and w1822;
w1824 <= w1818 and w1823;
w1825 <= w1812 and w1824;
w1826 <= not w1812 and w1824;
w1827 <= w1812 and not w1824;
w1828 <= not w1826 and not w1827;
w1829 <= not w236 and not w645;
w1830 <= not w1828 and w1829;
w1831 <= not w1825 and not w1830;
w1832 <= not w1707 and w1724;
w1833 <= not w1725 and not w1832;
w1834 <= not w1831 and w1833;
w1835 <= w1831 and not w1833;
w1836 <= not w1834 and not w1835;
w1837 <= w1778 and w1790;
w1838 <= not w1791 and not w1837;
w1839 <= not w1836 and not w1838;
w1840 <= w1836 and w1838;
w1841 <= not w229 and w983;
w1842 <= w229 and w818;
w1843 <= w236 and w986;
w1844 <= not w236 and w816;
w1845 <= not w1843 and not w1844;
w1846 <= not w1842 and w1845;
w1847 <= not w1841 and w1846;
w1848 <= not w971 and w1318;
w1849 <= w971 and w1267;
w1850 <= w963 and w1321;
w1851 <= not w963 and w1265;
w1852 <= not w1850 and not w1851;
w1853 <= not w1849 and w1852;
w1854 <= not w1848 and w1853;
w1855 <= not w1133 and w1191;
w1856 <= w1133 and w1149;
w1857 <= w225 and w1194;
w1858 <= not w225 and w1147;
w1859 <= not w1857 and not w1858;
w1860 <= not w1856 and w1859;
w1861 <= not w1855 and w1860;
w1862 <= w1854 and not w1861;
w1863 <= not w1854 and w1861;
w1864 <= not w1862 and not w1863;
w1865 <= w1847 and not w1864;
w1866 <= w1854 and w1861;
w1867 <= not w1865 and not w1866;
w1868 <= not w1773 and w1776;
w1869 <= not w1777 and not w1868;
w1870 <= not w1867 and w1869;
w1871 <= w1828 and not w1829;
w1872 <= not w1830 and not w1871;
w1873 <= not w1867 and not w1870;
w1874 <= w1869 and not w1870;
w1875 <= not w1873 and not w1874;
w1876 <= w1872 and not w1875;
w1877 <= not w1870 and not w1876;
w1878 <= not w778 and not w1822;
w1879 <= not w971 and w1500;
w1880 <= w971 and w1499;
w1881 <= w963 and not w1080;
w1882 <= w1437 and not w1881;
w1883 <= not w1880 and not w1882;
w1884 <= not w1879 and w1883;
w1885 <= not w236 and w1191;
w1886 <= w236 and not w959;
w1887 <= not w1194 and not w1886;
w1888 <= not w1885 and w1887;
w1889 <= w959 and w1888;
w1890 <= w1884 and w1889;
w1891 <= not w1823 and w1890;
w1892 <= not w1878 and w1891;
w1893 <= not w1133 and w1318;
w1894 <= w1133 and w1267;
w1895 <= w225 and w1321;
w1896 <= not w225 and w1265;
w1897 <= not w1895 and not w1896;
w1898 <= not w1894 and w1897;
w1899 <= not w1893 and w1898;
w1900 <= not w229 and w1191;
w1901 <= w229 and w1149;
w1902 <= w236 and w1194;
w1903 <= not w236 and w1147;
w1904 <= not w1902 and not w1903;
w1905 <= not w1901 and w1904;
w1906 <= not w1900 and w1905;
w1907 <= w1899 and w1906;
w1908 <= not w1884 and not w1889;
w1909 <= not w1890 and not w1908;
w1910 <= not w1899 and not w1906;
w1911 <= not w1907 and not w1910;
w1912 <= w1909 and w1911;
w1913 <= not w1907 and not w1912;
w1914 <= w1890 and not w1892;
w1915 <= not w1823 and not w1892;
w1916 <= not w1878 and w1915;
w1917 <= not w1914 and not w1916;
w1918 <= not w1913 and not w1917;
w1919 <= not w1892 and not w1918;
w1920 <= not w225 and w1191;
w1921 <= w225 and w1149;
w1922 <= w229 and w1194;
w1923 <= not w229 and w1147;
w1924 <= not w1922 and not w1923;
w1925 <= not w1921 and w1924;
w1926 <= not w1920 and w1925;
w1927 <= not w963 and w1318;
w1928 <= w963 and w1267;
w1929 <= w1133 and w1321;
w1930 <= not w1133 and w1265;
w1931 <= not w1929 and not w1930;
w1932 <= not w1928 and w1931;
w1933 <= not w1927 and w1932;
w1934 <= not w782 and w1500;
w1935 <= w782 and w1499;
w1936 <= w971 and not w1080;
w1937 <= w1437 and not w1936;
w1938 <= not w1935 and not w1937;
w1939 <= not w1934 and w1938;
w1940 <= not w1933 and w1939;
w1941 <= w1933 and not w1939;
w1942 <= not w1940 and not w1941;
w1943 <= not w1926 and w1942;
w1944 <= w1926 and not w1942;
w1945 <= not w963 and w1500;
w1946 <= w963 and w1499;
w1947 <= not w1080 and w1133;
w1948 <= w1437 and not w1947;
w1949 <= not w1946 and not w1948;
w1950 <= not w1945 and w1949;
w1951 <= not w225 and w1318;
w1952 <= w225 and w1267;
w1953 <= w229 and w1321;
w1954 <= not w229 and w1265;
w1955 <= not w1953 and not w1954;
w1956 <= not w1952 and w1955;
w1957 <= not w1951 and w1956;
w1958 <= w1950 and not w1957;
w1959 <= not w1950 and w1957;
w1960 <= not w1958 and not w1959;
w1961 <= not w1133 and w1500;
w1962 <= w1133 and w1499;
w1963 <= w225 and not w1080;
w1964 <= w1437 and not w1963;
w1965 <= not w1962 and not w1964;
w1966 <= not w1961 and w1965;
w1967 <= not w236 and w1318;
w1968 <= w236 and not w1127;
w1969 <= not w1321 and not w1968;
w1970 <= not w1967 and w1969;
w1971 <= w1127 and w1970;
w1972 <= w1966 and w1971;
w1973 <= w1960 and not w1972;
w1974 <= not w1960 and w1972;
w1975 <= not w229 and w1318;
w1976 <= w229 and w1267;
w1977 <= not w236 and w1265;
w1978 <= not w1127 and not w1970;
w1979 <= not w225 and w1500;
w1980 <= w225 and w1499;
w1981 <= not w229 and not w1437;
w1982 <= w1080 and w1437;
w1983 <= w229 and not w1982;
w1984 <= not w1981 and not w1983;
w1985 <= not w1980 and not w1984;
w1986 <= not w1979 and w1985;
w1987 <= w236 and not w1080;
w1988 <= not w1981 and w1987;
w1989 <= not w1986 and not w1988;
w1990 <= not w1971 and not w1989;
w1991 <= not w1978 and w1990;
w1992 <= w1986 and w1988;
w1993 <= not w1991 and not w1992;
w1994 <= not w1966 and not w1971;
w1995 <= not w1972 and not w1994;
w1996 <= w1993 and not w1995;
w1997 <= w236 and w1321;
w1998 <= not w1996 and not w1997;
w1999 <= not w1977 and w1998;
w2000 <= not w1976 and w1999;
w2001 <= not w1975 and w2000;
w2002 <= not w1993 and w1995;
w2003 <= not w2001 and not w2002;
w2004 <= not w236 and not w1144;
w2005 <= w2003 and not w2004;
w2006 <= not w1974 and not w2005;
w2007 <= not w1973 and w2006;
w2008 <= not w2003 and w2004;
w2009 <= not w2007 and not w2008;
w2010 <= w1909 and not w1912;
w2011 <= not w1910 and w1913;
w2012 <= not w2010 and not w2011;
w2013 <= w2009 and w2012;
w2014 <= w1950 and w1957;
w2015 <= not w1974 and not w2014;
w2016 <= not w2013 and not w2015;
w2017 <= not w2009 and not w2012;
w2018 <= not w2016 and not w2017;
w2019 <= not w1913 and not w1918;
w2020 <= not w1917 and not w1918;
w2021 <= not w2019 and not w2020;
w2022 <= w2018 and w2021;
w2023 <= not w1944 and not w2022;
w2024 <= not w1943 and w2023;
w2025 <= not w2018 and not w2021;
w2026 <= not w2024 and not w2025;
w2027 <= not w1919 and not w2026;
w2028 <= w1919 and w2026;
w2029 <= w1847 and not w1865;
w2030 <= not w1864 and not w1865;
w2031 <= not w2029 and not w2030;
w2032 <= not w1818 and not w1823;
w2033 <= not w1824 and not w2032;
w2034 <= w1933 and w1939;
w2035 <= not w1944 and not w2034;
w2036 <= w2033 and not w2035;
w2037 <= not w2033 and w2035;
w2038 <= not w2036 and not w2037;
w2039 <= not w2031 and w2038;
w2040 <= w2031 and not w2038;
w2041 <= not w2039 and not w2040;
w2042 <= not w2028 and w2041;
w2043 <= not w2027 and not w2042;
w2044 <= not w2036 and not w2039;
w2045 <= not w2043 and not w2044;
w2046 <= w2043 and w2044;
w2047 <= not w1872 and w1875;
w2048 <= not w1876 and not w2047;
w2049 <= not w2046 and w2048;
w2050 <= not w2045 and not w2049;
w2051 <= w1877 and w2050;
w2052 <= not w1840 and not w2051;
w2053 <= not w1839 and w2052;
w2054 <= not w1877 and not w2050;
w2055 <= not w2053 and not w2054;
w2056 <= not w1834 and not w1840;
w2057 <= not w2055 and not w2056;
w2058 <= w2055 and w2056;
w2059 <= w1800 and w1803;
w2060 <= not w1804 and not w2059;
w2061 <= not w2058 and w2060;
w2062 <= not w2057 and not w2061;
w2063 <= w1805 and w2062;
w2064 <= w1743 and w1746;
w2065 <= not w2063 and not w2064;
w2066 <= not w1747 and w2065;
w2067 <= not w1805 and not w2062;
w2068 <= not w2066 and not w2067;
w2069 <= w1749 and not w1751;
w2070 <= not w1752 and not w2069;
w2071 <= not w2068 and w2070;
w2072 <= not w1752 and not w2071;
w2073 <= w1696 and not w1698;
w2074 <= not w1699 and not w2073;
w2075 <= not w2072 and w2074;
w2076 <= not w1699 and not w2075;
w2077 <= w1616 and not w1618;
w2078 <= not w1619 and not w2077;
w2079 <= not w2076 and w2078;
w2080 <= not w1619 and not w2079;
w2081 <= w1573 and not w1575;
w2082 <= not w1576 and not w2081;
w2083 <= not w2080 and w2082;
w2084 <= not w1576 and not w2083;
w2085 <= not w1498 and not w2084;
w2086 <= not w1495 and not w2085;
w2087 <= w1374 and w1377;
w2088 <= not w1378 and not w2087;
w2089 <= not w2086 and w2088;
w2090 <= not w1378 and not w2089;
w2091 <= not w1245 and not w2090;
w2092 <= not w1242 and not w2091;
w2093 <= w1184 and not w1186;
w2094 <= not w1187 and not w2093;
w2095 <= not w2092 and w2094;
w2096 <= not w1187 and not w2095;
w2097 <= not w1024 and not w2096;
w2098 <= not w1018 and not w1021;
w2099 <= not w2097 and not w2098;
w2100 <= w845 and not w847;
w2101 <= not w848 and not w2100;
w2102 <= not w2099 and w2101;
w2103 <= not w848 and not w2102;
w2104 <= not w678 and not w2103;
w2105 <= not w672 and not w675;
w2106 <= not w2104 and not w2105;
w2107 <= w633 and not w2106;
w2108 <= not w633 and w2106;
w2109 <= not w2107 and not w2108;
w2110 <= w486 and w2109;
w2111 <= not w486 and not w2109;
w2112 <= not w2110 and not w2111;
w2113 <= not w343 and not w2112;
w2114 <= w343 and w2112;
w2115 <= not w84 and not w418;
w2116 <= not w169 and w2115;
w2117 <= not w204 and not w279;
w2118 <= not w308 and w2117;
w2119 <= not w276 and w2118;
w2120 <= not w292 and w2119;
w2121 <= w710 and w2120;
w2122 <= not w176 and w2121;
w2123 <= not w168 and w2122;
w2124 <= not w117 and w2123;
w2125 <= not w156 and w2124;
w2126 <= not w140 and w2125;
w2127 <= not w539 and w2126;
w2128 <= not w686 and w2127;
w2129 <= not w365 and w576;
w2130 <= not w247 and w2129;
w2131 <= not w306 and w2130;
w2132 <= not w311 and w918;
w2133 <= not w92 and w2132;
w2134 <= w505 and w2133;
w2135 <= w426 and w2134;
w2136 <= w1041 and w2135;
w2137 <= w2131 and w2136;
w2138 <= w936 and w2137;
w2139 <= w703 and w2138;
w2140 <= not w104 and w2139;
w2141 <= not w90 and w742;
w2142 <= not w249 and w2141;
w2143 <= not w408 and w2142;
w2144 <= not w307 and w2143;
w2145 <= not w98 and w2144;
w2146 <= not w503 and w2145;
w2147 <= w103 and w758;
w2148 <= w347 and w2147;
w2149 <= w723 and w2148;
w2150 <= w2146 and w2149;
w2151 <= w2140 and w2150;
w2152 <= w2128 and w2151;
w2153 <= w2116 and w2152;
w2154 <= not w278 and w2153;
w2155 <= not w178 and w2154;
w2156 <= not w127 and w2155;
w2157 <= not w454 and w2156;
w2158 <= not w317 and w2157;
w2159 <= not w165 and w2158;
w2160 <= w678 and w2103;
w2161 <= not w2104 and not w2160;
w2162 <= not w2159 and not w2161;
w2163 <= w95 and w744;
w2164 <= w269 and w2163;
w2165 <= w424 and w2164;
w2166 <= w587 and w2165;
w2167 <= w689 and w2166;
w2168 <= w917 and w2167;
w2169 <= w556 and w2168;
w2170 <= w1054 and w2169;
w2171 <= not w408 and w2170;
w2172 <= not w247 and w2171;
w2173 <= not w308 and w2172;
w2174 <= not w118 and w2173;
w2175 <= not w187 and w2174;
w2176 <= w2099 and not w2101;
w2177 <= not w2102 and not w2176;
w2178 <= not w2175 and not w2177;
w2179 <= w2175 and w2177;
w2180 <= w281 and w2133;
w2181 <= w186 and w2180;
w2182 <= w251 and w2181;
w2183 <= w587 and w2182;
w2184 <= w2116 and w2183;
w2185 <= w305 and w2184;
w2186 <= not w171 and w2185;
w2187 <= not w344 and w2186;
w2188 <= not w175 and w2187;
w2189 <= not w156 and w2188;
w2190 <= not w204 and w856;
w2191 <= not w397 and w2190;
w2192 <= not w98 and w2191;
w2193 <= not w61 and w2192;
w2194 <= not w188 and w2193;
w2195 <= w531 and w578;
w2196 <= w2194 and w2195;
w2197 <= not w177 and w2196;
w2198 <= not w367 and w2197;
w2199 <= not w73 and w2198;
w2200 <= not w686 and w2199;
w2201 <= not w128 and not w456;
w2202 <= not w421 and w2201;
w2203 <= not w252 and not w263;
w2204 <= not w395 and w2203;
w2205 <= w428 and w2204;
w2206 <= w2202 and w2205;
w2207 <= w106 and w2206;
w2208 <= w527 and w2207;
w2209 <= w594 and w2208;
w2210 <= w2200 and w2209;
w2211 <= w2189 and w2210;
w2212 <= not w267 and w2211;
w2213 <= not w286 and w2212;
w2214 <= not w504 and w2213;
w2215 <= w1024 and w2096;
w2216 <= not w2097 and not w2215;
w2217 <= not w2214 and not w2216;
w2218 <= w346 and w2202;
w2219 <= w401 and w2218;
w2220 <= not w89 and w2219;
w2221 <= not w138 and w2220;
w2222 <= not w79 and w2221;
w2223 <= not w309 and w2222;
w2224 <= not w285 and w2223;
w2225 <= not w317 and w2224;
w2226 <= not w549 and w2225;
w2227 <= not w397 and not w502;
w2228 <= not w187 and w2227;
w2229 <= not w102 and w2189;
w2230 <= not w246 and w2229;
w2231 <= not w165 and w2230;
w2232 <= w1409 and w2231;
w2233 <= w2228 and w2232;
w2234 <= w275 and w2233;
w2235 <= w2146 and w2234;
w2236 <= w2226 and w2235;
w2237 <= w930 and w2236;
w2238 <= not w126 and w2237;
w2239 <= not w293 and w2238;
w2240 <= not w117 and w2239;
w2241 <= not w310 and w2240;
w2242 <= not w263 and w2241;
w2243 <= w2092 and not w2094;
w2244 <= not w2095 and not w2243;
w2245 <= not w2242 and not w2244;
w2246 <= w2242 and w2244;
w2247 <= not w88 and not w177;
w2248 <= not w73 and w2247;
w2249 <= not w122 and w2248;
w2250 <= not w184 and w2249;
w2251 <= not w307 and w2250;
w2252 <= not w166 and w2251;
w2253 <= not w118 and w2252;
w2254 <= w91 and w1066;
w2255 <= w894 and w2254;
w2256 <= w594 and w2255;
w2257 <= w319 and w2256;
w2258 <= not w287 and w2257;
w2259 <= not w408 and w2258;
w2260 <= not w397 and w2259;
w2261 <= not w297 and w2260;
w2262 <= not w56 and w873;
w2263 <= not w276 and w2262;
w2264 <= not w167 and not w178;
w2265 <= not w96 and w2264;
w2266 <= not w161 and w2265;
w2267 <= not w419 and w2266;
w2268 <= w2263 and w2267;
w2269 <= w2261 and w2268;
w2270 <= w2253 and w2269;
w2271 <= not w278 and w2270;
w2272 <= not w358 and w2271;
w2273 <= not w144 and w2272;
w2274 <= not w169 and w2273;
w2275 <= not w248 and w2274;
w2276 <= w400 and w2275;
w2277 <= not w395 and w2276;
w2278 <= w1245 and w2090;
w2279 <= not w2091 and not w2278;
w2280 <= not w2277 and not w2279;
w2281 <= not w163 and w458;
w2282 <= not w686 and w2281;
w2283 <= not w295 and w2282;
w2284 <= w253 and w709;
w2285 <= w881 and w2284;
w2286 <= not w119 and w2285;
w2287 <= not w64 and w2286;
w2288 <= not w276 and w2287;
w2289 <= not w419 and w2288;
w2290 <= not w88 and not w96;
w2291 <= not w56 and not w298;
w2292 <= not w188 and w2291;
w2293 <= w382 and w2292;
w2294 <= w2290 and w2293;
w2295 <= w1056 and w2294;
w2296 <= w294 and w2295;
w2297 <= w264 and w2296;
w2298 <= w2289 and w2297;
w2299 <= w945 and w2298;
w2300 <= w880 and w2299;
w2301 <= w2283 and w2300;
w2302 <= not w102 and w2301;
w2303 <= not w167 and w2302;
w2304 <= not w445 and w2303;
w2305 <= w2086 and not w2088;
w2306 <= not w2089 and not w2305;
w2307 <= not w2304 and not w2306;
w2308 <= w2304 and w2306;
w2309 <= w91 and not w262;
w2310 <= not w367 and w2309;
w2311 <= not w263 and w2310;
w2312 <= not w174 and w2311;
w2313 <= not w503 and w2312;
w2314 <= not w185 and w2313;
w2315 <= not w205 and not w399;
w2316 <= not w504 and w2315;
w2317 <= not w144 and not w187;
w2318 <= w2316 and w2317;
w2319 <= w860 and w2318;
w2320 <= not w138 and w2319;
w2321 <= not w277 and w2320;
w2322 <= not w298 and w2321;
w2323 <= not w279 and w2322;
w2324 <= not w141 and w2323;
w2325 <= not w453 and w2324;
w2326 <= w332 and w398;
w2327 <= w2325 and w2326;
w2328 <= w703 and w2327;
w2329 <= w2314 and w2328;
w2330 <= not w146 and w2329;
w2331 <= not w171 and w2330;
w2332 <= not w344 and w2331;
w2333 <= not w117 and w2332;
w2334 <= not w297 and w2333;
w2335 <= not w422 and w2334;
w2336 <= w1498 and w2084;
w2337 <= not w2085 and not w2336;
w2338 <= not w2335 and not w2337;
w2339 <= w514 and w2204;
w2340 <= w856 and w2339;
w2341 <= w361 and w2340;
w2342 <= not w310 and w2341;
w2343 <= not w64 and w2342;
w2344 <= not w276 and w2343;
w2345 <= not w173 and w2344;
w2346 <= w366 and w423;
w2347 <= not w248 and w2346;
w2348 <= not w68 and w2347;
w2349 <= not w174 and w2348;
w2350 <= not w317 and w2349;
w2351 <= w540 and w2350;
w2352 <= w2345 and w2351;
w2353 <= w702 and w2352;
w2354 <= w936 and w2353;
w2355 <= w99 and w2354;
w2356 <= not w178 and w2355;
w2357 <= not w169 and w2356;
w2358 <= not w176 and w2357;
w2359 <= not w286 and w2358;
w2360 <= not w184 and w2359;
w2361 <= not w208 and w2360;
w2362 <= not w504 and w2361;
w2363 <= not w292 and w2362;
w2364 <= not w246 and w2363;
w2365 <= w2080 and not w2082;
w2366 <= not w2083 and not w2365;
w2367 <= not w2364 and not w2366;
w2368 <= not w503 and not w549;
w2369 <= not w285 and w2368;
w2370 <= not w61 and w2369;
w2371 <= not w427 and w2370;
w2372 <= not w246 and not w399;
w2373 <= w920 and w2372;
w2374 <= w2371 and w2373;
w2375 <= w2228 and w2374;
w2376 <= w323 and w2375;
w2377 <= w2283 and w2376;
w2378 <= w876 and w2377;
w2379 <= not w309 and w2378;
w2380 <= not w308 and w2379;
w2381 <= not w422 and w2380;
w2382 <= not w173 and w2381;
w2383 <= not w301 and not w454;
w2384 <= w346 and w756;
w2385 <= w2383 and w2384;
w2386 <= w2350 and w2385;
w2387 <= w275 and w2386;
w2388 <= w273 and w2387;
w2389 <= w933 and w2388;
w2390 <= w2382 and w2389;
w2391 <= w115 and w2390;
w2392 <= not w278 and w2391;
w2393 <= not w164 and w2392;
w2394 <= not w207 and w2393;
w2395 <= not w310 and w2394;
w2396 <= not w188 and w2395;
w2397 <= w2076 and not w2078;
w2398 <= not w2079 and not w2397;
w2399 <= not w2396 and not w2398;
w2400 <= w2396 and w2398;
w2401 <= not w102 and w1067;
w2402 <= not w177 and w2401;
w2403 <= not w297 and w2402;
w2404 <= not w504 and w2403;
w2405 <= not w126 and not w262;
w2406 <= not w320 and w2405;
w2407 <= not w311 and w2406;
w2408 <= not w82 and w2407;
w2409 <= w2404 and w2408;
w2410 <= not w293 and w2409;
w2411 <= not w408 and w2410;
w2412 <= not w309 and w2411;
w2413 <= not w502 and w2412;
w2414 <= not w104 and w2413;
w2415 <= w206 and w2372;
w2416 <= w424 and w2415;
w2417 <= w2289 and w2416;
w2418 <= w2414 and w2417;
w2419 <= w739 and w2418;
w2420 <= not w287 and w2419;
w2421 <= not w158 and w2420;
w2422 <= not w84 and w2421;
w2423 <= not w142 and w2422;
w2424 <= not w73 and w2423;
w2425 <= not w174 and w2424;
w2426 <= not w307 and w2425;
w2427 <= not w395 and w2426;
w2428 <= w2072 and not w2074;
w2429 <= not w2075 and not w2428;
w2430 <= not w2427 and not w2429;
w2431 <= w2427 and w2429;
w2432 <= not w2068 and not w2071;
w2433 <= w2070 and not w2071;
w2434 <= not w2432 and not w2433;
w2435 <= w727 and w1046;
w2436 <= w864 and w2435;
w2437 <= w323 and w2436;
w2438 <= w2345 and w2437;
w2439 <= w689 and w2438;
w2440 <= w2140 and w2439;
w2441 <= not w367 and w2440;
w2442 <= not w142 and w2441;
w2443 <= not w308 and w2442;
w2444 <= not w140 and w2443;
w2445 <= not w549 and w2444;
w2446 <= not w2434 and w2445;
w2447 <= not w2430 and not w2446;
w2448 <= not w2431 and w2447;
w2449 <= not w2430 and not w2448;
w2450 <= not w2399 and not w2449;
w2451 <= not w2400 and w2450;
w2452 <= not w2399 and not w2451;
w2453 <= w2364 and w2366;
w2454 <= not w2367 and not w2453;
w2455 <= not w2452 and w2454;
w2456 <= not w2367 and not w2455;
w2457 <= w2335 and w2337;
w2458 <= not w2338 and not w2457;
w2459 <= not w2456 and w2458;
w2460 <= not w2338 and not w2459;
w2461 <= not w2307 and not w2460;
w2462 <= not w2308 and w2461;
w2463 <= not w2307 and not w2462;
w2464 <= not w2277 and not w2280;
w2465 <= not w2279 and not w2280;
w2466 <= not w2464 and not w2465;
w2467 <= not w2463 and not w2466;
w2468 <= not w2280 and not w2467;
w2469 <= not w2245 and not w2468;
w2470 <= not w2246 and w2469;
w2471 <= not w2245 and not w2470;
w2472 <= w2214 and w2216;
w2473 <= not w2217 and not w2472;
w2474 <= not w2471 and w2473;
w2475 <= not w2217 and not w2474;
w2476 <= not w2178 and not w2475;
w2477 <= not w2179 and w2476;
w2478 <= not w2178 and not w2477;
w2479 <= w2159 and w2161;
w2480 <= not w2162 and not w2479;
w2481 <= not w2478 and w2480;
w2482 <= not w2162 and not w2481;
w2483 <= not w2113 and not w2482;
w2484 <= not w2114 and w2483;
w2485 <= not w2113 and not w2484;
w2486 <= not w358 and w746;
w2487 <= not w138 and w2486;
w2488 <= not w177 and w2487;
w2489 <= not w124 and w2488;
w2490 <= not w318 and w2489;
w2491 <= w428 and w1041;
w2492 <= w2289 and w2491;
w2493 <= w1418 and w2492;
w2494 <= w2490 and w2493;
w2495 <= w603 and w2494;
w2496 <= w99 and w2495;
w2497 <= not w249 and w2496;
w2498 <= w895 and w2497;
w2499 <= not w502 and w2498;
w2500 <= not w504 and w2499;
w2501 <= not w173 and w2500;
w2502 <= w2485 and w2501;
w2503 <= not w2485 and not w2501;
w2504 <= not w2502 and not w2503;
w2505 <= w245 and not w2504;
w2506 <= not w229 and w236;
w2507 <= w229 and not w236;
w2508 <= not w2506 and not w2507;
w2509 <= not w232 and w244;
w2510 <= w2508 and w2509;
w2511 <= w2478 and not w2480;
w2512 <= not w2481 and not w2511;
w2513 <= w2510 and w2512;
w2514 <= not w2482 and not w2484;
w2515 <= not w2114 and w2485;
w2516 <= not w2514 and not w2515;
w2517 <= w244 and not w2508;
w2518 <= not w2516 and w2517;
w2519 <= not w2513 and not w2518;
w2520 <= not w2505 and w2519;
w2521 <= not w232 and not w244;
w2522 <= w2512 and not w2516;
w2523 <= not w2475 and not w2477;
w2524 <= not w2179 and w2478;
w2525 <= not w2523 and not w2524;
w2526 <= w2512 and not w2525;
w2527 <= w2471 and not w2473;
w2528 <= not w2474 and not w2527;
w2529 <= not w2525 and w2528;
w2530 <= not w2468 and not w2470;
w2531 <= not w2246 and w2471;
w2532 <= not w2530 and not w2531;
w2533 <= w2528 and not w2532;
w2534 <= not w2463 and not w2467;
w2535 <= not w2466 and not w2467;
w2536 <= not w2534 and not w2535;
w2537 <= not w2532 and not w2536;
w2538 <= not w2460 and not w2462;
w2539 <= not w2308 and w2463;
w2540 <= not w2538 and not w2539;
w2541 <= not w2536 and not w2540;
w2542 <= w2456 and not w2458;
w2543 <= not w2459 and not w2542;
w2544 <= not w2540 and w2543;
w2545 <= w2452 and not w2454;
w2546 <= not w2455 and not w2545;
w2547 <= w2543 and w2546;
w2548 <= not w2449 and not w2451;
w2549 <= not w2400 and w2452;
w2550 <= not w2548 and not w2549;
w2551 <= w2546 and not w2550;
w2552 <= not w2446 and not w2448;
w2553 <= not w2431 and w2449;
w2554 <= not w2552 and not w2553;
w2555 <= not w2550 and not w2554;
w2556 <= w2434 and not w2445;
w2557 <= not w2446 and not w2556;
w2558 <= not w2554 and not w2557;
w2559 <= w2550 and w2558;
w2560 <= not w2555 and not w2559;
w2561 <= not w2546 and w2550;
w2562 <= not w2560 and not w2561;
w2563 <= not w2551 and w2562;
w2564 <= not w2551 and not w2563;
w2565 <= not w2543 and not w2546;
w2566 <= not w2564 and not w2565;
w2567 <= not w2547 and w2566;
w2568 <= not w2547 and not w2567;
w2569 <= w2540 and not w2543;
w2570 <= not w2544 and not w2569;
w2571 <= not w2568 and w2570;
w2572 <= not w2544 and not w2571;
w2573 <= w2536 and w2540;
w2574 <= not w2541 and not w2573;
w2575 <= not w2572 and w2574;
w2576 <= not w2541 and not w2575;
w2577 <= w2532 and w2536;
w2578 <= not w2537 and not w2577;
w2579 <= not w2576 and w2578;
w2580 <= not w2537 and not w2579;
w2581 <= not w2528 and w2532;
w2582 <= not w2533 and not w2581;
w2583 <= not w2580 and w2582;
w2584 <= not w2533 and not w2583;
w2585 <= w2525 and not w2528;
w2586 <= not w2529 and not w2585;
w2587 <= not w2584 and w2586;
w2588 <= not w2529 and not w2587;
w2589 <= not w2512 and w2525;
w2590 <= not w2526 and not w2589;
w2591 <= not w2588 and w2590;
w2592 <= not w2526 and not w2591;
w2593 <= not w2512 and w2516;
w2594 <= not w2522 and not w2593;
w2595 <= not w2592 and w2594;
w2596 <= not w2522 and not w2595;
w2597 <= not w2504 and not w2516;
w2598 <= w2504 and w2516;
w2599 <= not w2597 and not w2598;
w2600 <= not w2596 and w2599;
w2601 <= w2596 and not w2599;
w2602 <= not w2600 and not w2601;
w2603 <= w2521 and w2602;
w2604 <= w2520 and not w2603;
w2605 <= not w225 and not w2604;
w2606 <= w225 and w2604;
w2607 <= not w2605 and not w2606;
w2608 <= w619 and not w627;
w2609 <= not w619 and w627;
w2610 <= not w2608 and not w2609;
w2611 <= not w2557 and not w2610;
w2612 <= not w475 and not w2611;
w2613 <= w479 and not w627;
w2614 <= not w479 and w627;
w2615 <= not w2613 and not w2614;
w2616 <= w2610 and not w2615;
w2617 <= not w2557 and w2616;
w2618 <= w482 and not w2610;
w2619 <= not w2554 and w2618;
w2620 <= not w2617 and not w2619;
w2621 <= w2554 and not w2557;
w2622 <= not w2554 and w2557;
w2623 <= not w2621 and not w2622;
w2624 <= not w482 and not w2610;
w2625 <= not w2623 and w2624;
w2626 <= w2620 and not w2625;
w2627 <= not w475 and not w2626;
w2628 <= not w475 and not w2627;
w2629 <= not w2626 and not w2627;
w2630 <= not w2628 and not w2629;
w2631 <= w2612 and not w2630;
w2632 <= not w2612 and w2630;
w2633 <= not w2631 and not w2632;
w2634 <= w782 and not w971;
w2635 <= not w782 and w971;
w2636 <= not w2634 and not w2635;
w2637 <= w619 and not w790;
w2638 <= not w619 and w790;
w2639 <= not w2637 and not w2638;
w2640 <= not w2636 and not w2639;
w2641 <= w782 and not w790;
w2642 <= not w782 and w790;
w2643 <= not w2641 and not w2642;
w2644 <= w2636 and not w2639;
w2645 <= w2643 and w2644;
w2646 <= not w2550 and w2645;
w2647 <= w2636 and not w2643;
w2648 <= w2546 and w2647;
w2649 <= not w2636 and w2639;
w2650 <= w2543 and w2649;
w2651 <= not w2648 and not w2650;
w2652 <= not w2646 and w2651;
w2653 <= not w2640 and w2652;
w2654 <= not w2564 and not w2567;
w2655 <= not w2565 and w2568;
w2656 <= not w2654 and not w2655;
w2657 <= w2652 and w2656;
w2658 <= not w2653 and not w2657;
w2659 <= w619 and not w2658;
w2660 <= not w619 and w2658;
w2661 <= not w2659 and not w2660;
w2662 <= w2633 and w2661;
w2663 <= not w2557 and not w2636;
w2664 <= not w619 and not w2663;
w2665 <= not w2557 and w2647;
w2666 <= not w2554 and w2649;
w2667 <= not w2665 and not w2666;
w2668 <= not w2623 and w2640;
w2669 <= w2667 and not w2668;
w2670 <= not w619 and not w2669;
w2671 <= w619 and w2669;
w2672 <= not w2670 and not w2671;
w2673 <= w2664 and w2672;
w2674 <= not w2550 and w2649;
w2675 <= not w2557 and w2645;
w2676 <= not w2554 and w2647;
w2677 <= not w2675 and not w2676;
w2678 <= not w2674 and w2677;
w2679 <= not w2640 and w2678;
w2680 <= w2550 and not w2622;
w2681 <= not w2550 and w2622;
w2682 <= not w2680 and not w2681;
w2683 <= w2678 and not w2682;
w2684 <= not w2679 and not w2683;
w2685 <= w619 and not w2684;
w2686 <= not w619 and w2684;
w2687 <= not w2685 and not w2686;
w2688 <= w2673 and w2687;
w2689 <= w2611 and w2688;
w2690 <= w2688 and not w2689;
w2691 <= w2611 and not w2689;
w2692 <= not w2690 and not w2691;
w2693 <= not w2550 and w2647;
w2694 <= w2546 and w2649;
w2695 <= not w2554 and w2645;
w2696 <= not w2694 and not w2695;
w2697 <= not w2693 and w2696;
w2698 <= not w2560 and not w2563;
w2699 <= not w2561 and w2564;
w2700 <= not w2698 and not w2699;
w2701 <= w2640 and not w2700;
w2702 <= w2697 and not w2701;
w2703 <= not w619 and not w2702;
w2704 <= w619 and w2702;
w2705 <= not w2703 and not w2704;
w2706 <= not w2692 and w2705;
w2707 <= not w2689 and not w2706;
w2708 <= not w2633 and not w2661;
w2709 <= not w2662 and not w2708;
w2710 <= not w2707 and w2709;
w2711 <= not w2662 and not w2710;
w2712 <= not w2540 and w2649;
w2713 <= w2546 and w2645;
w2714 <= w2543 and w2647;
w2715 <= not w2713 and not w2714;
w2716 <= not w2712 and w2715;
w2717 <= w2568 and not w2570;
w2718 <= not w2571 and not w2717;
w2719 <= w2640 and w2718;
w2720 <= w2716 and not w2719;
w2721 <= not w619 and not w2720;
w2722 <= w619 and w2720;
w2723 <= not w2721 and not w2722;
w2724 <= not w2550 and w2618;
w2725 <= not w482 and w2610;
w2726 <= w2615 and w2725;
w2727 <= not w2557 and w2726;
w2728 <= not w2554 and w2616;
w2729 <= not w2727 and not w2728;
w2730 <= not w2724 and w2729;
w2731 <= not w2624 and w2730;
w2732 <= not w2682 and w2730;
w2733 <= not w2731 and not w2732;
w2734 <= w475 and not w2733;
w2735 <= not w475 and w2733;
w2736 <= not w2734 and not w2735;
w2737 <= w2631 and w2736;
w2738 <= not w2631 and not w2736;
w2739 <= not w2737 and not w2738;
w2740 <= w2723 and w2739;
w2741 <= not w2723 and not w2739;
w2742 <= not w2740 and not w2741;
w2743 <= w2711 and not w2742;
w2744 <= not w2711 and w2742;
w2745 <= not w2743 and not w2744;
w2746 <= w963 and not w971;
w2747 <= not w963 and w971;
w2748 <= not w2746 and not w2747;
w2749 <= w225 and not w1133;
w2750 <= not w225 and w1133;
w2751 <= not w2749 and not w2750;
w2752 <= w2748 and not w2751;
w2753 <= w2528 and w2752;
w2754 <= w963 and not w1133;
w2755 <= not w963 and w1133;
w2756 <= not w2754 and not w2755;
w2757 <= not w2748 and w2751;
w2758 <= w2756 and w2757;
w2759 <= not w2536 and w2758;
w2760 <= w2751 and not w2756;
w2761 <= not w2532 and w2760;
w2762 <= not w2759 and not w2761;
w2763 <= not w2753 and w2762;
w2764 <= w2580 and not w2582;
w2765 <= not w2583 and not w2764;
w2766 <= w2763 and not w2765;
w2767 <= not w2748 and not w2751;
w2768 <= w2763 and not w2767;
w2769 <= not w2766 and not w2768;
w2770 <= w971 and not w2769;
w2771 <= not w971 and w2769;
w2772 <= not w2770 and not w2771;
w2773 <= w2745 and w2772;
w2774 <= not w2532 and w2752;
w2775 <= not w2540 and w2758;
w2776 <= not w2536 and w2760;
w2777 <= not w2775 and not w2776;
w2778 <= not w2774 and w2777;
w2779 <= w2576 and not w2578;
w2780 <= not w2579 and not w2779;
w2781 <= w2767 and w2780;
w2782 <= w2778 and not w2781;
w2783 <= not w971 and not w2782;
w2784 <= not w2782 and not w2783;
w2785 <= not w971 and not w2783;
w2786 <= not w2784 and not w2785;
w2787 <= w2707 and not w2709;
w2788 <= not w2710 and not w2787;
w2789 <= not w2786 and w2788;
w2790 <= not w2692 and not w2706;
w2791 <= w2705 and not w2706;
w2792 <= not w2790 and not w2791;
w2793 <= not w2536 and w2752;
w2794 <= w2543 and w2758;
w2795 <= not w2540 and w2760;
w2796 <= not w2794 and not w2795;
w2797 <= not w2793 and w2796;
w2798 <= w2572 and not w2574;
w2799 <= not w2575 and not w2798;
w2800 <= w2797 and not w2799;
w2801 <= not w2767 and w2797;
w2802 <= not w2800 and not w2801;
w2803 <= w971 and not w2802;
w2804 <= not w971 and w2802;
w2805 <= not w2803 and not w2804;
w2806 <= not w2792 and w2805;
w2807 <= not w2540 and w2752;
w2808 <= w2546 and w2758;
w2809 <= w2543 and w2760;
w2810 <= not w2808 and not w2809;
w2811 <= not w2807 and w2810;
w2812 <= w2718 and w2767;
w2813 <= w2811 and not w2812;
w2814 <= not w971 and not w2813;
w2815 <= not w2813 and not w2814;
w2816 <= not w971 and not w2814;
w2817 <= not w2815 and not w2816;
w2818 <= not w2673 and not w2687;
w2819 <= not w2688 and not w2818;
w2820 <= not w2817 and w2819;
w2821 <= not w2664 and not w2672;
w2822 <= not w2673 and not w2821;
w2823 <= not w2550 and w2758;
w2824 <= w2546 and w2760;
w2825 <= w2543 and w2752;
w2826 <= not w2824 and not w2825;
w2827 <= not w2823 and w2826;
w2828 <= not w2767 and w2827;
w2829 <= w2656 and w2827;
w2830 <= not w2828 and not w2829;
w2831 <= w971 and not w2830;
w2832 <= not w971 and w2830;
w2833 <= not w2831 and not w2832;
w2834 <= w2822 and w2833;
w2835 <= not w2557 and w2760;
w2836 <= not w2554 and w2752;
w2837 <= not w2835 and not w2836;
w2838 <= not w2623 and w2767;
w2839 <= w2837 and not w2838;
w2840 <= not w971 and not w2839;
w2841 <= not w971 and not w2840;
w2842 <= not w2839 and not w2840;
w2843 <= not w2841 and not w2842;
w2844 <= not w2557 and not w2751;
w2845 <= not w971 and not w2844;
w2846 <= not w2843 and w2845;
w2847 <= not w2550 and w2752;
w2848 <= not w2557 and w2758;
w2849 <= not w2554 and w2760;
w2850 <= not w2848 and not w2849;
w2851 <= not w2847 and w2850;
w2852 <= not w2682 and w2851;
w2853 <= not w2767 and w2851;
w2854 <= not w2852 and not w2853;
w2855 <= w971 and not w2854;
w2856 <= not w971 and w2854;
w2857 <= not w2855 and not w2856;
w2858 <= w2846 and w2857;
w2859 <= w2663 and w2858;
w2860 <= w2858 and not w2859;
w2861 <= w2663 and not w2859;
w2862 <= not w2860 and not w2861;
w2863 <= not w2550 and w2760;
w2864 <= w2546 and w2752;
w2865 <= not w2554 and w2758;
w2866 <= not w2864 and not w2865;
w2867 <= not w2863 and w2866;
w2868 <= not w2700 and w2767;
w2869 <= w2867 and not w2868;
w2870 <= not w971 and not w2869;
w2871 <= not w971 and not w2870;
w2872 <= not w2869 and not w2870;
w2873 <= not w2871 and not w2872;
w2874 <= not w2862 and not w2873;
w2875 <= not w2859 and not w2874;
w2876 <= not w2822 and not w2833;
w2877 <= not w2834 and not w2876;
w2878 <= not w2875 and w2877;
w2879 <= not w2834 and not w2878;
w2880 <= not w2817 and not w2820;
w2881 <= w2819 and not w2820;
w2882 <= not w2880 and not w2881;
w2883 <= not w2879 and not w2882;
w2884 <= not w2820 and not w2883;
w2885 <= not w2792 and not w2806;
w2886 <= w2805 and not w2806;
w2887 <= not w2885 and not w2886;
w2888 <= not w2884 and not w2887;
w2889 <= not w2806 and not w2888;
w2890 <= not w2786 and not w2789;
w2891 <= w2788 and not w2789;
w2892 <= not w2890 and not w2891;
w2893 <= not w2889 and not w2892;
w2894 <= not w2789 and not w2893;
w2895 <= w2745 and not w2773;
w2896 <= w2772 and not w2773;
w2897 <= not w2895 and not w2896;
w2898 <= not w2894 and not w2897;
w2899 <= not w2773 and not w2898;
w2900 <= not w2536 and w2649;
w2901 <= w2543 and w2645;
w2902 <= not w2540 and w2647;
w2903 <= not w2901 and not w2902;
w2904 <= not w2900 and w2903;
w2905 <= w2640 and w2799;
w2906 <= w2904 and not w2905;
w2907 <= not w619 and not w2906;
w2908 <= w619 and w2906;
w2909 <= not w2907 and not w2908;
w2910 <= not w2550 and w2616;
w2911 <= w2546 and w2618;
w2912 <= not w2554 and w2726;
w2913 <= not w2911 and not w2912;
w2914 <= not w2910 and w2913;
w2915 <= w2624 and not w2700;
w2916 <= w2914 and not w2915;
w2917 <= not w475 and not w2916;
w2918 <= not w2916 and not w2917;
w2919 <= not w475 and not w2917;
w2920 <= not w2918 and not w2919;
w2921 <= not w475 and not w2557;
w2922 <= not w2737 and not w2921;
w2923 <= w2737 and w2921;
w2924 <= not w2920 and not w2923;
w2925 <= not w2922 and w2924;
w2926 <= not w2920 and not w2925;
w2927 <= not w2923 and not w2925;
w2928 <= not w2922 and w2927;
w2929 <= not w2926 and not w2928;
w2930 <= w2909 and not w2929;
w2931 <= w2909 and not w2930;
w2932 <= not w2929 and not w2930;
w2933 <= not w2931 and not w2932;
w2934 <= not w2740 and not w2744;
w2935 <= w2933 and w2934;
w2936 <= not w2933 and not w2934;
w2937 <= not w2935 and not w2936;
w2938 <= w2584 and not w2586;
w2939 <= not w2587 and not w2938;
w2940 <= not w2525 and w2752;
w2941 <= not w2532 and w2758;
w2942 <= w2528 and w2760;
w2943 <= not w2941 and not w2942;
w2944 <= not w2940 and w2943;
w2945 <= not w2939 and w2944;
w2946 <= not w2767 and w2944;
w2947 <= not w2945 and not w2946;
w2948 <= w971 and not w2947;
w2949 <= not w971 and w2947;
w2950 <= not w2948 and not w2949;
w2951 <= w2937 and w2950;
w2952 <= w2937 and not w2951;
w2953 <= w2950 and not w2951;
w2954 <= not w2952 and not w2953;
w2955 <= not w2899 and not w2954;
w2956 <= not w2899 and not w2955;
w2957 <= not w2954 and not w2955;
w2958 <= not w2956 and not w2957;
w2959 <= w2607 and not w2958;
w2960 <= w2607 and not w2959;
w2961 <= not w2958 and not w2959;
w2962 <= not w2960 and not w2961;
w2963 <= not w2894 and not w2898;
w2964 <= not w2897 and not w2898;
w2965 <= not w2963 and not w2964;
w2966 <= w245 and not w2516;
w2967 <= w2510 and not w2525;
w2968 <= w2512 and w2517;
w2969 <= not w2967 and not w2968;
w2970 <= not w2966 and w2969;
w2971 <= w2592 and not w2594;
w2972 <= not w2595 and not w2971;
w2973 <= w2521 and w2972;
w2974 <= w2970 and not w2973;
w2975 <= not w225 and not w2974;
w2976 <= w225 and w2974;
w2977 <= not w2975 and not w2976;
w2978 <= not w2965 and w2977;
w2979 <= w2977 and not w2978;
w2980 <= not w2965 and not w2978;
w2981 <= not w2979 and not w2980;
w2982 <= not w2889 and w2892;
w2983 <= w2889 and not w2892;
w2984 <= not w2982 and not w2983;
w2985 <= w245 and w2512;
w2986 <= w2510 and w2528;
w2987 <= w2517 and not w2525;
w2988 <= not w2986 and not w2987;
w2989 <= not w2985 and w2988;
w2990 <= not w2521 and w2989;
w2991 <= w2588 and not w2590;
w2992 <= not w2591 and not w2991;
w2993 <= w2989 and not w2992;
w2994 <= not w2990 and not w2993;
w2995 <= w225 and not w2994;
w2996 <= not w225 and w2994;
w2997 <= not w2995 and not w2996;
w2998 <= not w2984 and w2997;
w2999 <= not w2884 and not w2888;
w3000 <= not w2887 and not w2888;
w3001 <= not w2999 and not w3000;
w3002 <= w245 and not w2525;
w3003 <= w2510 and not w2532;
w3004 <= w2517 and w2528;
w3005 <= not w3003 and not w3004;
w3006 <= not w3002 and w3005;
w3007 <= not w2521 and w3006;
w3008 <= not w2939 and w3006;
w3009 <= not w3007 and not w3008;
w3010 <= w225 and not w3009;
w3011 <= not w225 and w3009;
w3012 <= not w3010 and not w3011;
w3013 <= not w3001 and w3012;
w3014 <= not w2879 and w2882;
w3015 <= w2879 and not w2882;
w3016 <= not w3014 and not w3015;
w3017 <= w245 and w2528;
w3018 <= w2510 and not w2536;
w3019 <= w2517 and not w2532;
w3020 <= not w3018 and not w3019;
w3021 <= not w3017 and w3020;
w3022 <= not w2521 and w3021;
w3023 <= not w2765 and w3021;
w3024 <= not w3022 and not w3023;
w3025 <= w225 and not w3024;
w3026 <= not w225 and w3024;
w3027 <= not w3025 and not w3026;
w3028 <= not w3016 and w3027;
w3029 <= w245 and not w2532;
w3030 <= w2510 and not w2540;
w3031 <= w2517 and not w2536;
w3032 <= not w3030 and not w3031;
w3033 <= not w3029 and w3032;
w3034 <= w2521 and w2780;
w3035 <= w3033 and not w3034;
w3036 <= not w225 and not w3035;
w3037 <= w225 and w3035;
w3038 <= not w3036 and not w3037;
w3039 <= w2875 and not w2877;
w3040 <= not w2878 and not w3039;
w3041 <= w3038 and w3040;
w3042 <= not w2862 and not w2874;
w3043 <= not w2873 and not w2874;
w3044 <= not w3042 and not w3043;
w3045 <= w245 and not w2536;
w3046 <= w2510 and w2543;
w3047 <= w2517 and not w2540;
w3048 <= not w3046 and not w3047;
w3049 <= not w3045 and w3048;
w3050 <= not w2521 and w3049;
w3051 <= not w2799 and w3049;
w3052 <= not w3050 and not w3051;
w3053 <= w225 and not w3052;
w3054 <= not w225 and w3052;
w3055 <= not w3053 and not w3054;
w3056 <= not w3044 and w3055;
w3057 <= w245 and not w2540;
w3058 <= w2510 and w2546;
w3059 <= w2517 and w2543;
w3060 <= not w3058 and not w3059;
w3061 <= not w3057 and w3060;
w3062 <= w2521 and w2718;
w3063 <= w3061 and not w3062;
w3064 <= not w225 and not w3063;
w3065 <= w225 and w3063;
w3066 <= not w3064 and not w3065;
w3067 <= not w2846 and not w2857;
w3068 <= not w2858 and not w3067;
w3069 <= w3066 and w3068;
w3070 <= w2843 and not w2845;
w3071 <= not w2846 and not w3070;
w3072 <= w2510 and not w2550;
w3073 <= w2517 and w2546;
w3074 <= w245 and w2543;
w3075 <= not w3073 and not w3074;
w3076 <= not w3072 and w3075;
w3077 <= not w2521 and w3076;
w3078 <= w2656 and w3076;
w3079 <= not w3077 and not w3078;
w3080 <= w225 and not w3079;
w3081 <= not w225 and w3079;
w3082 <= not w3080 and not w3081;
w3083 <= w3071 and w3082;
w3084 <= not w244 and not w2557;
w3085 <= not w225 and not w3084;
w3086 <= w2517 and not w2557;
w3087 <= w245 and not w2554;
w3088 <= not w3086 and not w3087;
w3089 <= w2521 and not w2623;
w3090 <= w3088 and not w3089;
w3091 <= not w225 and not w3090;
w3092 <= w225 and w3090;
w3093 <= not w3091 and not w3092;
w3094 <= w3085 and w3093;
w3095 <= w245 and not w2550;
w3096 <= w2510 and not w2557;
w3097 <= w2517 and not w2554;
w3098 <= not w3096 and not w3097;
w3099 <= not w3095 and w3098;
w3100 <= not w2521 and w3099;
w3101 <= not w2682 and w3099;
w3102 <= not w3100 and not w3101;
w3103 <= w225 and not w3102;
w3104 <= not w225 and w3102;
w3105 <= not w3103 and not w3104;
w3106 <= w3094 and w3105;
w3107 <= w2844 and w3106;
w3108 <= w3106 and not w3107;
w3109 <= w2844 and not w3107;
w3110 <= not w3108 and not w3109;
w3111 <= w2517 and not w2550;
w3112 <= w245 and w2546;
w3113 <= w2510 and not w2554;
w3114 <= not w3112 and not w3113;
w3115 <= not w3111 and w3114;
w3116 <= w2521 and not w2700;
w3117 <= w3115 and not w3116;
w3118 <= not w225 and not w3117;
w3119 <= w225 and w3117;
w3120 <= not w3118 and not w3119;
w3121 <= not w3110 and w3120;
w3122 <= not w3107 and not w3121;
w3123 <= not w3071 and not w3082;
w3124 <= not w3083 and not w3123;
w3125 <= not w3122 and w3124;
w3126 <= not w3083 and not w3125;
w3127 <= not w3066 and not w3068;
w3128 <= not w3069 and not w3127;
w3129 <= not w3126 and w3128;
w3130 <= not w3069 and not w3129;
w3131 <= not w3044 and not w3056;
w3132 <= w3055 and not w3056;
w3133 <= not w3131 and not w3132;
w3134 <= not w3130 and not w3133;
w3135 <= not w3056 and not w3134;
w3136 <= not w3038 and not w3040;
w3137 <= not w3041 and not w3136;
w3138 <= not w3135 and w3137;
w3139 <= not w3041 and not w3138;
w3140 <= not w3016 and not w3028;
w3141 <= w3027 and not w3028;
w3142 <= not w3140 and not w3141;
w3143 <= not w3139 and not w3142;
w3144 <= not w3028 and not w3143;
w3145 <= not w3001 and not w3013;
w3146 <= w3012 and not w3013;
w3147 <= not w3145 and not w3146;
w3148 <= not w3144 and not w3147;
w3149 <= not w3013 and not w3148;
w3150 <= w2984 and not w2997;
w3151 <= not w2998 and not w3150;
w3152 <= not w3149 and w3151;
w3153 <= not w2998 and not w3152;
w3154 <= not w2981 and not w3153;
w3155 <= not w2978 and not w3154;
w3156 <= w2962 and w3155;
w3157 <= not w2962 and not w3155;
w3158 <= not w3156 and not w3157;
w3159 <= a(0) and not a(22);
w3160 <= a(1) and not w3159;
w3161 <= not a(1) and w3159;
w3162 <= not w3160 and not w3161;
w3163 <= not w241 and w3162;
w3164 <= w241 and not w3162;
w3165 <= not w3163 and not w3164;
w3166 <= a(0) and not w3165;
w3167 <= a(0) and w3165;
w3168 <= not w274 and w759;
w3169 <= w435 and w3168;
w3170 <= w381 and w3169;
w3171 <= w2194 and w3170;
w3172 <= w2283 and w3171;
w3173 <= w2368 and w3172;
w3174 <= w926 and w3173;
w3175 <= not w454 and w3174;
w3176 <= not w247 and w3175;
w3177 <= not w162 and w3176;
w3178 <= not w208 and w3177;
w3179 <= not w187 and w3178;
w3180 <= not w250 and w758;
w3181 <= not w276 and w3180;
w3182 <= w150 and w3181;
w3183 <= w2116 and w3182;
w3184 <= not w365 and w3183;
w3185 <= not w176 and w3184;
w3186 <= not w163 and w3185;
w3187 <= not w320 and w3186;
w3188 <= not w397 and w3187;
w3189 <= not w285 and w3188;
w3190 <= not w64 and w3189;
w3191 <= not w308 and w3190;
w3192 <= not w56 and w3191;
w3193 <= not w292 and w3192;
w3194 <= w694 and w2316;
w3195 <= w106 and w3194;
w3196 <= w718 and w3195;
w3197 <= w3193 and w3196;
w3198 <= w160 and w3197;
w3199 <= not w100 and w3198;
w3200 <= not w126 and w3199;
w3201 <= not w170 and w3200;
w3202 <= not w177 and w3201;
w3203 <= not w136 and w3202;
w3204 <= not w396 and w3203;
w3205 <= not w311 and w3204;
w3206 <= not w427 and w3205;
w3207 <= w2502 and w3206;
w3208 <= w3179 and w3207;
w3209 <= not w84 and not w355;
w3210 <= w299 and w373;
w3211 <= w1115 and w3210;
w3212 <= w347 and w3211;
w3213 <= w387 and w3212;
w3214 <= w264 and w3213;
w3215 <= w435 and w3214;
w3216 <= w452 and w3215;
w3217 <= w403 and w3216;
w3218 <= w3209 and w3217;
w3219 <= not w90 and w3218;
w3220 <= not w3208 and w3219;
w3221 <= w3208 and not w3219;
w3222 <= not w3220 and not w3221;
w3223 <= w3167 and w3222;
w3224 <= w238 and not w3165;
w3225 <= not w2502 and w3206;
w3226 <= w2502 and not w3206;
w3227 <= not w3225 and not w3226;
w3228 <= w3224 and w3227;
w3229 <= not w3179 and not w3207;
w3230 <= not w3208 and not w3229;
w3231 <= not a(0) and not w3162;
w3232 <= not w3230 and w3231;
w3233 <= not w3228 and not w3232;
w3234 <= not w3223 and w3233;
w3235 <= not w3166 and w3234;
w3236 <= w3227 and not w3230;
w3237 <= not w2504 and w3227;
w3238 <= not w2597 and not w2600;
w3239 <= w2504 and not w3227;
w3240 <= not w3237 and not w3239;
w3241 <= not w3238 and w3240;
w3242 <= not w3237 and not w3241;
w3243 <= not w3227 and w3230;
w3244 <= not w3236 and not w3243;
w3245 <= not w3242 and w3244;
w3246 <= not w3236 and not w3245;
w3247 <= not w3222 and w3230;
w3248 <= w3222 and not w3230;
w3249 <= not w3247 and not w3248;
w3250 <= not w3246 and w3249;
w3251 <= w3246 and not w3249;
w3252 <= not w3250 and not w3251;
w3253 <= w3234 and not w3252;
w3254 <= not w3235 and not w3253;
w3255 <= w241 and not w3254;
w3256 <= not w241 and w3254;
w3257 <= not w3255 and not w3256;
w3258 <= w3158 and w3257;
w3259 <= w2981 and w3153;
w3260 <= not w3154 and not w3259;
w3261 <= w3167 and not w3230;
w3262 <= not w2504 and w3224;
w3263 <= w3227 and w3231;
w3264 <= not w3262 and not w3263;
w3265 <= not w3261 and w3264;
w3266 <= not w3166 and w3265;
w3267 <= w3242 and not w3244;
w3268 <= not w3245 and not w3267;
w3269 <= w3265 and not w3268;
w3270 <= not w3266 and not w3269;
w3271 <= w241 and not w3270;
w3272 <= not w241 and w3270;
w3273 <= not w3271 and not w3272;
w3274 <= w3260 and w3273;
w3275 <= w3149 and not w3151;
w3276 <= w3167 and w3227;
w3277 <= not w2516 and w3224;
w3278 <= not w2504 and w3231;
w3279 <= not w3277 and not w3278;
w3280 <= not w3276 and w3279;
w3281 <= w3238 and not w3240;
w3282 <= not w3241 and not w3281;
w3283 <= w3166 and w3282;
w3284 <= w3280 and not w3283;
w3285 <= not w241 and not w3284;
w3286 <= not w3284 and not w3285;
w3287 <= not w241 and not w3285;
w3288 <= not w3286 and not w3287;
w3289 <= w2512 and w3167;
w3290 <= w2528 and w3224;
w3291 <= not w2525 and w3231;
w3292 <= not w3290 and not w3291;
w3293 <= not w3289 and w3292;
w3294 <= not w241 and not w3293;
w3295 <= w2992 and w3166;
w3296 <= w3293 and not w3295;
w3297 <= w241 and w3296;
w3298 <= not w241 and w3166;
w3299 <= w2992 and w3298;
w3300 <= not w2525 and w3167;
w3301 <= not w2532 and w3224;
w3302 <= w2528 and w3231;
w3303 <= not w3301 and not w3302;
w3304 <= not w3300 and w3303;
w3305 <= not w241 and not w3304;
w3306 <= w2939 and w3166;
w3307 <= w3304 and not w3306;
w3308 <= w241 and w3307;
w3309 <= w2939 and w3298;
w3310 <= w2528 and w3167;
w3311 <= not w2536 and w3224;
w3312 <= not w2532 and w3231;
w3313 <= not w3311 and not w3312;
w3314 <= not w3310 and w3313;
w3315 <= not w241 and not w3314;
w3316 <= w2765 and w3166;
w3317 <= w3314 and not w3316;
w3318 <= w241 and w3317;
w3319 <= w2765 and w3298;
w3320 <= w3122 and not w3124;
w3321 <= not w2536 and w3167;
w3322 <= w2543 and w3224;
w3323 <= not w2540 and w3231;
w3324 <= not w3322 and not w3323;
w3325 <= not w3321 and w3324;
w3326 <= not w241 and not w3325;
w3327 <= w2799 and w3166;
w3328 <= w3325 and not w3327;
w3329 <= w241 and w3328;
w3330 <= w2799 and w3298;
w3331 <= not w3094 and not w3105;
w3332 <= not w2550 and w3224;
w3333 <= w2546 and w3231;
w3334 <= w2543 and w3167;
w3335 <= not w3333 and not w3334;
w3336 <= not w3332 and w3335;
w3337 <= not w241 and not w3336;
w3338 <= not w2656 and w3166;
w3339 <= w3336 and not w3338;
w3340 <= w241 and w3339;
w3341 <= not w2656 and w3298;
w3342 <= a(0) and not w2557;
w3343 <= w2682 and w3298;
w3344 <= not w2550 and w3167;
w3345 <= not w2557 and w3224;
w3346 <= not w2554 and w3231;
w3347 <= not w3345 and not w3346;
w3348 <= not w3344 and w3347;
w3349 <= not w241 and not w3348;
w3350 <= not w2623 and w3298;
w3351 <= not w2554 and w3167;
w3352 <= not w2557 and w3231;
w3353 <= not w241 and not w3352;
w3354 <= not w3351 and w3353;
w3355 <= not w3350 and w3354;
w3356 <= not w3349 and w3355;
w3357 <= not w3343 and w3356;
w3358 <= not w3342 and w3357;
w3359 <= not w3084 and not w3358;
w3360 <= not w2550 and w3231;
w3361 <= w2546 and w3167;
w3362 <= not w2554 and w3224;
w3363 <= not w3361 and not w3362;
w3364 <= not w3360 and w3363;
w3365 <= not w2700 and w3166;
w3366 <= w3364 and not w3365;
w3367 <= not w241 and not w3366;
w3368 <= w241 and w3366;
w3369 <= not w3367 and not w3368;
w3370 <= not w3359 and w3369;
w3371 <= w3084 and w3358;
w3372 <= not w3370 and not w3371;
w3373 <= not w3085 and not w3093;
w3374 <= not w3094 and not w3373;
w3375 <= w3372 and not w3374;
w3376 <= not w3341 and not w3375;
w3377 <= not w3340 and w3376;
w3378 <= not w3337 and w3377;
w3379 <= not w3372 and w3374;
w3380 <= not w3378 and not w3379;
w3381 <= not w2540 and w3167;
w3382 <= w2546 and w3224;
w3383 <= w2543 and w3231;
w3384 <= not w3382 and not w3383;
w3385 <= not w3381 and w3384;
w3386 <= w2718 and w3166;
w3387 <= w3385 and not w3386;
w3388 <= not w241 and not w3387;
w3389 <= not w3387 and not w3388;
w3390 <= not w241 and not w3388;
w3391 <= not w3389 and not w3390;
w3392 <= w3380 and w3391;
w3393 <= not w3106 and not w3392;
w3394 <= not w3331 and w3393;
w3395 <= not w3380 and not w3391;
w3396 <= not w3394 and not w3395;
w3397 <= not w3110 and not w3121;
w3398 <= w3120 and not w3121;
w3399 <= not w3397 and not w3398;
w3400 <= w3396 and w3399;
w3401 <= not w3330 and not w3400;
w3402 <= not w3329 and w3401;
w3403 <= not w3326 and w3402;
w3404 <= not w3396 and not w3399;
w3405 <= not w3403 and not w3404;
w3406 <= not w2532 and w3167;
w3407 <= not w2540 and w3224;
w3408 <= not w2536 and w3231;
w3409 <= not w3407 and not w3408;
w3410 <= not w3406 and w3409;
w3411 <= w2780 and w3166;
w3412 <= w3410 and not w3411;
w3413 <= not w241 and not w3412;
w3414 <= not w3412 and not w3413;
w3415 <= not w241 and not w3413;
w3416 <= not w3414 and not w3415;
w3417 <= w3405 and w3416;
w3418 <= not w3125 and not w3417;
w3419 <= not w3320 and w3418;
w3420 <= not w3405 and not w3416;
w3421 <= not w3419 and not w3420;
w3422 <= w3126 and not w3128;
w3423 <= not w3129 and not w3422;
w3424 <= w3421 and not w3423;
w3425 <= not w3319 and not w3424;
w3426 <= not w3318 and w3425;
w3427 <= not w3315 and w3426;
w3428 <= not w3421 and w3423;
w3429 <= not w3427 and not w3428;
w3430 <= not w3130 and not w3134;
w3431 <= not w3133 and not w3134;
w3432 <= not w3430 and not w3431;
w3433 <= w3429 and w3432;
w3434 <= not w3309 and not w3433;
w3435 <= not w3308 and w3434;
w3436 <= not w3305 and w3435;
w3437 <= not w3429 and not w3432;
w3438 <= not w3436 and not w3437;
w3439 <= w3135 and not w3137;
w3440 <= not w3138 and not w3439;
w3441 <= w3438 and not w3440;
w3442 <= not w3299 and not w3441;
w3443 <= not w3297 and w3442;
w3444 <= not w3294 and w3443;
w3445 <= not w3438 and w3440;
w3446 <= not w3444 and not w3445;
w3447 <= w3139 and w3142;
w3448 <= not w3143 and not w3447;
w3449 <= not w3446 and w3448;
w3450 <= not w2516 and w3167;
w3451 <= not w2525 and w3224;
w3452 <= w2512 and w3231;
w3453 <= not w3451 and not w3452;
w3454 <= not w3450 and w3453;
w3455 <= w2972 and w3166;
w3456 <= w3454 and not w3455;
w3457 <= w241 and not w3456;
w3458 <= not w241 and w3456;
w3459 <= not w3457 and not w3458;
w3460 <= not w3449 and w3459;
w3461 <= w3446 and not w3448;
w3462 <= not w3460 and not w3461;
w3463 <= w3144 and w3147;
w3464 <= not w3148 and not w3463;
w3465 <= not w3462 and not w3464;
w3466 <= not w2504 and w3167;
w3467 <= w2512 and w3224;
w3468 <= not w2516 and w3231;
w3469 <= not w3467 and not w3468;
w3470 <= not w3466 and w3469;
w3471 <= w2602 and w3166;
w3472 <= w3470 and not w3471;
w3473 <= not w241 and not w3472;
w3474 <= w241 and w3472;
w3475 <= not w3473 and not w3474;
w3476 <= not w3465 and w3475;
w3477 <= w3462 and w3464;
w3478 <= not w3476 and not w3477;
w3479 <= w3288 and w3478;
w3480 <= not w3152 and not w3479;
w3481 <= not w3275 and w3480;
w3482 <= not w3288 and not w3478;
w3483 <= not w3481 and not w3482;
w3484 <= w3260 and not w3274;
w3485 <= w3273 and not w3274;
w3486 <= not w3484 and not w3485;
w3487 <= not w3483 and not w3486;
w3488 <= not w3274 and not w3487;
w3489 <= w3158 and not w3258;
w3490 <= w3257 and not w3258;
w3491 <= not w3489 and not w3490;
w3492 <= not w3488 and not w3491;
w3493 <= not w3258 and not w3492;
w3494 <= not w2959 and not w3157;
w3495 <= w245 and w3227;
w3496 <= w2510 and not w2516;
w3497 <= not w2504 and w2517;
w3498 <= not w3496 and not w3497;
w3499 <= not w3495 and w3498;
w3500 <= w2521 and w3282;
w3501 <= w3499 and not w3500;
w3502 <= not w225 and not w3501;
w3503 <= w225 and w3501;
w3504 <= not w3502 and not w3503;
w3505 <= not w2951 and not w2955;
w3506 <= not w2930 and not w2936;
w3507 <= not w2532 and w2649;
w3508 <= not w2540 and w2645;
w3509 <= not w2536 and w2647;
w3510 <= not w3508 and not w3509;
w3511 <= not w3507 and w3510;
w3512 <= w2640 and w2780;
w3513 <= w3511 and not w3512;
w3514 <= not w619 and not w3513;
w3515 <= w619 and w3513;
w3516 <= not w3514 and not w3515;
w3517 <= not w475 and not w2554;
w3518 <= not w2550 and w2726;
w3519 <= w2546 and w2616;
w3520 <= w2543 and w2618;
w3521 <= not w3519 and not w3520;
w3522 <= not w3518 and w3521;
w3523 <= w2624 and not w2656;
w3524 <= w3522 and not w3523;
w3525 <= not w475 and not w3524;
w3526 <= w3517 and not w3525;
w3527 <= w3517 and not w3526;
w3528 <= w475 and w3524;
w3529 <= not w3525 and not w3528;
w3530 <= not w3526 and w3529;
w3531 <= not w3527 and not w3530;
w3532 <= not w2927 and not w3531;
w3533 <= not w2927 and not w3532;
w3534 <= not w3531 and not w3532;
w3535 <= not w3533 and not w3534;
w3536 <= w3516 and not w3535;
w3537 <= w3516 and not w3536;
w3538 <= not w3535 and not w3536;
w3539 <= not w3537 and not w3538;
w3540 <= not w3506 and w3539;
w3541 <= w3506 and not w3539;
w3542 <= not w3540 and not w3541;
w3543 <= w2512 and w2752;
w3544 <= w2528 and w2758;
w3545 <= not w2525 and w2760;
w3546 <= not w3544 and not w3545;
w3547 <= not w3543 and w3546;
w3548 <= not w2992 and w3547;
w3549 <= not w2767 and w3547;
w3550 <= not w3548 and not w3549;
w3551 <= w971 and not w3550;
w3552 <= not w971 and w3550;
w3553 <= not w3551 and not w3552;
w3554 <= not w3542 and w3553;
w3555 <= w3542 and not w3553;
w3556 <= not w3554 and not w3555;
w3557 <= not w3505 and w3556;
w3558 <= w3505 and not w3556;
w3559 <= not w3557 and not w3558;
w3560 <= w3504 and w3559;
w3561 <= not w3504 and not w3559;
w3562 <= not w3560 and not w3561;
w3563 <= not w3494 and w3562;
w3564 <= w3494 and not w3562;
w3565 <= not w3563 and not w3564;
w3566 <= not w298 and w452;
w3567 <= not w98 and w3566;
w3568 <= w464 and w3567;
w3569 <= w435 and w3568;
w3570 <= w364 and w3569;
w3571 <= w354 and w3570;
w3572 <= not w138 and w3571;
w3573 <= not w169 and w3572;
w3574 <= not w174 and w3573;
w3575 <= w3208 and w3219;
w3576 <= not w3574 and not w3575;
w3577 <= w3574 and w3575;
w3578 <= not w3576 and not w3577;
w3579 <= w3167 and not w3578;
w3580 <= w3224 and not w3230;
w3581 <= w3222 and w3231;
w3582 <= not w3580 and not w3581;
w3583 <= not w3579 and w3582;
w3584 <= not w3166 and w3583;
w3585 <= not w3248 and not w3250;
w3586 <= not w3222 and w3578;
w3587 <= w3222 and not w3578;
w3588 <= not w3586 and not w3587;
w3589 <= not w3585 and w3588;
w3590 <= w3585 and not w3588;
w3591 <= not w3589 and not w3590;
w3592 <= w3583 and not w3591;
w3593 <= not w3584 and not w3592;
w3594 <= w241 and not w3593;
w3595 <= not w241 and w3593;
w3596 <= not w3594 and not w3595;
w3597 <= w3565 and w3596;
w3598 <= not w3565 and not w3596;
w3599 <= not w3597 and not w3598;
w3600 <= not w3493 and w3599;
w3601 <= w3493 and not w3599;
w3602 <= not w3600 and not w3601;
w3603 <= not w221 and w3602;
w3604 <= not w64 and not w456;
w3605 <= not w686 and w3604;
w3606 <= not w246 and w3605;
w3607 <= not w104 and w3606;
w3608 <= w756 and w3607;
w3609 <= not w89 and w3608;
w3610 <= not w100 and w3609;
w3611 <= not w136 and w3610;
w3612 <= not w263 and w3611;
w3613 <= not w83 and w3612;
w3614 <= not w309 and w3613;
w3615 <= not w92 and w3614;
w3616 <= not w56 and w3615;
w3617 <= w322 and w455;
w3618 <= w1084 and w3617;
w3619 <= not w167 and w3618;
w3620 <= not w205 and w3619;
w3621 <= not w445 and w3620;
w3622 <= not w503 and w3621;
w3623 <= not w395 and w3622;
w3624 <= not w421 and w3623;
w3625 <= not w165 and w3624;
w3626 <= w739 and w3625;
w3627 <= not w367 and w3626;
w3628 <= not w248 and w3627;
w3629 <= w2404 and w3628;
w3630 <= w3616 and w3629;
w3631 <= w930 and w3630;
w3632 <= not w87 and w3631;
w3633 <= not w204 and w3632;
w3634 <= not w277 and w3633;
w3635 <= not w396 and w3634;
w3636 <= not w96 and w3635;
w3637 <= not w247 and w3636;
w3638 <= not w285 and w3637;
w3639 <= not w420 and w3638;
w3640 <= not w292 and w3639;
w3641 <= w3488 and not w3490;
w3642 <= not w3489 and w3641;
w3643 <= not w3492 and not w3642;
w3644 <= w347 and w2228;
w3645 <= w2253 and w3644;
w3646 <= not w94 and w3645;
w3647 <= not w453 and w3646;
w3648 <= not w306 and w3647;
w3649 <= not w427 and w3648;
w3650 <= w291 and w763;
w3651 <= not w87 and w3650;
w3652 <= not w105 and w3651;
w3653 <= w410 and w2372;
w3654 <= w2383 and w3653;
w3655 <= w294 and w3654;
w3656 <= w3652 and w3655;
w3657 <= w3649 and w3656;
w3658 <= w2314 and w3657;
w3659 <= not w365 and w3658;
w3660 <= not w100 and w3659;
w3661 <= not w267 and w3660;
w3662 <= not w169 and w3661;
w3663 <= not w124 and w3662;
w3664 <= not w168 and w3663;
w3665 <= not w252 and w3664;
w3666 <= w3483 and w3486;
w3667 <= not w3487 and not w3666;
w3668 <= not w3665 and w3667;
w3669 <= not w3643 and not w3668;
w3670 <= not w3640 and not w3669;
w3671 <= w3643 and w3668;
w3672 <= not w3670 and not w3671;
w3673 <= not w221 and not w3603;
w3674 <= w3602 and not w3603;
w3675 <= not w3673 and not w3674;
w3676 <= not w3672 and not w3675;
w3677 <= not w3603 and not w3676;
w3678 <= w189 and w540;
w3679 <= not w300 and w3678;
w3680 <= not w73 and w3679;
w3681 <= not w263 and w3680;
w3682 <= not w157 and w3681;
w3683 <= not w395 and w3682;
w3684 <= not w419 and w3683;
w3685 <= w303 and not w418;
w3686 <= w284 and w3685;
w3687 <= w1112 and w3686;
w3688 <= w3684 and w3687;
w3689 <= w2368 and w3688;
w3690 <= not w172 and w3689;
w3691 <= not w267 and w3690;
w3692 <= not w127 and w3691;
w3693 <= not w168 and w3692;
w3694 <= not w504 and w3693;
w3695 <= not w161 and w3694;
w3696 <= not w82 and w3695;
w3697 <= not w173 and w3696;
w3698 <= not w3577 and w3697;
w3699 <= w3577 and not w3697;
w3700 <= not w3698 and not w3699;
w3701 <= w3167 and w3700;
w3702 <= w3222 and w3224;
w3703 <= w3231 and not w3578;
w3704 <= not w3702 and not w3703;
w3705 <= not w3701 and w3704;
w3706 <= not w3587 and not w3589;
w3707 <= w3578 and not w3700;
w3708 <= not w3578 and w3700;
w3709 <= not w3707 and not w3708;
w3710 <= not w3706 and w3709;
w3711 <= w3706 and not w3709;
w3712 <= not w3710 and not w3711;
w3713 <= w3166 and w3712;
w3714 <= w3705 and not w3713;
w3715 <= not w241 and not w3714;
w3716 <= not w3714 and not w3715;
w3717 <= not w241 and not w3715;
w3718 <= not w3716 and not w3717;
w3719 <= not w3560 and not w3563;
w3720 <= not w2516 and w2752;
w3721 <= not w2525 and w2758;
w3722 <= w2512 and w2760;
w3723 <= not w3721 and not w3722;
w3724 <= not w3720 and w3723;
w3725 <= w2767 and w2972;
w3726 <= w3724 and not w3725;
w3727 <= not w971 and not w3726;
w3728 <= not w3726 and not w3727;
w3729 <= not w971 and not w3727;
w3730 <= not w3728 and not w3729;
w3731 <= not w3506 and not w3539;
w3732 <= not w3536 and not w3731;
w3733 <= not w3526 and not w3532;
w3734 <= not w2540 and w2618;
w3735 <= w2546 and w2726;
w3736 <= w2543 and w2616;
w3737 <= not w3735 and not w3736;
w3738 <= not w3734 and w3737;
w3739 <= w2624 and w2718;
w3740 <= w3738 and not w3739;
w3741 <= not w475 and w2550;
w3742 <= not w3740 and w3741;
w3743 <= w3740 and not w3741;
w3744 <= not w3742 and not w3743;
w3745 <= not w3733 and w3744;
w3746 <= w3733 and not w3744;
w3747 <= not w3745 and not w3746;
w3748 <= w2528 and w2649;
w3749 <= not w2536 and w2645;
w3750 <= not w2532 and w2647;
w3751 <= not w3749 and not w3750;
w3752 <= not w3748 and w3751;
w3753 <= not w2640 and w3752;
w3754 <= not w2765 and w3752;
w3755 <= not w3753 and not w3754;
w3756 <= w619 and not w3755;
w3757 <= not w619 and w3755;
w3758 <= not w3756 and not w3757;
w3759 <= w3747 and w3758;
w3760 <= w3747 and not w3759;
w3761 <= w3758 and not w3759;
w3762 <= not w3760 and not w3761;
w3763 <= not w3732 and not w3762;
w3764 <= not w3732 and not w3763;
w3765 <= not w3762 and not w3763;
w3766 <= not w3764 and not w3765;
w3767 <= not w3730 and not w3766;
w3768 <= not w3730 and not w3767;
w3769 <= not w3766 and not w3767;
w3770 <= not w3768 and not w3769;
w3771 <= not w3554 and not w3557;
w3772 <= w3770 and w3771;
w3773 <= not w3770 and not w3771;
w3774 <= not w3772 and not w3773;
w3775 <= w245 and not w3230;
w3776 <= not w2504 and w2510;
w3777 <= w2517 and w3227;
w3778 <= not w3776 and not w3777;
w3779 <= not w3775 and w3778;
w3780 <= not w2521 and w3779;
w3781 <= not w3268 and w3779;
w3782 <= not w3780 and not w3781;
w3783 <= w225 and not w3782;
w3784 <= not w225 and w3782;
w3785 <= not w3783 and not w3784;
w3786 <= w3774 and w3785;
w3787 <= w3774 and not w3786;
w3788 <= w3785 and not w3786;
w3789 <= not w3787 and not w3788;
w3790 <= not w3719 and not w3789;
w3791 <= not w3719 and not w3790;
w3792 <= not w3789 and not w3790;
w3793 <= not w3791 and not w3792;
w3794 <= not w3718 and not w3793;
w3795 <= not w3718 and not w3794;
w3796 <= not w3793 and not w3794;
w3797 <= not w3795 and not w3796;
w3798 <= not w3597 and not w3600;
w3799 <= w3797 and w3798;
w3800 <= not w3797 and not w3798;
w3801 <= not w3799 and not w3800;
w3802 <= w189 and w1043;
w3803 <= w756 and w3802;
w3804 <= w1409 and w3803;
w3805 <= w2261 and w3804;
w3806 <= w593 and w3805;
w3807 <= w573 and w3806;
w3808 <= w160 and w3807;
w3809 <= not w205 and w3808;
w3810 <= not w98 and w3809;
w3811 <= not w295 and w3810;
w3812 <= not w3801 and w3811;
w3813 <= w3801 and not w3811;
w3814 <= not w3812 and not w3813;
w3815 <= not w3677 and w3814;
w3816 <= w3677 and not w3814;
w3817 <= not w3815 and not w3816;
w3818 <= not w3672 and not w3676;
w3819 <= not w3675 and not w3676;
w3820 <= not w3818 and not w3819;
w3821 <= w3817 and not w3820;
w3822 <= w3817 and not w3821;
w3823 <= not w3820 and not w3821;
w3824 <= not w3822 and not w3823;
w3825 <= not w3813 and not w3815;
w3826 <= w3577 and w3697;
w3827 <= w186 and w2383;
w3828 <= w407 and w3827;
w3829 <= w703 and w3828;
w3830 <= not w119 and w3829;
w3831 <= not w68 and w3830;
w3832 <= not w116 and w3831;
w3833 <= not w118 and w3832;
w3834 <= w266 and w505;
w3835 <= w765 and w3834;
w3836 <= w1426 and w3835;
w3837 <= w3833 and w3836;
w3838 <= w2382 and w3837;
w3839 <= w926 and w3838;
w3840 <= not w445 and w3839;
w3841 <= not w420 and w3840;
w3842 <= not w317 and w3841;
w3843 <= not w276 and w3842;
w3844 <= not w3826 and w3843;
w3845 <= w3826 and not w3843;
w3846 <= not w3844 and not w3845;
w3847 <= w3167 and w3846;
w3848 <= w3224 and not w3578;
w3849 <= w3231 and w3700;
w3850 <= not w3848 and not w3849;
w3851 <= not w3847 and w3850;
w3852 <= not w3708 and not w3710;
w3853 <= not w3700 and not w3846;
w3854 <= w3700 and w3846;
w3855 <= not w3853 and not w3854;
w3856 <= not w3852 and w3855;
w3857 <= w3852 and not w3855;
w3858 <= not w3856 and not w3857;
w3859 <= w3166 and w3858;
w3860 <= w3851 and not w3859;
w3861 <= not w241 and not w3860;
w3862 <= not w3860 and not w3861;
w3863 <= not w241 and not w3861;
w3864 <= not w3862 and not w3863;
w3865 <= not w3786 and not w3790;
w3866 <= not w2504 and w2752;
w3867 <= w2512 and w2758;
w3868 <= not w2516 and w2760;
w3869 <= not w3867 and not w3868;
w3870 <= not w3866 and w3869;
w3871 <= w2602 and w2767;
w3872 <= w3870 and not w3871;
w3873 <= not w971 and not w3872;
w3874 <= not w3872 and not w3873;
w3875 <= not w971 and not w3873;
w3876 <= not w3874 and not w3875;
w3877 <= not w3759 and not w3763;
w3878 <= not w475 and not w2550;
w3879 <= w3740 and w3878;
w3880 <= not w3745 and not w3879;
w3881 <= not w2536 and w2618;
w3882 <= w2543 and w2726;
w3883 <= not w2540 and w2616;
w3884 <= not w3882 and not w3883;
w3885 <= not w3881 and w3884;
w3886 <= w2624 and w2799;
w3887 <= w3885 and not w3886;
w3888 <= not w475 and not w2546;
w3889 <= not w3887 and w3888;
w3890 <= w3887 and not w3888;
w3891 <= not w3889 and not w3890;
w3892 <= not w3880 and w3891;
w3893 <= not w3880 and not w3892;
w3894 <= w3891 and not w3892;
w3895 <= not w3893 and not w3894;
w3896 <= not w2525 and w2649;
w3897 <= not w2532 and w2645;
w3898 <= w2528 and w2647;
w3899 <= not w3897 and not w3898;
w3900 <= not w3896 and w3899;
w3901 <= not w2640 and w3900;
w3902 <= not w2939 and w3900;
w3903 <= not w3901 and not w3902;
w3904 <= w619 and not w3903;
w3905 <= not w619 and w3903;
w3906 <= not w3904 and not w3905;
w3907 <= not w3895 and w3906;
w3908 <= not w3895 and not w3907;
w3909 <= w3906 and not w3907;
w3910 <= not w3908 and not w3909;
w3911 <= not w3877 and not w3910;
w3912 <= not w3877 and not w3911;
w3913 <= not w3910 and not w3911;
w3914 <= not w3912 and not w3913;
w3915 <= not w3876 and not w3914;
w3916 <= not w3876 and not w3915;
w3917 <= not w3914 and not w3915;
w3918 <= not w3916 and not w3917;
w3919 <= not w3767 and not w3773;
w3920 <= w3918 and w3919;
w3921 <= not w3918 and not w3919;
w3922 <= not w3920 and not w3921;
w3923 <= w245 and w3222;
w3924 <= w2510 and w3227;
w3925 <= w2517 and not w3230;
w3926 <= not w3924 and not w3925;
w3927 <= not w3923 and w3926;
w3928 <= not w2521 and w3927;
w3929 <= not w3252 and w3927;
w3930 <= not w3928 and not w3929;
w3931 <= w225 and not w3930;
w3932 <= not w225 and w3930;
w3933 <= not w3931 and not w3932;
w3934 <= w3922 and w3933;
w3935 <= w3922 and not w3934;
w3936 <= w3933 and not w3934;
w3937 <= not w3935 and not w3936;
w3938 <= not w3865 and not w3937;
w3939 <= not w3865 and not w3938;
w3940 <= not w3937 and not w3938;
w3941 <= not w3939 and not w3940;
w3942 <= not w3864 and not w3941;
w3943 <= not w3864 and not w3942;
w3944 <= not w3941 and not w3942;
w3945 <= not w3943 and not w3944;
w3946 <= not w3794 and not w3800;
w3947 <= w3945 and w3946;
w3948 <= not w3945 and not w3946;
w3949 <= not w3947 and not w3948;
w3950 <= not w90 and not w355;
w3951 <= not w311 and w3950;
w3952 <= not w208 and w3951;
w3953 <= w587 and w2290;
w3954 <= w2226 and w3953;
w3955 <= w199 and w3954;
w3956 <= w703 and w3955;
w3957 <= w3952 and w3956;
w3958 <= w160 and w3957;
w3959 <= w3181 and w3958;
w3960 <= not w125 and w3959;
w3961 <= not w105 and w3960;
w3962 <= not w277 and w3961;
w3963 <= not w141 and w3962;
w3964 <= not w68 and w3963;
w3965 <= not w395 and w3964;
w3966 <= not w3949 and w3965;
w3967 <= w3949 and not w3965;
w3968 <= not w3966 and not w3967;
w3969 <= not w3825 and w3968;
w3970 <= w3825 and not w3968;
w3971 <= not w3969 and not w3970;
w3972 <= w3821 and w3971;
w3973 <= not w3821 and not w3971;
w3974 <= not w3972 and not w3973;
w3975 <= a(22) and not a(23);
w3976 <= not a(22) and a(23);
w3977 <= not w3975 and not w3976;
w3978 <= not w3824 and not w3977;
w3979 <= not w3974 and w3978;
w3980 <= w3974 and not w3978;
w3981 <= not w3979 and not w3980;
w3982 <= not w3967 and not w3969;
w3983 <= w296 and not w358;
w3984 <= not w79 and w3983;
w3985 <= not w178 and w3984;
w3986 <= not w92 and w3985;
w3987 <= not w82 and w3986;
w3988 <= w366 and w558;
w3989 <= w755 and w3988;
w3990 <= w3987 and w3989;
w3991 <= w3649 and w3990;
w3992 <= not w263 and w3991;
w3993 <= not w408 and w3992;
w3994 <= not w454 and w3993;
w3995 <= not w248 and w3994;
w3996 <= not w96 and w3995;
w3997 <= not w456 and w3996;
w3998 <= not w276 and w3997;
w3999 <= not w3942 and not w3948;
w4000 <= w3224 and w3700;
w4001 <= w3231 and w3846;
w4002 <= not w4000 and not w4001;
w4003 <= not w3700 and not w3856;
w4004 <= w3846 and not w4003;
w4005 <= not w3846 and not w3856;
w4006 <= not w4004 and not w4005;
w4007 <= w3166 and w4006;
w4008 <= w4002 and not w4007;
w4009 <= not w241 and not w4008;
w4010 <= not w4008 and not w4009;
w4011 <= not w241 and not w4009;
w4012 <= not w4010 and not w4011;
w4013 <= not w3934 and not w3938;
w4014 <= w2752 and w3227;
w4015 <= not w2516 and w2758;
w4016 <= not w2504 and w2760;
w4017 <= not w4015 and not w4016;
w4018 <= not w4014 and w4017;
w4019 <= w2767 and w3282;
w4020 <= w4018 and not w4019;
w4021 <= not w971 and not w4020;
w4022 <= not w4020 and not w4021;
w4023 <= not w971 and not w4021;
w4024 <= not w4022 and not w4023;
w4025 <= not w3907 and not w3911;
w4026 <= not w475 and w3887;
w4027 <= w2546 and w4026;
w4028 <= not w3892 and not w4027;
w4029 <= not w2532 and w2618;
w4030 <= not w2540 and w2726;
w4031 <= not w2536 and w2616;
w4032 <= not w4030 and not w4031;
w4033 <= not w4029 and w4032;
w4034 <= w2624 and w2780;
w4035 <= w4033 and not w4034;
w4036 <= not w475 and not w2543;
w4037 <= not w4035 and w4036;
w4038 <= w4035 and not w4036;
w4039 <= not w4037 and not w4038;
w4040 <= not w4028 and w4039;
w4041 <= not w4028 and not w4040;
w4042 <= w4039 and not w4040;
w4043 <= not w4041 and not w4042;
w4044 <= w2512 and w2649;
w4045 <= w2528 and w2645;
w4046 <= not w2525 and w2647;
w4047 <= not w4045 and not w4046;
w4048 <= not w4044 and w4047;
w4049 <= not w2640 and w4048;
w4050 <= not w2992 and w4048;
w4051 <= not w4049 and not w4050;
w4052 <= w619 and not w4051;
w4053 <= not w619 and w4051;
w4054 <= not w4052 and not w4053;
w4055 <= not w4043 and w4054;
w4056 <= not w4043 and not w4055;
w4057 <= w4054 and not w4055;
w4058 <= not w4056 and not w4057;
w4059 <= not w4025 and not w4058;
w4060 <= not w4025 and not w4059;
w4061 <= not w4058 and not w4059;
w4062 <= not w4060 and not w4061;
w4063 <= not w4024 and not w4062;
w4064 <= not w4024 and not w4063;
w4065 <= not w4062 and not w4063;
w4066 <= not w4064 and not w4065;
w4067 <= not w3915 and not w3921;
w4068 <= w4066 and w4067;
w4069 <= not w4066 and not w4067;
w4070 <= not w4068 and not w4069;
w4071 <= w245 and not w3578;
w4072 <= w2510 and not w3230;
w4073 <= w2517 and w3222;
w4074 <= not w4072 and not w4073;
w4075 <= not w4071 and w4074;
w4076 <= not w2521 and w4075;
w4077 <= not w3591 and w4075;
w4078 <= not w4076 and not w4077;
w4079 <= w225 and not w4078;
w4080 <= not w225 and w4078;
w4081 <= not w4079 and not w4080;
w4082 <= w4070 and w4081;
w4083 <= w4070 and not w4082;
w4084 <= w4081 and not w4082;
w4085 <= not w4083 and not w4084;
w4086 <= not w4013 and not w4085;
w4087 <= not w4013 and not w4086;
w4088 <= not w4085 and not w4086;
w4089 <= not w4087 and not w4088;
w4090 <= not w4012 and not w4089;
w4091 <= not w4012 and not w4090;
w4092 <= not w4089 and not w4090;
w4093 <= not w4091 and not w4092;
w4094 <= not w3999 and w4093;
w4095 <= w3999 and not w4093;
w4096 <= not w4094 and not w4095;
w4097 <= not w3998 and not w4096;
w4098 <= w3998 and w4096;
w4099 <= not w3982 and not w4098;
w4100 <= not w4097 and w4099;
w4101 <= not w3982 and not w4100;
w4102 <= not w4097 and not w4100;
w4103 <= not w4098 and w4102;
w4104 <= not w4101 and not w4103;
w4105 <= not w3972 and w4104;
w4106 <= w3972 and not w4104;
w4107 <= not w4105 and not w4106;
w4108 <= w3824 and not w3974;
w4109 <= not w3977 and not w4108;
w4110 <= not w4107 and w4109;
w4111 <= w4107 and not w4109;
w4112 <= not w4110 and not w4111;
w4113 <= w2290 and w3607;
w4114 <= w347 and w4113;
w4115 <= w896 and w4114;
w4116 <= w2146 and w4115;
w4117 <= w1418 and w4116;
w4118 <= w685 and w4117;
w4119 <= w305 and w4118;
w4120 <= not w267 and w4119;
w4121 <= not w125 and w4120;
w4122 <= not w320 and w4121;
w4123 <= not w61 and w4122;
w4124 <= not w208 and w4123;
w4125 <= not w188 and w4124;
w4126 <= not w3999 and not w4093;
w4127 <= not w4090 and not w4126;
w4128 <= not w4082 and not w4086;
w4129 <= w3224 and w3846;
w4130 <= w3166 and w4004;
w4131 <= not w4129 and not w4130;
w4132 <= not w241 and not w4131;
w4133 <= not w4131 and not w4132;
w4134 <= not w241 and not w4132;
w4135 <= not w4133 and not w4134;
w4136 <= w2752 and not w3230;
w4137 <= not w2504 and w2758;
w4138 <= w2760 and w3227;
w4139 <= not w4137 and not w4138;
w4140 <= not w4136 and w4139;
w4141 <= w2767 and w3268;
w4142 <= w4140 and not w4141;
w4143 <= not w971 and not w4142;
w4144 <= not w4142 and not w4143;
w4145 <= not w971 and not w4143;
w4146 <= not w4144 and not w4145;
w4147 <= not w4055 and not w4059;
w4148 <= not w475 and w4035;
w4149 <= w2543 and w4148;
w4150 <= not w4040 and not w4149;
w4151 <= w2528 and w2618;
w4152 <= not w2536 and w2726;
w4153 <= not w2532 and w2616;
w4154 <= not w4152 and not w4153;
w4155 <= not w4151 and w4154;
w4156 <= w2624 and w2765;
w4157 <= w4155 and not w4156;
w4158 <= not w475 and w2540;
w4159 <= not w4157 and w4158;
w4160 <= w4157 and not w4158;
w4161 <= not w4159 and not w4160;
w4162 <= not w4150 and w4161;
w4163 <= not w4150 and not w4162;
w4164 <= w4161 and not w4162;
w4165 <= not w4163 and not w4164;
w4166 <= not w2516 and w2649;
w4167 <= not w2525 and w2645;
w4168 <= w2512 and w2647;
w4169 <= not w4167 and not w4168;
w4170 <= not w4166 and w4169;
w4171 <= not w2640 and w4170;
w4172 <= not w2972 and w4170;
w4173 <= not w4171 and not w4172;
w4174 <= w619 and not w4173;
w4175 <= not w619 and w4173;
w4176 <= not w4174 and not w4175;
w4177 <= not w4165 and w4176;
w4178 <= w4165 and not w4176;
w4179 <= not w4177 and not w4178;
w4180 <= not w4147 and w4179;
w4181 <= w4147 and not w4179;
w4182 <= not w4180 and not w4181;
w4183 <= not w4146 and w4182;
w4184 <= not w4146 and not w4183;
w4185 <= w4182 and not w4183;
w4186 <= not w4184 and not w4185;
w4187 <= not w4063 and not w4069;
w4188 <= w4186 and w4187;
w4189 <= not w4186 and not w4187;
w4190 <= not w4188 and not w4189;
w4191 <= w245 and w3700;
w4192 <= w2510 and w3222;
w4193 <= w2517 and not w3578;
w4194 <= not w4192 and not w4193;
w4195 <= not w4191 and w4194;
w4196 <= not w2521 and w4195;
w4197 <= not w3712 and w4195;
w4198 <= not w4196 and not w4197;
w4199 <= w225 and not w4198;
w4200 <= not w225 and w4198;
w4201 <= not w4199 and not w4200;
w4202 <= w4190 and w4201;
w4203 <= not w4190 and not w4201;
w4204 <= not w4202 and not w4203;
w4205 <= not w4135 and w4204;
w4206 <= w4135 and not w4204;
w4207 <= not w4205 and not w4206;
w4208 <= not w4128 and w4207;
w4209 <= w4128 and not w4207;
w4210 <= not w4208 and not w4209;
w4211 <= not w4127 and w4210;
w4212 <= w4127 and not w4210;
w4213 <= not w4211 and not w4212;
w4214 <= not w4125 and w4213;
w4215 <= not w4125 and not w4214;
w4216 <= w4213 and not w4214;
w4217 <= not w4215 and not w4216;
w4218 <= not w4102 and not w4217;
w4219 <= w4102 and not w4216;
w4220 <= not w4215 and w4219;
w4221 <= not w4218 and not w4220;
w4222 <= w4106 and w4221;
w4223 <= w4221 and not w4222;
w4224 <= w4106 and not w4222;
w4225 <= not w4223 and not w4224;
w4226 <= not w4107 and w4108;
w4227 <= not w3977 and not w4226;
w4228 <= not w4225 and w4227;
w4229 <= w4225 and not w4227;
w4230 <= not w4228 and not w4229;
w4231 <= not w4214 and not w4218;
w4232 <= w296 and w446;
w4233 <= w251 and w4232;
w4234 <= w2414 and w4233;
w4235 <= w925 and w4234;
w4236 <= w702 and w4235;
w4237 <= w594 and w4236;
w4238 <= w2368 and w4237;
w4239 <= not w128 and w4238;
w4240 <= not w144 and w4239;
w4241 <= not w539 and w4240;
w4242 <= not w4208 and not w4211;
w4243 <= not w4202 and not w4205;
w4244 <= not w4183 and not w4189;
w4245 <= not w4177 and not w4180;
w4246 <= not w2525 and w2618;
w4247 <= not w2532 and w2726;
w4248 <= w2528 and w2616;
w4249 <= not w4247 and not w4248;
w4250 <= not w4246 and w4249;
w4251 <= w2624 and w2939;
w4252 <= w4250 and not w4251;
w4253 <= not w475 and not w4252;
w4254 <= not w4252 and not w4253;
w4255 <= not w475 and not w4253;
w4256 <= not w4254 and not w4255;
w4257 <= not w241 and not w475;
w4258 <= not w2536 and w4257;
w4259 <= not w241 and not w4258;
w4260 <= not w2536 and not w4258;
w4261 <= not w475 and w4260;
w4262 <= not w4259 and not w4261;
w4263 <= not w4256 and not w4262;
w4264 <= not w4256 and not w4263;
w4265 <= not w4262 and not w4263;
w4266 <= not w4264 and not w4265;
w4267 <= not w475 and not w2540;
w4268 <= w4157 and w4267;
w4269 <= not w4162 and not w4268;
w4270 <= w4266 and not w4269;
w4271 <= not w4266 and w4269;
w4272 <= not w4270 and not w4271;
w4273 <= not w2504 and w2649;
w4274 <= w2512 and w2645;
w4275 <= not w2516 and w2647;
w4276 <= not w4274 and not w4275;
w4277 <= not w4273 and w4276;
w4278 <= w2602 and w2640;
w4279 <= w4277 and not w4278;
w4280 <= not w619 and not w4279;
w4281 <= w619 and w4279;
w4282 <= not w4280 and not w4281;
w4283 <= not w4272 and w4282;
w4284 <= not w4272 and not w4283;
w4285 <= w4282 and not w4283;
w4286 <= not w4284 and not w4285;
w4287 <= not w4245 and w4286;
w4288 <= w4245 and not w4286;
w4289 <= not w4287 and not w4288;
w4290 <= w2752 and w3222;
w4291 <= w2758 and w3227;
w4292 <= w2760 and not w3230;
w4293 <= not w4291 and not w4292;
w4294 <= not w4290 and w4293;
w4295 <= w2767 and w3252;
w4296 <= w4294 and not w4295;
w4297 <= not w971 and not w4296;
w4298 <= not w971 and not w4297;
w4299 <= not w4296 and not w4297;
w4300 <= not w4298 and not w4299;
w4301 <= not w4289 and not w4300;
w4302 <= w4289 and w4300;
w4303 <= not w4301 and not w4302;
w4304 <= not w4244 and w4303;
w4305 <= w4244 and not w4303;
w4306 <= not w4304 and not w4305;
w4307 <= w245 and w3846;
w4308 <= w2510 and not w3578;
w4309 <= w2517 and w3700;
w4310 <= not w4308 and not w4309;
w4311 <= not w4307 and w4310;
w4312 <= w2521 and w3858;
w4313 <= w4311 and not w4312;
w4314 <= not w225 and not w4313;
w4315 <= w225 and w4313;
w4316 <= not w4314 and not w4315;
w4317 <= w4306 and w4316;
w4318 <= not w4306 and not w4316;
w4319 <= not w4317 and not w4318;
w4320 <= not w4243 and w4319;
w4321 <= w4243 and not w4319;
w4322 <= not w4320 and not w4321;
w4323 <= w4242 and not w4322;
w4324 <= not w4242 and w4322;
w4325 <= not w4323 and not w4324;
w4326 <= w4241 and not w4325;
w4327 <= not w4241 and w4325;
w4328 <= not w4326 and not w4327;
w4329 <= not w4231 and w4328;
w4330 <= w4231 and not w4328;
w4331 <= not w4329 and not w4330;
w4332 <= not w4222 and not w4331;
w4333 <= w4222 and w4331;
w4334 <= not w4332 and not w4333;
w4335 <= w4225 and w4226;
w4336 <= not w3977 and not w4335;
w4337 <= not w4334 and w4336;
w4338 <= w4334 and not w4336;
w4339 <= not w4337 and not w4338;
w4340 <= not w4327 and not w4329;
w4341 <= not w267 and not w309;
w4342 <= not w422 and w4341;
w4343 <= w139 and w757;
w4344 <= w4342 and w4343;
w4345 <= w2267 and w4344;
w4346 <= w264 and w4345;
w4347 <= w3833 and w4346;
w4348 <= w3193 and w4347;
w4349 <= w3952 and w4348;
w4350 <= w319 and w4349;
w4351 <= not w128 and w4350;
w4352 <= not w367 and w4351;
w4353 <= not w249 and w4352;
w4354 <= not w187 and w4353;
w4355 <= not w4320 and not w4324;
w4356 <= not w4304 and not w4317;
w4357 <= not w4245 and not w4286;
w4358 <= not w4301 and not w4357;
w4359 <= w2752 and not w3578;
w4360 <= w2758 and not w3230;
w4361 <= w2760 and w3222;
w4362 <= not w4360 and not w4361;
w4363 <= not w4359 and w4362;
w4364 <= w2767 and w3591;
w4365 <= w4363 and not w4364;
w4366 <= not w971 and not w4365;
w4367 <= not w4365 and not w4366;
w4368 <= not w971 and not w4366;
w4369 <= not w4367 and not w4368;
w4370 <= not w4266 and not w4269;
w4371 <= not w4283 and not w4370;
w4372 <= not w4258 and not w4263;
w4373 <= not w2532 and w4257;
w4374 <= not w241 and not w4373;
w4375 <= not w2532 and not w4373;
w4376 <= not w475 and w4375;
w4377 <= not w4374 and not w4376;
w4378 <= not w4372 and not w4377;
w4379 <= not w4372 and not w4378;
w4380 <= not w4377 and not w4378;
w4381 <= not w4379 and not w4380;
w4382 <= w2512 and w2618;
w4383 <= w2528 and w2726;
w4384 <= not w2525 and w2616;
w4385 <= not w4383 and not w4384;
w4386 <= not w4382 and w4385;
w4387 <= not w2624 and w4386;
w4388 <= not w2992 and w4386;
w4389 <= not w4387 and not w4388;
w4390 <= w475 and not w4389;
w4391 <= not w475 and w4389;
w4392 <= not w4390 and not w4391;
w4393 <= not w4381 and w4392;
w4394 <= not w4381 and not w4393;
w4395 <= w4392 and not w4393;
w4396 <= not w4394 and not w4395;
w4397 <= w2649 and w3227;
w4398 <= not w2516 and w2645;
w4399 <= not w2504 and w2647;
w4400 <= not w4398 and not w4399;
w4401 <= not w4397 and w4400;
w4402 <= w2640 and w3282;
w4403 <= w4401 and not w4402;
w4404 <= not w619 and not w4403;
w4405 <= w619 and w4403;
w4406 <= not w4404 and not w4405;
w4407 <= not w4396 and w4406;
w4408 <= not w4395 and not w4406;
w4409 <= not w4394 and w4408;
w4410 <= not w4407 and not w4409;
w4411 <= not w4371 and w4410;
w4412 <= not w4371 and not w4411;
w4413 <= w4410 and not w4411;
w4414 <= not w4412 and not w4413;
w4415 <= not w4369 and not w4414;
w4416 <= w4369 and not w4413;
w4417 <= not w4412 and w4416;
w4418 <= not w4415 and not w4417;
w4419 <= not w4358 and w4418;
w4420 <= not w4358 and not w4419;
w4421 <= w4418 and not w4419;
w4422 <= not w4420 and not w4421;
w4423 <= w2510 and w3700;
w4424 <= w2517 and w3846;
w4425 <= not w4423 and not w4424;
w4426 <= w2521 and w4006;
w4427 <= w4425 and not w4426;
w4428 <= not w225 and not w4427;
w4429 <= w225 and w4427;
w4430 <= not w4428 and not w4429;
w4431 <= not w4422 and w4430;
w4432 <= not w4421 and not w4430;
w4433 <= not w4420 and w4432;
w4434 <= not w4431 and not w4433;
w4435 <= not w4356 and w4434;
w4436 <= w4356 and not w4434;
w4437 <= not w4435 and not w4436;
w4438 <= not w4355 and w4437;
w4439 <= w4355 and not w4437;
w4440 <= not w4438 and not w4439;
w4441 <= w4354 and not w4440;
w4442 <= not w4354 and w4440;
w4443 <= not w4441 and not w4442;
w4444 <= not w4340 and w4443;
w4445 <= w4340 and not w4443;
w4446 <= not w4444 and not w4445;
w4447 <= not w4333 and not w4446;
w4448 <= w4333 and w4446;
w4449 <= not w4447 and not w4448;
w4450 <= not w4334 and w4335;
w4451 <= not w3977 and not w4450;
w4452 <= not w4449 and w4451;
w4453 <= w4449 and not w4451;
w4454 <= not w4452 and not w4453;
w4455 <= not w4442 and not w4444;
w4456 <= w266 and w1067;
w4457 <= w536 and w4456;
w4458 <= w2371 and w4457;
w4459 <= w2290 and w4458;
w4460 <= w106 and w4459;
w4461 <= w319 and w4460;
w4462 <= w926 and w4461;
w4463 <= not w307 and w4462;
w4464 <= w203 and w920;
w4465 <= w2408 and w4464;
w4466 <= w3209 and w4465;
w4467 <= w4463 and w4466;
w4468 <= not w287 and w4467;
w4469 <= not w100 and w4468;
w4470 <= not w122 and w4469;
w4471 <= not w119 and w4470;
w4472 <= not w397 and w4471;
w4473 <= not w98 and w4472;
w4474 <= not w4435 and not w4438;
w4475 <= not w4419 and not w4431;
w4476 <= not w4411 and not w4415;
w4477 <= w2510 and w3846;
w4478 <= w2521 and w4004;
w4479 <= not w4477 and not w4478;
w4480 <= w225 and not w4479;
w4481 <= not w225 and w4479;
w4482 <= not w4480 and not w4481;
w4483 <= not w4476 and not w4482;
w4484 <= w4476 and w4482;
w4485 <= not w4483 and not w4484;
w4486 <= w2752 and w3700;
w4487 <= w2758 and w3222;
w4488 <= w2760 and not w3578;
w4489 <= not w4487 and not w4488;
w4490 <= not w4486 and w4489;
w4491 <= w2767 and w3712;
w4492 <= w4490 and not w4491;
w4493 <= not w971 and not w4492;
w4494 <= not w4492 and not w4493;
w4495 <= not w971 and not w4493;
w4496 <= not w4494 and not w4495;
w4497 <= not w4393 and not w4407;
w4498 <= not w4373 and not w4378;
w4499 <= w2528 and w4257;
w4500 <= not w241 and not w4499;
w4501 <= w2528 and not w4499;
w4502 <= not w475 and w4501;
w4503 <= not w4500 and not w4502;
w4504 <= not w4498 and not w4503;
w4505 <= not w4498 and not w4504;
w4506 <= not w4503 and not w4504;
w4507 <= not w4505 and not w4506;
w4508 <= not w2516 and w2618;
w4509 <= not w2525 and w2726;
w4510 <= w2512 and w2616;
w4511 <= not w4509 and not w4510;
w4512 <= not w4508 and w4511;
w4513 <= not w2624 and w4512;
w4514 <= not w2972 and w4512;
w4515 <= not w4513 and not w4514;
w4516 <= w475 and not w4515;
w4517 <= not w475 and w4515;
w4518 <= not w4516 and not w4517;
w4519 <= not w4507 and w4518;
w4520 <= not w4507 and not w4519;
w4521 <= w4518 and not w4519;
w4522 <= not w4520 and not w4521;
w4523 <= w2649 and not w3230;
w4524 <= not w2504 and w2645;
w4525 <= w2647 and w3227;
w4526 <= not w4524 and not w4525;
w4527 <= not w4523 and w4526;
w4528 <= w2640 and w3268;
w4529 <= w4527 and not w4528;
w4530 <= not w619 and not w4529;
w4531 <= w619 and w4529;
w4532 <= not w4530 and not w4531;
w4533 <= not w4522 and w4532;
w4534 <= not w4521 and not w4532;
w4535 <= not w4520 and w4534;
w4536 <= not w4533 and not w4535;
w4537 <= not w4497 and w4536;
w4538 <= not w4497 and not w4537;
w4539 <= w4536 and not w4537;
w4540 <= not w4538 and not w4539;
w4541 <= not w4496 and not w4540;
w4542 <= w4496 and not w4539;
w4543 <= not w4538 and w4542;
w4544 <= not w4541 and not w4543;
w4545 <= w4485 and w4544;
w4546 <= not w4485 and not w4544;
w4547 <= not w4545 and not w4546;
w4548 <= not w4475 and w4547;
w4549 <= w4475 and not w4547;
w4550 <= not w4548 and not w4549;
w4551 <= not w4474 and w4550;
w4552 <= w4474 and not w4550;
w4553 <= not w4551 and not w4552;
w4554 <= w4473 and not w4553;
w4555 <= not w4473 and w4553;
w4556 <= not w4554 and not w4555;
w4557 <= not w4455 and w4556;
w4558 <= w4455 and not w4556;
w4559 <= not w4557 and not w4558;
w4560 <= not w4448 and not w4559;
w4561 <= w4448 and w4559;
w4562 <= not w4560 and not w4561;
w4563 <= not w4449 and w4450;
w4564 <= not w3977 and not w4563;
w4565 <= not w4562 and w4564;
w4566 <= w4562 and not w4564;
w4567 <= not w4565 and not w4566;
w4568 <= not w4555 and not w4557;
w4569 <= not w4483 and not w4545;
w4570 <= not w4537 and not w4541;
w4571 <= w2752 and w3846;
w4572 <= w2758 and not w3578;
w4573 <= w2760 and w3700;
w4574 <= not w4572 and not w4573;
w4575 <= not w4571 and w4574;
w4576 <= not w3858 and w4575;
w4577 <= not w2767 and w4575;
w4578 <= not w4576 and not w4577;
w4579 <= w971 and not w4578;
w4580 <= not w971 and w4578;
w4581 <= not w4579 and not w4580;
w4582 <= not w4570 and w4581;
w4583 <= w4570 and not w4581;
w4584 <= not w4582 and not w4583;
w4585 <= not w4519 and not w4533;
w4586 <= not w4499 and not w4504;
w4587 <= not w2504 and w2618;
w4588 <= w2512 and w2726;
w4589 <= not w2516 and w2616;
w4590 <= not w4588 and not w4589;
w4591 <= not w4587 and w4590;
w4592 <= w2602 and w2624;
w4593 <= w4591 and not w4592;
w4594 <= not w475 and not w4593;
w4595 <= not w4593 and not w4594;
w4596 <= not w475 and not w4594;
w4597 <= not w4595 and not w4596;
w4598 <= not w475 and not w2525;
w4599 <= w225 and w241;
w4600 <= not w225 and not w241;
w4601 <= not w4599 and not w4600;
w4602 <= w4598 and w4601;
w4603 <= not w4598 and not w4601;
w4604 <= not w4602 and not w4603;
w4605 <= not w4597 and w4604;
w4606 <= not w4597 and not w4605;
w4607 <= w4604 and not w4605;
w4608 <= not w4606 and not w4607;
w4609 <= not w4586 and w4608;
w4610 <= w4586 and not w4608;
w4611 <= not w4609 and not w4610;
w4612 <= w2649 and w3222;
w4613 <= w2645 and w3227;
w4614 <= w2647 and not w3230;
w4615 <= not w4613 and not w4614;
w4616 <= not w4612 and w4615;
w4617 <= not w2640 and w4616;
w4618 <= not w3252 and w4616;
w4619 <= not w4617 and not w4618;
w4620 <= w619 and not w4619;
w4621 <= not w619 and w4619;
w4622 <= not w4620 and not w4621;
w4623 <= not w4611 and w4622;
w4624 <= not w4611 and not w4623;
w4625 <= w4622 and not w4623;
w4626 <= not w4624 and not w4625;
w4627 <= not w4585 and not w4626;
w4628 <= not w4585 and not w4627;
w4629 <= not w4626 and not w4627;
w4630 <= not w4628 and not w4629;
w4631 <= w4584 and not w4630;
w4632 <= w4584 and not w4631;
w4633 <= not w4630 and not w4631;
w4634 <= not w4632 and not w4633;
w4635 <= not w4569 and w4634;
w4636 <= w4569 and not w4634;
w4637 <= not w4635 and not w4636;
w4638 <= not w4548 and not w4551;
w4639 <= w4637 and w4638;
w4640 <= not w4637 and not w4638;
w4641 <= not w4639 and not w4640;
w4642 <= w881 and w2231;
w4643 <= w4342 and w4642;
w4644 <= w759 and w4643;
w4645 <= w4463 and w4644;
w4646 <= not w79 and w4645;
w4647 <= not w144 and w4646;
w4648 <= not w87 and w4647;
w4649 <= not w168 and w4648;
w4650 <= w1040 and w4649;
w4651 <= not w118 and w4650;
w4652 <= not w395 and w4651;
w4653 <= w4641 and not w4652;
w4654 <= not w4641 and w4652;
w4655 <= not w4653 and not w4654;
w4656 <= not w4568 and w4655;
w4657 <= w4568 and not w4655;
w4658 <= not w4656 and not w4657;
w4659 <= w4561 and w4658;
w4660 <= not w4561 and not w4658;
w4661 <= not w4659 and not w4660;
w4662 <= not w4562 and w4563;
w4663 <= not w3977 and not w4662;
w4664 <= not w4661 and w4663;
w4665 <= w4661 and not w4663;
w4666 <= not w4664 and not w4665;
w4667 <= not w4653 and not w4656;
w4668 <= w559 and w2131;
w4669 <= w115 and w4668;
w4670 <= not w171 and w4669;
w4671 <= not w169 and w4670;
w4672 <= not w117 and w4671;
w4673 <= not w175 and w4672;
w4674 <= not w396 and w4673;
w4675 <= not w61 and w4674;
w4676 <= not w161 and w4675;
w4677 <= w911 and w2292;
w4678 <= w929 and w4677;
w4679 <= w3628 and w4678;
w4680 <= w4676 and w4679;
w4681 <= not w358 and w4680;
w4682 <= not w207 and w4681;
w4683 <= not w157 and w4682;
w4684 <= not w311 and w4683;
w4685 <= not w174 and w4684;
w4686 <= not w276 and w4685;
w4687 <= not w419 and w4686;
w4688 <= not w4569 and not w4634;
w4689 <= not w4640 and not w4688;
w4690 <= not w4582 and not w4631;
w4691 <= w2758 and w3700;
w4692 <= w2760 and w3846;
w4693 <= not w4691 and not w4692;
w4694 <= w2767 and w4006;
w4695 <= w4693 and not w4694;
w4696 <= not w971 and not w4695;
w4697 <= not w4695 and not w4696;
w4698 <= not w971 and not w4696;
w4699 <= not w4697 and not w4698;
w4700 <= not w4623 and not w4627;
w4701 <= not w4586 and not w4608;
w4702 <= not w4605 and not w4701;
w4703 <= not w475 and w2512;
w4704 <= not w4599 and not w4602;
w4705 <= not w4703 and not w4704;
w4706 <= not w4703 and not w4705;
w4707 <= not w4704 and not w4705;
w4708 <= not w4706 and not w4707;
w4709 <= w2618 and w3227;
w4710 <= not w2516 and w2726;
w4711 <= not w2504 and w2616;
w4712 <= not w4710 and not w4711;
w4713 <= not w4709 and w4712;
w4714 <= not w2624 and w4713;
w4715 <= not w3282 and w4713;
w4716 <= not w4714 and not w4715;
w4717 <= w475 and not w4716;
w4718 <= not w475 and w4716;
w4719 <= not w4717 and not w4718;
w4720 <= not w4708 and w4719;
w4721 <= w4708 and not w4719;
w4722 <= not w4720 and not w4721;
w4723 <= not w4702 and w4722;
w4724 <= not w4702 and not w4723;
w4725 <= w4722 and not w4723;
w4726 <= not w4724 and not w4725;
w4727 <= w2649 and not w3578;
w4728 <= w2645 and not w3230;
w4729 <= w2647 and w3222;
w4730 <= not w4728 and not w4729;
w4731 <= not w4727 and w4730;
w4732 <= w2640 and w3591;
w4733 <= w4731 and not w4732;
w4734 <= not w619 and not w4733;
w4735 <= w619 and w4733;
w4736 <= not w4734 and not w4735;
w4737 <= not w4726 and w4736;
w4738 <= not w4725 and not w4736;
w4739 <= not w4724 and w4738;
w4740 <= not w4737 and not w4739;
w4741 <= not w4700 and w4740;
w4742 <= w4700 and not w4740;
w4743 <= not w4741 and not w4742;
w4744 <= not w4699 and w4743;
w4745 <= w4699 and not w4743;
w4746 <= not w4744 and not w4745;
w4747 <= not w4690 and w4746;
w4748 <= w4690 and not w4746;
w4749 <= not w4747 and not w4748;
w4750 <= not w4689 and w4749;
w4751 <= w4689 and not w4749;
w4752 <= not w4750 and not w4751;
w4753 <= w4687 and not w4752;
w4754 <= not w4687 and w4752;
w4755 <= not w4753 and not w4754;
w4756 <= not w4667 and w4755;
w4757 <= w4667 and not w4755;
w4758 <= not w4756 and not w4757;
w4759 <= not w4659 and not w4758;
w4760 <= w4659 and w4758;
w4761 <= not w4759 and not w4760;
w4762 <= not w4661 and w4662;
w4763 <= not w3977 and not w4762;
w4764 <= not w4761 and w4763;
w4765 <= w4761 and not w4763;
w4766 <= not w4764 and not w4765;
w4767 <= not w4754 and not w4756;
w4768 <= w707 and w759;
w4769 <= w154 and w4768;
w4770 <= w3181 and w4769;
w4771 <= w2382 and w4770;
w4772 <= w3209 and w4771;
w4773 <= not w287 and w4772;
w4774 <= not w277 and w4773;
w4775 <= not w175 and w4774;
w4776 <= not w83 and w4775;
w4777 <= not w184 and w4776;
w4778 <= not w306 and w4777;
w4779 <= not w166 and w4778;
w4780 <= not w4741 and not w4744;
w4781 <= not w4705 and not w4720;
w4782 <= w2618 and not w3230;
w4783 <= not w2504 and w2726;
w4784 <= w2616 and w3227;
w4785 <= not w4783 and not w4784;
w4786 <= not w4782 and w4785;
w4787 <= w2624 and w3268;
w4788 <= w4786 and not w4787;
w4789 <= not w475 and not w4788;
w4790 <= not w4788 and not w4789;
w4791 <= not w475 and not w4789;
w4792 <= not w4790 and not w4791;
w4793 <= not w475 and w2594;
w4794 <= not w4792 and not w4793;
w4795 <= not w4792 and not w4794;
w4796 <= not w4793 and not w4794;
w4797 <= not w4795 and not w4796;
w4798 <= not w4781 and w4797;
w4799 <= w4781 and not w4797;
w4800 <= not w4798 and not w4799;
w4801 <= w2649 and w3700;
w4802 <= w2645 and w3222;
w4803 <= w2647 and not w3578;
w4804 <= not w4802 and not w4803;
w4805 <= not w4801 and w4804;
w4806 <= w2640 and w3712;
w4807 <= w4805 and not w4806;
w4808 <= not w619 and not w4807;
w4809 <= w619 and w4807;
w4810 <= not w4808 and not w4809;
w4811 <= not w4800 and w4810;
w4812 <= not w4800 and not w4811;
w4813 <= w4810 and not w4811;
w4814 <= not w4812 and not w4813;
w4815 <= not w4723 and not w4737;
w4816 <= w2758 and w3846;
w4817 <= w2767 and w4004;
w4818 <= not w4816 and not w4817;
w4819 <= not w971 and w4818;
w4820 <= w971 and not w4818;
w4821 <= not w4819 and not w4820;
w4822 <= not w4815 and not w4821;
w4823 <= w4815 and w4821;
w4824 <= not w4822 and not w4823;
w4825 <= not w4814 and w4824;
w4826 <= not w4814 and not w4825;
w4827 <= w4824 and not w4825;
w4828 <= not w4826 and not w4827;
w4829 <= not w4780 and w4828;
w4830 <= w4780 and not w4828;
w4831 <= not w4829 and not w4830;
w4832 <= not w4747 and not w4750;
w4833 <= w4831 and w4832;
w4834 <= not w4831 and not w4832;
w4835 <= not w4833 and not w4834;
w4836 <= w4779 and not w4835;
w4837 <= not w4779 and w4835;
w4838 <= not w4836 and not w4837;
w4839 <= not w4767 and w4838;
w4840 <= w4767 and not w4838;
w4841 <= not w4839 and not w4840;
w4842 <= not w4760 and not w4841;
w4843 <= w4760 and w4841;
w4844 <= not w4842 and not w4843;
w4845 <= not w4761 and w4762;
w4846 <= not w3977 and not w4845;
w4847 <= not w4844 and w4846;
w4848 <= w4844 and not w4846;
w4849 <= not w4847 and not w4848;
w4850 <= not w4837 and not w4839;
w4851 <= w209 and w605;
w4852 <= w426 and w4851;
w4853 <= w455 and w4852;
w4854 <= w160 and w4853;
w4855 <= w3616 and w4854;
w4856 <= w1054 and w4855;
w4857 <= w3209 and w4856;
w4858 <= w927 and w4857;
w4859 <= not w262 and w4858;
w4860 <= not w142 and w4859;
w4861 <= not w265 and w4860;
w4862 <= not w4780 and not w4828;
w4863 <= not w4834 and not w4862;
w4864 <= not w4822 and not w4825;
w4865 <= not w2516 and not w4703;
w4866 <= not w475 and w4865;
w4867 <= not w4794 and not w4866;
w4868 <= not w475 and not w2504;
w4869 <= not w971 and not w4868;
w4870 <= w971 and w4868;
w4871 <= w4703 and not w4870;
w4872 <= not w4869 and w4871;
w4873 <= w4703 and not w4872;
w4874 <= not w4870 and not w4872;
w4875 <= not w4869 and w4874;
w4876 <= not w4873 and not w4875;
w4877 <= not w4867 and not w4876;
w4878 <= not w4867 and not w4877;
w4879 <= not w4876 and not w4877;
w4880 <= not w4878 and not w4879;
w4881 <= w2618 and w3222;
w4882 <= w2726 and w3227;
w4883 <= w2616 and not w3230;
w4884 <= not w4882 and not w4883;
w4885 <= not w4881 and w4884;
w4886 <= w2624 and w3252;
w4887 <= w4885 and not w4886;
w4888 <= not w475 and not w4887;
w4889 <= not w475 and not w4888;
w4890 <= not w4887 and not w4888;
w4891 <= not w4889 and not w4890;
w4892 <= not w4880 and not w4891;
w4893 <= not w4880 and not w4892;
w4894 <= not w4891 and not w4892;
w4895 <= not w4893 and not w4894;
w4896 <= not w4781 and not w4797;
w4897 <= not w4811 and not w4896;
w4898 <= w2649 and w3846;
w4899 <= w2645 and not w3578;
w4900 <= w2647 and w3700;
w4901 <= not w4899 and not w4900;
w4902 <= not w4898 and w4901;
w4903 <= not w2640 and w4902;
w4904 <= not w3858 and w4902;
w4905 <= not w4903 and not w4904;
w4906 <= w619 and not w4905;
w4907 <= not w619 and w4905;
w4908 <= not w4906 and not w4907;
w4909 <= not w4897 and w4908;
w4910 <= not w4897 and not w4909;
w4911 <= w4908 and not w4909;
w4912 <= not w4910 and not w4911;
w4913 <= not w4895 and not w4912;
w4914 <= w4895 and not w4911;
w4915 <= not w4910 and w4914;
w4916 <= not w4913 and not w4915;
w4917 <= not w4864 and w4916;
w4918 <= w4864 and not w4916;
w4919 <= not w4917 and not w4918;
w4920 <= not w4863 and w4919;
w4921 <= w4863 and not w4919;
w4922 <= not w4920 and not w4921;
w4923 <= w4861 and not w4922;
w4924 <= not w4861 and w4922;
w4925 <= not w4923 and not w4924;
w4926 <= not w4850 and w4925;
w4927 <= w4850 and not w4925;
w4928 <= not w4926 and not w4927;
w4929 <= not w4843 and not w4928;
w4930 <= w4843 and w4928;
w4931 <= not w4929 and not w4930;
w4932 <= not w4844 and w4845;
w4933 <= not w3977 and not w4932;
w4934 <= not w4931 and w4933;
w4935 <= w4931 and not w4933;
w4936 <= not w4934 and not w4935;
w4937 <= not w4924 and not w4926;
w4938 <= w861 and w919;
w4939 <= w449 and w4938;
w4940 <= w3684 and w4939;
w4941 <= w586 and w4940;
w4942 <= w403 and w4941;
w4943 <= not w286 and w4942;
w4944 <= not w4917 and not w4920;
w4945 <= not w4909 and not w4913;
w4946 <= not w4877 and not w4892;
w4947 <= not w475 and w3227;
w4948 <= not w4874 and w4947;
w4949 <= w4874 and not w4947;
w4950 <= not w4948 and not w4949;
w4951 <= w2618 and not w3578;
w4952 <= w2726 and not w3230;
w4953 <= w2616 and w3222;
w4954 <= not w4952 and not w4953;
w4955 <= not w4951 and w4954;
w4956 <= not w2624 and w4955;
w4957 <= not w3591 and w4955;
w4958 <= not w4956 and not w4957;
w4959 <= w475 and not w4958;
w4960 <= not w475 and w4958;
w4961 <= not w4959 and not w4960;
w4962 <= not w4950 and w4961;
w4963 <= w4950 and not w4961;
w4964 <= not w4962 and not w4963;
w4965 <= not w4946 and w4964;
w4966 <= not w4946 and not w4965;
w4967 <= w4964 and not w4965;
w4968 <= not w4966 and not w4967;
w4969 <= w2645 and w3700;
w4970 <= w2647 and w3846;
w4971 <= not w4969 and not w4970;
w4972 <= w2640 and w4006;
w4973 <= w4971 and not w4972;
w4974 <= not w619 and not w4973;
w4975 <= w619 and w4973;
w4976 <= not w4974 and not w4975;
w4977 <= not w4968 and w4976;
w4978 <= not w4967 and not w4976;
w4979 <= not w4966 and w4978;
w4980 <= not w4977 and not w4979;
w4981 <= not w4945 and w4980;
w4982 <= w4945 and not w4980;
w4983 <= not w4981 and not w4982;
w4984 <= not w4944 and w4983;
w4985 <= w4944 and not w4983;
w4986 <= not w4984 and not w4985;
w4987 <= w4943 and not w4986;
w4988 <= not w4943 and w4986;
w4989 <= not w4987 and not w4988;
w4990 <= not w4937 and w4989;
w4991 <= w4937 and not w4989;
w4992 <= not w4990 and not w4991;
w4993 <= not w4930 and not w4992;
w4994 <= w4930 and w4992;
w4995 <= not w4993 and not w4994;
w4996 <= not w4931 and w4932;
w4997 <= not w3977 and not w4996;
w4998 <= not w4995 and w4997;
w4999 <= w4995 and not w4997;
w5000 <= not w4998 and not w4999;
w5001 <= not w4988 and not w4990;
w5002 <= not w127 and not w136;
w5003 <= not w157 and w5002;
w5004 <= not w184 and w5003;
w5005 <= not w285 and w5004;
w5006 <= w2317 and w5005;
w5007 <= w896 and w5006;
w5008 <= w3987 and w5007;
w5009 <= w2200 and w5008;
w5010 <= w330 and w5009;
w5011 <= not w89 and w5010;
w5012 <= not w84 and w5011;
w5013 <= not w161 and w5012;
w5014 <= not w4981 and not w4984;
w5015 <= not w4965 and not w4977;
w5016 <= w2645 and w3846;
w5017 <= w2640 and w4004;
w5018 <= not w5016 and not w5017;
w5019 <= not w619 and not w5018;
w5020 <= w619 and w5018;
w5021 <= not w5019 and not w5020;
w5022 <= w2618 and w3700;
w5023 <= w2726 and w3222;
w5024 <= w2616 and not w3578;
w5025 <= not w5023 and not w5024;
w5026 <= not w5022 and w5025;
w5027 <= w2624 and w3712;
w5028 <= w5026 and not w5027;
w5029 <= not w475 and not w5028;
w5030 <= not w475 and not w5029;
w5031 <= not w5028 and not w5029;
w5032 <= not w5030 and not w5031;
w5033 <= w5021 and not w5032;
w5034 <= w5021 and not w5033;
w5035 <= not w5032 and not w5033;
w5036 <= not w5034 and not w5035;
w5037 <= not w4874 and not w4947;
w5038 <= not w4962 and not w5037;
w5039 <= not w475 and not w3230;
w5040 <= not w4947 and w5039;
w5041 <= w4947 and not w5039;
w5042 <= not w5038 and not w5041;
w5043 <= not w5040 and w5042;
w5044 <= not w5038 and not w5043;
w5045 <= not w5041 and not w5043;
w5046 <= not w5040 and w5045;
w5047 <= not w5044 and not w5046;
w5048 <= not w5036 and w5047;
w5049 <= w5036 and not w5047;
w5050 <= not w5048 and not w5049;
w5051 <= not w5015 and not w5050;
w5052 <= w5015 and w5050;
w5053 <= not w5051 and not w5052;
w5054 <= not w5014 and w5053;
w5055 <= w5014 and not w5053;
w5056 <= not w5054 and not w5055;
w5057 <= w5013 and not w5056;
w5058 <= not w5013 and w5056;
w5059 <= not w5057 and not w5058;
w5060 <= not w5001 and w5059;
w5061 <= w5001 and not w5059;
w5062 <= not w5060 and not w5061;
w5063 <= not w4994 and not w5062;
w5064 <= w4994 and w5062;
w5065 <= not w5063 and not w5064;
w5066 <= not w4995 and w4996;
w5067 <= not w3977 and not w5066;
w5068 <= not w5065 and w5067;
w5069 <= w5065 and not w5067;
w5070 <= not w5068 and not w5069;
w5071 <= not w5058 and not w5060;
w5072 <= not w144 and not w344;
w5073 <= not w205 and w5072;
w5074 <= not w310 and w5073;
w5075 <= not w68 and w5074;
w5076 <= w106 and w5075;
w5077 <= w3952 and w5076;
w5078 <= w261 and w5077;
w5079 <= w2128 and w5078;
w5080 <= w930 and w5079;
w5081 <= w3649 and w5080;
w5082 <= not w146 and w5081;
w5083 <= not w293 and w5082;
w5084 <= not w207 and w5083;
w5085 <= not w119 and w5084;
w5086 <= not w92 and w5085;
w5087 <= not w420 and w5086;
w5088 <= not w301 and w5087;
w5089 <= not w5051 and not w5054;
w5090 <= w2618 and w3846;
w5091 <= w2726 and not w3578;
w5092 <= w2616 and w3700;
w5093 <= not w5091 and not w5092;
w5094 <= not w5090 and w5093;
w5095 <= w2624 and w3858;
w5096 <= w5094 and not w5095;
w5097 <= not w475 and not w5096;
w5098 <= not w5096 and not w5097;
w5099 <= not w475 and not w5097;
w5100 <= not w5098 and not w5099;
w5101 <= w619 and w5039;
w5102 <= not w619 and not w5039;
w5103 <= not w5101 and not w5102;
w5104 <= not w475 and w3222;
w5105 <= w5103 and w5104;
w5106 <= not w5103 and not w5104;
w5107 <= not w5105 and not w5106;
w5108 <= not w5100 and w5107;
w5109 <= not w5100 and not w5108;
w5110 <= w5107 and not w5108;
w5111 <= not w5109 and not w5110;
w5112 <= not w5045 and w5111;
w5113 <= w5045 and not w5111;
w5114 <= not w5112 and not w5113;
w5115 <= not w5036 and not w5047;
w5116 <= not w5033 and not w5115;
w5117 <= not w5114 and not w5116;
w5118 <= w5114 and w5116;
w5119 <= not w5117 and not w5118;
w5120 <= not w5089 and w5119;
w5121 <= w5089 and not w5119;
w5122 <= not w5120 and not w5121;
w5123 <= not w5088 and w5122;
w5124 <= w5088 and not w5122;
w5125 <= not w5071 and not w5124;
w5126 <= not w5123 and w5125;
w5127 <= not w5071 and not w5126;
w5128 <= not w5123 and not w5126;
w5129 <= not w5124 and w5128;
w5130 <= not w5127 and not w5129;
w5131 <= not w5064 and w5130;
w5132 <= w5064 and not w5130;
w5133 <= not w5131 and not w5132;
w5134 <= not w5065 and w5066;
w5135 <= not w3977 and not w5134;
w5136 <= not w5133 and w5135;
w5137 <= w5133 and not w5135;
w5138 <= not w5136 and not w5137;
w5139 <= w2317 and w2383;
w5140 <= w423 and w5139;
w5141 <= w917 and w5140;
w5142 <= w2140 and w5141;
w5143 <= w1407 and w5142;
w5144 <= w933 and w5143;
w5145 <= w3209 and w5144;
w5146 <= not w88 and w5145;
w5147 <= not w126 and w5146;
w5148 <= not w77 and w5147;
w5149 <= not w293 and w5148;
w5150 <= not w320 and w5149;
w5151 <= not w286 and w5150;
w5152 <= not w456 and w5151;
w5153 <= not w5117 and not w5120;
w5154 <= not w5045 and not w5111;
w5155 <= not w5108 and not w5154;
w5156 <= not w475 and not w3578;
w5157 <= not w5101 and not w5105;
w5158 <= not w5156 and not w5157;
w5159 <= not w5156 and not w5158;
w5160 <= not w5157 and not w5158;
w5161 <= not w5159 and not w5160;
w5162 <= w2726 and w3700;
w5163 <= w2616 and w3846;
w5164 <= not w5162 and not w5163;
w5165 <= not w2624 and w5164;
w5166 <= not w4006 and w5164;
w5167 <= not w5165 and not w5166;
w5168 <= w475 and not w5167;
w5169 <= not w475 and w5167;
w5170 <= not w5168 and not w5169;
w5171 <= not w5161 and w5170;
w5172 <= w5161 and not w5170;
w5173 <= not w5171 and not w5172;
w5174 <= not w5155 and w5173;
w5175 <= w5155 and not w5173;
w5176 <= not w5174 and not w5175;
w5177 <= not w5153 and w5176;
w5178 <= w5153 and not w5176;
w5179 <= not w5177 and not w5178;
w5180 <= w5152 and not w5179;
w5181 <= not w5152 and w5179;
w5182 <= not w5180 and not w5181;
w5183 <= not w5128 and w5182;
w5184 <= w5128 and not w5182;
w5185 <= not w5183 and not w5184;
w5186 <= not w5132 and not w5185;
w5187 <= w5132 and w5185;
w5188 <= not w5186 and not w5187;
w5189 <= not w5133 and w5134;
w5190 <= not w3977 and not w5189;
w5191 <= not w5188 and w5190;
w5192 <= w5188 and not w5190;
w5193 <= not w5191 and not w5192;
w5194 <= not w5181 and not w5183;
w5195 <= not w287 and w1095;
w5196 <= not w278 and w5195;
w5197 <= not w204 and w5196;
w5198 <= w920 and w5197;
w5199 <= w294 and w5198;
w5200 <= w5005 and w5199;
w5201 <= w2325 and w5200;
w5202 <= w1065 and w5201;
w5203 <= not w77 and w5202;
w5204 <= not w176 and w5203;
w5205 <= not w167 and w5204;
w5206 <= not w306 and w5205;
w5207 <= not w456 and w5206;
w5208 <= not w686 and w5207;
w5209 <= w2726 and w3846;
w5210 <= w2624 and w4004;
w5211 <= not w5209 and not w5210;
w5212 <= not w475 and not w5211;
w5213 <= not w5211 and not w5212;
w5214 <= not w475 and not w5212;
w5215 <= not w5213 and not w5214;
w5216 <= not w475 and w3709;
w5217 <= not w5215 and not w5216;
w5218 <= not w5215 and not w5217;
w5219 <= not w5216 and not w5217;
w5220 <= not w5218 and not w5219;
w5221 <= not w5158 and not w5171;
w5222 <= w5220 and w5221;
w5223 <= not w5220 and not w5221;
w5224 <= not w5222 and not w5223;
w5225 <= not w5174 and not w5177;
w5226 <= not w5224 and w5225;
w5227 <= w5224 and not w5225;
w5228 <= not w5226 and not w5227;
w5229 <= not w5208 and w5228;
w5230 <= w5208 and not w5228;
w5231 <= not w5194 and not w5230;
w5232 <= not w5229 and w5231;
w5233 <= not w5194 and not w5232;
w5234 <= not w5229 and not w5232;
w5235 <= not w5230 and w5234;
w5236 <= not w5233 and not w5235;
w5237 <= not w5187 and w5236;
w5238 <= w5187 and not w5236;
w5239 <= not w5237 and not w5238;
w5240 <= not w5188 and w5189;
w5241 <= not w3977 and not w5240;
w5242 <= not w5239 and w5241;
w5243 <= w5239 and not w5241;
w5244 <= not w5242 and not w5243;
w5245 <= w588 and w2263;
w5246 <= w2202 and w5245;
w5247 <= w5075 and w5246;
w5248 <= w183 and w5247;
w5249 <= w425 and w5248;
w5250 <= w3652 and w5249;
w5251 <= not w158 and w5250;
w5252 <= not w397 and w5251;
w5253 <= not w427 and w5252;
w5254 <= not w5223 and not w5227;
w5255 <= w3700 and not w5156;
w5256 <= not w475 and w5255;
w5257 <= not w5217 and not w5256;
w5258 <= not w5254 and w5257;
w5259 <= w5254 and not w5257;
w5260 <= not w5258 and not w5259;
w5261 <= w3846 and not w5156;
w5262 <= not w3846 and w5156;
w5263 <= not w5261 and not w5262;
w5264 <= not w475 and w5263;
w5265 <= w5260 and not w5264;
w5266 <= not w5260 and w5264;
w5267 <= not w5265 and not w5266;
w5268 <= not w5253 and not w5267;
w5269 <= w5253 and w5267;
w5270 <= not w5234 and not w5269;
w5271 <= not w5268 and w5270;
w5272 <= not w5234 and not w5271;
w5273 <= not w5268 and not w5271;
w5274 <= not w5269 and w5273;
w5275 <= not w5272 and not w5274;
w5276 <= not w5238 and w5275;
w5277 <= w5238 and not w5275;
w5278 <= not w5276 and not w5277;
w5279 <= not w5239 and w5240;
w5280 <= not w3977 and not w5279;
w5281 <= not w5278 and w5280;
w5282 <= w5278 and not w5280;
w5283 <= not w5281 and not w5282;
w5284 <= w108 and w725;
w5285 <= w856 and w5284;
w5286 <= w209 and w5285;
w5287 <= w3193 and w5286;
w5288 <= w521 and w5287;
w5289 <= w930 and w5288;
w5290 <= not w89 and w5289;
w5291 <= not w157 and w5290;
w5292 <= not w247 and w5291;
w5293 <= not w318 and w5292;
w5294 <= not w165 and w5293;
w5295 <= not w5273 and not w5294;
w5296 <= w5273 and w5294;
w5297 <= not w5295 and not w5296;
w5298 <= not w5277 and w5297;
w5299 <= w5277 and not w5297;
w5300 <= not w5298 and not w5299;
w5301 <= not w5278 and w5279;
w5302 <= not w3977 and not w5301;
w5303 <= not w5300 and w5302;
w5304 <= w5300 and not w5302;
w5305 <= not w5303 and not w5304;
w5306 <= w5277 and w5297;
w5307 <= w538 and w2120;
w5308 <= w558 and w5307;
w5309 <= w1102 and w5308;
w5310 <= w1058 and w5309;
w5311 <= w936 and w5310;
w5312 <= w3625 and w5311;
w5313 <= not w126 and w5312;
w5314 <= not w177 and w5313;
w5315 <= not w157 and w5314;
w5316 <= not w307 and w5315;
w5317 <= not w188 and w5316;
w5318 <= w5295 and not w5317;
w5319 <= not w5295 and w5317;
w5320 <= not w5318 and not w5319;
w5321 <= not w5306 and not w5320;
w5322 <= w5306 and not w5319;
w5323 <= not w5321 and not w5322;
w5324 <= w5300 and w5301;
w5325 <= not w3977 and not w5324;
w5326 <= not w5323 and w5325;
w5327 <= w5323 and not w5325;
w5328 <= not w5326 and not w5327;
w5329 <= w4342 and w5197;
w5330 <= w323 and w5329;
w5331 <= w2490 and w5330;
w5332 <= w888 and w5331;
w5333 <= not w94 and w5332;
w5334 <= not w102 and w5333;
w5335 <= not w158 and w5334;
w5336 <= not w90 and w5335;
w5337 <= not w396 and w5336;
w5338 <= not w248 and w5337;
w5339 <= not w156 and w5338;
w5340 <= not w5318 and w5339;
w5341 <= w5318 and not w5339;
w5342 <= not w5340 and not w5341;
w5343 <= not w5322 and not w5342;
w5344 <= w5322 and w5342;
w5345 <= not w5343 and not w5344;
w5346 <= not w5323 and w5324;
w5347 <= not w3977 and not w5346;
w5348 <= not w5345 and w5347;
w5349 <= w5345 and not w5347;
w5350 <= not w5348 and not w5349;
w5351 <= w139 and w409;
w5352 <= w949 and w5351;
w5353 <= w452 and w5352;
w5354 <= w4676 and w5353;
w5355 <= w319 and w5354;
w5356 <= not w144 and w5355;
w5357 <= not w177 and w5356;
w5358 <= not w262 and w5357;
w5359 <= not w168 and w5358;
w5360 <= not w163 and w5359;
w5361 <= not w162 and w5360;
w5362 <= not w504 and w5361;
w5363 <= w5341 and not w5362;
w5364 <= not w5341 and w5362;
w5365 <= not w5363 and not w5364;
w5366 <= not w5344 and not w5365;
w5367 <= w5344 and not w5364;
w5368 <= not w5366 and not w5367;
w5369 <= not w5345 and w5346;
w5370 <= not w3977 and not w5369;
w5371 <= not w5368 and w5370;
w5372 <= w5368 and not w5370;
w5373 <= not w5371 and not w5372;
w5374 <= w439 and w3567;
w5375 <= w394 and w5374;
w5376 <= not w293 and w5375;
w5377 <= not w310 and w5376;
w5378 <= not w5363 and w5377;
w5379 <= w5363 and not w5377;
w5380 <= not w5378 and not w5379;
w5381 <= not w5367 and not w5380;
w5382 <= w5367 and w5380;
w5383 <= not w5381 and not w5382;
w5384 <= not w5368 and w5369;
w5385 <= not w3977 and not w5384;
w5386 <= not w5383 and w5385;
w5387 <= w5383 and not w5385;
w5388 <= not w5386 and not w5387;
w5389 <= w394 and w467;
w5390 <= w5379 and not w5389;
w5391 <= not w5379 and w5389;
w5392 <= not w5390 and not w5391;
w5393 <= not w5382 and not w5392;
w5394 <= w5382 and not w5391;
w5395 <= not w5393 and not w5394;
w5396 <= not w5383 and w5384;
w5397 <= not w3977 and not w5396;
w5398 <= not w5395 and w5397;
w5399 <= w5395 and not w5397;
w5400 <= not w5398 and not w5399;
w5401 <= not a(22) and w21;
w5402 <= not w5390 and not w5394;
w5403 <= w5390 and w5394;
w5404 <= not w5402 and not w5403;
w5405 <= not w5395 and w5396;
w5406 <= not w3977 and not w5405;
w5407 <= w5404 and not w5406;
w5408 <= not w5404 and w5406;
w5409 <= not w5407 and not w5408;
w5410 <= not w5401 and w5409;
w5411 <= not w5402 and w5405;
w5412 <= not w5403 and not w5405;
w5413 <= not w5411 and not w5412;
w5414 <= not w5401 and w5413;
w5415 <= not w3977 and not w5414;
one <= '1';
sin(0) <= not w3824;-- level 177
sin(1) <= not w3981;-- level 180
sin(2) <= not w4112;-- level 185
sin(3) <= w4230;-- level 187
sin(4) <= not w4339;-- level 189
sin(5) <= not w4454;-- level 190
sin(6) <= not w4567;-- level 191
sin(7) <= not w4666;-- level 193
sin(8) <= not w4766;-- level 195
sin(9) <= not w4849;-- level 197
sin(10) <= not w4936;-- level 199
sin(11) <= not w5000;-- level 201
sin(12) <= not w5070;-- level 203
sin(13) <= not w5138;-- level 208
sin(14) <= not w5193;-- level 210
sin(15) <= not w5244;-- level 213
sin(16) <= not w5283;-- level 216
sin(17) <= w5305;-- level 218
sin(18) <= not w5328;-- level 219
sin(19) <= not w5350;-- level 220
sin(20) <= not w5373;-- level 221
sin(21) <= not w5388;-- level 222
sin(22) <= not w5400;-- level 223
sin(23) <= not w5410;-- level 225
sin(24) <= w5415;-- level 225
end Behavioral;