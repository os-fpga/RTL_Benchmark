//
// Exhibits situation where design has a very small number of inputs.
// Here 9 inputs : theoritically we should map on maximum 11 Lut6 with BDD/mux
// decomposition.
//

module top ( 
    ys__n17, ys__n27, ys__n30, ys__n45, ys__n50, ys__n65, ys__n74, ys__n77,
    ys__n119,
    ys__n2841  );
  input  ys__n17, ys__n27, ys__n30, ys__n45, ys__n50, ys__n65, ys__n74,
    ys__n77, ys__n119;
  output ys__n2841;
  wire new_ys__n136_, new_new_new_ys__n11___, new_new_new_ys__n15___,
    new_new_new_ys__n0___, new_new_new_ys__n4___, new_new_new_ys__n5___,
    new_new_new_ys__n6___, new_new_new_ys__n7___, new_new_new_ys__n8___,
    new_new_new_ys__n12___, new_new_new_ys__n13___, new_new_new_ys__n14___,
    new_new_new_ys__n16___, new_new_new_ys__n18___, new_new_new_ys__n19___,
    new_new_new_ys__n20___, new_new_new_ys__n21___, new_new_new_ys__n22___,
    new_new_new_ys__n23___, new_new_new_ys__n24___, new_new_new_ys__n25___,
    new_new_new_ys__n26___, new_new_new_ys__n28___, new_new_new_ys__n29___,
    new_new_new_ys__n31___, new_new_new_ys__n33___, new_new_new_ys__n35___,
    new_new_new_ys__n36___, new_new_new_ys__n38___, new_new_new_ys__n39___,
    new_new_new_ys__n40___, new_new_new_ys__n41___, new_new_new_ys__n42___,
    new_new_new_ys__n43___, new_new_new_ys__n44___, new_new_new_ys__n47___,
    new_new_new_ys__n52___, new_new_new_ys__n54___, new_new_new_ys__n56___,
    new_new_new_ys__n59___, new_new_new_ys__n61___, new_new_new_ys__n63___,
    new_new_new_ys__n64___, new_new_new_ys__n68___, new_new_new_ys__n71___,
    new_new_new_ys__n73___, new_new_new_ys__n76___, new_new_new_ys__n88___,
    new_new_new_ys__n96___, new_new_new_ys__n98___,
    new_new_new_ys__n100___, new_new_new_ys__n104___,
    new_new_new_ys__n114___, new_new_new_ys__n121___,
    new_new_new_ys__n123___, new_new_new_ys__n124___,
    new_new_new_ys__n126___, new_new_new_ys__n132___,
    new_new_new_ys__n140___, new_new_new_ys__n141___,
    new_new_new_ys__n148___, new_new_new_ys__n149___,
    new_new_new_ys__n150___, new_new_new_ys__n161___,
    new_new_new_ys__n179___, new_new_new_ys__n185___,
    new_new_new_ys__n186___, new_new_new_ys__n188___,
    new_new_new_ys__n190___, new_new_new_ys__n194___,
    new_new_new_ys__n196___, new_new_new_ys__n203___,
    new_new_new_ys__n205___, new_new_new_ys__n208___,
    new_new_new_ys__n209___, new_new_new_ys__n210___,
    new_new_new_ys__n211___, new_new_new_ys__n212___,
    new_new_new_ys__n213___, new_new_new_ys__n214___,
    new_new_new_ys__n215___, new_new_new_ys__n216___,
    new_new_new_ys__n217___, new_new_new_ys__n218___,
    new_new_new_ys__n219___, new_new_new_ys__n220___,
    new_new_new_ys__n221___, new_new_new_ys__n231___,
    new_new_new_ys__n232___, new_new_new_ys__n233___,
    new_new_new_ys__n234___, new_new_new_ys__n235___,
    new_new_new_ys__n236___, new_new_new_ys__n237___,
    new_new_new_ys__n238___, new_new_new_ys__n239___,
    new_new_new_ys__n240___, new_new_new_ys__n249___,
    new_new_new_ys__n250___, new_new_new_ys__n252___,
    new_new_new_ys__n253___, new_new_new_ys__n254___,
    new_new_new_ys__n255___, new_new_new_ys__n256___,
    new_new_new_ys__n257___, new_new_new_ys__n258___,
    new_new_new_ys__n259___, new_new_new_ys__n260___,
    new_new_new_ys__n261___, new_new_new_ys__n262___,
    new_new_new_ys__n263___, new_new_new_ys__n264___,
    new_new_new_ys__n265___, new_new_new_ys__n266___,
    new_new_new_ys__n267___, new_new_new_ys__n268___,
    new_new_new_ys__n269___, new_new_new_ys__n270___,
    new_new_new_ys__n271___, new_new_new_ys__n272___,
    new_new_new_ys__n273___, new_new_new_ys__n286___,
    new_new_new_ys__n297___, new_new_new_ys__n309___,
    new_new_new_ys__n319___, new_new_new_ys__n331___,
    new_new_new_ys__n337___, new_new_new_ys__n348___,
    new_new_new_ys__n356___, new_new_new_ys__n357___,
    new_new_new_ys__n366___, new_new_new_ys__n389___,
    new_new_new_ys__n396___, new_new_new_ys__n398___,
    new_new_new_ys__n402___, new_new_new_ys__n403___,
    new_new_new_ys__n404___, new_new_new_ys__n405___,
    new_new_new_ys__n406___, new_new_new_ys__n407___,
    new_new_new_ys__n408___, new_new_new_ys__n409___,
    new_new_new_ys__n410___, new_new_new_ys__n414___,
    new_new_new_ys__n416___, new_new_new_ys__n417___,
    new_new_new_ys__n418___, new_new_new_ys__n419___,
    new_new_new_ys__n420___, new_new_new_ys__n421___,
    new_new_new_ys__n422___, new_new_new_ys__n423___,
    new_new_new_ys__n424___, new_new_new_ys__n425___,
    new_new_new_ys__n426___, new_new_new_ys__n427___,
    new_new_new_ys__n428___, new_new_new_ys__n429___,
    new_new_new_ys__n430___, new_new_new_ys__n431___,
    new_new_new_ys__n432___, new_new_new_ys__n449___,
    new_new_new_ys__n452___, new_new_new_ys__n455___,
    new_new_new_ys__n456___, new_new_new_ys__n457___,
    new_new_new_ys__n458___, new_new_new_ys__n459___,
    new_new_new_ys__n460___, new_new_new_ys__n461___,
    new_new_new_ys__n462___, new_new_new_ys__n470___,
    new_new_new_ys__n474___, new_new_new_ys__n475___,
    new_new_new_ys__n476___, new_new_new_ys__n487___,
    new_new_new_ys__n488___, new_new_new_ys__n495___,
    new_new_new_ys__n507___, new_new_new_ys__n517___,
    new_new_new_ys__n518___, new_new_new_ys__n519___,
    new_new_new_ys__n520___, new_new_new_ys__n521___,
    new_new_new_ys__n522___, new_new_new_ys__n523___,
    new_new_new_ys__n524___, new_new_new_ys__n525___,
    new_new_new_ys__n526___, new_new_new_ys__n527___,
    new_new_new_ys__n528___, new_new_new_ys__n529___,
    new_new_new_ys__n530___, new_new_new_ys__n531___,
    new_new_new_ys__n532___, new_new_new_ys__n533___,
    new_new_new_ys__n534___, new_new_new_ys__n535___,
    new_new_new_ys__n536___, new_new_new_ys__n537___,
    new_new_new_ys__n538___, new_new_new_ys__n539___,
    new_new_new_ys__n540___, new_new_new_ys__n541___,
    new_new_new_ys__n542___, new_new_new_ys__n543___,
    new_new_new_ys__n544___, new_new_new_ys__n545___,
    new_new_new_ys__n546___, new_new_new_ys__n547___,
    new_new_new_ys__n548___, new_new_new_ys__n549___,
    new_new_new_ys__n561___, new_new_new_ys__n562___,
    new_new_new_ys__n563___, new_new_new_ys__n564___,
    new_new_new_ys__n565___, new_new_new_ys__n566___,
    new_new_new_ys__n567___, new_new_new_ys__n568___,
    new_new_new_ys__n569___, new_new_new_ys__n570___,
    new_new_new_ys__n571___, new_new_new_ys__n572___,
    new_new_new_ys__n573___, new_new_new_ys__n574___,
    new_new_new_ys__n575___, new_new_new_ys__n576___,
    new_new_new_ys__n577___, new_new_new_ys__n578___,
    new_new_new_ys__n579___, new_new_new_ys__n580___,
    new_new_new_ys__n581___, new_new_new_ys__n582___,
    new_new_new_ys__n583___, new_new_new_ys__n584___,
    new_new_new_ys__n585___, new_new_new_ys__n586___,
    new_new_new_ys__n587___, new_new_new_ys__n588___,
    new_new_new_ys__n589___, new_new_new_ys__n590___,
    new_new_new_ys__n591___, new_new_new_ys__n592___,
    new_new_new_ys__n593___, new_new_new_ys__n594___,
    new_new_new_ys__n595___, new_new_new_ys__n596___,
    new_new_new_ys__n597___, new_new_new_ys__n598___,
    new_new_new_ys__n599___, new_new_new_ys__n600___,
    new_new_new_ys__n601___, new_new_new_ys__n602___,
    new_new_new_ys__n603___, new_new_new_ys__n604___,
    new_new_new_ys__n605___, new_new_new_ys__n606___,
    new_new_new_ys__n607___, new_new_new_ys__n608___,
    new_new_new_ys__n609___, new_new_new_ys__n610___,
    new_new_new_ys__n611___, new_new_new_ys__n612___,
    new_new_new_ys__n613___, new_new_new_ys__n614___,
    new_new_new_ys__n615___, new_new_new_ys__n616___,
    new_new_new_ys__n617___, new_new_new_ys__n618___,
    new_new_new_ys__n619___, new_new_new_ys__n642___,
    new_new_new_ys__n643___, new_new_new_ys__n644___,
    new_new_new_ys__n645___, new_new_new_ys__n646___,
    new_new_new_ys__n647___, new_new_new_ys__n648___,
    new_new_new_ys__n649___, new_new_new_ys__n650___,
    new_new_new_ys__n651___, new_new_new_ys__n652___,
    new_new_new_ys__n665___, new_new_new_ys__n666___,
    new_new_new_ys__n667___, new_new_new_ys__n668___,
    new_new_new_ys__n669___, new_new_new_ys__n670___,
    new_new_new_ys__n683___, new_new_new_ys__n690___,
    new_new_new_ys__n691___, new_new_new_ys__n692___,
    new_new_new_ys__n693___, new_new_new_ys__n694___,
    new_new_new_ys__n695___, new_new_new_ys__n696___,
    new_new_new_ys__n697___, new_new_new_ys__n698___,
    new_new_new_ys__n699___, new_new_new_ys__n700___,
    new_new_new_ys__n728___, new_new_new_ys__n729___,
    new_new_new_ys__n730___, new_new_new_ys__n731___,
    new_new_new_ys__n732___, new_new_new_ys__n733___,
    new_new_new_ys__n734___, new_new_new_ys__n735___,
    new_new_new_ys__n745___, new_new_new_ys__n746___,
    new_new_new_ys__n747___, new_new_new_ys__n748___,
    new_new_new_ys__n749___, new_new_new_ys__n750___,
    new_new_new_ys__n751___, new_new_new_ys__n752___,
    new_new_new_ys__n753___, new_new_new_ys__n754___,
    new_new_new_ys__n755___, new_new_new_ys__n756___,
    new_new_new_ys__n757___, new_new_new_ys__n773___,
    new_new_new_ys__n813___, new_new_new_ys__n826___,
    new_new_new_ys__n827___, new_new_new_ys__n828___,
    new_new_new_ys__n829___, new_new_new_ys__n830___,
    new_new_new_ys__n831___, new_new_new_ys__n832___,
    new_new_new_ys__n833___, new_new_new_ys__n834___,
    new_new_new_ys__n835___, new_new_new_ys__n871___,
    new_new_new_ys__n872___, new_new_new_ys__n873___,
    new_new_new_ys__n874___, new_new_new_ys__n875___,
    new_new_new_ys__n876___, new_new_new_ys__n877___,
    new_new_new_ys__n878___, new_new_new_ys__n879___,
    new_new_new_ys__n880___, new_new_new_ys__n881___,
    new_new_new_ys__n882___, new_new_new_ys__n883___,
    new_new_new_ys__n884___, new_new_new_ys__n902___,
    new_new_new_ys__n903___, new_new_new_ys__n1039___,
    new_new_new_ys__n1040___, new_new_new_ys__n1041___,
    new_new_new_ys__n1042___, new_new_new_ys__n1043___,
    new_new_new_ys__n1044___, new_new_new_ys__n1045___,
    new_new_new_ys__n1046___, new_new_new_ys__n1047___,
    new_new_new_ys__n1048___, new_new_new_ys__n1049___,
    new_new_new_ys__n1050___, new_new_new_ys__n1051___,
    new_new_new_ys__n1052___, new_new_new_ys__n1053___,
    new_new_new_ys__n1054___, new_new_new_ys__n1064___,
    new_new_new_ys__n1067___, new_new_new_ys__n1068___,
    new_new_new_ys__n1069___, new_new_new_ys__n1070___,
    new_new_new_ys__n1071___, new_new_new_ys__n1072___,
    new_new_new_ys__n1073___, new_new_new_ys__n1074___,
    new_new_new_ys__n1148___, new_new_new_ys__n1149___,
    new_new_new_ys__n1150___, new_new_new_ys__n1151___,
    new_new_new_ys__n1152___, new_new_new_ys__n1153___,
    new_new_new_ys__n1154___, new_new_new_ys__n1155___,
    new_new_new_ys__n1156___, new_new_new_ys__n1157___,
    new_new_new_ys__n1158___, new_new_new_ys__n1159___,
    new_new_new_ys__n1161___, new_new_new_ys__n1171___,
    new_new_new_ys__n1172___, new_new_new_ys__n1173___,
    new_new_new_ys__n1174___, new_new_new_ys__n1175___,
    new_new_new_ys__n1176___, new_new_new_ys__n1177___,
    new_new_new_ys__n1184___, new_new_new_ys__n1197___,
    new_new_new_ys__n1324___, new_new_new_ys__n1363___,
    new_new_new_ys__n1364___, new_new_new_ys__n1403___,
    new_new_new_ys__n1406___, new_new_new_ys__n1628___,
    new_new_new_ys__n1630___, new_new_new_ys__n1643___,
    new_new_new_ys__n1644___, new_new_new_ys__n1645___,
    new_new_new_ys__n1646___, new_new_new_ys__n1647___,
    new_new_new_ys__n1648___, new_new_new_ys__n1663___,
    new_new_new_ys__n1672___, new_new_new_ys__n1709___,
    new_new_new_ys__n1759___, new_new_new_ys__n1760___,
    new_new_new_ys__n1761___, new_new_new_ys__n1762___,
    new_new_new_ys__n1786___, new_new_new_ys__n1788___,
    new_new_new_ys__n1798___, new_new_new_ys__n1817___,
    new_new_new_ys__n1980___, new_new_new_ys__n1981___,
    new_new_new_ys__n1982___, new_new_new_ys__n1983___,
    new_new_new_ys__n1984___, new_new_new_ys__n1985___,
    new_new_new_ys__n1986___, new_new_new_ys__n1991___,
    new_new_new_ys__n1992___, new_new_new_ys__n1993___,
    new_new_new_ys__n1994___, new_new_new_ys__n1995___,
    new_new_new_ys__n1996___, new_new_new_ys__n1997___,
    new_new_new_ys__n1998___, new_new_new_ys__n1999___,
    new_new_new_ys__n2000___, new_new_new_ys__n2009___,
    new_new_new_ys__n2010___, new_new_new_ys__n2011___,
    new_new_new_ys__n2029___, new_new_new_ys__n2030___,
    new_new_new_ys__n2031___, new_new_new_ys__n2032___,
    new_new_new_ys__n2033___, new_new_new_ys__n2037___,
    new_new_new_ys__n2038___, new_new_new_ys__n2039___,
    new_new_new_ys__n2040___, new_new_new_ys__n2041___,
    new_new_new_ys__n2042___, new_new_new_ys__n2043___,
    new_new_new_ys__n2044___, new_new_new_ys__n2045___,
    new_new_new_ys__n2046___, new_new_new_ys__n2047___,
    new_new_new_ys__n2048___, new_new_new_ys__n2049___,
    new_new_new_ys__n2050___, new_new_new_ys__n2051___,
    new_new_new_ys__n2052___, new_new_new_ys__n2053___,
    new_new_new_ys__n2054___, new_new_new_ys__n2055___,
    new_new_new_ys__n2056___, new_new_new_ys__n2100___,
    new_new_new_ys__n2101___, new_new_new_ys__n2102___,
    new_new_new_ys__n2103___, new_new_new_ys__n2104___,
    new_new_new_ys__n2105___, new_new_new_ys__n2106___,
    new_new_new_ys__n2107___, new_new_new_ys__n2108___,
    new_new_new_ys__n2109___, new_new_new_ys__n2110___,
    new_new_new_ys__n2111___, new_new_new_ys__n2112___,
    new_new_new_ys__n2113___, new_new_new_ys__n2114___,
    new_new_new_ys__n2115___, new_new_new_ys__n2116___,
    new_new_new_ys__n2117___, new_new_new_ys__n2118___,
    new_new_new_ys__n2119___, new_new_new_ys__n2120___,
    new_new_new_ys__n2121___, new_new_new_ys__n2122___,
    new_new_new_ys__n2123___, new_new_new_ys__n2124___,
    new_new_new_ys__n2125___, new_new_new_ys__n2126___,
    new_new_new_ys__n2154___, new_new_new_ys__n2155___,
    new_new_new_ys__n2156___, new_new_new_ys__n2157___,
    new_new_new_ys__n2158___, new_new_new_ys__n2159___,
    new_new_new_ys__n2160___, new_new_new_ys__n2161___,
    new_new_new_ys__n2162___, new_new_new_ys__n2163___,
    new_new_new_ys__n2164___, new_new_new_ys__n2165___,
    new_new_new_ys__n2166___, new_new_new_ys__n2175___,
    new_new_new_ys__n2176___, new_new_new_ys__n2177___,
    new_new_new_ys__n2178___, new_new_new_ys__n2179___,
    new_new_new_ys__n2180___, new_new_new_ys__n2181___,
    new_new_new_ys__n2182___, new_new_new_ys__n2183___,
    new_new_new_ys__n2184___, new_new_new_ys__n2185___,
    new_new_new_ys__n2186___, new_new_new_ys__n2187___,
    new_new_new_ys__n2188___, new_new_new_ys__n2189___,
    new_new_new_ys__n2190___, new_new_new_ys__n2191___,
    new_new_new_ys__n2192___, new_new_new_ys__n2193___,
    new_new_new_ys__n2194___, new_new_new_ys__n2195___,
    new_new_new_ys__n2196___, new_new_new_ys__n2197___,
    new_new_new_ys__n2198___, new_new_new_ys__n2199___,
    new_new_new_ys__n2200___, new_new_new_ys__n2201___,
    new_new_new_ys__n2202___, new_new_new_ys__n2203___,
    new_new_new_ys__n2204___, new_new_new_ys__n2205___,
    new_new_new_ys__n2206___, new_new_new_ys__n2375___,
    new_new_new_ys__n2376___, new_new_new_ys__n2377___,
    new_new_new_ys__n2378___, new_new_new_ys__n2379___,
    new_new_new_ys__n2380___, new_new_new_ys__n2381___,
    new_new_new_ys__n2382___, new_new_new_ys__n2383___,
    new_new_new_ys__n2384___, new_new_new_ys__n2385___,
    new_new_new_ys__n2386___, new_new_new_ys__n2390___,
    new_new_new_ys__n2393___, new_new_new_ys__n2394___,
    new_new_new_ys__n2395___, new_new_new_ys__n2396___,
    new_new_new_ys__n2397___, new_new_new_ys__n2398___,
    new_new_new_ys__n2399___, new_new_new_ys__n2400___,
    new_new_new_ys__n2423___, new_new_new_ys__n2518___,
    new_new_new_ys__n2552___, new_new_new_ys__n2553___,
    new_new_new_ys__n2554___, new_new_new_ys__n2555___,
    new_new_new_ys__n2568___, new_new_new_ys__n2668___,
    new_new_new_ys__n2719___, new_new_new_ys__n2720___,
    new_new_new_ys__n2721___, new_new_new_ys__n2722___,
    new_new_new_ys__n2778___, new_new_new_ys__n2779___,
    new_new_new_ys__n2788___, new_new_new_ys__n2791___,
    new_new_new_ys__n2821___, new_new_new_ys__n2822___,
    new_new_new_ys__n2823___, new_new_new_ys__n2824___,
    new_new_new_ys__n2825___, new_new_new_ys__n2826___,
    new_new_new_ys__n2827___, new_new_new_ys__n2828___,
    new_new_new_ys__n2829___, new_new_new_ys__n2830___,
    new_new_new_ys__n2831___, new_new_new_ys__n2832___,
    new_new_new_ys__n2833___, new_new_new_ys__n2834___,
    new_new_new_ys__n2835___, new_new_new_ys__n2836___,
    new_new_new_ys__n2837___, new_new_new_ys__n2838___,
    new_new_new_ys__n2839___, new_new_new_ys__n2840___,
    new_new_new_ys__n2848___, new_new_new_ys__n2866___,
    new_new_new_ys__n2867___, new_new_new_ys__n2868___,
    new_new_new_ys__n2869___, new_new_new_ys__n2882___,
    new_new_new_ys__n2883___, new_new_new_ys__n2884___,
    new_new_new_ys__n2894___, new_new_new_ys__n2895___,
    new_new_new_ys__n2896___, new_new_new_ys__n2897___,
    new_new_new_ys__n2898___, new_new_new_ys__n2899___,
    new_new_new_ys__n2900___, new_new_new_ys__n2901___,
    new_new_new_ys__n2902___, new_new_new_ys__n2903___,
    new_new_new_ys__n2904___, new_new_new_ys__n2905___,
    new_new_new_ys__n2906___, new_new_new_ys__n2918___,
    new_new_new_ys__n2919___, new_new_new_ys__n2920___,
    new_new_new_ys__n2921___, new_new_new_ys__n2922___,
    new_new_new_ys__n2923___, new_new_new_ys__n2924___,
    new_new_new_ys__n2945___, new_new_new_ys__n2946___,
    new_new_new_ys__n2960___, new_new_new_ys__n2961___,
    new_new_new_ys__n2962___, new_new_new_ys__n2963___,
    new_new_new_ys__n2964___, new_new_new_ys__n2965___,
    new_new_new_ys__n2966___, new_new_new_ys__n2967___,
    new_new_new_ys__n2972___, new_new_new_ys__n2973___,
    new_new_new_ys__n2974___, new_new_new_ys__n2975___,
    new_new_new_ys__n2976___, new_new_new_ys__n2981___,
    new_new_new_ys__n2982___, new_new_new_ys__n2983___,
    new_new_new_ys__n2984___, new_new_new_ys__n2985___,
    new_new_new_ys__n2992___, new_new_new_ys__n2993___,
    new_new_new_ys__n2994___, new_new_new_ys__n2995___,
    new_new_new_ys__n2996___, new_new_new_ys__n2997___,
    new_new_new_ys__n2998___, new_new_new_ys__n2999___,
    new_new_new_ys__n3000___, new_new_new_ys__n3029___,
    new_new_new_ys__n3030___, new_new_new_ys__n3031___,
    new_new_new_ys__n3032___, new_new_new_ys__n3033___,
    new_new_new_ys__n3034___, new_new_new_ys__n3035___,
    new_new_new_ys__n3040___, new_new_new_ys__n3041___,
    new_new_new_ys__n3042___, new_new_new_ys__n3043___,
    new_new_new_ys__n3075___, new_new_new_ys__n3076___,
    new_new_new_ys__n3077___;
  assign new_ys__n136_ = 1'b1;
  assign new_new_new_ys__n11___ = 1'b0;
  assign new_new_new_ys__n15___ = 1'b1;
  assign new_new_new_ys__n0___ = ys__n77 ? new_new_new_ys__n11___ : new_new_new_ys__n8___;
  assign new_new_new_ys__n4___ = ys__n74 ? new_ys__n136_ : new_new_new_ys__n15___;
  assign new_new_new_ys__n5___ = ys__n74 ? new_ys__n136_ : new_new_new_ys__n8___;
  assign new_new_new_ys__n6___ = new_new_new_ys__n487___ ? new_new_new_ys__n33___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n7___ = new_new_new_ys__n6___ ? new_new_new_ys__n5___ : new_new_new_ys__n4___;
  assign new_new_new_ys__n8___ = ~new_ys__n136_;
  assign new_new_new_ys__n12___ = ~new_new_new_ys__n96___;
  assign new_new_new_ys__n13___ = ys__n50 ? new_new_new_ys__n2568___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n14___ = new_new_new_ys__n13___ ? new_new_new_ys__n12___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n16___ = new_new_new_ys__n13___ ? new_new_new_ys__n12___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n18___ = ys__n17 ? new_new_new_ys__n11___ : new_new_new_ys__n12___;
  assign new_new_new_ys__n19___ = ~new_new_new_ys__n13___;
  assign new_new_new_ys__n20___ = ys__n17 ? new_new_new_ys__n11___ : new_new_new_ys__n19___;
  assign new_new_new_ys__n21___ = ys__n17 ? new_new_new_ys__n14___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n22___ = ys__n17 ? new_new_new_ys__n16___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n23___ = ys__n17 ? new_new_new_ys__n2113___ : new_new_new_ys__n2112___;
  assign new_new_new_ys__n24___ = new_new_new_ys__n23___ ? new_new_new_ys__n15___ : new_new_new_ys__n18___;
  assign new_new_new_ys__n25___ = new_new_new_ys__n23___ ? new_new_new_ys__n15___ : new_new_new_ys__n20___;
  assign new_new_new_ys__n26___ = new_new_new_ys__n23___ ? new_new_new_ys__n22___ : new_new_new_ys__n21___;
  assign new_new_new_ys__n28___ = ys__n27 ? new_new_new_ys__n15___ : new_new_new_ys__n24___;
  assign new_new_new_ys__n29___ = ys__n27 ? new_new_new_ys__n26___ : new_new_new_ys__n25___;
  assign new_new_new_ys__n31___ = ys__n30 ? new_new_new_ys__n29___ : new_new_new_ys__n28___;
  assign new_new_new_ys__n33___ = ys__n17 ? new_new_new_ys__n11___ : new_new_new_ys__n1363___;
  assign new_new_new_ys__n35___ = ~new_new_new_ys__n813___;
  assign new_new_new_ys__n36___ = new_ys__n136_ ? new_new_new_ys__n2779___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n38___ = new_new_new_ys__n460___ ? new_new_new_ys__n459___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n39___ = ys__n50 ? new_new_new_ys__n2000___ : new_new_new_ys__n1999___;
  assign new_new_new_ys__n40___ = new_new_new_ys__n190___ ? ys__n119 : new_new_new_ys__n11___;
  assign new_new_new_ys__n41___ = new_new_new_ys__n40___ ? new_new_new_ys__n39___ : new_new_new_ys__n38___;
  assign new_new_new_ys__n42___ = new_new_new_ys__n357___ ? new_new_new_ys__n2011___ : new_new_new_ys__n2009___;
  assign new_new_new_ys__n43___ = new_new_new_ys__n42___ ? new_new_new_ys__n41___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n44___ = ~new_new_new_ys__n190___;
  assign new_new_new_ys__n47___ = ~new_new_new_ys__n488___;
  assign new_new_new_ys__n52___ = new_new_new_ys__n331___ ? new_new_new_ys__n73___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n54___ = ys__n77 ? new_new_new_ys__n1064___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n56___ = new_new_new_ys__n309___ ? new_new_new_ys__n73___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n59___ = ys__n30 ? new_new_new_ys__n2518___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n61___ = ~new_new_new_ys__n205___;
  assign new_new_new_ys__n63___ = ~new_new_new_ys__n188___;
  assign new_new_new_ys__n64___ = ys__n30 ? new_new_new_ys__n15___ : new_new_new_ys__n63___;
  assign new_new_new_ys__n68___ = new_ys__n136_ ? new_new_new_ys__n1403___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n71___ = new_new_new_ys__n59___ ? ys__n119 : new_new_new_ys__n11___;
  assign new_new_new_ys__n73___ = ~ys__n65;
  assign new_new_new_ys__n76___ = ~ys__n74;
  assign new_new_new_ys__n88___ = new_new_new_ys__n527___ ? new_new_new_ys__n903___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n96___ = new_new_new_ys__n452___ ? new_new_new_ys__n132___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n98___ = new_new_new_ys__n54___ ? new_new_new_ys__n132___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n100___ = ys__n17 ? new_new_new_ys__n690___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n104___ = ~new_new_new_ys__n357___;
  assign new_new_new_ys__n114___ = ~new_new_new_ys__n56___;
  assign new_new_new_ys__n121___ = ys__n74 ? new_new_new_ys__n2924___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n123___ = ys__n30 ? new_new_new_ys__n249___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n124___ = ys__n27 ? new_new_new_ys__n461___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n126___ = new_new_new_ys__n521___ ? new_new_new_ys__n132___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n132___ = ~ys__n119;
  assign new_new_new_ys__n140___ = ~new_new_new_ys__n179___;
  assign new_new_new_ys__n141___ = ys__n27 ? new_new_new_ys__n2206___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n148___ = ~new_new_new_ys__n40___;
  assign new_new_new_ys__n149___ = new_new_new_ys__n309___ ? ys__n65 : new_new_new_ys__n11___;
  assign new_new_new_ys__n150___ = new_new_new_ys__n149___ ? new_new_new_ys__n148___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n161___ = ys__n45 ? new_new_new_ys__n1628___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n179___ = new_new_new_ys__n331___ ? ys__n65 : new_new_new_ys__n11___;
  assign new_new_new_ys__n185___ = ~new_new_new_ys__n149___;
  assign new_new_new_ys__n186___ = new_new_new_ys__n414___ ? ys__n119 : new_new_new_ys__n11___;
  assign new_new_new_ys__n188___ = ys__n77 ? new_new_new_ys__n1817___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n190___ = ys__n17 ? new_new_new_ys__n1324___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n194___ = ~new_new_new_ys__n405___;
  assign new_new_new_ys__n196___ = new_new_new_ys__n0___ ? ys__n74 : new_new_new_ys__n11___;
  assign new_new_new_ys__n203___ = ys__n65 ? new_new_new_ys__n2848___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n205___ = new_ys__n136_ ? new_new_new_ys__n2423___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n208___ = ys__n77 ? ys__n119 : new_new_new_ys__n15___;
  assign new_new_new_ys__n209___ = ys__n77 ? new_new_new_ys__n132___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n210___ = ys__n77 ? new_new_new_ys__n15___ : ys__n119;
  assign new_new_new_ys__n211___ = ys__n74 ? new_new_new_ys__n208___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n212___ = ys__n74 ? new_new_new_ys__n15___ : new_new_new_ys__n209___;
  assign new_new_new_ys__n213___ = ys__n74 ? new_new_new_ys__n210___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n214___ = ys__n74 ? new_new_new_ys__n15___ : new_new_new_ys__n210___;
  assign new_new_new_ys__n215___ = ys__n17 ? new_new_new_ys__n15___ : new_new_new_ys__n211___;
  assign new_new_new_ys__n216___ = ys__n17 ? new_new_new_ys__n212___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n217___ = ys__n17 ? new_new_new_ys__n15___ : new_new_new_ys__n213___;
  assign new_new_new_ys__n218___ = ys__n17 ? new_new_new_ys__n214___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n219___ = ys__n30 ? new_new_new_ys__n216___ : new_new_new_ys__n215___;
  assign new_new_new_ys__n220___ = ys__n30 ? new_new_new_ys__n218___ : new_new_new_ys__n217___;
  assign new_new_new_ys__n221___ = new_ys__n136_ ? new_new_new_ys__n220___ : new_new_new_ys__n219___;
  assign new_new_new_ys__n231___ = new_new_new_ys__n68___ ? new_new_new_ys__n35___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n232___ = ys__n27 ? new_new_new_ys__n1761___ : new_new_new_ys__n1760___;
  assign new_new_new_ys__n233___ = new_new_new_ys__n232___ ? new_new_new_ys__n11___ : new_new_new_ys__n231___;
  assign new_new_new_ys__n234___ = ~new_new_new_ys__n232___;
  assign new_new_new_ys__n235___ = new_new_new_ys__n190___ ? new_new_new_ys__n1788___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n236___ = new_new_new_ys__n235___ ? new_new_new_ys__n11___ : new_new_new_ys__n233___;
  assign new_new_new_ys__n237___ = new_new_new_ys__n235___ ? new_new_new_ys__n11___ : new_new_new_ys__n234___;
  assign new_new_new_ys__n238___ = ys__n119 ? new_new_new_ys__n234___ : new_new_new_ys__n237___;
  assign new_new_new_ys__n239___ = ys__n119 ? new_new_new_ys__n237___ : new_new_new_ys__n236___;
  assign new_new_new_ys__n240___ = new_new_new_ys__n13___ ? new_new_new_ys__n239___ : new_new_new_ys__n238___;
  assign new_new_new_ys__n249___ = ys__n17 ? new_new_new_ys__n11___ : new_new_new_ys__n297___;
  assign new_new_new_ys__n250___ = new_new_new_ys__n188___ ? new_new_new_ys__n132___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n252___ = ~ys__n77;
  assign new_new_new_ys__n253___ = ys__n50 ? new_new_new_ys__n252___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n254___ = ys__n50 ? new_new_new_ys__n15___ : ys__n77;
  assign new_new_new_ys__n255___ = ys__n50 ? ys__n77 : new_new_new_ys__n15___;
  assign new_new_new_ys__n256___ = ys__n45 ? new_new_new_ys__n255___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n257___ = ys__n45 ? new_new_new_ys__n253___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n258___ = ys__n45 ? new_new_new_ys__n15___ : new_new_new_ys__n254___;
  assign new_new_new_ys__n259___ = ys__n74 ? new_new_new_ys__n15___ : new_new_new_ys__n256___;
  assign new_new_new_ys__n260___ = ys__n74 ? new_new_new_ys__n258___ : new_new_new_ys__n257___;
  assign new_new_new_ys__n261___ = ys__n65 ? new_new_new_ys__n260___ : new_new_new_ys__n259___;
  assign new_new_new_ys__n262___ = new_new_new_ys__n6___ ? new_new_new_ys__n11___ : new_new_new_ys__n2160___;
  assign new_new_new_ys__n263___ = new_new_new_ys__n521___ ? new_new_new_ys__n2123___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n264___ = new_new_new_ys__n263___ ? new_new_new_ys__n11___ : new_new_new_ys__n262___;
  assign new_new_new_ys__n265___ = ~new_new_new_ys__n263___;
  assign new_new_new_ys__n266___ = new_new_new_ys__n13___ ? new_new_new_ys__n2126___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n267___ = new_new_new_ys__n266___ ? new_new_new_ys__n11___ : new_new_new_ys__n264___;
  assign new_new_new_ys__n268___ = new_new_new_ys__n266___ ? new_new_new_ys__n11___ : new_new_new_ys__n265___;
  assign new_new_new_ys__n269___ = ys__n119 ? new_new_new_ys__n265___ : new_new_new_ys__n267___;
  assign new_new_new_ys__n270___ = ys__n119 ? new_new_new_ys__n265___ : new_new_new_ys__n268___;
  assign new_new_new_ys__n271___ = ys__n74 ? new_new_new_ys__n268___ : new_new_new_ys__n270___;
  assign new_new_new_ys__n272___ = ys__n74 ? new_new_new_ys__n270___ : new_new_new_ys__n269___;
  assign new_new_new_ys__n273___ = new_ys__n136_ ? new_new_new_ys__n272___ : new_new_new_ys__n271___;
  assign new_new_new_ys__n286___ = ~new_new_new_ys__n98___;
  assign new_new_new_ys__n297___ = ~ys__n27;
  assign new_new_new_ys__n309___ = ys__n45 ? new_new_new_ys__n11___ : new_new_new_ys__n581___;
  assign new_new_new_ys__n319___ = ~new_new_new_ys__n141___;
  assign new_new_new_ys__n331___ = ys__n45 ? ys__n50 : new_new_new_ys__n11___;
  assign new_new_new_ys__n337___ = ~ys__n30;
  assign new_new_new_ys__n348___ = ~new_new_new_ys__n71___;
  assign new_new_new_ys__n356___ = ~new_new_new_ys__n100___;
  assign new_new_new_ys__n357___ = new_new_new_ys__n68___ ? new_new_new_ys__n132___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n366___ = ~ys__n45;
  assign new_new_new_ys__n389___ = ~new_new_new_ys__n124___;
  assign new_new_new_ys__n396___ = ~new_new_new_ys__n68___;
  assign new_new_new_ys__n398___ = ~new_new_new_ys__n54___;
  assign new_new_new_ys__n402___ = new_new_new_ys__n123___ ? ys__n119 : new_new_new_ys__n15___;
  assign new_new_new_ys__n403___ = new_new_new_ys__n52___ ? new_new_new_ys__n11___ : new_new_new_ys__n402___;
  assign new_new_new_ys__n404___ = ~new_new_new_ys__n52___;
  assign new_new_new_ys__n405___ = new_new_new_ys__n33___ ? ys__n119 : new_new_new_ys__n11___;
  assign new_new_new_ys__n406___ = new_new_new_ys__n405___ ? new_new_new_ys__n404___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n407___ = new_new_new_ys__n405___ ? new_new_new_ys__n403___ : new_new_new_ys__n402___;
  assign new_new_new_ys__n408___ = new_new_new_ys__n203___ ? new_new_new_ys__n194___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n409___ = new_new_new_ys__n203___ ? new_new_new_ys__n407___ : new_new_new_ys__n406___;
  assign new_new_new_ys__n410___ = ys__n77 ? new_new_new_ys__n409___ : new_new_new_ys__n408___;
  assign new_new_new_ys__n414___ = ys__n27 ? new_new_new_ys__n1630___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n416___ = ys__n45 ? new_new_new_ys__n11___ : new_new_new_ys__n104___;
  assign new_new_new_ys__n417___ = ys__n45 ? new_new_new_ys__n15___ : new_new_new_ys__n104___;
  assign new_new_new_ys__n418___ = ys__n45 ? new_new_new_ys__n15___ : new_new_new_ys__n286___;
  assign new_new_new_ys__n419___ = ys__n50 ? new_new_new_ys__n416___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n420___ = ys__n50 ? new_new_new_ys__n418___ : new_new_new_ys__n417___;
  assign new_new_new_ys__n421___ = ys__n65 ? new_new_new_ys__n420___ : new_new_new_ys__n419___;
  assign new_new_new_ys__n422___ = new_new_new_ys__n240___ ? new_new_new_ys__n1054___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n423___ = new_new_new_ys__n603___ ? new_new_new_ys__n602___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n424___ = new_new_new_ys__n423___ ? new_new_new_ys__n422___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n425___ = ys__n45 ? new_new_new_ys__n2400___ : new_new_new_ys__n2399___;
  assign new_new_new_ys__n426___ = new_new_new_ys__n425___ ? new_new_new_ys__n424___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n427___ = ys__n74 ? new_new_new_ys__n2380___ : new_new_new_ys__n2376___;
  assign new_new_new_ys__n428___ = new_new_new_ys__n427___ ? new_new_new_ys__n426___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n429___ = ys__n50 ? new_new_new_ys__n1159___ : new_new_new_ys__n1158___;
  assign new_new_new_ys__n430___ = new_new_new_ys__n429___ ? new_new_new_ys__n428___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n431___ = new_new_new_ys__n124___ ? new_new_new_ys__n1648___ : new_new_new_ys__n1647___;
  assign new_new_new_ys__n432___ = new_new_new_ys__n431___ ? new_new_new_ys__n430___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n449___ = new_new_new_ys__n54___ ? new_new_new_ys__n537___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n452___ = new_new_new_ys__n0___ ? new_new_new_ys__n76___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n455___ = ~new_new_new_ys__n59___;
  assign new_new_new_ys__n456___ = new_new_new_ys__n421___ ? new_new_new_ys__n15___ : new_new_new_ys__n455___;
  assign new_new_new_ys__n457___ = new_new_new_ys__n488___ ? new_new_new_ys__n585___ : new_new_new_ys__n584___;
  assign new_new_new_ys__n458___ = new_new_new_ys__n421___ ? new_new_new_ys__n15___ : new_new_new_ys__n457___;
  assign new_new_new_ys__n459___ = ys__n45 ? new_new_new_ys__n458___ : new_new_new_ys__n456___;
  assign new_new_new_ys__n460___ = new_new_new_ys__n141___ ? new_new_new_ys__n3077___ : new_new_new_ys__n3075___;
  assign new_new_new_ys__n461___ = ys__n17 ? new_new_new_ys__n11___ : new_new_new_ys__n337___;
  assign new_new_new_ys__n462___ = ~new_new_new_ys__n203___;
  assign new_new_new_ys__n470___ = new_new_new_ys__n196___ ? new_new_new_ys__n132___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n474___ = new_new_new_ys__n121___ ? new_new_new_ys__n132___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n475___ = new_new_new_ys__n474___ ? new_new_new_ys__n124___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n476___ = new_new_new_ys__n13___ ? new_new_new_ys__n475___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n487___ = ys__n65 ? new_new_new_ys__n1364___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n488___ = new_new_new_ys__n813___ ? ys__n119 : new_new_new_ys__n11___;
  assign new_new_new_ys__n495___ = ~new_new_new_ys__n121___;
  assign new_new_new_ys__n507___ = new_new_new_ys__n533___ ? new_new_new_ys__n532___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n517___ = new_new_new_ys__n54___ ? new_new_new_ys__n194___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n518___ = new_new_new_ys__n56___ ? new_new_new_ys__n517___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n519___ = new_new_new_ys__n52___ ? new_new_new_ys__n2555___ : new_new_new_ys__n2553___;
  assign new_new_new_ys__n520___ = new_new_new_ys__n519___ ? new_new_new_ys__n518___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n521___ = ys__n74 ? new_new_new_ys__n773___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n522___ = new_new_new_ys__n521___ ? new_new_new_ys__n140___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n523___ = new_new_new_ys__n100___ ? ys__n119 : new_new_new_ys__n11___;
  assign new_new_new_ys__n524___ = new_new_new_ys__n523___ ? new_new_new_ys__n522___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n525___ = new_new_new_ys__n56___ ? new_new_new_ys__n11___ : new_new_new_ys__n524___;
  assign new_new_new_ys__n526___ = new_new_new_ys__n36___ ? new_new_new_ys__n525___ : new_new_new_ys__n524___;
  assign new_new_new_ys__n527___ = new_new_new_ys__n123___ ? new_new_new_ys__n526___ : new_new_new_ys__n524___;
  assign new_new_new_ys__n528___ = ys__n30 ? new_new_new_ys__n652___ : new_new_new_ys__n651___;
  assign new_new_new_ys__n529___ = new_ys__n136_ ? new_new_new_ys__n528___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n530___ = new_ys__n136_ ? new_new_new_ys__n735___ : new_new_new_ys__n734___;
  assign new_new_new_ys__n531___ = new_new_new_ys__n530___ ? new_new_new_ys__n11___ : new_new_new_ys__n529___;
  assign new_new_new_ys__n532___ = new_new_new_ys__n59___ ? new_new_new_ys__n531___ : new_new_new_ys__n529___;
  assign new_new_new_ys__n533___ = ys__n50 ? new_new_new_ys__n570___ : new_new_new_ys__n569___;
  assign new_new_new_ys__n534___ = new_new_new_ys__n523___ ? new_new_new_ys__n11___ : new_new_new_ys__n348___;
  assign new_new_new_ys__n535___ = new_new_new_ys__n123___ ? ys__n119 : new_new_new_ys__n11___;
  assign new_new_new_ys__n536___ = new_new_new_ys__n535___ ? new_new_new_ys__n11___ : new_new_new_ys__n534___;
  assign new_new_new_ys__n537___ = ~new_new_new_ys__n535___;
  assign new_new_new_ys__n538___ = new_new_new_ys__n54___ ? new_new_new_ys__n536___ : new_new_new_ys__n534___;
  assign new_new_new_ys__n539___ = new_new_new_ys__n121___ ? new_new_new_ys__n538___ : new_new_new_ys__n449___;
  assign new_new_new_ys__n540___ = ~new_new_new_ys__n123___;
  assign new_new_new_ys__n541___ = new_new_new_ys__n52___ ? new_new_new_ys__n540___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n542___ = new_new_new_ys__n36___ ? new_new_new_ys__n541___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n543___ = ~new_new_new_ys__n36___;
  assign new_new_new_ys__n544___ = new_new_new_ys__n13___ ? new_new_new_ys__n813___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n545___ = new_new_new_ys__n544___ ? new_new_new_ys__n543___ : new_new_new_ys__n542___;
  assign new_new_new_ys__n546___ = new_new_new_ys__n523___ ? new_new_new_ys__n1070___ : new_new_new_ys__n1068___;
  assign new_new_new_ys__n547___ = new_new_new_ys__n546___ ? new_new_new_ys__n545___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n548___ = new_new_new_ys__n203___ ? new_new_new_ys__n1074___ : new_new_new_ys__n1072___;
  assign new_new_new_ys__n549___ = new_new_new_ys__n548___ ? new_new_new_ys__n547___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n561___ = new_new_new_ys__n405___ ? new_new_new_ys__n11___ : new_new_new_ys__n47___;
  assign new_new_new_ys__n562___ = new_new_new_ys__n523___ ? new_new_new_ys__n605___ : new_new_new_ys__n604___;
  assign new_new_new_ys__n563___ = new_new_new_ys__n405___ ? new_new_new_ys__n11___ : new_new_new_ys__n562___;
  assign new_new_new_ys__n564___ = ys__n50 ? new_new_new_ys__n594___ : new_new_new_ys__n593___;
  assign new_new_new_ys__n565___ = new_new_new_ys__n564___ ? new_new_new_ys__n47___ : new_new_new_ys__n561___;
  assign new_new_new_ys__n566___ = new_new_new_ys__n564___ ? new_new_new_ys__n562___ : new_new_new_ys__n563___;
  assign new_new_new_ys__n567___ = new_new_new_ys__n564___ ? new_new_new_ys__n15___ : new_new_new_ys__n194___;
  assign new_new_new_ys__n568___ = ys__n65 ? new_new_new_ys__n582___ : new_new_new_ys__n580___;
  assign new_new_new_ys__n569___ = new_new_new_ys__n568___ ? new_new_new_ys__n567___ : new_new_new_ys__n565___;
  assign new_new_new_ys__n570___ = new_new_new_ys__n568___ ? new_new_new_ys__n567___ : new_new_new_ys__n566___;
  assign new_new_new_ys__n571___ = new_ys__n136_ ? new_new_new_ys__n252___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n572___ = new_ys__n136_ ? new_new_new_ys__n15___ : ys__n77;
  assign new_new_new_ys__n573___ = ys__n74 ? new_new_new_ys__n572___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n574___ = new_ys__n136_ ? ys__n77 : new_new_new_ys__n15___;
  assign new_new_new_ys__n575___ = ys__n74 ? new_new_new_ys__n15___ : new_new_new_ys__n574___;
  assign new_new_new_ys__n576___ = ys__n74 ? new_new_new_ys__n571___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n577___ = ys__n50 ? new_new_new_ys__n15___ : new_new_new_ys__n573___;
  assign new_new_new_ys__n578___ = ys__n50 ? new_new_new_ys__n15___ : new_new_new_ys__n575___;
  assign new_new_new_ys__n579___ = ys__n50 ? new_new_new_ys__n15___ : new_new_new_ys__n576___;
  assign new_new_new_ys__n580___ = ys__n45 ? new_new_new_ys__n578___ : new_new_new_ys__n577___;
  assign new_new_new_ys__n581___ = ~ys__n50;
  assign new_new_new_ys__n582___ = ys__n45 ? new_new_new_ys__n581___ : new_new_new_ys__n579___;
  assign new_new_new_ys__n583___ = ys__n27 ? ys__n30 : new_new_new_ys__n15___;
  assign new_new_new_ys__n584___ = new_new_new_ys__n470___ ? new_new_new_ys__n583___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n585___ = new_new_new_ys__n205___ ? new_new_new_ys__n11___ : new_new_new_ys__n584___;
  assign new_new_new_ys__n586___ = ys__n65 ? new_new_new_ys__n15___ : ys__n45;
  assign new_new_new_ys__n587___ = ys__n65 ? new_new_new_ys__n366___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n588___ = ys__n77 ? new_new_new_ys__n586___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n589___ = ys__n77 ? new_new_new_ys__n15___ : new_new_new_ys__n586___;
  assign new_new_new_ys__n590___ = ys__n77 ? new_new_new_ys__n587___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n591___ = ys__n74 ? new_new_new_ys__n588___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n592___ = ys__n74 ? new_new_new_ys__n590___ : new_new_new_ys__n589___;
  assign new_new_new_ys__n593___ = new_ys__n136_ ? new_new_new_ys__n15___ : new_new_new_ys__n591___;
  assign new_new_new_ys__n594___ = new_ys__n136_ ? new_new_new_ys__n592___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n595___ = new_new_new_ys__n250___ ? new_new_new_ys__n2946___ : new_new_new_ys__n2945___;
  assign new_new_new_ys__n596___ = new_new_new_ys__n179___ ? new_new_new_ys__n595___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n597___ = new_new_new_ys__n884___ ? new_new_new_ys__n883___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n598___ = new_new_new_ys__n597___ ? new_new_new_ys__n596___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n599___ = new_new_new_ys__n757___ ? new_new_new_ys__n756___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n600___ = new_new_new_ys__n599___ ? new_new_new_ys__n598___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n601___ = ys__n119 ? new_new_new_ys__n2967___ : new_new_new_ys__n2966___;
  assign new_new_new_ys__n602___ = new_new_new_ys__n601___ ? new_new_new_ys__n600___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n603___ = new_new_new_ys__n203___ ? new_new_new_ys__n3043___ : new_new_new_ys__n871___;
  assign new_new_new_ys__n604___ = new_new_new_ys__n470___ ? new_new_new_ys__n44___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n605___ = new_new_new_ys__n452___ ? new_new_new_ys__n11___ : new_new_new_ys__n604___;
  assign new_new_new_ys__n606___ = ys__n27 ? new_new_new_ys__n2106___ : new_new_new_ys__n2105___;
  assign new_new_new_ys__n607___ = new_new_new_ys__n606___ ? new_new_new_ys__n15___ : new_new_new_ys__n114___;
  assign new_new_new_ys__n608___ = new_new_new_ys__n606___ ? new_new_new_ys__n15___ : new_new_new_ys__n462___;
  assign new_new_new_ys__n609___ = ys__n30 ? new_new_new_ys__n608___ : new_new_new_ys__n607___;
  assign new_new_new_ys__n610___ = new_new_new_ys__n521___ ? new_new_new_ys__n2108___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n611___ = new_new_new_ys__n610___ ? new_new_new_ys__n11___ : new_new_new_ys__n609___;
  assign new_new_new_ys__n612___ = new_new_new_ys__n31___ ? new_new_new_ys__n611___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n613___ = new_new_new_ys__n149___ ? ys__n74 : new_new_new_ys__n15___;
  assign new_new_new_ys__n614___ = ys__n119 ? new_new_new_ys__n2178___ : new_new_new_ys__n2177___;
  assign new_new_new_ys__n615___ = new_new_new_ys__n614___ ? new_new_new_ys__n15___ : new_new_new_ys__n613___;
  assign new_new_new_ys__n616___ = new_new_new_ys__n2158___ ? new_new_new_ys__n11___ : new_new_new_ys__n2157___;
  assign new_new_new_ys__n617___ = new_new_new_ys__n616___ ? new_new_new_ys__n11___ : new_new_new_ys__n615___;
  assign new_new_new_ys__n618___ = new_new_new_ys__n273___ ? new_new_new_ys__n617___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n619___ = new_new_new_ys__n612___ ? new_new_new_ys__n618___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n642___ = ys__n17 ? new_new_new_ys__n700___ : new_new_new_ys__n699___;
  assign new_new_new_ys__n643___ = new_new_new_ys__n642___ ? new_new_new_ys__n15___ : new_new_new_ys__n404___;
  assign new_new_new_ys__n644___ = ~new_new_new_ys__n642___;
  assign new_new_new_ys__n645___ = ys__n17 ? new_new_new_ys__n642___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n646___ = ys__n17 ? new_new_new_ys__n15___ : new_new_new_ys__n642___;
  assign new_new_new_ys__n647___ = ys__n17 ? new_new_new_ys__n644___ : new_new_new_ys__n643___;
  assign new_new_new_ys__n648___ = ys__n27 ? new_new_new_ys__n645___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n649___ = ys__n27 ? new_new_new_ys__n646___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n650___ = ys__n27 ? new_new_new_ys__n15___ : new_new_new_ys__n647___;
  assign new_new_new_ys__n651___ = ys__n119 ? new_new_new_ys__n648___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n652___ = ys__n119 ? new_new_new_ys__n650___ : new_new_new_ys__n649___;
  assign new_new_new_ys__n665___ = new_new_new_ys__n205___ ? new_new_new_ys__n535___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n666___ = ~new_new_new_ys__n186___;
  assign new_new_new_ys__n667___ = new_new_new_ys__n205___ ? new_new_new_ys__n666___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n668___ = ys__n65 ? new_new_new_ys__n44___ : new_new_new_ys__n665___;
  assign new_new_new_ys__n669___ = ys__n65 ? new_new_new_ys__n15___ : new_new_new_ys__n667___;
  assign new_new_new_ys__n670___ = ys__n50 ? new_new_new_ys__n669___ : new_new_new_ys__n668___;
  assign new_new_new_ys__n683___ = ~ys__n17;
  assign new_new_new_ys__n690___ = ys__n30 ? new_new_new_ys__n297___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n691___ = ys__n27 ? new_new_new_ys__n462___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n692___ = ys__n27 ? new_new_new_ys__n15___ : new_new_new_ys__n203___;
  assign new_new_new_ys__n693___ = ~new_new_new_ys__n487___;
  assign new_new_new_ys__n694___ = ys__n27 ? new_new_new_ys__n693___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n695___ = ys__n27 ? new_new_new_ys__n462___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n696___ = ys__n74 ? new_new_new_ys__n694___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n697___ = ys__n74 ? new_new_new_ys__n694___ : new_new_new_ys__n692___;
  assign new_new_new_ys__n698___ = ys__n74 ? ys__n27 : new_new_new_ys__n695___;
  assign new_new_new_ys__n699___ = ys__n77 ? new_new_new_ys__n696___ : new_new_new_ys__n691___;
  assign new_new_new_ys__n700___ = ys__n77 ? new_new_new_ys__n698___ : new_new_new_ys__n697___;
  assign new_new_new_ys__n728___ = ys__n119 ? new_new_new_ys__n15___ : new_new_new_ys__n56___;
  assign new_new_new_ys__n729___ = ys__n119 ? new_new_new_ys__n11___ : new_new_new_ys__n52___;
  assign new_new_new_ys__n730___ = ys__n74 ? new_new_new_ys__n11___ : new_new_new_ys__n729___;
  assign new_new_new_ys__n731___ = ys__n74 ? new_new_new_ys__n11___ : ys__n119;
  assign new_new_new_ys__n732___ = ys__n74 ? new_new_new_ys__n11___ : new_new_new_ys__n728___;
  assign new_new_new_ys__n733___ = ys__n119 ? new_new_new_ys__n752___ : new_new_new_ys__n252___;
  assign new_new_new_ys__n734___ = new_new_new_ys__n733___ ? new_new_new_ys__n731___ : new_new_new_ys__n730___;
  assign new_new_new_ys__n735___ = new_new_new_ys__n733___ ? new_new_new_ys__n11___ : new_new_new_ys__n732___;
  assign new_new_new_ys__n745___ = ys__n50 ? new_new_new_ys__n11___ : ys__n45;
  assign new_new_new_ys__n746___ = ys__n65 ? new_new_new_ys__n11___ : new_new_new_ys__n745___;
  assign new_new_new_ys__n747___ = ys__n65 ? new_new_new_ys__n745___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n748___ = ys__n50 ? ys__n45 : new_new_new_ys__n15___;
  assign new_new_new_ys__n749___ = ys__n65 ? new_new_new_ys__n748___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n750___ = new_ys__n136_ ? new_new_new_ys__n15___ : new_new_new_ys__n746___;
  assign new_new_new_ys__n751___ = new_ys__n136_ ? new_new_new_ys__n749___ : new_new_new_ys__n747___;
  assign new_new_new_ys__n752___ = ys__n77 ? new_new_new_ys__n751___ : new_new_new_ys__n750___;
  assign new_new_new_ys__n753___ = ys__n77 ? new_new_new_ys__n835___ : new_new_new_ys__n834___;
  assign new_new_new_ys__n754___ = new_new_new_ys__n186___ ? new_new_new_ys__n753___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n755___ = new_new_new_ys__n520___ ? new_new_new_ys__n754___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n756___ = new_new_new_ys__n88___ ? new_new_new_ys__n755___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n757___ = new_new_new_ys__n3031___ ? new_new_new_ys__n3030___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n773___ = new_ys__n136_ ? new_new_new_ys__n252___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n813___ = ys__n17 ? new_new_new_ys__n1363___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n826___ = ys__n50 ? new_new_new_ys__n15___ : new_new_new_ys__n366___;
  assign new_new_new_ys__n827___ = ys__n65 ? new_new_new_ys__n826___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n828___ = ys__n65 ? new_new_new_ys__n15___ : new_new_new_ys__n748___;
  assign new_new_new_ys__n829___ = ys__n65 ? new_new_new_ys__n15___ : ys__n50;
  assign new_new_new_ys__n830___ = ys__n65 ? new_new_new_ys__n15___ : new_new_new_ys__n826___;
  assign new_new_new_ys__n831___ = ys__n74 ? new_new_new_ys__n827___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n832___ = ys__n74 ? new_new_new_ys__n829___ : new_new_new_ys__n828___;
  assign new_new_new_ys__n833___ = ys__n74 ? new_new_new_ys__n15___ : new_new_new_ys__n830___;
  assign new_new_new_ys__n834___ = new_ys__n136_ ? new_new_new_ys__n15___ : new_new_new_ys__n831___;
  assign new_new_new_ys__n835___ = new_ys__n136_ ? new_new_new_ys__n833___ : new_new_new_ys__n832___;
  assign new_new_new_ys__n871___ = new_new_new_ys__n250___ ? new_new_new_ys__n875___ : new_new_new_ys__n873___;
  assign new_new_new_ys__n872___ = new_new_new_ys__n71___ ? new_new_new_ys__n140___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n873___ = new_new_new_ys__n54___ ? new_new_new_ys__n872___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n874___ = new_new_new_ys__n190___ ? new_new_new_ys__n11___ : new_new_new_ys__n873___;
  assign new_new_new_ys__n875___ = new_new_new_ys__n13___ ? new_new_new_ys__n874___ : new_new_new_ys__n873___;
  assign new_new_new_ys__n876___ = new_new_new_ys__n205___ ? new_new_new_ys__n1986___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n877___ = ~new_new_new_ys__n876___;
  assign new_new_new_ys__n878___ = ys__n119 ? new_new_new_ys__n877___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n879___ = ys__n45 ? new_new_new_ys__n878___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n880___ = new_new_new_ys__n149___ ? new_new_new_ys__n2976___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n881___ = new_new_new_ys__n880___ ? new_new_new_ys__n11___ : new_new_new_ys__n879___;
  assign new_new_new_ys__n882___ = new_new_new_ys__n126___ ? new_new_new_ys__n2722___ : new_new_new_ys__n2720___;
  assign new_new_new_ys__n883___ = new_new_new_ys__n882___ ? new_new_new_ys__n881___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n884___ = new_new_new_ys__n487___ ? new_new_new_ys__n3000___ : new_new_new_ys__n2999___;
  assign new_new_new_ys__n902___ = new_new_new_ys__n196___ ? new_new_new_ys__n150___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n903___ = new_new_new_ys__n476___ ? new_new_new_ys__n11___ : new_new_new_ys__n902___;
  assign new_new_new_ys__n1039___ = ys__n30 ? new_new_new_ys__n581___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1040___ = ys__n30 ? ys__n50 : new_new_new_ys__n15___;
  assign new_new_new_ys__n1041___ = ys__n30 ? new_new_new_ys__n15___ : ys__n50;
  assign new_new_new_ys__n1042___ = ys__n17 ? new_new_new_ys__n15___ : new_new_new_ys__n1041___;
  assign new_new_new_ys__n1043___ = ys__n17 ? new_new_new_ys__n1039___ : new_new_new_ys__n581___;
  assign new_new_new_ys__n1044___ = ys__n17 ? new_new_new_ys__n1040___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1045___ = ys__n17 ? new_new_new_ys__n1041___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1046___ = ys__n27 ? new_new_new_ys__n1042___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1047___ = ys__n27 ? new_new_new_ys__n1043___ : new_new_new_ys__n581___;
  assign new_new_new_ys__n1048___ = ys__n27 ? new_new_new_ys__n1045___ : new_new_new_ys__n1044___;
  assign new_new_new_ys__n1049___ = ys__n65 ? new_new_new_ys__n1047___ : new_new_new_ys__n1046___;
  assign new_new_new_ys__n1050___ = ys__n65 ? new_new_new_ys__n15___ : new_new_new_ys__n1048___;
  assign new_new_new_ys__n1051___ = ys__n45 ? new_new_new_ys__n1050___ : new_new_new_ys__n1049___;
  assign new_new_new_ys__n1052___ = new_new_new_ys__n1051___ ? new_new_new_ys__n15___ : new_new_new_ys__n543___;
  assign new_new_new_ys__n1053___ = new_new_new_ys__n1051___ ? new_new_new_ys__n15___ : new_new_new_ys__n539___;
  assign new_new_new_ys__n1054___ = ys__n50 ? new_new_new_ys__n1053___ : new_new_new_ys__n1052___;
  assign new_new_new_ys__n1064___ = ys__n74 ? new_new_new_ys__n11___ : new_new_new_ys__n8___;
  assign new_new_new_ys__n1067___ = new_new_new_ys__n121___ ? new_new_new_ys__n19___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1068___ = new_new_new_ys__n40___ ? new_new_new_ys__n1067___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1069___ = new_new_new_ys__n487___ ? new_new_new_ys__n11___ : new_new_new_ys__n1068___;
  assign new_new_new_ys__n1070___ = new_new_new_ys__n68___ ? new_new_new_ys__n1069___ : new_new_new_ys__n1068___;
  assign new_new_new_ys__n1071___ = new_new_new_ys__n54___ ? new_new_new_ys__n319___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1072___ = new_new_new_ys__n161___ ? new_new_new_ys__n1071___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1073___ = new_new_new_ys__n488___ ? new_new_new_ys__n11___ : new_new_new_ys__n1072___;
  assign new_new_new_ys__n1074___ = new_new_new_ys__n452___ ? new_new_new_ys__n1073___ : new_new_new_ys__n1072___;
  assign new_new_new_ys__n1148___ = ys__n65 ? new_new_new_ys__n540___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1149___ = ys__n65 ? new_new_new_ys__n123___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1150___ = new_new_new_ys__n470___ ? new_new_new_ys__n73___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1151___ = new_new_new_ys__n470___ ? new_new_new_ys__n1148___ : ys__n65;
  assign new_new_new_ys__n1152___ = new_new_new_ys__n470___ ? ys__n65 : new_new_new_ys__n1148___;
  assign new_new_new_ys__n1153___ = new_new_new_ys__n470___ ? new_new_new_ys__n540___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1154___ = new_new_new_ys__n470___ ? new_new_new_ys__n15___ : new_new_new_ys__n1149___;
  assign new_new_new_ys__n1155___ = new_new_new_ys__n670___ ? new_new_new_ys__n1151___ : new_new_new_ys__n1150___;
  assign new_new_new_ys__n1156___ = new_new_new_ys__n670___ ? new_new_new_ys__n1153___ : new_new_new_ys__n1152___;
  assign new_new_new_ys__n1157___ = new_new_new_ys__n670___ ? new_new_new_ys__n15___ : new_new_new_ys__n1154___;
  assign new_new_new_ys__n1158___ = ys__n45 ? new_new_new_ys__n1155___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1159___ = ys__n45 ? new_new_new_ys__n1157___ : new_new_new_ys__n1156___;
  assign new_new_new_ys__n1161___ = ~new_new_new_ys__n470___;
  assign new_new_new_ys__n1171___ = ys__n119 ? new_new_new_ys__n185___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1172___ = ys__n119 ? new_new_new_ys__n15___ : new_new_new_ys__n140___;
  assign new_new_new_ys__n1173___ = ys__n77 ? new_new_new_ys__n1171___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1174___ = ys__n77 ? new_new_new_ys__n1172___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1175___ = new_new_new_ys__n33___ ? new_new_new_ys__n1173___ : ys__n77;
  assign new_new_new_ys__n1176___ = new_new_new_ys__n33___ ? new_new_new_ys__n1174___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1177___ = new_ys__n136_ ? new_new_new_ys__n1176___ : new_new_new_ys__n1175___;
  assign new_new_new_ys__n1184___ = new_new_new_ys__n196___ ? new_new_new_ys__n148___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1197___ = ~new_new_new_ys__n250___;
  assign new_new_new_ys__n1324___ = ys__n27 ? new_new_new_ys__n337___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1363___ = ys__n27 ? new_new_new_ys__n11___ : new_new_new_ys__n337___;
  assign new_new_new_ys__n1364___ = ys__n45 ? new_new_new_ys__n581___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1403___ = ys__n77 ? new_new_new_ys__n76___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1406___ = new_new_new_ys__n452___ ? new_new_new_ys__n537___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1628___ = ys__n65 ? new_new_new_ys__n11___ : new_new_new_ys__n581___;
  assign new_new_new_ys__n1630___ = ys__n30 ? ys__n17 : new_new_new_ys__n11___;
  assign new_new_new_ys__n1643___ = new_new_new_ys__n203___ ? new_new_new_ys__n1161___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1644___ = new_new_new_ys__n98___ ? new_new_new_ys__n11___ : new_new_new_ys__n1643___;
  assign new_new_new_ys__n1645___ = new_new_new_ys__n161___ ? new_new_new_ys__n1644___ : new_new_new_ys__n1643___;
  assign new_new_new_ys__n1646___ = new_new_new_ys__n179___ ? new_new_new_ys__n1663___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1647___ = ~new_new_new_ys__n1646___;
  assign new_new_new_ys__n1648___ = new_new_new_ys__n1646___ ? new_new_new_ys__n11___ : new_new_new_ys__n1645___;
  assign new_new_new_ys__n1663___ = new_new_new_ys__n121___ ? new_new_new_ys__n535___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1672___ = new_new_new_ys__n161___ ? new_new_new_ys__n123___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1709___ = new_new_new_ys__n124___ ? new_new_new_ys__n179___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1759___ = new_new_new_ys__n52___ ? new_new_new_ys__n521___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1760___ = new_new_new_ys__n221___ ? new_new_new_ys__n11___ : new_new_new_ys__n203___;
  assign new_new_new_ys__n1761___ = new_new_new_ys__n221___ ? new_new_new_ys__n11___ : new_new_new_ys__n1759___;
  assign new_new_new_ys__n1762___ = new_new_new_ys__n71___ ? new_new_new_ys__n396___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1786___ = new_new_new_ys__n149___ ? new_new_new_ys__n452___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1788___ = ys__n119 ? new_new_new_ys__n521___ : new_new_new_ys__n1786___;
  assign new_new_new_ys__n1798___ = ~new_new_new_ys__n196___;
  assign new_new_new_ys__n1817___ = new_ys__n136_ ? ys__n74 : new_new_new_ys__n11___;
  assign new_new_new_ys__n1980___ = ys__n65 ? ys__n30 : new_new_new_ys__n11___;
  assign new_new_new_ys__n1981___ = ys__n65 ? new_new_new_ys__n11___ : new_new_new_ys__n337___;
  assign new_new_new_ys__n1982___ = ys__n17 ? new_new_new_ys__n11___ : new_new_new_ys__n1980___;
  assign new_new_new_ys__n1983___ = ys__n17 ? new_new_new_ys__n1981___ : new_new_new_ys__n1980___;
  assign new_new_new_ys__n1984___ = ys__n50 ? new_new_new_ys__n11___ : new_new_new_ys__n1982___;
  assign new_new_new_ys__n1985___ = ys__n50 ? new_new_new_ys__n1983___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n1986___ = ys__n27 ? new_new_new_ys__n1985___ : new_new_new_ys__n1984___;
  assign new_new_new_ys__n1991___ = ys__n74 ? new_new_new_ys__n73___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1992___ = ys__n74 ? new_new_new_ys__n15___ : ys__n65;
  assign new_new_new_ys__n1993___ = new_ys__n136_ ? new_new_new_ys__n1991___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1994___ = new_ys__n136_ ? new_new_new_ys__n1992___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1995___ = new_ys__n136_ ? new_new_new_ys__n15___ : new_new_new_ys__n1992___;
  assign new_new_new_ys__n1996___ = ys__n45 ? new_new_new_ys__n15___ : new_new_new_ys__n1993___;
  assign new_new_new_ys__n1997___ = ys__n45 ? new_new_new_ys__n15___ : new_new_new_ys__n1994___;
  assign new_new_new_ys__n1998___ = ys__n45 ? new_new_new_ys__n1995___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n1999___ = ys__n77 ? new_new_new_ys__n15___ : new_new_new_ys__n1996___;
  assign new_new_new_ys__n2000___ = ys__n77 ? new_new_new_ys__n1998___ : new_new_new_ys__n1997___;
  assign new_new_new_ys__n2009___ = new_new_new_ys__n487___ ? new_new_new_ys__n1184___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2010___ = new_new_new_ys__n56___ ? new_new_new_ys__n11___ : new_new_new_ys__n2009___;
  assign new_new_new_ys__n2011___ = new_new_new_ys__n100___ ? new_new_new_ys__n2010___ : new_new_new_ys__n2009___;
  assign new_new_new_ys__n2029___ = ys__n77 ? new_new_new_ys__n319___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2030___ = new_new_new_ys__n71___ ? new_new_new_ys__n11___ : new_new_new_ys__n2029___;
  assign new_new_new_ys__n2031___ = new_new_new_ys__n549___ ? new_new_new_ys__n2030___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2032___ = new_new_new_ys__n261___ ? new_new_new_ys__n549___ : new_new_new_ys__n2031___;
  assign new_new_new_ys__n2033___ = new_ys__n136_ ? new_new_new_ys__n2032___ : new_new_new_ys__n549___;
  assign new_new_new_ys__n2037___ = ys__n17 ? new_new_new_ys__n8___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2038___ = ys__n17 ? new_new_new_ys__n11___ : new_ys__n136_;
  assign new_new_new_ys__n2039___ = ys__n17 ? new_new_new_ys__n15___ : new_ys__n136_;
  assign new_new_new_ys__n2040___ = ys__n17 ? new_new_new_ys__n15___ : new_new_new_ys__n8___;
  assign new_new_new_ys__n2041___ = ys__n50 ? new_new_new_ys__n15___ : new_new_new_ys__n2040___;
  assign new_new_new_ys__n2042___ = ys__n50 ? new_new_new_ys__n8___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2043___ = ys__n17 ? new_ys__n136_ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2044___ = ys__n50 ? new_new_new_ys__n2043___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2045___ = ys__n50 ? new_new_new_ys__n11___ : new_new_new_ys__n2037___;
  assign new_new_new_ys__n2046___ = ys__n50 ? new_new_new_ys__n11___ : new_new_new_ys__n2038___;
  assign new_new_new_ys__n2047___ = ys__n50 ? new_new_new_ys__n15___ : new_new_new_ys__n2039___;
  assign new_new_new_ys__n2048___ = ys__n50 ? new_new_new_ys__n2040___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2049___ = ys__n50 ? new_new_new_ys__n15___ : new_new_new_ys__n2043___;
  assign new_new_new_ys__n2050___ = ys__n119 ? new_new_new_ys__n2042___ : new_new_new_ys__n2041___;
  assign new_new_new_ys__n2051___ = ys__n119 ? new_new_new_ys__n2045___ : new_new_new_ys__n2044___;
  assign new_new_new_ys__n2052___ = ys__n119 ? new_new_new_ys__n2047___ : new_new_new_ys__n2046___;
  assign new_new_new_ys__n2053___ = ys__n119 ? new_new_new_ys__n2049___ : new_new_new_ys__n2048___;
  assign new_new_new_ys__n2054___ = ys__n45 ? new_new_new_ys__n2051___ : new_new_new_ys__n2050___;
  assign new_new_new_ys__n2055___ = ys__n45 ? new_new_new_ys__n2053___ : new_new_new_ys__n2052___;
  assign new_new_new_ys__n2056___ = ys__n65 ? new_new_new_ys__n2055___ : new_new_new_ys__n2054___;
  assign new_new_new_ys__n2100___ = ys__n30 ? new_new_new_ys__n63___ : new_new_new_ys__n398___;
  assign new_new_new_ys__n2101___ = ys__n30 ? new_new_new_ys__n15___ : new_new_new_ys__n398___;
  assign new_new_new_ys__n2102___ = ys__n119 ? new_new_new_ys__n15___ : new_new_new_ys__n64___;
  assign new_new_new_ys__n2103___ = ys__n119 ? new_new_new_ys__n15___ : new_new_new_ys__n2100___;
  assign new_new_new_ys__n2104___ = ys__n119 ? new_new_new_ys__n2101___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2105___ = ys__n17 ? new_new_new_ys__n2102___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2106___ = ys__n17 ? new_new_new_ys__n2104___ : new_new_new_ys__n2103___;
  assign new_new_new_ys__n2107___ = new_new_new_ys__n414___ ? new_new_new_ys__n203___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2108___ = ys__n119 ? new_new_new_ys__n1709___ : new_new_new_ys__n2107___;
  assign new_new_new_ys__n2109___ = ys__n119 ? new_new_new_ys__n15___ : new_new_new_ys__n185___;
  assign new_new_new_ys__n2110___ = new_new_new_ys__n196___ ? new_new_new_ys__n132___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2111___ = new_new_new_ys__n196___ ? new_new_new_ys__n2109___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2112___ = ys__n30 ? new_new_new_ys__n2110___ : new_new_new_ys__n693___;
  assign new_new_new_ys__n2113___ = ys__n30 ? new_new_new_ys__n15___ : new_new_new_ys__n2111___;
  assign new_new_new_ys__n2114___ = ys__n65 ? new_new_new_ys__n2166___ : new_new_new_ys__n2165___;
  assign new_new_new_ys__n2115___ = new_new_new_ys__n2114___ ? new_new_new_ys__n11___ : ys__n27;
  assign new_new_new_ys__n2116___ = ~new_new_new_ys__n2114___;
  assign new_new_new_ys__n2117___ = new_new_new_ys__n2114___ ? new_new_new_ys__n11___ : new_new_new_ys__n297___;
  assign new_new_new_ys__n2118___ = ys__n119 ? new_new_new_ys__n11___ : new_new_new_ys__n2115___;
  assign new_new_new_ys__n2119___ = ys__n119 ? new_new_new_ys__n2116___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2120___ = ys__n119 ? new_new_new_ys__n11___ : new_new_new_ys__n2117___;
  assign new_new_new_ys__n2121___ = ys__n45 ? new_new_new_ys__n11___ : new_new_new_ys__n2118___;
  assign new_new_new_ys__n2122___ = ys__n45 ? new_new_new_ys__n2120___ : new_new_new_ys__n2119___;
  assign new_new_new_ys__n2123___ = ys__n17 ? new_new_new_ys__n2122___ : new_new_new_ys__n2121___;
  assign new_new_new_ys__n2124___ = new_new_new_ys__n7___ ? ys__n119 : new_new_new_ys__n15___;
  assign new_new_new_ys__n2125___ = ys__n77 ? new_new_new_ys__n11___ : new_new_new_ys__n2124___;
  assign new_new_new_ys__n2126___ = new_new_new_ys__n59___ ? new_new_new_ys__n2125___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2154___ = new_new_new_ys__n203___ ? new_new_new_ys__n405___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2155___ = ys__n77 ? new_new_new_ys__n15___ : new_new_new_ys__n2154___;
  assign new_new_new_ys__n2156___ = new_new_new_ys__n1672___ ? new_new_new_ys__n15___ : new_new_new_ys__n2155___;
  assign new_new_new_ys__n2157___ = new_ys__n136_ ? new_new_new_ys__n11___ : new_new_new_ys__n2156___;
  assign new_new_new_ys__n2158___ = ys__n74 ? new_new_new_ys__n2205___ : new_new_new_ys__n2204___;
  assign new_new_new_ys__n2159___ = new_new_new_ys__n331___ ? new_new_new_ys__n252___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2160___ = new_new_new_ys__n414___ ? new_new_new_ys__n2159___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2161___ = ys__n30 ? new_new_new_ys__n15___ : new_new_new_ys__n132___;
  assign new_new_new_ys__n2162___ = ys__n30 ? new_new_new_ys__n15___ : ys__n119;
  assign new_new_new_ys__n2163___ = ys__n27 ? new_new_new_ys__n15___ : new_new_new_ys__n2161___;
  assign new_new_new_ys__n2164___ = ys__n27 ? new_new_new_ys__n337___ : new_new_new_ys__n2162___;
  assign new_new_new_ys__n2165___ = ys__n50 ? new_new_new_ys__n2163___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2166___ = ys__n50 ? new_new_new_ys__n15___ : new_new_new_ys__n2164___;
  assign new_new_new_ys__n2175___ = ys__n77 ? new_new_new_ys__n15___ : new_new_new_ys__n356___;
  assign new_new_new_ys__n2176___ = ys__n77 ? new_new_new_ys__n389___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2177___ = new_ys__n136_ ? new_new_new_ys__n389___ : new_new_new_ys__n2175___;
  assign new_new_new_ys__n2178___ = new_ys__n136_ ? new_new_new_ys__n15___ : new_new_new_ys__n2176___;
  assign new_new_new_ys__n2179___ = ys__n50 ? new_new_new_ys__n15___ : ys__n17;
  assign new_new_new_ys__n2180___ = ys__n50 ? ys__n17 : new_new_new_ys__n11___;
  assign new_new_new_ys__n2181___ = ys__n50 ? new_new_new_ys__n11___ : ys__n17;
  assign new_new_new_ys__n2182___ = ys__n119 ? new_new_new_ys__n2179___ : ys__n17;
  assign new_new_new_ys__n2183___ = ys__n119 ? new_new_new_ys__n2180___ : ys__n17;
  assign new_new_new_ys__n2184___ = ys__n119 ? new_new_new_ys__n2181___ : new_new_new_ys__n581___;
  assign new_new_new_ys__n2185___ = ys__n119 ? ys__n17 : new_new_new_ys__n2180___;
  assign new_new_new_ys__n2186___ = ys__n65 ? new_new_new_ys__n2182___ : new_new_new_ys__n2185___;
  assign new_new_new_ys__n2187___ = ys__n65 ? new_new_new_ys__n2183___ : ys__n17;
  assign new_new_new_ys__n2188___ = ys__n65 ? new_new_new_ys__n2184___ : ys__n17;
  assign new_new_new_ys__n2189___ = ys__n65 ? ys__n17 : new_new_new_ys__n2185___;
  assign new_new_new_ys__n2190___ = ys__n27 ? new_new_new_ys__n2187___ : new_new_new_ys__n2186___;
  assign new_new_new_ys__n2191___ = ys__n27 ? new_new_new_ys__n2189___ : new_new_new_ys__n2188___;
  assign new_new_new_ys__n2192___ = ys__n30 ? new_new_new_ys__n2191___ : new_new_new_ys__n2190___;
  assign new_new_new_ys__n2193___ = ys__n45 ? new_new_new_ys__n252___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2194___ = ys__n45 ? ys__n77 : new_new_new_ys__n11___;
  assign new_new_new_ys__n2195___ = ys__n45 ? new_new_new_ys__n11___ : ys__n77;
  assign new_new_new_ys__n2196___ = new_new_new_ys__n2192___ ? new_new_new_ys__n252___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2197___ = new_new_new_ys__n2192___ ? new_new_new_ys__n15___ : new_new_new_ys__n2193___;
  assign new_new_new_ys__n2198___ = new_new_new_ys__n2192___ ? new_new_new_ys__n2194___ : ys__n77;
  assign new_new_new_ys__n2199___ = new_new_new_ys__n2192___ ? ys__n77 : new_new_new_ys__n2195___;
  assign new_new_new_ys__n2200___ = ys__n119 ? new_new_new_ys__n2196___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2201___ = ys__n119 ? new_new_new_ys__n2197___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2202___ = ys__n119 ? ys__n77 : new_new_new_ys__n2198___;
  assign new_new_new_ys__n2203___ = ys__n119 ? ys__n77 : new_new_new_ys__n2199___;
  assign new_new_new_ys__n2204___ = ys__n17 ? new_new_new_ys__n2201___ : new_new_new_ys__n2200___;
  assign new_new_new_ys__n2205___ = ys__n17 ? new_new_new_ys__n2203___ : new_new_new_ys__n2202___;
  assign new_new_new_ys__n2206___ = ys__n119 ? new_new_new_ys__n461___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2375___ = new_new_new_ys__n488___ ? new_new_new_ys__n114___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2376___ = new_new_new_ys__n71___ ? new_new_new_ys__n2869___ : new_new_new_ys__n2867___;
  assign new_new_new_ys__n2377___ = new_new_new_ys__n2376___ ? new_new_new_ys__n2375___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2378___ = ys__n77 ? new_new_new_ys__n11___ : new_new_new_ys__n2376___;
  assign new_new_new_ys__n2379___ = ys__n77 ? new_new_new_ys__n2376___ : new_new_new_ys__n2377___;
  assign new_new_new_ys__n2380___ = new_new_new_ys__n1177___ ? new_new_new_ys__n2379___ : new_new_new_ys__n2378___;
  assign new_new_new_ys__n2381___ = ys__n30 ? new_new_new_ys__n414___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2382___ = new_new_new_ys__n126___ ? new_new_new_ys__n2381___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2383___ = new_new_new_ys__n126___ ? ys__n30 : new_new_new_ys__n15___;
  assign new_new_new_ys__n2384___ = ys__n50 ? new_new_new_ys__n1197___ : new_new_new_ys__n250___;
  assign new_new_new_ys__n2385___ = ys__n50 ? new_new_new_ys__n2383___ : new_new_new_ys__n2382___;
  assign new_new_new_ys__n2386___ = ys__n65 ? new_new_new_ys__n2385___ : new_new_new_ys__n2384___;
  assign new_new_new_ys__n2390___ = new_new_new_ys__n2827___ ? new_new_new_ys__n2835___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2393___ = new_new_new_ys__n59___ ? new_new_new_ys__n12___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2394___ = ys__n50 ? new_new_new_ys__n455___ : new_new_new_ys__n2393___;
  assign new_new_new_ys__n2395___ = ys__n50 ? new_new_new_ys__n15___ : new_new_new_ys__n455___;
  assign new_new_new_ys__n2396___ = ys__n65 ? new_new_new_ys__n581___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2397___ = ys__n65 ? new_new_new_ys__n15___ : new_new_new_ys__n2394___;
  assign new_new_new_ys__n2398___ = ys__n65 ? ys__n50 : new_new_new_ys__n2395___;
  assign new_new_new_ys__n2399___ = new_new_new_ys__n2386___ ? new_new_new_ys__n15___ : new_new_new_ys__n2396___;
  assign new_new_new_ys__n2400___ = new_new_new_ys__n2386___ ? new_new_new_ys__n2398___ : new_new_new_ys__n2397___;
  assign new_new_new_ys__n2423___ = ys__n74 ? new_new_new_ys__n11___ : new_new_new_ys__n252___;
  assign new_new_new_ys__n2518___ = ys__n27 ? new_new_new_ys__n683___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2552___ = new_new_new_ys__n161___ ? new_new_new_ys__n1197___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2553___ = new_new_new_ys__n124___ ? new_new_new_ys__n2552___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2554___ = new_new_new_ys__n100___ ? new_new_new_ys__n11___ : new_new_new_ys__n2553___;
  assign new_new_new_ys__n2555___ = new_new_new_ys__n36___ ? new_new_new_ys__n2554___ : new_new_new_ys__n2553___;
  assign new_new_new_ys__n2568___ = ys__n65 ? new_new_new_ys__n11___ : new_new_new_ys__n366___;
  assign new_new_new_ys__n2668___ = new_new_new_ys__n149___ ? new_new_new_ys__n495___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2719___ = new_new_new_ys__n188___ ? new_new_new_ys__n140___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2720___ = new_new_new_ys__n40___ ? new_new_new_ys__n2719___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2721___ = new_new_new_ys__n33___ ? new_new_new_ys__n11___ : new_new_new_ys__n2720___;
  assign new_new_new_ys__n2722___ = new_new_new_ys__n161___ ? new_new_new_ys__n2721___ : new_new_new_ys__n2720___;
  assign new_new_new_ys__n2778___ = ys__n77 ? new_new_new_ys__n11___ : new_new_new_ys__n132___;
  assign new_new_new_ys__n2779___ = ys__n74 ? new_new_new_ys__n11___ : new_new_new_ys__n2778___;
  assign new_new_new_ys__n2788___ = ys__n45 ? new_new_new_ys__n15___ : ys__n65;
  assign new_new_new_ys__n2791___ = ys__n45 ? new_new_new_ys__n73___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2821___ = new_new_new_ys__n161___ ? new_new_new_ys__n319___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2822___ = ys__n77 ? new_new_new_ys__n15___ : new_new_new_ys__n2821___;
  assign new_new_new_ys__n2823___ = ys__n77 ? new_new_new_ys__n410___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2824___ = ys__n77 ? new_new_new_ys__n15___ : new_new_new_ys__n410___;
  assign new_new_new_ys__n2825___ = new_ys__n136_ ? new_new_new_ys__n15___ : new_new_new_ys__n2822___;
  assign new_new_new_ys__n2826___ = new_ys__n136_ ? new_new_new_ys__n2824___ : new_new_new_ys__n2823___;
  assign new_new_new_ys__n2827___ = ys__n74 ? new_new_new_ys__n2826___ : new_new_new_ys__n2825___;
  assign new_new_new_ys__n2828___ = ys__n17 ? new_new_new_ys__n11___ : new_new_new_ys__n2884___;
  assign new_new_new_ys__n2829___ = ~new_new_new_ys__n2828___;
  assign new_new_new_ys__n2830___ = ys__n74 ? new_new_new_ys__n2906___ : new_new_new_ys__n2905___;
  assign new_new_new_ys__n2831___ = ys__n30 ? new_new_new_ys__n2830___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2832___ = ys__n30 ? new_new_new_ys__n2829___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2833___ = ys__n27 ? new_new_new_ys__n2832___ : new_new_new_ys__n2831___;
  assign new_new_new_ys__n2834___ = new_new_new_ys__n331___ ? new_new_new_ys__n2923___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2835___ = new_new_new_ys__n2834___ ? new_new_new_ys__n11___ : new_new_new_ys__n2833___;
  assign new_new_new_ys__n2836___ = ~new_new_new_ys__n2390___;
  assign new_new_new_ys__n2837___ = new_new_new_ys__n2033___ ? new_new_new_ys__n2836___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2838___ = new_new_new_ys__n619___ ? new_new_new_ys__n2837___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2839___ = new_new_new_ys__n432___ ? new_new_new_ys__n2838___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2840___ = new_new_new_ys__n43___ ? new_new_new_ys__n2839___ : new_new_new_ys__n15___;
  assign ys__n2841 = new_new_new_ys__n507___ ? new_new_new_ys__n2840___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2848___ = ys__n50 ? new_new_new_ys__n366___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2866___ = new_new_new_ys__n535___ ? new_new_new_ys__n61___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2867___ = new_new_new_ys__n203___ ? new_new_new_ys__n2866___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2868___ = new_new_new_ys__n487___ ? new_new_new_ys__n11___ : new_new_new_ys__n2867___;
  assign new_new_new_ys__n2869___ = new_new_new_ys__n196___ ? new_new_new_ys__n2868___ : new_new_new_ys__n2867___;
  assign new_new_new_ys__n2882___ = new_new_new_ys__n98___ ? new_new_new_ys__n56___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2883___ = new_new_new_ys__n179___ ? new_new_new_ys__n15___ : new_new_new_ys__n2882___;
  assign new_new_new_ys__n2884___ = new_new_new_ys__n96___ ? new_new_new_ys__n2883___ : new_new_new_ys__n2882___;
  assign new_new_new_ys__n2894___ = ys__n45 ? ys__n65 : new_new_new_ys__n15___;
  assign new_new_new_ys__n2895___ = ys__n45 ? new_new_new_ys__n73___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2896___ = ys__n45 ? new_new_new_ys__n15___ : new_new_new_ys__n73___;
  assign new_new_new_ys__n2897___ = ys__n119 ? new_new_new_ys__n15___ : new_new_new_ys__n2791___;
  assign new_new_new_ys__n2898___ = ys__n119 ? new_new_new_ys__n15___ : new_new_new_ys__n2788___;
  assign new_new_new_ys__n2899___ = ys__n119 ? new_new_new_ys__n2895___ : new_new_new_ys__n2894___;
  assign new_new_new_ys__n2900___ = ys__n119 ? new_new_new_ys__n15___ : new_new_new_ys__n2896___;
  assign new_new_new_ys__n2901___ = new_new_new_ys__n2056___ ? new_new_new_ys__n15___ : new_new_new_ys__n2897___;
  assign new_new_new_ys__n2902___ = new_new_new_ys__n2056___ ? new_new_new_ys__n15___ : new_new_new_ys__n2898___;
  assign new_new_new_ys__n2903___ = new_new_new_ys__n2056___ ? new_new_new_ys__n15___ : new_new_new_ys__n2899___;
  assign new_new_new_ys__n2904___ = new_new_new_ys__n2056___ ? new_new_new_ys__n2900___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2905___ = ys__n77 ? new_new_new_ys__n2902___ : new_new_new_ys__n2901___;
  assign new_new_new_ys__n2906___ = ys__n77 ? new_new_new_ys__n2904___ : new_new_new_ys__n2903___;
  assign new_new_new_ys__n2918___ = new_new_new_ys__n474___ ? new_new_new_ys__n15___ : new_new_new_ys__n813___;
  assign new_new_new_ys__n2919___ = new_new_new_ys__n414___ ? new_new_new_ys__n474___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2920___ = new_new_new_ys__n414___ ? new_new_new_ys__n2918___ : new_new_new_ys__n813___;
  assign new_new_new_ys__n2921___ = new_new_new_ys__n126___ ? new_new_new_ys__n414___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2922___ = new_new_new_ys__n126___ ? new_new_new_ys__n2920___ : new_new_new_ys__n2919___;
  assign new_new_new_ys__n2923___ = ys__n65 ? new_new_new_ys__n2922___ : new_new_new_ys__n2921___;
  assign new_new_new_ys__n2924___ = ys__n77 ? new_new_new_ys__n8___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2945___ = new_new_new_ys__n141___ ? new_new_new_ys__n1798___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2946___ = new_new_new_ys__n59___ ? new_new_new_ys__n11___ : new_new_new_ys__n2945___;
  assign new_new_new_ys__n2960___ = ys__n74 ? new_new_new_ys__n11___ : new_new_new_ys__n693___;
  assign new_new_new_ys__n2961___ = new_new_new_ys__n813___ ? new_new_new_ys__n2960___ : new_new_new_ys__n76___;
  assign new_new_new_ys__n2962___ = new_new_new_ys__n0___ ? new_new_new_ys__n2961___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2963___ = ys__n119 ? new_new_new_ys__n813___ : new_new_new_ys__n2962___;
  assign new_new_new_ys__n2964___ = new_new_new_ys__n121___ ? new_new_new_ys__n114___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2965___ = new_new_new_ys__n1672___ ? new_new_new_ys__n11___ : ys__n74;
  assign new_new_new_ys__n2966___ = new_new_new_ys__n2963___ ? new_new_new_ys__n15___ : new_new_new_ys__n2965___;
  assign new_new_new_ys__n2967___ = new_new_new_ys__n2963___ ? new_new_new_ys__n2964___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2972___ = new_new_new_ys__n68___ ? new_new_new_ys__n15___ : new_new_new_ys__n452___;
  assign new_new_new_ys__n2973___ = new_new_new_ys__n100___ ? new_new_new_ys__n15___ : new_new_new_ys__n2972___;
  assign new_new_new_ys__n2974___ = new_new_new_ys__n470___ ? new_new_new_ys__n100___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2975___ = new_new_new_ys__n470___ ? new_new_new_ys__n2973___ : new_new_new_ys__n2972___;
  assign new_new_new_ys__n2976___ = new_new_new_ys__n40___ ? new_new_new_ys__n2975___ : new_new_new_ys__n2974___;
  assign new_new_new_ys__n2981___ = new_new_new_ys__n179___ ? new_new_new_ys__n44___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2982___ = new_new_new_ys__n98___ ? new_new_new_ys__n2981___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2983___ = new_new_new_ys__n56___ ? new_new_new_ys__n11___ : new_new_new_ys__n2982___;
  assign new_new_new_ys__n2984___ = new_new_new_ys__n535___ ? new_new_new_ys__n2983___ : new_new_new_ys__n2982___;
  assign new_new_new_ys__n2985___ = new_new_new_ys__n521___ ? new_new_new_ys__n2984___ : new_new_new_ys__n2982___;
  assign new_new_new_ys__n2992___ = new_new_new_ys__n813___ ? new_new_new_ys__n2668___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n2993___ = new_new_new_ys__n813___ ? new_new_new_ys__n452___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2994___ = ys__n119 ? new_new_new_ys__n2993___ : new_new_new_ys__n2992___;
  assign new_new_new_ys__n2995___ = new_new_new_ys__n2985___ ? new_new_new_ys__n1762___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2996___ = ys__n119 ? new_new_new_ys__n2985___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2997___ = ys__n119 ? new_new_new_ys__n2995___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n2998___ = ys__n119 ? new_new_new_ys__n11___ : new_new_new_ys__n2995___;
  assign new_new_new_ys__n2999___ = new_new_new_ys__n2994___ ? new_new_new_ys__n2985___ : new_new_new_ys__n2996___;
  assign new_new_new_ys__n3000___ = new_new_new_ys__n2994___ ? new_new_new_ys__n2998___ : new_new_new_ys__n2997___;
  assign new_new_new_ys__n3029___ = new_new_new_ys__n124___ ? new_new_new_ys__n693___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n3030___ = new_new_new_ys__n96___ ? new_new_new_ys__n3029___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n3031___ = new_new_new_ys__n357___ ? new_new_new_ys__n3035___ : new_new_new_ys__n3033___;
  assign new_new_new_ys__n3032___ = new_new_new_ys__n405___ ? new_new_new_ys__n495___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n3033___ = new_new_new_ys__n161___ ? new_new_new_ys__n3032___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n3034___ = new_new_new_ys__n813___ ? new_new_new_ys__n11___ : new_new_new_ys__n3033___;
  assign new_new_new_ys__n3035___ = new_new_new_ys__n179___ ? new_new_new_ys__n3034___ : new_new_new_ys__n3033___;
  assign new_new_new_ys__n3040___ = new_new_new_ys__n40___ ? new_new_new_ys__n63___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n3041___ = new_new_new_ys__n124___ ? new_new_new_ys__n11___ : new_new_new_ys__n3040___;
  assign new_new_new_ys__n3042___ = new_new_new_ys__n98___ ? new_new_new_ys__n3041___ : new_new_new_ys__n3040___;
  assign new_new_new_ys__n3043___ = new_new_new_ys__n871___ ? new_new_new_ys__n3042___ : new_new_new_ys__n11___;
  assign new_new_new_ys__n3075___ = new_new_new_ys__n161___ ? new_new_new_ys__n1406___ : new_new_new_ys__n15___;
  assign new_new_new_ys__n3076___ = new_new_new_ys__n487___ ? new_new_new_ys__n11___ : new_new_new_ys__n3075___;
  assign new_new_new_ys__n3077___ = new_new_new_ys__n188___ ? new_new_new_ys__n3076___ : new_new_new_ys__n3075___;
endmodule


