library ieee;
use ieee.std_logic_1164.all;

entity top is
 port(B: in std_logic_vector(10 downto 0);
 M: out std_logic_vector(3 downto 0);
 E: out std_logic_vector(2 downto 0));
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259: std_logic;

begin

w0 <= not B(1) and B(4);
w1 <= not B(4) and not B(8);
w2 <= not w0 and not w1;
w3 <= B(0) and not w2;
w4 <= B(1) and B(4);
w5 <= not B(0) and w4;
w6 <= not w3 and not w5;
w7 <= not B(6) and not w6;
w8 <= not B(7) and w7;
w9 <= B(4) and B(8);
w10 <= not w8 and not w9;
w11 <= not B(5) and not w10;
w12 <= not B(4) and B(7);
w13 <= B(1) and not B(2);
w14 <= B(5) and not B(7);
w15 <= w13 and w14;
w16 <= not w12 and not w15;
w17 <= B(3) and not w16;
w18 <= B(4) and B(7);
w19 <= not B(3) and w18;
w20 <= not w17 and not w19;
w21 <= not B(8) and not w20;
w22 <= B(5) and B(8);
w23 <= not B(4) and w22;
w24 <= not w21 and not w23;
w25 <= not w11 and w24;
w26 <= not B(9) and not w25;
w27 <= B(4) and not B(8);
w28 <= not B(3) and w27;
w29 <= not B(4) and not B(7);
w30 <= not w28 and not w29;
w31 <= not B(2) and not w30;
w32 <= B(1) and w31;
w33 <= not B(1) and B(2);
w34 <= not B(7) and not B(8);
w35 <= w33 and w34;
w36 <= not B(9) and not w35;
w37 <= not w32 and w36;
w38 <= not B(6) and not w37;
w39 <= B(5) and w38;
w40 <= B(6) and B(9);
w41 <= not B(5) and w40;
w42 <= not w39 and not w41;
w43 <= not w26 and w42;
w44 <= not B(10) and not w43;
w45 <= not B(2) and B(3);
w46 <= B(2) and not B(3);
w47 <= not w45 and not w46;
w48 <= not B(9) and not w47;
w49 <= not B(8) and w48;
w50 <= not B(10) and not w49;
w51 <= not B(7) and not w50;
w52 <= B(9) and B(10);
w53 <= B(8) and w52;
w54 <= not w51 and not w53;
w55 <= B(6) and not w54;
w56 <= not B(6) and B(10);
w57 <= B(7) and w56;
w58 <= not w55 and not w57;
w59 <= not w44 and w58;
w60 <= not B(4) and not B(9);
w61 <= not B(2) and not B(7);
w62 <= not w60 and not w61;
w63 <= not B(1) and not w62;
w64 <= B(1) and B(2);
w65 <= B(0) and w64;
w66 <= not B(0) and not B(2);
w67 <= not w65 and not w66;
w68 <= not B(7) and not w67;
w69 <= B(4) and w68;
w70 <= B(8) and not B(9);
w71 <= not w69 and not w70;
w72 <= not w63 and w71;
w73 <= not B(6) and not w72;
w74 <= B(3) and B(4);
w75 <= B(7) and not w74;
w76 <= not B(9) and w75;
w77 <= not B(8) and w76;
w78 <= not B(7) and B(9);
w79 <= not w77 and not w78;
w80 <= not w73 and w79;
w81 <= not B(5) and not w80;
w82 <= not B(8) and not B(9);
w83 <= B(4) and w82;
w84 <= not B(6) and not B(7);
w85 <= not B(4) and w84;
w86 <= not w83 and not w85;
w87 <= B(2) and not w86;
w88 <= B(1) and w87;
w89 <= B(7) and not B(9);
w90 <= w27 and w89;
w91 <= not w88 and not w90;
w92 <= B(3) and not w91;
w93 <= B(4) and w70;
w94 <= B(7) and B(9);
w95 <= not w93 and not w94;
w96 <= B(6) and not w95;
w97 <= not w92 and not w96;
w98 <= B(5) and not w97;
w99 <= not B(4) and w70;
w100 <= not w78 and not w99;
w101 <= not B(6) and not w100;
w102 <= not w98 and not w101;
w103 <= not w81 and w102;
w104 <= not B(10) and not w103;
w105 <= B(6) and not B(9);
w106 <= not B(4) and w105;
w107 <= B(5) and not B(6);
w108 <= not B(3) and w107;
w109 <= not w106 and not w108;
w110 <= not B(2) and not w109;
w111 <= not B(1) and w107;
w112 <= not w106 and not w111;
w113 <= not B(3) and not w112;
w114 <= B(2) and B(3);
w115 <= B(4) and w105;
w116 <= w114 and w115;
w117 <= not B(10) and not w116;
w118 <= not w113 and w117;
w119 <= not w110 and w118;
w120 <= not B(7) and not w119;
w121 <= not w56 and not w120;
w122 <= not B(8) and not w121;
w123 <= B(6) and B(10);
w124 <= B(7) and w123;
w125 <= w70 and w124;
w126 <= not w122 and not w125;
w127 <= not w104 and w126;
w128 <= B(4) and not B(6);
w129 <= B(0) and not B(3);
w130 <= w128 and w129;
w131 <= not B(4) and B(5);
w132 <= B(3) and w131;
w133 <= not w130 and not w132;
w134 <= B(1) and not w133;
w135 <= not B(4) and not B(6);
w136 <= B(0) and B(1);
w137 <= B(4) and not w136;
w138 <= B(3) and w137;
w139 <= not w135 and not w138;
w140 <= not B(5) and not w139;
w141 <= not w134 and not w140;
w142 <= B(2) and not w141;
w143 <= B(3) and not B(6);
w144 <= not B(2) and w143;
w145 <= not B(3) and B(5);
w146 <= not w144 and not w145;
w147 <= B(4) and not w146;
w148 <= not w142 and not w147;
w149 <= not B(7) and not w148;
w150 <= not B(5) and B(6);
w151 <= B(2) and w150;
w152 <= not w111 and not w151;
w153 <= B(4) and not w152;
w154 <= B(3) and w153;
w155 <= B(5) and not w74;
w156 <= B(6) and w155;
w157 <= not w154 and not w156;
w158 <= not w149 and w157;
w159 <= not B(8) and not w158;
w160 <= not B(6) and B(7);
w161 <= B(3) and w160;
w162 <= B(6) and not B(7);
w163 <= not B(2) and w162;
w164 <= not w161 and not w163;
w165 <= B(5) and not w164;
w166 <= B(4) and w165;
w167 <= B(4) and B(5);
w168 <= B(7) and not w167;
w169 <= B(6) and w168;
w170 <= not w166 and not w169;
w171 <= not w159 and w170;
w172 <= not B(9) and not w171;
w173 <= B(4) and B(6);
w174 <= w14 and w173;
w175 <= not w160 and not w174;
w176 <= B(8) and not w175;
w177 <= not w172 and not w176;
w178 <= not B(10) and not w177;
w179 <= B(8) and B(10);
w180 <= not B(8) and B(9);
w181 <= B(5) and w180;
w182 <= not w179 and not w181;
w183 <= B(7) and not w182;
w184 <= B(6) and w183;
w185 <= B(5) and B(7);
w186 <= B(8) and not w185;
w187 <= not B(10) and not w186;
w188 <= B(9) and not w187;
w189 <= not w184 and not w188;
w190 <= not w178 and w189;
w191 <= B(6) and B(7);
w192 <= not B(2) and w191;
w193 <= B(5) and w9;
w194 <= w192 and w193;
w195 <= not B(5) and w1;
w196 <= w84 and w195;
w197 <= not w194 and not w196;
w198 <= not B(9) and not w197;
w199 <= not B(10) and w198;
w200 <= not B(3) and w199;
w201 <= B(5) and B(6);
w202 <= B(4) and not B(7);
w203 <= w201 and w202;
w204 <= not B(5) and not B(6);
w205 <= w136 and w204;
w206 <= not w203 and not w205;
w207 <= B(3) and not w206;
w208 <= B(2) and w207;
w209 <= not B(4) and not w162;
w210 <= not B(7) and not w107;
w211 <= not B(3) and not w210;
w212 <= B(7) and not w201;
w213 <= not B(6) and not w64;
w214 <= B(5) and w213;
w215 <= not B(9) and not w214;
w216 <= not w212 and w215;
w217 <= not w211 and w216;
w218 <= not w209 and w217;
w219 <= not w208 and w218;
w220 <= not B(8) and not w219;
w221 <= B(3) and B(8);
w222 <= not w46 and not w221;
w223 <= B(6) and not w222;
w224 <= B(5) and w223;
w225 <= B(7) and w224;
w226 <= not B(9) and w225;
w227 <= B(4) and w226;
w228 <= B(7) and w201;
w229 <= B(9) and not w228;
w230 <= not w227 and not w229;
w231 <= not w220 and w230;
w232 <= not B(10) and not w231;
w233 <= B(6) and B(8);
w234 <= w185 and w233;
w235 <= B(1) and B(3);
w236 <= B(0) and w235;
w237 <= not B(5) and not B(7);
w238 <= not B(8) and w237;
w239 <= w236 and w238;
w240 <= not w234 and not w239;
w241 <= B(2) and not w240;
w242 <= B(8) and w185;
w243 <= B(3) and B(6);
w244 <= w242 and w243;
w245 <= not w241 and not w244;
w246 <= B(4) and not w245;
w247 <= w114 and w173;
w248 <= B(5) and not w247;
w249 <= not w150 and not w248;
w250 <= not B(7) and not w249;
w251 <= not B(8) and w250;
w252 <= not B(9) and not B(10);
w253 <= not w251 and w252;
w254 <= not w246 and w253;
w255 <= B(2) and w74;
w256 <= w201 and w255;
w257 <= not B(9) and not w256;
w258 <= not B(10) and w257;
w259 <= w34 and w258;
one <= '1';
M(0) <= not w59;-- level 13
M(1) <= w127;-- level 13
M(2) <= not w190;-- level 16
M(3) <= not w200;-- level 7
E(0) <= not w232;-- level 11
E(1) <= not w254;-- level 8
E(2) <= not w259;-- level 6
end Behavioral;