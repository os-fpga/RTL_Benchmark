`ifndef _fft_w_
`define _fft_w_
`include "round32.sv"

module W_int32 #(parameter POW, W_WIDTH)(clk, k, W_Re, W_Im);
// N = 2**POW, Max POW = 10, Max W_WIDTH = 32
// File contains the rotate coefficients
// W(k, N) =  exp(-2i * pi * k / N)
// in the scale W * 2^30

   input wire clk;
   input wire [POW-2:0] k;
   output wire signed [W_WIDTH-1:0] W_Re, W_Im;

   generate
      if (POW == 1)
         begin
            localparam bit signed [31:0] W_Re_table = 32'sh40000000;
            localparam bit signed [31:0] W_Im_table = 32'sh00000000;

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_table, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_table, W_Im);
         end
      else if (POW == 2)
         begin
            reg signed [31:0] W_Re_table[2] = '{
               32'sh40000000, 32'sh00000000
            };

            reg signed [31:0] W_Im_table[2] = '{
               32'sh00000000, 32'shc0000000
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 3)
         begin
            reg signed [31:0] W_Re_table[4] = '{
               32'sh40000000, 32'sh2d413ccd, 32'sh00000000, 32'shd2bec333
            };

            reg signed [31:0] W_Im_table[4] = '{
               32'sh00000000, 32'shd2bec333, 32'shc0000000, 32'shd2bec333
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 4)
         begin
            reg signed [31:0] W_Re_table[8] = '{
               32'sh40000000, 32'sh3b20d79e, 32'sh2d413ccd, 32'sh187de2a7, 32'sh00000000, 32'she7821d59, 32'shd2bec333, 32'shc4df2862
            };

            reg signed [31:0] W_Im_table[8] = '{
               32'sh00000000, 32'she7821d59, 32'shd2bec333, 32'shc4df2862, 32'shc0000000, 32'shc4df2862, 32'shd2bec333, 32'she7821d59
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 5)
         begin
            reg signed [31:0] W_Re_table[16] = '{
               32'sh40000000, 32'sh3ec52fa0, 32'sh3b20d79e, 32'sh3536cc52, 32'sh2d413ccd, 32'sh238e7673, 32'sh187de2a7, 32'sh0c7c5c1e, 
               32'sh00000000, 32'shf383a3e2, 32'she7821d59, 32'shdc71898d, 32'shd2bec333, 32'shcac933ae, 32'shc4df2862, 32'shc13ad060
            };

            reg signed [31:0] W_Im_table[16] = '{
               32'sh00000000, 32'shf383a3e2, 32'she7821d59, 32'shdc71898d, 32'shd2bec333, 32'shcac933ae, 32'shc4df2862, 32'shc13ad060, 
               32'shc0000000, 32'shc13ad060, 32'shc4df2862, 32'shcac933ae, 32'shd2bec333, 32'shdc71898d, 32'she7821d59, 32'shf383a3e2
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 6)
         begin
            reg signed [31:0] W_Re_table[32] = '{
               32'sh40000000, 32'sh3fb11b48, 32'sh3ec52fa0, 32'sh3d3e82ae, 32'sh3b20d79e, 32'sh387165e3, 32'sh3536cc52, 32'sh317900d6, 
               32'sh2d413ccd, 32'sh2899e64a, 32'sh238e7673, 32'sh1e2b5d38, 32'sh187de2a7, 32'sh1294062f, 32'sh0c7c5c1e, 32'sh0645e9af, 
               32'sh00000000, 32'shf9ba1651, 32'shf383a3e2, 32'shed6bf9d1, 32'she7821d59, 32'she1d4a2c8, 32'shdc71898d, 32'shd76619b6, 
               32'shd2bec333, 32'shce86ff2a, 32'shcac933ae, 32'shc78e9a1d, 32'shc4df2862, 32'shc2c17d52, 32'shc13ad060, 32'shc04ee4b8
            };

            reg signed [31:0] W_Im_table[32] = '{
               32'sh00000000, 32'shf9ba1651, 32'shf383a3e2, 32'shed6bf9d1, 32'she7821d59, 32'she1d4a2c8, 32'shdc71898d, 32'shd76619b6, 
               32'shd2bec333, 32'shce86ff2a, 32'shcac933ae, 32'shc78e9a1d, 32'shc4df2862, 32'shc2c17d52, 32'shc13ad060, 32'shc04ee4b8, 
               32'shc0000000, 32'shc04ee4b8, 32'shc13ad060, 32'shc2c17d52, 32'shc4df2862, 32'shc78e9a1d, 32'shcac933ae, 32'shce86ff2a, 
               32'shd2bec333, 32'shd76619b6, 32'shdc71898d, 32'she1d4a2c8, 32'she7821d59, 32'shed6bf9d1, 32'shf383a3e2, 32'shf9ba1651
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 7)
         begin
            reg signed [31:0] W_Re_table[64] = '{
               32'sh40000000, 32'sh3fec43c7, 32'sh3fb11b48, 32'sh3f4eaafe, 32'sh3ec52fa0, 32'sh3e14fdf7, 32'sh3d3e82ae, 32'sh3c42420a, 
               32'sh3b20d79e, 32'sh39daf5e8, 32'sh387165e3, 32'sh36e5068a, 32'sh3536cc52, 32'sh3367c090, 32'sh317900d6, 32'sh2f6bbe45, 
               32'sh2d413ccd, 32'sh2afad269, 32'sh2899e64a, 32'sh261feffa, 32'sh238e7673, 32'sh20e70f32, 32'sh1e2b5d38, 32'sh1b5d100a, 
               32'sh187de2a7, 32'sh158f9a76, 32'sh1294062f, 32'sh0f8cfcbe, 32'sh0c7c5c1e, 32'sh09640837, 32'sh0645e9af, 32'sh0323ecbe, 
               32'sh00000000, 32'shfcdc1342, 32'shf9ba1651, 32'shf69bf7c9, 32'shf383a3e2, 32'shf0730342, 32'shed6bf9d1, 32'shea70658a, 
               32'she7821d59, 32'she4a2eff6, 32'she1d4a2c8, 32'shdf18f0ce, 32'shdc71898d, 32'shd9e01006, 32'shd76619b6, 32'shd5052d97, 
               32'shd2bec333, 32'shd09441bb, 32'shce86ff2a, 32'shcc983f70, 32'shcac933ae, 32'shc91af976, 32'shc78e9a1d, 32'shc6250a18, 
               32'shc4df2862, 32'shc3bdbdf6, 32'shc2c17d52, 32'shc1eb0209, 32'shc13ad060, 32'shc0b15502, 32'shc04ee4b8, 32'shc013bc39
            };

            reg signed [31:0] W_Im_table[64] = '{
               32'sh00000000, 32'shfcdc1342, 32'shf9ba1651, 32'shf69bf7c9, 32'shf383a3e2, 32'shf0730342, 32'shed6bf9d1, 32'shea70658a, 
               32'she7821d59, 32'she4a2eff6, 32'she1d4a2c8, 32'shdf18f0ce, 32'shdc71898d, 32'shd9e01006, 32'shd76619b6, 32'shd5052d97, 
               32'shd2bec333, 32'shd09441bb, 32'shce86ff2a, 32'shcc983f70, 32'shcac933ae, 32'shc91af976, 32'shc78e9a1d, 32'shc6250a18, 
               32'shc4df2862, 32'shc3bdbdf6, 32'shc2c17d52, 32'shc1eb0209, 32'shc13ad060, 32'shc0b15502, 32'shc04ee4b8, 32'shc013bc39, 
               32'shc0000000, 32'shc013bc39, 32'shc04ee4b8, 32'shc0b15502, 32'shc13ad060, 32'shc1eb0209, 32'shc2c17d52, 32'shc3bdbdf6, 
               32'shc4df2862, 32'shc6250a18, 32'shc78e9a1d, 32'shc91af976, 32'shcac933ae, 32'shcc983f70, 32'shce86ff2a, 32'shd09441bb, 
               32'shd2bec333, 32'shd5052d97, 32'shd76619b6, 32'shd9e01006, 32'shdc71898d, 32'shdf18f0ce, 32'she1d4a2c8, 32'she4a2eff6, 
               32'she7821d59, 32'shea70658a, 32'shed6bf9d1, 32'shf0730342, 32'shf383a3e2, 32'shf69bf7c9, 32'shf9ba1651, 32'shfcdc1342
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 8)
         begin
            reg signed [31:0] W_Re_table[128] = '{
               32'sh40000000, 32'sh3ffb10c1, 32'sh3fec43c7, 32'sh3fd39b5a, 32'sh3fb11b48, 32'sh3f84c8e2, 32'sh3f4eaafe, 32'sh3f0ec9f5, 
               32'sh3ec52fa0, 32'sh3e71e759, 32'sh3e14fdf7, 32'sh3dae81cf, 32'sh3d3e82ae, 32'sh3cc511d9, 32'sh3c42420a, 32'sh3bb6276e, 
               32'sh3b20d79e, 32'sh3a8269a3, 32'sh39daf5e8, 32'sh392a9642, 32'sh387165e3, 32'sh37af8159, 32'sh36e5068a, 32'sh361214b0, 
               32'sh3536cc52, 32'sh34534f41, 32'sh3367c090, 32'sh32744493, 32'sh317900d6, 32'sh30761c18, 32'sh2f6bbe45, 32'sh2e5a1070, 
               32'sh2d413ccd, 32'sh2c216eaa, 32'sh2afad269, 32'sh29cd9578, 32'sh2899e64a, 32'sh275ff452, 32'sh261feffa, 32'sh24da0a9a, 
               32'sh238e7673, 32'sh223d66a8, 32'sh20e70f32, 32'sh1f8ba4dc, 32'sh1e2b5d38, 32'sh1cc66e99, 32'sh1b5d100a, 32'sh19ef7944, 
               32'sh187de2a7, 32'sh17088531, 32'sh158f9a76, 32'sh14135c94, 32'sh1294062f, 32'sh1111d263, 32'sh0f8cfcbe, 32'sh0e05c135, 
               32'sh0c7c5c1e, 32'sh0af10a22, 32'sh09640837, 32'sh07d59396, 32'sh0645e9af, 32'sh04b54825, 32'sh0323ecbe, 32'sh0192155f, 
               32'sh00000000, 32'shfe6deaa1, 32'shfcdc1342, 32'shfb4ab7db, 32'shf9ba1651, 32'shf82a6c6a, 32'shf69bf7c9, 32'shf50ef5de, 
               32'shf383a3e2, 32'shf1fa3ecb, 32'shf0730342, 32'sheeee2d9d, 32'shed6bf9d1, 32'shebeca36c, 32'shea70658a, 32'she8f77acf, 
               32'she7821d59, 32'she61086bc, 32'she4a2eff6, 32'she3399167, 32'she1d4a2c8, 32'she0745b24, 32'shdf18f0ce, 32'shddc29958, 
               32'shdc71898d, 32'shdb25f566, 32'shd9e01006, 32'shd8a00bae, 32'shd76619b6, 32'shd6326a88, 32'shd5052d97, 32'shd3de9156, 
               32'shd2bec333, 32'shd1a5ef90, 32'shd09441bb, 32'shcf89e3e8, 32'shce86ff2a, 32'shcd8bbb6d, 32'shcc983f70, 32'shcbacb0bf, 
               32'shcac933ae, 32'shc9edeb50, 32'shc91af976, 32'shc8507ea7, 32'shc78e9a1d, 32'shc6d569be, 32'shc6250a18, 32'shc57d965d, 
               32'shc4df2862, 32'shc449d892, 32'shc3bdbdf6, 32'shc33aee27, 32'shc2c17d52, 32'shc2517e31, 32'shc1eb0209, 32'shc18e18a7, 
               32'shc13ad060, 32'shc0f1360b, 32'shc0b15502, 32'shc07b371e, 32'shc04ee4b8, 32'shc02c64a6, 32'shc013bc39, 32'shc004ef3f
            };

            reg signed [31:0] W_Im_table[128] = '{
               32'sh00000000, 32'shfe6deaa1, 32'shfcdc1342, 32'shfb4ab7db, 32'shf9ba1651, 32'shf82a6c6a, 32'shf69bf7c9, 32'shf50ef5de, 
               32'shf383a3e2, 32'shf1fa3ecb, 32'shf0730342, 32'sheeee2d9d, 32'shed6bf9d1, 32'shebeca36c, 32'shea70658a, 32'she8f77acf, 
               32'she7821d59, 32'she61086bc, 32'she4a2eff6, 32'she3399167, 32'she1d4a2c8, 32'she0745b24, 32'shdf18f0ce, 32'shddc29958, 
               32'shdc71898d, 32'shdb25f566, 32'shd9e01006, 32'shd8a00bae, 32'shd76619b6, 32'shd6326a88, 32'shd5052d97, 32'shd3de9156, 
               32'shd2bec333, 32'shd1a5ef90, 32'shd09441bb, 32'shcf89e3e8, 32'shce86ff2a, 32'shcd8bbb6d, 32'shcc983f70, 32'shcbacb0bf, 
               32'shcac933ae, 32'shc9edeb50, 32'shc91af976, 32'shc8507ea7, 32'shc78e9a1d, 32'shc6d569be, 32'shc6250a18, 32'shc57d965d, 
               32'shc4df2862, 32'shc449d892, 32'shc3bdbdf6, 32'shc33aee27, 32'shc2c17d52, 32'shc2517e31, 32'shc1eb0209, 32'shc18e18a7, 
               32'shc13ad060, 32'shc0f1360b, 32'shc0b15502, 32'shc07b371e, 32'shc04ee4b8, 32'shc02c64a6, 32'shc013bc39, 32'shc004ef3f, 
               32'shc0000000, 32'shc004ef3f, 32'shc013bc39, 32'shc02c64a6, 32'shc04ee4b8, 32'shc07b371e, 32'shc0b15502, 32'shc0f1360b, 
               32'shc13ad060, 32'shc18e18a7, 32'shc1eb0209, 32'shc2517e31, 32'shc2c17d52, 32'shc33aee27, 32'shc3bdbdf6, 32'shc449d892, 
               32'shc4df2862, 32'shc57d965d, 32'shc6250a18, 32'shc6d569be, 32'shc78e9a1d, 32'shc8507ea7, 32'shc91af976, 32'shc9edeb50, 
               32'shcac933ae, 32'shcbacb0bf, 32'shcc983f70, 32'shcd8bbb6d, 32'shce86ff2a, 32'shcf89e3e8, 32'shd09441bb, 32'shd1a5ef90, 
               32'shd2bec333, 32'shd3de9156, 32'shd5052d97, 32'shd6326a88, 32'shd76619b6, 32'shd8a00bae, 32'shd9e01006, 32'shdb25f566, 
               32'shdc71898d, 32'shddc29958, 32'shdf18f0ce, 32'she0745b24, 32'she1d4a2c8, 32'she3399167, 32'she4a2eff6, 32'she61086bc, 
               32'she7821d59, 32'she8f77acf, 32'shea70658a, 32'shebeca36c, 32'shed6bf9d1, 32'sheeee2d9d, 32'shf0730342, 32'shf1fa3ecb, 
               32'shf383a3e2, 32'shf50ef5de, 32'shf69bf7c9, 32'shf82a6c6a, 32'shf9ba1651, 32'shfb4ab7db, 32'shfcdc1342, 32'shfe6deaa1
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 9)
         begin
            reg signed [31:0] W_Re_table[256] = '{
               32'sh40000000, 32'sh3ffec42d, 32'sh3ffb10c1, 32'sh3ff4e5e0, 32'sh3fec43c7, 32'sh3fe12acb, 32'sh3fd39b5a, 32'sh3fc395f9, 
               32'sh3fb11b48, 32'sh3f9c2bfb, 32'sh3f84c8e2, 32'sh3f6af2e3, 32'sh3f4eaafe, 32'sh3f2ff24a, 32'sh3f0ec9f5, 32'sh3eeb3347, 
               32'sh3ec52fa0, 32'sh3e9cc076, 32'sh3e71e759, 32'sh3e44a5ef, 32'sh3e14fdf7, 32'sh3de2f148, 32'sh3dae81cf, 32'sh3d77b192, 
               32'sh3d3e82ae, 32'sh3d02f757, 32'sh3cc511d9, 32'sh3c84d496, 32'sh3c42420a, 32'sh3bfd5cc4, 32'sh3bb6276e, 32'sh3b6ca4c4, 
               32'sh3b20d79e, 32'sh3ad2c2e8, 32'sh3a8269a3, 32'sh3a2fcee8, 32'sh39daf5e8, 32'sh3983e1e8, 32'sh392a9642, 32'sh38cf1669, 
               32'sh387165e3, 32'sh3811884d, 32'sh37af8159, 32'sh374b54ce, 32'sh36e5068a, 32'sh367c9a7e, 32'sh361214b0, 32'sh35a5793c, 
               32'sh3536cc52, 32'sh34c61236, 32'sh34534f41, 32'sh33de87de, 32'sh3367c090, 32'sh32eefdea, 32'sh32744493, 32'sh31f79948, 
               32'sh317900d6, 32'sh30f8801f, 32'sh30761c18, 32'sh2ff1d9c7, 32'sh2f6bbe45, 32'sh2ee3cebe, 32'sh2e5a1070, 32'sh2dce88aa, 
               32'sh2d413ccd, 32'sh2cb2324c, 32'sh2c216eaa, 32'sh2b8ef77d, 32'sh2afad269, 32'sh2a650525, 32'sh29cd9578, 32'sh29348937, 
               32'sh2899e64a, 32'sh27fdb2a7, 32'sh275ff452, 32'sh26c0b162, 32'sh261feffa, 32'sh257db64c, 32'sh24da0a9a, 32'sh2434f332, 
               32'sh238e7673, 32'sh22e69ac8, 32'sh223d66a8, 32'sh2192e09b, 32'sh20e70f32, 32'sh2039f90f, 32'sh1f8ba4dc, 32'sh1edc1953, 
               32'sh1e2b5d38, 32'sh1d79775c, 32'sh1cc66e99, 32'sh1c1249d8, 32'sh1b5d100a, 32'sh1aa6c82b, 32'sh19ef7944, 32'sh19372a64, 
               32'sh187de2a7, 32'sh17c3a931, 32'sh17088531, 32'sh164c7ddd, 32'sh158f9a76, 32'sh14d1e242, 32'sh14135c94, 32'sh135410c3, 
               32'sh1294062f, 32'sh11d3443f, 32'sh1111d263, 32'sh104fb80e, 32'sh0f8cfcbe, 32'sh0ec9a7f3, 32'sh0e05c135, 32'sh0d415013, 
               32'sh0c7c5c1e, 32'sh0bb6ecef, 32'sh0af10a22, 32'sh0a2abb59, 32'sh09640837, 32'sh089cf867, 32'sh07d59396, 32'sh070de172, 
               32'sh0645e9af, 32'sh057db403, 32'sh04b54825, 32'sh03ecadcf, 32'sh0323ecbe, 32'sh025b0caf, 32'sh0192155f, 32'sh00c90e90, 
               32'sh00000000, 32'shff36f170, 32'shfe6deaa1, 32'shfda4f351, 32'shfcdc1342, 32'shfc135231, 32'shfb4ab7db, 32'shfa824bfd, 
               32'shf9ba1651, 32'shf8f21e8e, 32'shf82a6c6a, 32'shf7630799, 32'shf69bf7c9, 32'shf5d544a7, 32'shf50ef5de, 32'shf4491311, 
               32'shf383a3e2, 32'shf2beafed, 32'shf1fa3ecb, 32'shf136580d, 32'shf0730342, 32'shefb047f2, 32'sheeee2d9d, 32'shee2cbbc1, 
               32'shed6bf9d1, 32'shecabef3d, 32'shebeca36c, 32'sheb2e1dbe, 32'shea70658a, 32'she9b38223, 32'she8f77acf, 32'she83c56cf, 
               32'she7821d59, 32'she6c8d59c, 32'she61086bc, 32'she55937d5, 32'she4a2eff6, 32'she3edb628, 32'she3399167, 32'she28688a4, 
               32'she1d4a2c8, 32'she123e6ad, 32'she0745b24, 32'shdfc606f1, 32'shdf18f0ce, 32'shde6d1f65, 32'shddc29958, 32'shdd196538, 
               32'shdc71898d, 32'shdbcb0cce, 32'shdb25f566, 32'shda8249b4, 32'shd9e01006, 32'shd93f4e9e, 32'shd8a00bae, 32'shd8024d59, 
               32'shd76619b6, 32'shd6cb76c9, 32'shd6326a88, 32'shd59afadb, 32'shd5052d97, 32'shd4710883, 32'shd3de9156, 32'shd34dcdb4, 
               32'shd2bec333, 32'shd2317756, 32'shd1a5ef90, 32'shd11c3142, 32'shd09441bb, 32'shd00e2639, 32'shcf89e3e8, 32'shcf077fe1, 
               32'shce86ff2a, 32'shce0866b8, 32'shcd8bbb6d, 32'shcd110216, 32'shcc983f70, 32'shcc217822, 32'shcbacb0bf, 32'shcb39edca, 
               32'shcac933ae, 32'shca5a86c4, 32'shc9edeb50, 32'shc9836582, 32'shc91af976, 32'shc8b4ab32, 32'shc8507ea7, 32'shc7ee77b3, 
               32'shc78e9a1d, 32'shc730e997, 32'shc6d569be, 32'shc67c1e18, 32'shc6250a18, 32'shc5d03118, 32'shc57d965d, 32'shc52d3d18, 
               32'shc4df2862, 32'shc4935b3c, 32'shc449d892, 32'shc402a33c, 32'shc3bdbdf6, 32'shc37b2b6a, 32'shc33aee27, 32'shc2fd08a9, 
               32'shc2c17d52, 32'shc2884e6e, 32'shc2517e31, 32'shc21d0eb8, 32'shc1eb0209, 32'shc1bb5a11, 32'shc18e18a7, 32'shc1633f8a, 
               32'shc13ad060, 32'shc114ccb9, 32'shc0f1360b, 32'shc0d00db6, 32'shc0b15502, 32'shc0950d1d, 32'shc07b371e, 32'shc063d405, 
               32'shc04ee4b8, 32'shc03c6a07, 32'shc02c64a6, 32'shc01ed535, 32'shc013bc39, 32'shc00b1a20, 32'shc004ef3f, 32'shc0013bd3
            };

            reg signed [31:0] W_Im_table[256] = '{
               32'sh00000000, 32'shff36f170, 32'shfe6deaa1, 32'shfda4f351, 32'shfcdc1342, 32'shfc135231, 32'shfb4ab7db, 32'shfa824bfd, 
               32'shf9ba1651, 32'shf8f21e8e, 32'shf82a6c6a, 32'shf7630799, 32'shf69bf7c9, 32'shf5d544a7, 32'shf50ef5de, 32'shf4491311, 
               32'shf383a3e2, 32'shf2beafed, 32'shf1fa3ecb, 32'shf136580d, 32'shf0730342, 32'shefb047f2, 32'sheeee2d9d, 32'shee2cbbc1, 
               32'shed6bf9d1, 32'shecabef3d, 32'shebeca36c, 32'sheb2e1dbe, 32'shea70658a, 32'she9b38223, 32'she8f77acf, 32'she83c56cf, 
               32'she7821d59, 32'she6c8d59c, 32'she61086bc, 32'she55937d5, 32'she4a2eff6, 32'she3edb628, 32'she3399167, 32'she28688a4, 
               32'she1d4a2c8, 32'she123e6ad, 32'she0745b24, 32'shdfc606f1, 32'shdf18f0ce, 32'shde6d1f65, 32'shddc29958, 32'shdd196538, 
               32'shdc71898d, 32'shdbcb0cce, 32'shdb25f566, 32'shda8249b4, 32'shd9e01006, 32'shd93f4e9e, 32'shd8a00bae, 32'shd8024d59, 
               32'shd76619b6, 32'shd6cb76c9, 32'shd6326a88, 32'shd59afadb, 32'shd5052d97, 32'shd4710883, 32'shd3de9156, 32'shd34dcdb4, 
               32'shd2bec333, 32'shd2317756, 32'shd1a5ef90, 32'shd11c3142, 32'shd09441bb, 32'shd00e2639, 32'shcf89e3e8, 32'shcf077fe1, 
               32'shce86ff2a, 32'shce0866b8, 32'shcd8bbb6d, 32'shcd110216, 32'shcc983f70, 32'shcc217822, 32'shcbacb0bf, 32'shcb39edca, 
               32'shcac933ae, 32'shca5a86c4, 32'shc9edeb50, 32'shc9836582, 32'shc91af976, 32'shc8b4ab32, 32'shc8507ea7, 32'shc7ee77b3, 
               32'shc78e9a1d, 32'shc730e997, 32'shc6d569be, 32'shc67c1e18, 32'shc6250a18, 32'shc5d03118, 32'shc57d965d, 32'shc52d3d18, 
               32'shc4df2862, 32'shc4935b3c, 32'shc449d892, 32'shc402a33c, 32'shc3bdbdf6, 32'shc37b2b6a, 32'shc33aee27, 32'shc2fd08a9, 
               32'shc2c17d52, 32'shc2884e6e, 32'shc2517e31, 32'shc21d0eb8, 32'shc1eb0209, 32'shc1bb5a11, 32'shc18e18a7, 32'shc1633f8a, 
               32'shc13ad060, 32'shc114ccb9, 32'shc0f1360b, 32'shc0d00db6, 32'shc0b15502, 32'shc0950d1d, 32'shc07b371e, 32'shc063d405, 
               32'shc04ee4b8, 32'shc03c6a07, 32'shc02c64a6, 32'shc01ed535, 32'shc013bc39, 32'shc00b1a20, 32'shc004ef3f, 32'shc0013bd3, 
               32'shc0000000, 32'shc0013bd3, 32'shc004ef3f, 32'shc00b1a20, 32'shc013bc39, 32'shc01ed535, 32'shc02c64a6, 32'shc03c6a07, 
               32'shc04ee4b8, 32'shc063d405, 32'shc07b371e, 32'shc0950d1d, 32'shc0b15502, 32'shc0d00db6, 32'shc0f1360b, 32'shc114ccb9, 
               32'shc13ad060, 32'shc1633f8a, 32'shc18e18a7, 32'shc1bb5a11, 32'shc1eb0209, 32'shc21d0eb8, 32'shc2517e31, 32'shc2884e6e, 
               32'shc2c17d52, 32'shc2fd08a9, 32'shc33aee27, 32'shc37b2b6a, 32'shc3bdbdf6, 32'shc402a33c, 32'shc449d892, 32'shc4935b3c, 
               32'shc4df2862, 32'shc52d3d18, 32'shc57d965d, 32'shc5d03118, 32'shc6250a18, 32'shc67c1e18, 32'shc6d569be, 32'shc730e997, 
               32'shc78e9a1d, 32'shc7ee77b3, 32'shc8507ea7, 32'shc8b4ab32, 32'shc91af976, 32'shc9836582, 32'shc9edeb50, 32'shca5a86c4, 
               32'shcac933ae, 32'shcb39edca, 32'shcbacb0bf, 32'shcc217822, 32'shcc983f70, 32'shcd110216, 32'shcd8bbb6d, 32'shce0866b8, 
               32'shce86ff2a, 32'shcf077fe1, 32'shcf89e3e8, 32'shd00e2639, 32'shd09441bb, 32'shd11c3142, 32'shd1a5ef90, 32'shd2317756, 
               32'shd2bec333, 32'shd34dcdb4, 32'shd3de9156, 32'shd4710883, 32'shd5052d97, 32'shd59afadb, 32'shd6326a88, 32'shd6cb76c9, 
               32'shd76619b6, 32'shd8024d59, 32'shd8a00bae, 32'shd93f4e9e, 32'shd9e01006, 32'shda8249b4, 32'shdb25f566, 32'shdbcb0cce, 
               32'shdc71898d, 32'shdd196538, 32'shddc29958, 32'shde6d1f65, 32'shdf18f0ce, 32'shdfc606f1, 32'she0745b24, 32'she123e6ad, 
               32'she1d4a2c8, 32'she28688a4, 32'she3399167, 32'she3edb628, 32'she4a2eff6, 32'she55937d5, 32'she61086bc, 32'she6c8d59c, 
               32'she7821d59, 32'she83c56cf, 32'she8f77acf, 32'she9b38223, 32'shea70658a, 32'sheb2e1dbe, 32'shebeca36c, 32'shecabef3d, 
               32'shed6bf9d1, 32'shee2cbbc1, 32'sheeee2d9d, 32'shefb047f2, 32'shf0730342, 32'shf136580d, 32'shf1fa3ecb, 32'shf2beafed, 
               32'shf383a3e2, 32'shf4491311, 32'shf50ef5de, 32'shf5d544a7, 32'shf69bf7c9, 32'shf7630799, 32'shf82a6c6a, 32'shf8f21e8e, 
               32'shf9ba1651, 32'shfa824bfd, 32'shfb4ab7db, 32'shfc135231, 32'shfcdc1342, 32'shfda4f351, 32'shfe6deaa1, 32'shff36f170
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 10)
         begin
            reg signed [31:0] W_Re_table[512] = '{
               32'sh40000000, 32'sh3fffb10b, 32'sh3ffec42d, 32'sh3ffd3969, 32'sh3ffb10c1, 32'sh3ff84a3c, 32'sh3ff4e5e0, 32'sh3ff0e3b6, 
               32'sh3fec43c7, 32'sh3fe7061f, 32'sh3fe12acb, 32'sh3fdab1d9, 32'sh3fd39b5a, 32'sh3fcbe75e, 32'sh3fc395f9, 32'sh3fbaa740, 
               32'sh3fb11b48, 32'sh3fa6f228, 32'sh3f9c2bfb, 32'sh3f90c8da, 32'sh3f84c8e2, 32'sh3f782c30, 32'sh3f6af2e3, 32'sh3f5d1d1d, 
               32'sh3f4eaafe, 32'sh3f3f9cab, 32'sh3f2ff24a, 32'sh3f1fabff, 32'sh3f0ec9f5, 32'sh3efd4c54, 32'sh3eeb3347, 32'sh3ed87efc, 
               32'sh3ec52fa0, 32'sh3eb14563, 32'sh3e9cc076, 32'sh3e87a10c, 32'sh3e71e759, 32'sh3e5b9392, 32'sh3e44a5ef, 32'sh3e2d1ea8, 
               32'sh3e14fdf7, 32'sh3dfc4418, 32'sh3de2f148, 32'sh3dc905c5, 32'sh3dae81cf, 32'sh3d9365a8, 32'sh3d77b192, 32'sh3d5b65d2, 
               32'sh3d3e82ae, 32'sh3d21086c, 32'sh3d02f757, 32'sh3ce44fb7, 32'sh3cc511d9, 32'sh3ca53e09, 32'sh3c84d496, 32'sh3c63d5d1, 
               32'sh3c42420a, 32'sh3c201994, 32'sh3bfd5cc4, 32'sh3bda0bf0, 32'sh3bb6276e, 32'sh3b91af97, 32'sh3b6ca4c4, 32'sh3b470753, 
               32'sh3b20d79e, 32'sh3afa1605, 32'sh3ad2c2e8, 32'sh3aaadea6, 32'sh3a8269a3, 32'sh3a596442, 32'sh3a2fcee8, 32'sh3a05a9fd, 
               32'sh39daf5e8, 32'sh39afb313, 32'sh3983e1e8, 32'sh395782d3, 32'sh392a9642, 32'sh38fd1ca4, 32'sh38cf1669, 32'sh38a08402, 
               32'sh387165e3, 32'sh3841bc7f, 32'sh3811884d, 32'sh37e0c9c3, 32'sh37af8159, 32'sh377daf89, 32'sh374b54ce, 32'sh371871a5, 
               32'sh36e5068a, 32'sh36b113fd, 32'sh367c9a7e, 32'sh36479a8e, 32'sh361214b0, 32'sh35dc0968, 32'sh35a5793c, 32'sh356e64b2, 
               32'sh3536cc52, 32'sh34feb0a5, 32'sh34c61236, 32'sh348cf190, 32'sh34534f41, 32'sh34192bd5, 32'sh33de87de, 32'sh33a363ec, 
               32'sh3367c090, 32'sh332b9e5e, 32'sh32eefdea, 32'sh32b1dfc9, 32'sh32744493, 32'sh32362ce0, 32'sh31f79948, 32'sh31b88a66, 
               32'sh317900d6, 32'sh3138fd35, 32'sh30f8801f, 32'sh30b78a36, 32'sh30761c18, 32'sh30343667, 32'sh2ff1d9c7, 32'sh2faf06da, 
               32'sh2f6bbe45, 32'sh2f2800af, 32'sh2ee3cebe, 32'sh2e9f291b, 32'sh2e5a1070, 32'sh2e148566, 32'sh2dce88aa, 32'sh2d881ae8, 
               32'sh2d413ccd, 32'sh2cf9ef09, 32'sh2cb2324c, 32'sh2c6a0746, 32'sh2c216eaa, 32'sh2bd8692b, 32'sh2b8ef77d, 32'sh2b451a55, 
               32'sh2afad269, 32'sh2ab02071, 32'sh2a650525, 32'sh2a19813f, 32'sh29cd9578, 32'sh2981428c, 32'sh29348937, 32'sh28e76a37, 
               32'sh2899e64a, 32'sh284bfe2f, 32'sh27fdb2a7, 32'sh27af0472, 32'sh275ff452, 32'sh2710830c, 32'sh26c0b162, 32'sh2670801a, 
               32'sh261feffa, 32'sh25cf01c8, 32'sh257db64c, 32'sh252c0e4f, 32'sh24da0a9a, 32'sh2487abf7, 32'sh2434f332, 32'sh23e1e117, 
               32'sh238e7673, 32'sh233ab414, 32'sh22e69ac8, 32'sh22922b5e, 32'sh223d66a8, 32'sh21e84d76, 32'sh2192e09b, 32'sh213d20e8, 
               32'sh20e70f32, 32'sh2090ac4d, 32'sh2039f90f, 32'sh1fe2f64c, 32'sh1f8ba4dc, 32'sh1f340596, 32'sh1edc1953, 32'sh1e83e0eb, 
               32'sh1e2b5d38, 32'sh1dd28f15, 32'sh1d79775c, 32'sh1d2016e9, 32'sh1cc66e99, 32'sh1c6c7f4a, 32'sh1c1249d8, 32'sh1bb7cf23, 
               32'sh1b5d100a, 32'sh1b020d6c, 32'sh1aa6c82b, 32'sh1a4b4128, 32'sh19ef7944, 32'sh19937161, 32'sh19372a64, 32'sh18daa52f, 
               32'sh187de2a7, 32'sh1820e3b0, 32'sh17c3a931, 32'sh1766340f, 32'sh17088531, 32'sh16aa9d7e, 32'sh164c7ddd, 32'sh15ee2738, 
               32'sh158f9a76, 32'sh1530d881, 32'sh14d1e242, 32'sh1472b8a5, 32'sh14135c94, 32'sh13b3cefa, 32'sh135410c3, 32'sh12f422db, 
               32'sh1294062f, 32'sh1233bbac, 32'sh11d3443f, 32'sh1172a0d7, 32'sh1111d263, 32'sh10b0d9d0, 32'sh104fb80e, 32'sh0fee6e0d, 
               32'sh0f8cfcbe, 32'sh0f2b650f, 32'sh0ec9a7f3, 32'sh0e67c65a, 32'sh0e05c135, 32'sh0da39978, 32'sh0d415013, 32'sh0cdee5f9, 
               32'sh0c7c5c1e, 32'sh0c19b374, 32'sh0bb6ecef, 32'sh0b540982, 32'sh0af10a22, 32'sh0a8defc3, 32'sh0a2abb59, 32'sh09c76dd8, 
               32'sh09640837, 32'sh09008b6a, 32'sh089cf867, 32'sh08395024, 32'sh07d59396, 32'sh0771c3b3, 32'sh070de172, 32'sh06a9edc9, 
               32'sh0645e9af, 32'sh05e1d61b, 32'sh057db403, 32'sh0519845e, 32'sh04b54825, 32'sh0451004d, 32'sh03ecadcf, 32'sh038851a2, 
               32'sh0323ecbe, 32'sh02bf801a, 32'sh025b0caf, 32'sh01f69373, 32'sh0192155f, 32'sh012d936c, 32'sh00c90e90, 32'sh006487c4, 
               32'sh00000000, 32'shff9b783c, 32'shff36f170, 32'shfed26c94, 32'shfe6deaa1, 32'shfe096c8d, 32'shfda4f351, 32'shfd407fe6, 
               32'shfcdc1342, 32'shfc77ae5e, 32'shfc135231, 32'shfbaeffb3, 32'shfb4ab7db, 32'shfae67ba2, 32'shfa824bfd, 32'shfa1e29e5, 
               32'shf9ba1651, 32'shf9561237, 32'shf8f21e8e, 32'shf88e3c4d, 32'shf82a6c6a, 32'shf7c6afdc, 32'shf7630799, 32'shf6ff7496, 
               32'shf69bf7c9, 32'shf6389228, 32'shf5d544a7, 32'shf572103d, 32'shf50ef5de, 32'shf4abf67e, 32'shf4491311, 32'shf3e64c8c, 
               32'shf383a3e2, 32'shf3211a07, 32'shf2beafed, 32'shf25c6688, 32'shf1fa3ecb, 32'shf19839a6, 32'shf136580d, 32'shf0d49af1, 
               32'shf0730342, 32'shf01191f3, 32'shefb047f2, 32'shef4f2630, 32'sheeee2d9d, 32'shee8d5f29, 32'shee2cbbc1, 32'shedcc4454, 
               32'shed6bf9d1, 32'shed0bdd25, 32'shecabef3d, 32'shec4c3106, 32'shebeca36c, 32'sheb8d475b, 32'sheb2e1dbe, 32'sheacf277f, 
               32'shea70658a, 32'shea11d8c8, 32'she9b38223, 32'she9556282, 32'she8f77acf, 32'she899cbf1, 32'she83c56cf, 32'she7df1c50, 
               32'she7821d59, 32'she7255ad1, 32'she6c8d59c, 32'she66c8e9f, 32'she61086bc, 32'she5b4bed8, 32'she55937d5, 32'she4fdf294, 
               32'she4a2eff6, 32'she44830dd, 32'she3edb628, 32'she39380b6, 32'she3399167, 32'she2dfe917, 32'she28688a4, 32'she22d70eb, 
               32'she1d4a2c8, 32'she17c1f15, 32'she123e6ad, 32'she0cbfa6a, 32'she0745b24, 32'she01d09b4, 32'shdfc606f1, 32'shdf6f53b3, 
               32'shdf18f0ce, 32'shdec2df18, 32'shde6d1f65, 32'shde17b28a, 32'shddc29958, 32'shdd6dd4a2, 32'shdd196538, 32'shdcc54bec, 
               32'shdc71898d, 32'shdc1e1ee9, 32'shdbcb0cce, 32'shdb785409, 32'shdb25f566, 32'shdad3f1b1, 32'shda8249b4, 32'shda30fe38, 
               32'shd9e01006, 32'shd98f7fe6, 32'shd93f4e9e, 32'shd8ef7cf4, 32'shd8a00bae, 32'shd850fb8e, 32'shd8024d59, 32'shd7b401d1, 
               32'shd76619b6, 32'shd71895c9, 32'shd6cb76c9, 32'shd67ebd74, 32'shd6326a88, 32'shd5e67ec1, 32'shd59afadb, 32'shd54fdf8f, 
               32'shd5052d97, 32'shd4bae5ab, 32'shd4710883, 32'shd42796d5, 32'shd3de9156, 32'shd395f8ba, 32'shd34dcdb4, 32'shd30610f7, 
               32'shd2bec333, 32'shd277e518, 32'shd2317756, 32'shd1eb7a9a, 32'shd1a5ef90, 32'shd160d6e5, 32'shd11c3142, 32'shd0d7ff51, 
               32'shd09441bb, 32'shd050f926, 32'shd00e2639, 32'shcfcbc999, 32'shcf89e3e8, 32'shcf4875ca, 32'shcf077fe1, 32'shcec702cb, 
               32'shce86ff2a, 32'shce47759a, 32'shce0866b8, 32'shcdc9d320, 32'shcd8bbb6d, 32'shcd4e2037, 32'shcd110216, 32'shccd461a2, 
               32'shcc983f70, 32'shcc5c9c14, 32'shcc217822, 32'shcbe6d42b, 32'shcbacb0bf, 32'shcb730e70, 32'shcb39edca, 32'shcb014f5b, 
               32'shcac933ae, 32'shca919b4e, 32'shca5a86c4, 32'shca23f698, 32'shc9edeb50, 32'shc9b86572, 32'shc9836582, 32'shc94eec03, 
               32'shc91af976, 32'shc8e78e5b, 32'shc8b4ab32, 32'shc8825077, 32'shc8507ea7, 32'shc81f363d, 32'shc7ee77b3, 32'shc7be4381, 
               32'shc78e9a1d, 32'shc75f7bfe, 32'shc730e997, 32'shc702e35c, 32'shc6d569be, 32'shc6a87d2d, 32'shc67c1e18, 32'shc6504ced, 
               32'shc6250a18, 32'shc5fa5603, 32'shc5d03118, 32'shc5a69bbe, 32'shc57d965d, 32'shc555215a, 32'shc52d3d18, 32'shc505e9fb, 
               32'shc4df2862, 32'shc4b8f8ad, 32'shc4935b3c, 32'shc46e5069, 32'shc449d892, 32'shc425f410, 32'shc402a33c, 32'shc3dfe66c, 
               32'shc3bdbdf6, 32'shc39c2a2f, 32'shc37b2b6a, 32'shc35ac1f7, 32'shc33aee27, 32'shc31bb049, 32'shc2fd08a9, 32'shc2def794, 
               32'shc2c17d52, 32'shc2a49a2e, 32'shc2884e6e, 32'shc26c9a58, 32'shc2517e31, 32'shc236fa3b, 32'shc21d0eb8, 32'shc203bbe8, 
               32'shc1eb0209, 32'shc1d2e158, 32'shc1bb5a11, 32'shc1a46c6e, 32'shc18e18a7, 32'shc1785ef4, 32'shc1633f8a, 32'shc14eba9d, 
               32'shc13ad060, 32'shc1278104, 32'shc114ccb9, 32'shc102b3ac, 32'shc0f1360b, 32'shc0e05401, 32'shc0d00db6, 32'shc0c06355, 
               32'shc0b15502, 32'shc0a2e2e3, 32'shc0950d1d, 32'shc087d3d0, 32'shc07b371e, 32'shc06f3726, 32'shc063d405, 32'shc0590dd8, 
               32'shc04ee4b8, 32'shc04558c0, 32'shc03c6a07, 32'shc03418a2, 32'shc02c64a6, 32'shc0254e27, 32'shc01ed535, 32'shc018f9e1, 
               32'shc013bc39, 32'shc00f1c4a, 32'shc00b1a20, 32'shc007b5c4, 32'shc004ef3f, 32'shc002c697, 32'shc0013bd3, 32'shc0004ef5
            };

            reg signed [31:0] W_Im_table[512] = '{
               32'sh00000000, 32'shff9b783c, 32'shff36f170, 32'shfed26c94, 32'shfe6deaa1, 32'shfe096c8d, 32'shfda4f351, 32'shfd407fe6, 
               32'shfcdc1342, 32'shfc77ae5e, 32'shfc135231, 32'shfbaeffb3, 32'shfb4ab7db, 32'shfae67ba2, 32'shfa824bfd, 32'shfa1e29e5, 
               32'shf9ba1651, 32'shf9561237, 32'shf8f21e8e, 32'shf88e3c4d, 32'shf82a6c6a, 32'shf7c6afdc, 32'shf7630799, 32'shf6ff7496, 
               32'shf69bf7c9, 32'shf6389228, 32'shf5d544a7, 32'shf572103d, 32'shf50ef5de, 32'shf4abf67e, 32'shf4491311, 32'shf3e64c8c, 
               32'shf383a3e2, 32'shf3211a07, 32'shf2beafed, 32'shf25c6688, 32'shf1fa3ecb, 32'shf19839a6, 32'shf136580d, 32'shf0d49af1, 
               32'shf0730342, 32'shf01191f3, 32'shefb047f2, 32'shef4f2630, 32'sheeee2d9d, 32'shee8d5f29, 32'shee2cbbc1, 32'shedcc4454, 
               32'shed6bf9d1, 32'shed0bdd25, 32'shecabef3d, 32'shec4c3106, 32'shebeca36c, 32'sheb8d475b, 32'sheb2e1dbe, 32'sheacf277f, 
               32'shea70658a, 32'shea11d8c8, 32'she9b38223, 32'she9556282, 32'she8f77acf, 32'she899cbf1, 32'she83c56cf, 32'she7df1c50, 
               32'she7821d59, 32'she7255ad1, 32'she6c8d59c, 32'she66c8e9f, 32'she61086bc, 32'she5b4bed8, 32'she55937d5, 32'she4fdf294, 
               32'she4a2eff6, 32'she44830dd, 32'she3edb628, 32'she39380b6, 32'she3399167, 32'she2dfe917, 32'she28688a4, 32'she22d70eb, 
               32'she1d4a2c8, 32'she17c1f15, 32'she123e6ad, 32'she0cbfa6a, 32'she0745b24, 32'she01d09b4, 32'shdfc606f1, 32'shdf6f53b3, 
               32'shdf18f0ce, 32'shdec2df18, 32'shde6d1f65, 32'shde17b28a, 32'shddc29958, 32'shdd6dd4a2, 32'shdd196538, 32'shdcc54bec, 
               32'shdc71898d, 32'shdc1e1ee9, 32'shdbcb0cce, 32'shdb785409, 32'shdb25f566, 32'shdad3f1b1, 32'shda8249b4, 32'shda30fe38, 
               32'shd9e01006, 32'shd98f7fe6, 32'shd93f4e9e, 32'shd8ef7cf4, 32'shd8a00bae, 32'shd850fb8e, 32'shd8024d59, 32'shd7b401d1, 
               32'shd76619b6, 32'shd71895c9, 32'shd6cb76c9, 32'shd67ebd74, 32'shd6326a88, 32'shd5e67ec1, 32'shd59afadb, 32'shd54fdf8f, 
               32'shd5052d97, 32'shd4bae5ab, 32'shd4710883, 32'shd42796d5, 32'shd3de9156, 32'shd395f8ba, 32'shd34dcdb4, 32'shd30610f7, 
               32'shd2bec333, 32'shd277e518, 32'shd2317756, 32'shd1eb7a9a, 32'shd1a5ef90, 32'shd160d6e5, 32'shd11c3142, 32'shd0d7ff51, 
               32'shd09441bb, 32'shd050f926, 32'shd00e2639, 32'shcfcbc999, 32'shcf89e3e8, 32'shcf4875ca, 32'shcf077fe1, 32'shcec702cb, 
               32'shce86ff2a, 32'shce47759a, 32'shce0866b8, 32'shcdc9d320, 32'shcd8bbb6d, 32'shcd4e2037, 32'shcd110216, 32'shccd461a2, 
               32'shcc983f70, 32'shcc5c9c14, 32'shcc217822, 32'shcbe6d42b, 32'shcbacb0bf, 32'shcb730e70, 32'shcb39edca, 32'shcb014f5b, 
               32'shcac933ae, 32'shca919b4e, 32'shca5a86c4, 32'shca23f698, 32'shc9edeb50, 32'shc9b86572, 32'shc9836582, 32'shc94eec03, 
               32'shc91af976, 32'shc8e78e5b, 32'shc8b4ab32, 32'shc8825077, 32'shc8507ea7, 32'shc81f363d, 32'shc7ee77b3, 32'shc7be4381, 
               32'shc78e9a1d, 32'shc75f7bfe, 32'shc730e997, 32'shc702e35c, 32'shc6d569be, 32'shc6a87d2d, 32'shc67c1e18, 32'shc6504ced, 
               32'shc6250a18, 32'shc5fa5603, 32'shc5d03118, 32'shc5a69bbe, 32'shc57d965d, 32'shc555215a, 32'shc52d3d18, 32'shc505e9fb, 
               32'shc4df2862, 32'shc4b8f8ad, 32'shc4935b3c, 32'shc46e5069, 32'shc449d892, 32'shc425f410, 32'shc402a33c, 32'shc3dfe66c, 
               32'shc3bdbdf6, 32'shc39c2a2f, 32'shc37b2b6a, 32'shc35ac1f7, 32'shc33aee27, 32'shc31bb049, 32'shc2fd08a9, 32'shc2def794, 
               32'shc2c17d52, 32'shc2a49a2e, 32'shc2884e6e, 32'shc26c9a58, 32'shc2517e31, 32'shc236fa3b, 32'shc21d0eb8, 32'shc203bbe8, 
               32'shc1eb0209, 32'shc1d2e158, 32'shc1bb5a11, 32'shc1a46c6e, 32'shc18e18a7, 32'shc1785ef4, 32'shc1633f8a, 32'shc14eba9d, 
               32'shc13ad060, 32'shc1278104, 32'shc114ccb9, 32'shc102b3ac, 32'shc0f1360b, 32'shc0e05401, 32'shc0d00db6, 32'shc0c06355, 
               32'shc0b15502, 32'shc0a2e2e3, 32'shc0950d1d, 32'shc087d3d0, 32'shc07b371e, 32'shc06f3726, 32'shc063d405, 32'shc0590dd8, 
               32'shc04ee4b8, 32'shc04558c0, 32'shc03c6a07, 32'shc03418a2, 32'shc02c64a6, 32'shc0254e27, 32'shc01ed535, 32'shc018f9e1, 
               32'shc013bc39, 32'shc00f1c4a, 32'shc00b1a20, 32'shc007b5c4, 32'shc004ef3f, 32'shc002c697, 32'shc0013bd3, 32'shc0004ef5, 
               32'shc0000000, 32'shc0004ef5, 32'shc0013bd3, 32'shc002c697, 32'shc004ef3f, 32'shc007b5c4, 32'shc00b1a20, 32'shc00f1c4a, 
               32'shc013bc39, 32'shc018f9e1, 32'shc01ed535, 32'shc0254e27, 32'shc02c64a6, 32'shc03418a2, 32'shc03c6a07, 32'shc04558c0, 
               32'shc04ee4b8, 32'shc0590dd8, 32'shc063d405, 32'shc06f3726, 32'shc07b371e, 32'shc087d3d0, 32'shc0950d1d, 32'shc0a2e2e3, 
               32'shc0b15502, 32'shc0c06355, 32'shc0d00db6, 32'shc0e05401, 32'shc0f1360b, 32'shc102b3ac, 32'shc114ccb9, 32'shc1278104, 
               32'shc13ad060, 32'shc14eba9d, 32'shc1633f8a, 32'shc1785ef4, 32'shc18e18a7, 32'shc1a46c6e, 32'shc1bb5a11, 32'shc1d2e158, 
               32'shc1eb0209, 32'shc203bbe8, 32'shc21d0eb8, 32'shc236fa3b, 32'shc2517e31, 32'shc26c9a58, 32'shc2884e6e, 32'shc2a49a2e, 
               32'shc2c17d52, 32'shc2def794, 32'shc2fd08a9, 32'shc31bb049, 32'shc33aee27, 32'shc35ac1f7, 32'shc37b2b6a, 32'shc39c2a2f, 
               32'shc3bdbdf6, 32'shc3dfe66c, 32'shc402a33c, 32'shc425f410, 32'shc449d892, 32'shc46e5069, 32'shc4935b3c, 32'shc4b8f8ad, 
               32'shc4df2862, 32'shc505e9fb, 32'shc52d3d18, 32'shc555215a, 32'shc57d965d, 32'shc5a69bbe, 32'shc5d03118, 32'shc5fa5603, 
               32'shc6250a18, 32'shc6504ced, 32'shc67c1e18, 32'shc6a87d2d, 32'shc6d569be, 32'shc702e35c, 32'shc730e997, 32'shc75f7bfe, 
               32'shc78e9a1d, 32'shc7be4381, 32'shc7ee77b3, 32'shc81f363d, 32'shc8507ea7, 32'shc8825077, 32'shc8b4ab32, 32'shc8e78e5b, 
               32'shc91af976, 32'shc94eec03, 32'shc9836582, 32'shc9b86572, 32'shc9edeb50, 32'shca23f698, 32'shca5a86c4, 32'shca919b4e, 
               32'shcac933ae, 32'shcb014f5b, 32'shcb39edca, 32'shcb730e70, 32'shcbacb0bf, 32'shcbe6d42b, 32'shcc217822, 32'shcc5c9c14, 
               32'shcc983f70, 32'shccd461a2, 32'shcd110216, 32'shcd4e2037, 32'shcd8bbb6d, 32'shcdc9d320, 32'shce0866b8, 32'shce47759a, 
               32'shce86ff2a, 32'shcec702cb, 32'shcf077fe1, 32'shcf4875ca, 32'shcf89e3e8, 32'shcfcbc999, 32'shd00e2639, 32'shd050f926, 
               32'shd09441bb, 32'shd0d7ff51, 32'shd11c3142, 32'shd160d6e5, 32'shd1a5ef90, 32'shd1eb7a9a, 32'shd2317756, 32'shd277e518, 
               32'shd2bec333, 32'shd30610f7, 32'shd34dcdb4, 32'shd395f8ba, 32'shd3de9156, 32'shd42796d5, 32'shd4710883, 32'shd4bae5ab, 
               32'shd5052d97, 32'shd54fdf8f, 32'shd59afadb, 32'shd5e67ec1, 32'shd6326a88, 32'shd67ebd74, 32'shd6cb76c9, 32'shd71895c9, 
               32'shd76619b6, 32'shd7b401d1, 32'shd8024d59, 32'shd850fb8e, 32'shd8a00bae, 32'shd8ef7cf4, 32'shd93f4e9e, 32'shd98f7fe6, 
               32'shd9e01006, 32'shda30fe38, 32'shda8249b4, 32'shdad3f1b1, 32'shdb25f566, 32'shdb785409, 32'shdbcb0cce, 32'shdc1e1ee9, 
               32'shdc71898d, 32'shdcc54bec, 32'shdd196538, 32'shdd6dd4a2, 32'shddc29958, 32'shde17b28a, 32'shde6d1f65, 32'shdec2df18, 
               32'shdf18f0ce, 32'shdf6f53b3, 32'shdfc606f1, 32'she01d09b4, 32'she0745b24, 32'she0cbfa6a, 32'she123e6ad, 32'she17c1f15, 
               32'she1d4a2c8, 32'she22d70eb, 32'she28688a4, 32'she2dfe917, 32'she3399167, 32'she39380b6, 32'she3edb628, 32'she44830dd, 
               32'she4a2eff6, 32'she4fdf294, 32'she55937d5, 32'she5b4bed8, 32'she61086bc, 32'she66c8e9f, 32'she6c8d59c, 32'she7255ad1, 
               32'she7821d59, 32'she7df1c50, 32'she83c56cf, 32'she899cbf1, 32'she8f77acf, 32'she9556282, 32'she9b38223, 32'shea11d8c8, 
               32'shea70658a, 32'sheacf277f, 32'sheb2e1dbe, 32'sheb8d475b, 32'shebeca36c, 32'shec4c3106, 32'shecabef3d, 32'shed0bdd25, 
               32'shed6bf9d1, 32'shedcc4454, 32'shee2cbbc1, 32'shee8d5f29, 32'sheeee2d9d, 32'shef4f2630, 32'shefb047f2, 32'shf01191f3, 
               32'shf0730342, 32'shf0d49af1, 32'shf136580d, 32'shf19839a6, 32'shf1fa3ecb, 32'shf25c6688, 32'shf2beafed, 32'shf3211a07, 
               32'shf383a3e2, 32'shf3e64c8c, 32'shf4491311, 32'shf4abf67e, 32'shf50ef5de, 32'shf572103d, 32'shf5d544a7, 32'shf6389228, 
               32'shf69bf7c9, 32'shf6ff7496, 32'shf7630799, 32'shf7c6afdc, 32'shf82a6c6a, 32'shf88e3c4d, 32'shf8f21e8e, 32'shf9561237, 
               32'shf9ba1651, 32'shfa1e29e5, 32'shfa824bfd, 32'shfae67ba2, 32'shfb4ab7db, 32'shfbaeffb3, 32'shfc135231, 32'shfc77ae5e, 
               32'shfcdc1342, 32'shfd407fe6, 32'shfda4f351, 32'shfe096c8d, 32'shfe6deaa1, 32'shfed26c94, 32'shff36f170, 32'shff9b783c
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 11)
         begin
            reg signed [31:0] W_Re_table[1024] = '{
               32'sh40000000, 32'sh3fffec43, 32'sh3fffb10b, 32'sh3fff4e59, 32'sh3ffec42d, 32'sh3ffe1288, 32'sh3ffd3969, 32'sh3ffc38d1, 
               32'sh3ffb10c1, 32'sh3ff9c13a, 32'sh3ff84a3c, 32'sh3ff6abc8, 32'sh3ff4e5e0, 32'sh3ff2f884, 32'sh3ff0e3b6, 32'sh3feea776, 
               32'sh3fec43c7, 32'sh3fe9b8a9, 32'sh3fe7061f, 32'sh3fe42c2a, 32'sh3fe12acb, 32'sh3fde0205, 32'sh3fdab1d9, 32'sh3fd73a4a, 
               32'sh3fd39b5a, 32'sh3fcfd50b, 32'sh3fcbe75e, 32'sh3fc7d258, 32'sh3fc395f9, 32'sh3fbf3246, 32'sh3fbaa740, 32'sh3fb5f4ea, 
               32'sh3fb11b48, 32'sh3fac1a5b, 32'sh3fa6f228, 32'sh3fa1a2b2, 32'sh3f9c2bfb, 32'sh3f968e07, 32'sh3f90c8da, 32'sh3f8adc77, 
               32'sh3f84c8e2, 32'sh3f7e8e1e, 32'sh3f782c30, 32'sh3f71a31b, 32'sh3f6af2e3, 32'sh3f641b8d, 32'sh3f5d1d1d, 32'sh3f55f796, 
               32'sh3f4eaafe, 32'sh3f473759, 32'sh3f3f9cab, 32'sh3f37dafa, 32'sh3f2ff24a, 32'sh3f27e29f, 32'sh3f1fabff, 32'sh3f174e70, 
               32'sh3f0ec9f5, 32'sh3f061e95, 32'sh3efd4c54, 32'sh3ef45338, 32'sh3eeb3347, 32'sh3ee1ec87, 32'sh3ed87efc, 32'sh3eceeaad, 
               32'sh3ec52fa0, 32'sh3ebb4ddb, 32'sh3eb14563, 32'sh3ea7163f, 32'sh3e9cc076, 32'sh3e92440d, 32'sh3e87a10c, 32'sh3e7cd778, 
               32'sh3e71e759, 32'sh3e66d0b4, 32'sh3e5b9392, 32'sh3e502ff9, 32'sh3e44a5ef, 32'sh3e38f57c, 32'sh3e2d1ea8, 32'sh3e212179, 
               32'sh3e14fdf7, 32'sh3e08b42a, 32'sh3dfc4418, 32'sh3defadca, 32'sh3de2f148, 32'sh3dd60e99, 32'sh3dc905c5, 32'sh3dbbd6d4, 
               32'sh3dae81cf, 32'sh3da106bd, 32'sh3d9365a8, 32'sh3d859e96, 32'sh3d77b192, 32'sh3d699ea3, 32'sh3d5b65d2, 32'sh3d4d0728, 
               32'sh3d3e82ae, 32'sh3d2fd86c, 32'sh3d21086c, 32'sh3d1212b7, 32'sh3d02f757, 32'sh3cf3b653, 32'sh3ce44fb7, 32'sh3cd4c38b, 
               32'sh3cc511d9, 32'sh3cb53aaa, 32'sh3ca53e09, 32'sh3c951bff, 32'sh3c84d496, 32'sh3c7467d9, 32'sh3c63d5d1, 32'sh3c531e88, 
               32'sh3c42420a, 32'sh3c314060, 32'sh3c201994, 32'sh3c0ecdb2, 32'sh3bfd5cc4, 32'sh3bebc6d5, 32'sh3bda0bf0, 32'sh3bc82c1f, 
               32'sh3bb6276e, 32'sh3ba3fde7, 32'sh3b91af97, 32'sh3b7f3c87, 32'sh3b6ca4c4, 32'sh3b59e85a, 32'sh3b470753, 32'sh3b3401bb, 
               32'sh3b20d79e, 32'sh3b0d8909, 32'sh3afa1605, 32'sh3ae67ea1, 32'sh3ad2c2e8, 32'sh3abee2e5, 32'sh3aaadea6, 32'sh3a96b636, 
               32'sh3a8269a3, 32'sh3a6df8f8, 32'sh3a596442, 32'sh3a44ab8e, 32'sh3a2fcee8, 32'sh3a1ace5f, 32'sh3a05a9fd, 32'sh39f061d2, 
               32'sh39daf5e8, 32'sh39c5664f, 32'sh39afb313, 32'sh3999dc42, 32'sh3983e1e8, 32'sh396dc414, 32'sh395782d3, 32'sh39411e33, 
               32'sh392a9642, 32'sh3913eb0e, 32'sh38fd1ca4, 32'sh38e62b13, 32'sh38cf1669, 32'sh38b7deb4, 32'sh38a08402, 32'sh38890663, 
               32'sh387165e3, 32'sh3859a292, 32'sh3841bc7f, 32'sh3829b3b9, 32'sh3811884d, 32'sh37f93a4b, 32'sh37e0c9c3, 32'sh37c836c2, 
               32'sh37af8159, 32'sh3796a996, 32'sh377daf89, 32'sh37649341, 32'sh374b54ce, 32'sh3731f440, 32'sh371871a5, 32'sh36fecd0e, 
               32'sh36e5068a, 32'sh36cb1e2a, 32'sh36b113fd, 32'sh3696e814, 32'sh367c9a7e, 32'sh36622b4c, 32'sh36479a8e, 32'sh362ce855, 
               32'sh361214b0, 32'sh35f71fb1, 32'sh35dc0968, 32'sh35c0d1e7, 32'sh35a5793c, 32'sh3589ff7a, 32'sh356e64b2, 32'sh3552a8f4, 
               32'sh3536cc52, 32'sh351acedd, 32'sh34feb0a5, 32'sh34e271bd, 32'sh34c61236, 32'sh34a99221, 32'sh348cf190, 32'sh34703095, 
               32'sh34534f41, 32'sh34364da6, 32'sh34192bd5, 32'sh33fbe9e2, 32'sh33de87de, 32'sh33c105db, 32'sh33a363ec, 32'sh3385a222, 
               32'sh3367c090, 32'sh3349bf48, 32'sh332b9e5e, 32'sh330d5de3, 32'sh32eefdea, 32'sh32d07e85, 32'sh32b1dfc9, 32'sh329321c7, 
               32'sh32744493, 32'sh32554840, 32'sh32362ce0, 32'sh3216f287, 32'sh31f79948, 32'sh31d82137, 32'sh31b88a66, 32'sh3198d4ea, 
               32'sh317900d6, 32'sh31590e3e, 32'sh3138fd35, 32'sh3118cdcf, 32'sh30f8801f, 32'sh30d8143b, 32'sh30b78a36, 32'sh3096e223, 
               32'sh30761c18, 32'sh30553828, 32'sh30343667, 32'sh301316eb, 32'sh2ff1d9c7, 32'sh2fd07f0f, 32'sh2faf06da, 32'sh2f8d713a, 
               32'sh2f6bbe45, 32'sh2f49ee0f, 32'sh2f2800af, 32'sh2f05f637, 32'sh2ee3cebe, 32'sh2ec18a58, 32'sh2e9f291b, 32'sh2e7cab1c, 
               32'sh2e5a1070, 32'sh2e37592c, 32'sh2e148566, 32'sh2df19534, 32'sh2dce88aa, 32'sh2dab5fdf, 32'sh2d881ae8, 32'sh2d64b9da, 
               32'sh2d413ccd, 32'sh2d1da3d5, 32'sh2cf9ef09, 32'sh2cd61e7f, 32'sh2cb2324c, 32'sh2c8e2a87, 32'sh2c6a0746, 32'sh2c45c8a0, 
               32'sh2c216eaa, 32'sh2bfcf97c, 32'sh2bd8692b, 32'sh2bb3bdce, 32'sh2b8ef77d, 32'sh2b6a164d, 32'sh2b451a55, 32'sh2b2003ac, 
               32'sh2afad269, 32'sh2ad586a3, 32'sh2ab02071, 32'sh2a8a9fea, 32'sh2a650525, 32'sh2a3f503a, 32'sh2a19813f, 32'sh29f3984c, 
               32'sh29cd9578, 32'sh29a778db, 32'sh2981428c, 32'sh295af2a3, 32'sh29348937, 32'sh290e0661, 32'sh28e76a37, 32'sh28c0b4d2, 
               32'sh2899e64a, 32'sh2872feb6, 32'sh284bfe2f, 32'sh2824e4cc, 32'sh27fdb2a7, 32'sh27d667d5, 32'sh27af0472, 32'sh27878893, 
               32'sh275ff452, 32'sh273847c8, 32'sh2710830c, 32'sh26e8a637, 32'sh26c0b162, 32'sh2698a4a6, 32'sh2670801a, 32'sh264843d9, 
               32'sh261feffa, 32'sh25f78497, 32'sh25cf01c8, 32'sh25a667a7, 32'sh257db64c, 32'sh2554edd1, 32'sh252c0e4f, 32'sh250317df, 
               32'sh24da0a9a, 32'sh24b0e699, 32'sh2487abf7, 32'sh245e5acc, 32'sh2434f332, 32'sh240b7543, 32'sh23e1e117, 32'sh23b836ca, 
               32'sh238e7673, 32'sh2364a02e, 32'sh233ab414, 32'sh2310b23e, 32'sh22e69ac8, 32'sh22bc6dca, 32'sh22922b5e, 32'sh2267d3a0, 
               32'sh223d66a8, 32'sh2212e492, 32'sh21e84d76, 32'sh21bda171, 32'sh2192e09b, 32'sh21680b0f, 32'sh213d20e8, 32'sh21122240, 
               32'sh20e70f32, 32'sh20bbe7d8, 32'sh2090ac4d, 32'sh20655cac, 32'sh2039f90f, 32'sh200e8190, 32'sh1fe2f64c, 32'sh1fb7575c, 
               32'sh1f8ba4dc, 32'sh1f5fdee6, 32'sh1f340596, 32'sh1f081907, 32'sh1edc1953, 32'sh1eb00696, 32'sh1e83e0eb, 32'sh1e57a86d, 
               32'sh1e2b5d38, 32'sh1dfeff67, 32'sh1dd28f15, 32'sh1da60c5d, 32'sh1d79775c, 32'sh1d4cd02c, 32'sh1d2016e9, 32'sh1cf34baf, 
               32'sh1cc66e99, 32'sh1c997fc4, 32'sh1c6c7f4a, 32'sh1c3f6d47, 32'sh1c1249d8, 32'sh1be51518, 32'sh1bb7cf23, 32'sh1b8a7815, 
               32'sh1b5d100a, 32'sh1b2f971e, 32'sh1b020d6c, 32'sh1ad47312, 32'sh1aa6c82b, 32'sh1a790cd4, 32'sh1a4b4128, 32'sh1a1d6544, 
               32'sh19ef7944, 32'sh19c17d44, 32'sh19937161, 32'sh196555b8, 32'sh19372a64, 32'sh1908ef82, 32'sh18daa52f, 32'sh18ac4b87, 
               32'sh187de2a7, 32'sh184f6aab, 32'sh1820e3b0, 32'sh17f24dd3, 32'sh17c3a931, 32'sh1794f5e6, 32'sh1766340f, 32'sh173763c9, 
               32'sh17088531, 32'sh16d99864, 32'sh16aa9d7e, 32'sh167b949d, 32'sh164c7ddd, 32'sh161d595d, 32'sh15ee2738, 32'sh15bee78c, 
               32'sh158f9a76, 32'sh15604013, 32'sh1530d881, 32'sh150163dc, 32'sh14d1e242, 32'sh14a253d1, 32'sh1472b8a5, 32'sh144310dd, 
               32'sh14135c94, 32'sh13e39be9, 32'sh13b3cefa, 32'sh1383f5e3, 32'sh135410c3, 32'sh13241fb6, 32'sh12f422db, 32'sh12c41a4f, 
               32'sh1294062f, 32'sh1263e699, 32'sh1233bbac, 32'sh12038584, 32'sh11d3443f, 32'sh11a2f7fc, 32'sh1172a0d7, 32'sh11423ef0, 
               32'sh1111d263, 32'sh10e15b4e, 32'sh10b0d9d0, 32'sh10804e06, 32'sh104fb80e, 32'sh101f1807, 32'sh0fee6e0d, 32'sh0fbdba40, 
               32'sh0f8cfcbe, 32'sh0f5c35a3, 32'sh0f2b650f, 32'sh0efa8b20, 32'sh0ec9a7f3, 32'sh0e98bba7, 32'sh0e67c65a, 32'sh0e36c82a, 
               32'sh0e05c135, 32'sh0dd4b19a, 32'sh0da39978, 32'sh0d7278eb, 32'sh0d415013, 32'sh0d101f0e, 32'sh0cdee5f9, 32'sh0cada4f5, 
               32'sh0c7c5c1e, 32'sh0c4b0b94, 32'sh0c19b374, 32'sh0be853de, 32'sh0bb6ecef, 32'sh0b857ec7, 32'sh0b540982, 32'sh0b228d42, 
               32'sh0af10a22, 32'sh0abf8043, 32'sh0a8defc3, 32'sh0a5c58c0, 32'sh0a2abb59, 32'sh09f917ac, 32'sh09c76dd8, 32'sh0995bdfd, 
               32'sh09640837, 32'sh09324ca7, 32'sh09008b6a, 32'sh08cec4a0, 32'sh089cf867, 32'sh086b26de, 32'sh08395024, 32'sh08077457, 
               32'sh07d59396, 32'sh07a3adff, 32'sh0771c3b3, 32'sh073fd4cf, 32'sh070de172, 32'sh06dbe9bb, 32'sh06a9edc9, 32'sh0677edbb, 
               32'sh0645e9af, 32'sh0613e1c5, 32'sh05e1d61b, 32'sh05afc6d0, 32'sh057db403, 32'sh054b9dd3, 32'sh0519845e, 32'sh04e767c5, 
               32'sh04b54825, 32'sh0483259d, 32'sh0451004d, 32'sh041ed854, 32'sh03ecadcf, 32'sh03ba80df, 32'sh038851a2, 32'sh03562038, 
               32'sh0323ecbe, 32'sh02f1b755, 32'sh02bf801a, 32'sh028d472e, 32'sh025b0caf, 32'sh0228d0bb, 32'sh01f69373, 32'sh01c454f5, 
               32'sh0192155f, 32'sh015fd4d2, 32'sh012d936c, 32'sh00fb514b, 32'sh00c90e90, 32'sh0096cb58, 32'sh006487c4, 32'sh003243f1, 
               32'sh00000000, 32'shffcdbc0f, 32'shff9b783c, 32'shff6934a8, 32'shff36f170, 32'shff04aeb5, 32'shfed26c94, 32'shfea02b2e, 
               32'shfe6deaa1, 32'shfe3bab0b, 32'shfe096c8d, 32'shfdd72f45, 32'shfda4f351, 32'shfd72b8d2, 32'shfd407fe6, 32'shfd0e48ab, 
               32'shfcdc1342, 32'shfca9dfc8, 32'shfc77ae5e, 32'shfc457f21, 32'shfc135231, 32'shfbe127ac, 32'shfbaeffb3, 32'shfb7cda63, 
               32'shfb4ab7db, 32'shfb18983b, 32'shfae67ba2, 32'shfab4622d, 32'shfa824bfd, 32'shfa503930, 32'shfa1e29e5, 32'shf9ec1e3b, 
               32'shf9ba1651, 32'shf9881245, 32'shf9561237, 32'shf9241645, 32'shf8f21e8e, 32'shf8c02b31, 32'shf88e3c4d, 32'shf85c5201, 
               32'shf82a6c6a, 32'shf7f88ba9, 32'shf7c6afdc, 32'shf794d922, 32'shf7630799, 32'shf7313b60, 32'shf6ff7496, 32'shf6cdb359, 
               32'shf69bf7c9, 32'shf66a4203, 32'shf6389228, 32'shf606e854, 32'shf5d544a7, 32'shf5a3a740, 32'shf572103d, 32'shf5407fbd, 
               32'shf50ef5de, 32'shf4dd72be, 32'shf4abf67e, 32'shf47a8139, 32'shf4491311, 32'shf417ac22, 32'shf3e64c8c, 32'shf3b4f46c, 
               32'shf383a3e2, 32'shf3525b0b, 32'shf3211a07, 32'shf2efe0f2, 32'shf2beafed, 32'shf28d8715, 32'shf25c6688, 32'shf22b4e66, 
               32'shf1fa3ecb, 32'shf1c937d6, 32'shf19839a6, 32'shf1674459, 32'shf136580d, 32'shf10574e0, 32'shf0d49af1, 32'shf0a3ca5d, 
               32'shf0730342, 32'shf04245c0, 32'shf01191f3, 32'shefe0e7f9, 32'shefb047f2, 32'shef7fb1fa, 32'shef4f2630, 32'shef1ea4b2, 
               32'sheeee2d9d, 32'sheebdc110, 32'shee8d5f29, 32'shee5d0804, 32'shee2cbbc1, 32'shedfc7a7c, 32'shedcc4454, 32'shed9c1967, 
               32'shed6bf9d1, 32'shed3be5b1, 32'shed0bdd25, 32'shecdbe04a, 32'shecabef3d, 32'shec7c0a1d, 32'shec4c3106, 32'shec1c6417, 
               32'shebeca36c, 32'shebbcef23, 32'sheb8d475b, 32'sheb5dac2f, 32'sheb2e1dbe, 32'sheafe9c24, 32'sheacf277f, 32'shea9fbfed, 
               32'shea70658a, 32'shea411874, 32'shea11d8c8, 32'she9e2a6a3, 32'she9b38223, 32'she9846b63, 32'she9556282, 32'she926679c, 
               32'she8f77acf, 32'she8c89c37, 32'she899cbf1, 32'she86b0a1a, 32'she83c56cf, 32'she80db22d, 32'she7df1c50, 32'she7b09555, 
               32'she7821d59, 32'she753b479, 32'she7255ad1, 32'she6f7107e, 32'she6c8d59c, 32'she69aaa48, 32'she66c8e9f, 32'she63e82bc, 
               32'she61086bc, 32'she5e29abc, 32'she5b4bed8, 32'she586f32c, 32'she55937d5, 32'she52b8cee, 32'she4fdf294, 32'she4d068e2, 
               32'she4a2eff6, 32'she47587eb, 32'she44830dd, 32'she41aeae8, 32'she3edb628, 32'she3c092b9, 32'she39380b6, 32'she366803c, 
               32'she3399167, 32'she30cb451, 32'she2dfe917, 32'she2b32fd4, 32'she28688a4, 32'she259f3a3, 32'she22d70eb, 32'she2010099, 
               32'she1d4a2c8, 32'she1a85793, 32'she17c1f15, 32'she14ff96a, 32'she123e6ad, 32'she0f7e6f9, 32'she0cbfa6a, 32'she0a0211a, 
               32'she0745b24, 32'she048a8a4, 32'she01d09b4, 32'shdff17e70, 32'shdfc606f1, 32'shdf9aa354, 32'shdf6f53b3, 32'shdf441828, 
               32'shdf18f0ce, 32'shdeedddc0, 32'shdec2df18, 32'shde97f4f1, 32'shde6d1f65, 32'shde425e8f, 32'shde17b28a, 32'shdded1b6e, 
               32'shddc29958, 32'shdd982c60, 32'shdd6dd4a2, 32'shdd439236, 32'shdd196538, 32'shdcef4dc2, 32'shdcc54bec, 32'shdc9b5fd2, 
               32'shdc71898d, 32'shdc47c936, 32'shdc1e1ee9, 32'shdbf48abd, 32'shdbcb0cce, 32'shdba1a534, 32'shdb785409, 32'shdb4f1967, 
               32'shdb25f566, 32'shdafce821, 32'shdad3f1b1, 32'shdaab122f, 32'shda8249b4, 32'shda599859, 32'shda30fe38, 32'shda087b69, 
               32'shd9e01006, 32'shd9b7bc27, 32'shd98f7fe6, 32'shd9675b5a, 32'shd93f4e9e, 32'shd91759c9, 32'shd8ef7cf4, 32'shd8c7b838, 
               32'shd8a00bae, 32'shd878776d, 32'shd850fb8e, 32'shd829982b, 32'shd8024d59, 32'shd7db1b34, 32'shd7b401d1, 32'shd78d014a, 
               32'shd76619b6, 32'shd73f4b2e, 32'shd71895c9, 32'shd6f1f99f, 32'shd6cb76c9, 32'shd6a50d5d, 32'shd67ebd74, 32'shd6588725, 
               32'shd6326a88, 32'shd60c67b4, 32'shd5e67ec1, 32'shd5c0afc6, 32'shd59afadb, 32'shd5756016, 32'shd54fdf8f, 32'shd52a795d, 
               32'shd5052d97, 32'shd4dffc54, 32'shd4bae5ab, 32'shd495e9b3, 32'shd4710883, 32'shd44c4232, 32'shd42796d5, 32'shd4030684, 
               32'shd3de9156, 32'shd3ba3760, 32'shd395f8ba, 32'shd371d579, 32'shd34dcdb4, 32'shd329e181, 32'shd30610f7, 32'shd2e25c2b, 
               32'shd2bec333, 32'shd29b4626, 32'shd277e518, 32'shd254a021, 32'shd2317756, 32'shd20e6acc, 32'shd1eb7a9a, 32'shd1c8a6d4, 
               32'shd1a5ef90, 32'shd18354e4, 32'shd160d6e5, 32'shd13e75a8, 32'shd11c3142, 32'shd0fa09c9, 32'shd0d7ff51, 32'shd0b611f1, 
               32'shd09441bb, 32'shd0728ec6, 32'shd050f926, 32'shd02f80f1, 32'shd00e2639, 32'shcfece915, 32'shcfcbc999, 32'shcfaac7d8, 
               32'shcf89e3e8, 32'shcf691ddd, 32'shcf4875ca, 32'shcf27ebc5, 32'shcf077fe1, 32'shcee73231, 32'shcec702cb, 32'shcea6f1c2, 
               32'shce86ff2a, 32'shce672b16, 32'shce47759a, 32'shce27dec9, 32'shce0866b8, 32'shcde90d79, 32'shcdc9d320, 32'shcdaab7c0, 
               32'shcd8bbb6d, 32'shcd6cde39, 32'shcd4e2037, 32'shcd2f817b, 32'shcd110216, 32'shccf2a21d, 32'shccd461a2, 32'shccb640b8, 
               32'shcc983f70, 32'shcc7a5dde, 32'shcc5c9c14, 32'shcc3efa25, 32'shcc217822, 32'shcc04161e, 32'shcbe6d42b, 32'shcbc9b25a, 
               32'shcbacb0bf, 32'shcb8fcf6b, 32'shcb730e70, 32'shcb566ddf, 32'shcb39edca, 32'shcb1d8e43, 32'shcb014f5b, 32'shcae53123, 
               32'shcac933ae, 32'shcaad570c, 32'shca919b4e, 32'shca760086, 32'shca5a86c4, 32'shca3f2e19, 32'shca23f698, 32'shca08e04f, 
               32'shc9edeb50, 32'shc9d317ab, 32'shc9b86572, 32'shc99dd4b4, 32'shc9836582, 32'shc96917ec, 32'shc94eec03, 32'shc934e1d6, 
               32'shc91af976, 32'shc90132f2, 32'shc8e78e5b, 32'shc8ce0bc0, 32'shc8b4ab32, 32'shc89b6cbf, 32'shc8825077, 32'shc869566a, 
               32'shc8507ea7, 32'shc837c93e, 32'shc81f363d, 32'shc806c5b5, 32'shc7ee77b3, 32'shc7d64c47, 32'shc7be4381, 32'shc7a65d6e, 
               32'shc78e9a1d, 32'shc776f99d, 32'shc75f7bfe, 32'shc748214c, 32'shc730e997, 32'shc719d4ed, 32'shc702e35c, 32'shc6ec14f2, 
               32'shc6d569be, 32'shc6bee1cd, 32'shc6a87d2d, 32'shc6923bec, 32'shc67c1e18, 32'shc66623be, 32'shc6504ced, 32'shc63a99b1, 
               32'shc6250a18, 32'shc60f9e2e, 32'shc5fa5603, 32'shc5e531a1, 32'shc5d03118, 32'shc5bb5472, 32'shc5a69bbe, 32'shc5920708, 
               32'shc57d965d, 32'shc56949ca, 32'shc555215a, 32'shc5411d1b, 32'shc52d3d18, 32'shc519815f, 32'shc505e9fb, 32'shc4f276f7, 
               32'shc4df2862, 32'shc4cbfe45, 32'shc4b8f8ad, 32'shc4a617a6, 32'shc4935b3c, 32'shc480c379, 32'shc46e5069, 32'shc45c0219, 
               32'shc449d892, 32'shc437d3e1, 32'shc425f410, 32'shc414392b, 32'shc402a33c, 32'shc3f1324e, 32'shc3dfe66c, 32'shc3cebfa0, 
               32'shc3bdbdf6, 32'shc3ace178, 32'shc39c2a2f, 32'shc38b9827, 32'shc37b2b6a, 32'shc36ae401, 32'shc35ac1f7, 32'shc34ac556, 
               32'shc33aee27, 32'shc32b3c75, 32'shc31bb049, 32'shc30c49ad, 32'shc2fd08a9, 32'shc2eded49, 32'shc2def794, 32'shc2d02794, 
               32'shc2c17d52, 32'shc2b2f8d8, 32'shc2a49a2e, 32'shc296615d, 32'shc2884e6e, 32'shc27a616a, 32'shc26c9a58, 32'shc25ef943, 
               32'shc2517e31, 32'shc244292c, 32'shc236fa3b, 32'shc229f167, 32'shc21d0eb8, 32'shc2105236, 32'shc203bbe8, 32'shc1f74bd6, 
               32'shc1eb0209, 32'shc1dede87, 32'shc1d2e158, 32'shc1c70a84, 32'shc1bb5a11, 32'shc1afd007, 32'shc1a46c6e, 32'shc1992f4c, 
               32'shc18e18a7, 32'shc1832888, 32'shc1785ef4, 32'shc16dbbf3, 32'shc1633f8a, 32'shc158e9c1, 32'shc14eba9d, 32'shc144b225, 
               32'shc13ad060, 32'shc1311553, 32'shc1278104, 32'shc11e1379, 32'shc114ccb9, 32'shc10bacc8, 32'shc102b3ac, 32'shc0f9e16b, 
               32'shc0f1360b, 32'shc0e8b190, 32'shc0e05401, 32'shc0d81d61, 32'shc0d00db6, 32'shc0c82506, 32'shc0c06355, 32'shc0b8c8a7, 
               32'shc0b15502, 32'shc0aa086a, 32'shc0a2e2e3, 32'shc09be473, 32'shc0950d1d, 32'shc08e5ce5, 32'shc087d3d0, 32'shc08171e2, 
               32'shc07b371e, 32'shc0752389, 32'shc06f3726, 32'shc06971f9, 32'shc063d405, 32'shc05e5d4e, 32'shc0590dd8, 32'shc053e5a5, 
               32'shc04ee4b8, 32'shc04a0b16, 32'shc04558c0, 32'shc040cdba, 32'shc03c6a07, 32'shc0382da8, 32'shc03418a2, 32'shc0302af5, 
               32'shc02c64a6, 32'shc028c5b6, 32'shc0254e27, 32'shc021fdfb, 32'shc01ed535, 32'shc01bd3d6, 32'shc018f9e1, 32'shc0164757, 
               32'shc013bc39, 32'shc011588a, 32'shc00f1c4a, 32'shc00d077c, 32'shc00b1a20, 32'shc0095438, 32'shc007b5c4, 32'shc0063ec6, 
               32'shc004ef3f, 32'shc003c72f, 32'shc002c697, 32'shc001ed78, 32'shc0013bd3, 32'shc000b1a7, 32'shc0004ef5, 32'shc00013bd
            };

            reg signed [31:0] W_Im_table[1024] = '{
               32'sh00000000, 32'shffcdbc0f, 32'shff9b783c, 32'shff6934a8, 32'shff36f170, 32'shff04aeb5, 32'shfed26c94, 32'shfea02b2e, 
               32'shfe6deaa1, 32'shfe3bab0b, 32'shfe096c8d, 32'shfdd72f45, 32'shfda4f351, 32'shfd72b8d2, 32'shfd407fe6, 32'shfd0e48ab, 
               32'shfcdc1342, 32'shfca9dfc8, 32'shfc77ae5e, 32'shfc457f21, 32'shfc135231, 32'shfbe127ac, 32'shfbaeffb3, 32'shfb7cda63, 
               32'shfb4ab7db, 32'shfb18983b, 32'shfae67ba2, 32'shfab4622d, 32'shfa824bfd, 32'shfa503930, 32'shfa1e29e5, 32'shf9ec1e3b, 
               32'shf9ba1651, 32'shf9881245, 32'shf9561237, 32'shf9241645, 32'shf8f21e8e, 32'shf8c02b31, 32'shf88e3c4d, 32'shf85c5201, 
               32'shf82a6c6a, 32'shf7f88ba9, 32'shf7c6afdc, 32'shf794d922, 32'shf7630799, 32'shf7313b60, 32'shf6ff7496, 32'shf6cdb359, 
               32'shf69bf7c9, 32'shf66a4203, 32'shf6389228, 32'shf606e854, 32'shf5d544a7, 32'shf5a3a740, 32'shf572103d, 32'shf5407fbd, 
               32'shf50ef5de, 32'shf4dd72be, 32'shf4abf67e, 32'shf47a8139, 32'shf4491311, 32'shf417ac22, 32'shf3e64c8c, 32'shf3b4f46c, 
               32'shf383a3e2, 32'shf3525b0b, 32'shf3211a07, 32'shf2efe0f2, 32'shf2beafed, 32'shf28d8715, 32'shf25c6688, 32'shf22b4e66, 
               32'shf1fa3ecb, 32'shf1c937d6, 32'shf19839a6, 32'shf1674459, 32'shf136580d, 32'shf10574e0, 32'shf0d49af1, 32'shf0a3ca5d, 
               32'shf0730342, 32'shf04245c0, 32'shf01191f3, 32'shefe0e7f9, 32'shefb047f2, 32'shef7fb1fa, 32'shef4f2630, 32'shef1ea4b2, 
               32'sheeee2d9d, 32'sheebdc110, 32'shee8d5f29, 32'shee5d0804, 32'shee2cbbc1, 32'shedfc7a7c, 32'shedcc4454, 32'shed9c1967, 
               32'shed6bf9d1, 32'shed3be5b1, 32'shed0bdd25, 32'shecdbe04a, 32'shecabef3d, 32'shec7c0a1d, 32'shec4c3106, 32'shec1c6417, 
               32'shebeca36c, 32'shebbcef23, 32'sheb8d475b, 32'sheb5dac2f, 32'sheb2e1dbe, 32'sheafe9c24, 32'sheacf277f, 32'shea9fbfed, 
               32'shea70658a, 32'shea411874, 32'shea11d8c8, 32'she9e2a6a3, 32'she9b38223, 32'she9846b63, 32'she9556282, 32'she926679c, 
               32'she8f77acf, 32'she8c89c37, 32'she899cbf1, 32'she86b0a1a, 32'she83c56cf, 32'she80db22d, 32'she7df1c50, 32'she7b09555, 
               32'she7821d59, 32'she753b479, 32'she7255ad1, 32'she6f7107e, 32'she6c8d59c, 32'she69aaa48, 32'she66c8e9f, 32'she63e82bc, 
               32'she61086bc, 32'she5e29abc, 32'she5b4bed8, 32'she586f32c, 32'she55937d5, 32'she52b8cee, 32'she4fdf294, 32'she4d068e2, 
               32'she4a2eff6, 32'she47587eb, 32'she44830dd, 32'she41aeae8, 32'she3edb628, 32'she3c092b9, 32'she39380b6, 32'she366803c, 
               32'she3399167, 32'she30cb451, 32'she2dfe917, 32'she2b32fd4, 32'she28688a4, 32'she259f3a3, 32'she22d70eb, 32'she2010099, 
               32'she1d4a2c8, 32'she1a85793, 32'she17c1f15, 32'she14ff96a, 32'she123e6ad, 32'she0f7e6f9, 32'she0cbfa6a, 32'she0a0211a, 
               32'she0745b24, 32'she048a8a4, 32'she01d09b4, 32'shdff17e70, 32'shdfc606f1, 32'shdf9aa354, 32'shdf6f53b3, 32'shdf441828, 
               32'shdf18f0ce, 32'shdeedddc0, 32'shdec2df18, 32'shde97f4f1, 32'shde6d1f65, 32'shde425e8f, 32'shde17b28a, 32'shdded1b6e, 
               32'shddc29958, 32'shdd982c60, 32'shdd6dd4a2, 32'shdd439236, 32'shdd196538, 32'shdcef4dc2, 32'shdcc54bec, 32'shdc9b5fd2, 
               32'shdc71898d, 32'shdc47c936, 32'shdc1e1ee9, 32'shdbf48abd, 32'shdbcb0cce, 32'shdba1a534, 32'shdb785409, 32'shdb4f1967, 
               32'shdb25f566, 32'shdafce821, 32'shdad3f1b1, 32'shdaab122f, 32'shda8249b4, 32'shda599859, 32'shda30fe38, 32'shda087b69, 
               32'shd9e01006, 32'shd9b7bc27, 32'shd98f7fe6, 32'shd9675b5a, 32'shd93f4e9e, 32'shd91759c9, 32'shd8ef7cf4, 32'shd8c7b838, 
               32'shd8a00bae, 32'shd878776d, 32'shd850fb8e, 32'shd829982b, 32'shd8024d59, 32'shd7db1b34, 32'shd7b401d1, 32'shd78d014a, 
               32'shd76619b6, 32'shd73f4b2e, 32'shd71895c9, 32'shd6f1f99f, 32'shd6cb76c9, 32'shd6a50d5d, 32'shd67ebd74, 32'shd6588725, 
               32'shd6326a88, 32'shd60c67b4, 32'shd5e67ec1, 32'shd5c0afc6, 32'shd59afadb, 32'shd5756016, 32'shd54fdf8f, 32'shd52a795d, 
               32'shd5052d97, 32'shd4dffc54, 32'shd4bae5ab, 32'shd495e9b3, 32'shd4710883, 32'shd44c4232, 32'shd42796d5, 32'shd4030684, 
               32'shd3de9156, 32'shd3ba3760, 32'shd395f8ba, 32'shd371d579, 32'shd34dcdb4, 32'shd329e181, 32'shd30610f7, 32'shd2e25c2b, 
               32'shd2bec333, 32'shd29b4626, 32'shd277e518, 32'shd254a021, 32'shd2317756, 32'shd20e6acc, 32'shd1eb7a9a, 32'shd1c8a6d4, 
               32'shd1a5ef90, 32'shd18354e4, 32'shd160d6e5, 32'shd13e75a8, 32'shd11c3142, 32'shd0fa09c9, 32'shd0d7ff51, 32'shd0b611f1, 
               32'shd09441bb, 32'shd0728ec6, 32'shd050f926, 32'shd02f80f1, 32'shd00e2639, 32'shcfece915, 32'shcfcbc999, 32'shcfaac7d8, 
               32'shcf89e3e8, 32'shcf691ddd, 32'shcf4875ca, 32'shcf27ebc5, 32'shcf077fe1, 32'shcee73231, 32'shcec702cb, 32'shcea6f1c2, 
               32'shce86ff2a, 32'shce672b16, 32'shce47759a, 32'shce27dec9, 32'shce0866b8, 32'shcde90d79, 32'shcdc9d320, 32'shcdaab7c0, 
               32'shcd8bbb6d, 32'shcd6cde39, 32'shcd4e2037, 32'shcd2f817b, 32'shcd110216, 32'shccf2a21d, 32'shccd461a2, 32'shccb640b8, 
               32'shcc983f70, 32'shcc7a5dde, 32'shcc5c9c14, 32'shcc3efa25, 32'shcc217822, 32'shcc04161e, 32'shcbe6d42b, 32'shcbc9b25a, 
               32'shcbacb0bf, 32'shcb8fcf6b, 32'shcb730e70, 32'shcb566ddf, 32'shcb39edca, 32'shcb1d8e43, 32'shcb014f5b, 32'shcae53123, 
               32'shcac933ae, 32'shcaad570c, 32'shca919b4e, 32'shca760086, 32'shca5a86c4, 32'shca3f2e19, 32'shca23f698, 32'shca08e04f, 
               32'shc9edeb50, 32'shc9d317ab, 32'shc9b86572, 32'shc99dd4b4, 32'shc9836582, 32'shc96917ec, 32'shc94eec03, 32'shc934e1d6, 
               32'shc91af976, 32'shc90132f2, 32'shc8e78e5b, 32'shc8ce0bc0, 32'shc8b4ab32, 32'shc89b6cbf, 32'shc8825077, 32'shc869566a, 
               32'shc8507ea7, 32'shc837c93e, 32'shc81f363d, 32'shc806c5b5, 32'shc7ee77b3, 32'shc7d64c47, 32'shc7be4381, 32'shc7a65d6e, 
               32'shc78e9a1d, 32'shc776f99d, 32'shc75f7bfe, 32'shc748214c, 32'shc730e997, 32'shc719d4ed, 32'shc702e35c, 32'shc6ec14f2, 
               32'shc6d569be, 32'shc6bee1cd, 32'shc6a87d2d, 32'shc6923bec, 32'shc67c1e18, 32'shc66623be, 32'shc6504ced, 32'shc63a99b1, 
               32'shc6250a18, 32'shc60f9e2e, 32'shc5fa5603, 32'shc5e531a1, 32'shc5d03118, 32'shc5bb5472, 32'shc5a69bbe, 32'shc5920708, 
               32'shc57d965d, 32'shc56949ca, 32'shc555215a, 32'shc5411d1b, 32'shc52d3d18, 32'shc519815f, 32'shc505e9fb, 32'shc4f276f7, 
               32'shc4df2862, 32'shc4cbfe45, 32'shc4b8f8ad, 32'shc4a617a6, 32'shc4935b3c, 32'shc480c379, 32'shc46e5069, 32'shc45c0219, 
               32'shc449d892, 32'shc437d3e1, 32'shc425f410, 32'shc414392b, 32'shc402a33c, 32'shc3f1324e, 32'shc3dfe66c, 32'shc3cebfa0, 
               32'shc3bdbdf6, 32'shc3ace178, 32'shc39c2a2f, 32'shc38b9827, 32'shc37b2b6a, 32'shc36ae401, 32'shc35ac1f7, 32'shc34ac556, 
               32'shc33aee27, 32'shc32b3c75, 32'shc31bb049, 32'shc30c49ad, 32'shc2fd08a9, 32'shc2eded49, 32'shc2def794, 32'shc2d02794, 
               32'shc2c17d52, 32'shc2b2f8d8, 32'shc2a49a2e, 32'shc296615d, 32'shc2884e6e, 32'shc27a616a, 32'shc26c9a58, 32'shc25ef943, 
               32'shc2517e31, 32'shc244292c, 32'shc236fa3b, 32'shc229f167, 32'shc21d0eb8, 32'shc2105236, 32'shc203bbe8, 32'shc1f74bd6, 
               32'shc1eb0209, 32'shc1dede87, 32'shc1d2e158, 32'shc1c70a84, 32'shc1bb5a11, 32'shc1afd007, 32'shc1a46c6e, 32'shc1992f4c, 
               32'shc18e18a7, 32'shc1832888, 32'shc1785ef4, 32'shc16dbbf3, 32'shc1633f8a, 32'shc158e9c1, 32'shc14eba9d, 32'shc144b225, 
               32'shc13ad060, 32'shc1311553, 32'shc1278104, 32'shc11e1379, 32'shc114ccb9, 32'shc10bacc8, 32'shc102b3ac, 32'shc0f9e16b, 
               32'shc0f1360b, 32'shc0e8b190, 32'shc0e05401, 32'shc0d81d61, 32'shc0d00db6, 32'shc0c82506, 32'shc0c06355, 32'shc0b8c8a7, 
               32'shc0b15502, 32'shc0aa086a, 32'shc0a2e2e3, 32'shc09be473, 32'shc0950d1d, 32'shc08e5ce5, 32'shc087d3d0, 32'shc08171e2, 
               32'shc07b371e, 32'shc0752389, 32'shc06f3726, 32'shc06971f9, 32'shc063d405, 32'shc05e5d4e, 32'shc0590dd8, 32'shc053e5a5, 
               32'shc04ee4b8, 32'shc04a0b16, 32'shc04558c0, 32'shc040cdba, 32'shc03c6a07, 32'shc0382da8, 32'shc03418a2, 32'shc0302af5, 
               32'shc02c64a6, 32'shc028c5b6, 32'shc0254e27, 32'shc021fdfb, 32'shc01ed535, 32'shc01bd3d6, 32'shc018f9e1, 32'shc0164757, 
               32'shc013bc39, 32'shc011588a, 32'shc00f1c4a, 32'shc00d077c, 32'shc00b1a20, 32'shc0095438, 32'shc007b5c4, 32'shc0063ec6, 
               32'shc004ef3f, 32'shc003c72f, 32'shc002c697, 32'shc001ed78, 32'shc0013bd3, 32'shc000b1a7, 32'shc0004ef5, 32'shc00013bd, 
               32'shc0000000, 32'shc00013bd, 32'shc0004ef5, 32'shc000b1a7, 32'shc0013bd3, 32'shc001ed78, 32'shc002c697, 32'shc003c72f, 
               32'shc004ef3f, 32'shc0063ec6, 32'shc007b5c4, 32'shc0095438, 32'shc00b1a20, 32'shc00d077c, 32'shc00f1c4a, 32'shc011588a, 
               32'shc013bc39, 32'shc0164757, 32'shc018f9e1, 32'shc01bd3d6, 32'shc01ed535, 32'shc021fdfb, 32'shc0254e27, 32'shc028c5b6, 
               32'shc02c64a6, 32'shc0302af5, 32'shc03418a2, 32'shc0382da8, 32'shc03c6a07, 32'shc040cdba, 32'shc04558c0, 32'shc04a0b16, 
               32'shc04ee4b8, 32'shc053e5a5, 32'shc0590dd8, 32'shc05e5d4e, 32'shc063d405, 32'shc06971f9, 32'shc06f3726, 32'shc0752389, 
               32'shc07b371e, 32'shc08171e2, 32'shc087d3d0, 32'shc08e5ce5, 32'shc0950d1d, 32'shc09be473, 32'shc0a2e2e3, 32'shc0aa086a, 
               32'shc0b15502, 32'shc0b8c8a7, 32'shc0c06355, 32'shc0c82506, 32'shc0d00db6, 32'shc0d81d61, 32'shc0e05401, 32'shc0e8b190, 
               32'shc0f1360b, 32'shc0f9e16b, 32'shc102b3ac, 32'shc10bacc8, 32'shc114ccb9, 32'shc11e1379, 32'shc1278104, 32'shc1311553, 
               32'shc13ad060, 32'shc144b225, 32'shc14eba9d, 32'shc158e9c1, 32'shc1633f8a, 32'shc16dbbf3, 32'shc1785ef4, 32'shc1832888, 
               32'shc18e18a7, 32'shc1992f4c, 32'shc1a46c6e, 32'shc1afd007, 32'shc1bb5a11, 32'shc1c70a84, 32'shc1d2e158, 32'shc1dede87, 
               32'shc1eb0209, 32'shc1f74bd6, 32'shc203bbe8, 32'shc2105236, 32'shc21d0eb8, 32'shc229f167, 32'shc236fa3b, 32'shc244292c, 
               32'shc2517e31, 32'shc25ef943, 32'shc26c9a58, 32'shc27a616a, 32'shc2884e6e, 32'shc296615d, 32'shc2a49a2e, 32'shc2b2f8d8, 
               32'shc2c17d52, 32'shc2d02794, 32'shc2def794, 32'shc2eded49, 32'shc2fd08a9, 32'shc30c49ad, 32'shc31bb049, 32'shc32b3c75, 
               32'shc33aee27, 32'shc34ac556, 32'shc35ac1f7, 32'shc36ae401, 32'shc37b2b6a, 32'shc38b9827, 32'shc39c2a2f, 32'shc3ace178, 
               32'shc3bdbdf6, 32'shc3cebfa0, 32'shc3dfe66c, 32'shc3f1324e, 32'shc402a33c, 32'shc414392b, 32'shc425f410, 32'shc437d3e1, 
               32'shc449d892, 32'shc45c0219, 32'shc46e5069, 32'shc480c379, 32'shc4935b3c, 32'shc4a617a6, 32'shc4b8f8ad, 32'shc4cbfe45, 
               32'shc4df2862, 32'shc4f276f7, 32'shc505e9fb, 32'shc519815f, 32'shc52d3d18, 32'shc5411d1b, 32'shc555215a, 32'shc56949ca, 
               32'shc57d965d, 32'shc5920708, 32'shc5a69bbe, 32'shc5bb5472, 32'shc5d03118, 32'shc5e531a1, 32'shc5fa5603, 32'shc60f9e2e, 
               32'shc6250a18, 32'shc63a99b1, 32'shc6504ced, 32'shc66623be, 32'shc67c1e18, 32'shc6923bec, 32'shc6a87d2d, 32'shc6bee1cd, 
               32'shc6d569be, 32'shc6ec14f2, 32'shc702e35c, 32'shc719d4ed, 32'shc730e997, 32'shc748214c, 32'shc75f7bfe, 32'shc776f99d, 
               32'shc78e9a1d, 32'shc7a65d6e, 32'shc7be4381, 32'shc7d64c47, 32'shc7ee77b3, 32'shc806c5b5, 32'shc81f363d, 32'shc837c93e, 
               32'shc8507ea7, 32'shc869566a, 32'shc8825077, 32'shc89b6cbf, 32'shc8b4ab32, 32'shc8ce0bc0, 32'shc8e78e5b, 32'shc90132f2, 
               32'shc91af976, 32'shc934e1d6, 32'shc94eec03, 32'shc96917ec, 32'shc9836582, 32'shc99dd4b4, 32'shc9b86572, 32'shc9d317ab, 
               32'shc9edeb50, 32'shca08e04f, 32'shca23f698, 32'shca3f2e19, 32'shca5a86c4, 32'shca760086, 32'shca919b4e, 32'shcaad570c, 
               32'shcac933ae, 32'shcae53123, 32'shcb014f5b, 32'shcb1d8e43, 32'shcb39edca, 32'shcb566ddf, 32'shcb730e70, 32'shcb8fcf6b, 
               32'shcbacb0bf, 32'shcbc9b25a, 32'shcbe6d42b, 32'shcc04161e, 32'shcc217822, 32'shcc3efa25, 32'shcc5c9c14, 32'shcc7a5dde, 
               32'shcc983f70, 32'shccb640b8, 32'shccd461a2, 32'shccf2a21d, 32'shcd110216, 32'shcd2f817b, 32'shcd4e2037, 32'shcd6cde39, 
               32'shcd8bbb6d, 32'shcdaab7c0, 32'shcdc9d320, 32'shcde90d79, 32'shce0866b8, 32'shce27dec9, 32'shce47759a, 32'shce672b16, 
               32'shce86ff2a, 32'shcea6f1c2, 32'shcec702cb, 32'shcee73231, 32'shcf077fe1, 32'shcf27ebc5, 32'shcf4875ca, 32'shcf691ddd, 
               32'shcf89e3e8, 32'shcfaac7d8, 32'shcfcbc999, 32'shcfece915, 32'shd00e2639, 32'shd02f80f1, 32'shd050f926, 32'shd0728ec6, 
               32'shd09441bb, 32'shd0b611f1, 32'shd0d7ff51, 32'shd0fa09c9, 32'shd11c3142, 32'shd13e75a8, 32'shd160d6e5, 32'shd18354e4, 
               32'shd1a5ef90, 32'shd1c8a6d4, 32'shd1eb7a9a, 32'shd20e6acc, 32'shd2317756, 32'shd254a021, 32'shd277e518, 32'shd29b4626, 
               32'shd2bec333, 32'shd2e25c2b, 32'shd30610f7, 32'shd329e181, 32'shd34dcdb4, 32'shd371d579, 32'shd395f8ba, 32'shd3ba3760, 
               32'shd3de9156, 32'shd4030684, 32'shd42796d5, 32'shd44c4232, 32'shd4710883, 32'shd495e9b3, 32'shd4bae5ab, 32'shd4dffc54, 
               32'shd5052d97, 32'shd52a795d, 32'shd54fdf8f, 32'shd5756016, 32'shd59afadb, 32'shd5c0afc6, 32'shd5e67ec1, 32'shd60c67b4, 
               32'shd6326a88, 32'shd6588725, 32'shd67ebd74, 32'shd6a50d5d, 32'shd6cb76c9, 32'shd6f1f99f, 32'shd71895c9, 32'shd73f4b2e, 
               32'shd76619b6, 32'shd78d014a, 32'shd7b401d1, 32'shd7db1b34, 32'shd8024d59, 32'shd829982b, 32'shd850fb8e, 32'shd878776d, 
               32'shd8a00bae, 32'shd8c7b838, 32'shd8ef7cf4, 32'shd91759c9, 32'shd93f4e9e, 32'shd9675b5a, 32'shd98f7fe6, 32'shd9b7bc27, 
               32'shd9e01006, 32'shda087b69, 32'shda30fe38, 32'shda599859, 32'shda8249b4, 32'shdaab122f, 32'shdad3f1b1, 32'shdafce821, 
               32'shdb25f566, 32'shdb4f1967, 32'shdb785409, 32'shdba1a534, 32'shdbcb0cce, 32'shdbf48abd, 32'shdc1e1ee9, 32'shdc47c936, 
               32'shdc71898d, 32'shdc9b5fd2, 32'shdcc54bec, 32'shdcef4dc2, 32'shdd196538, 32'shdd439236, 32'shdd6dd4a2, 32'shdd982c60, 
               32'shddc29958, 32'shdded1b6e, 32'shde17b28a, 32'shde425e8f, 32'shde6d1f65, 32'shde97f4f1, 32'shdec2df18, 32'shdeedddc0, 
               32'shdf18f0ce, 32'shdf441828, 32'shdf6f53b3, 32'shdf9aa354, 32'shdfc606f1, 32'shdff17e70, 32'she01d09b4, 32'she048a8a4, 
               32'she0745b24, 32'she0a0211a, 32'she0cbfa6a, 32'she0f7e6f9, 32'she123e6ad, 32'she14ff96a, 32'she17c1f15, 32'she1a85793, 
               32'she1d4a2c8, 32'she2010099, 32'she22d70eb, 32'she259f3a3, 32'she28688a4, 32'she2b32fd4, 32'she2dfe917, 32'she30cb451, 
               32'she3399167, 32'she366803c, 32'she39380b6, 32'she3c092b9, 32'she3edb628, 32'she41aeae8, 32'she44830dd, 32'she47587eb, 
               32'she4a2eff6, 32'she4d068e2, 32'she4fdf294, 32'she52b8cee, 32'she55937d5, 32'she586f32c, 32'she5b4bed8, 32'she5e29abc, 
               32'she61086bc, 32'she63e82bc, 32'she66c8e9f, 32'she69aaa48, 32'she6c8d59c, 32'she6f7107e, 32'she7255ad1, 32'she753b479, 
               32'she7821d59, 32'she7b09555, 32'she7df1c50, 32'she80db22d, 32'she83c56cf, 32'she86b0a1a, 32'she899cbf1, 32'she8c89c37, 
               32'she8f77acf, 32'she926679c, 32'she9556282, 32'she9846b63, 32'she9b38223, 32'she9e2a6a3, 32'shea11d8c8, 32'shea411874, 
               32'shea70658a, 32'shea9fbfed, 32'sheacf277f, 32'sheafe9c24, 32'sheb2e1dbe, 32'sheb5dac2f, 32'sheb8d475b, 32'shebbcef23, 
               32'shebeca36c, 32'shec1c6417, 32'shec4c3106, 32'shec7c0a1d, 32'shecabef3d, 32'shecdbe04a, 32'shed0bdd25, 32'shed3be5b1, 
               32'shed6bf9d1, 32'shed9c1967, 32'shedcc4454, 32'shedfc7a7c, 32'shee2cbbc1, 32'shee5d0804, 32'shee8d5f29, 32'sheebdc110, 
               32'sheeee2d9d, 32'shef1ea4b2, 32'shef4f2630, 32'shef7fb1fa, 32'shefb047f2, 32'shefe0e7f9, 32'shf01191f3, 32'shf04245c0, 
               32'shf0730342, 32'shf0a3ca5d, 32'shf0d49af1, 32'shf10574e0, 32'shf136580d, 32'shf1674459, 32'shf19839a6, 32'shf1c937d6, 
               32'shf1fa3ecb, 32'shf22b4e66, 32'shf25c6688, 32'shf28d8715, 32'shf2beafed, 32'shf2efe0f2, 32'shf3211a07, 32'shf3525b0b, 
               32'shf383a3e2, 32'shf3b4f46c, 32'shf3e64c8c, 32'shf417ac22, 32'shf4491311, 32'shf47a8139, 32'shf4abf67e, 32'shf4dd72be, 
               32'shf50ef5de, 32'shf5407fbd, 32'shf572103d, 32'shf5a3a740, 32'shf5d544a7, 32'shf606e854, 32'shf6389228, 32'shf66a4203, 
               32'shf69bf7c9, 32'shf6cdb359, 32'shf6ff7496, 32'shf7313b60, 32'shf7630799, 32'shf794d922, 32'shf7c6afdc, 32'shf7f88ba9, 
               32'shf82a6c6a, 32'shf85c5201, 32'shf88e3c4d, 32'shf8c02b31, 32'shf8f21e8e, 32'shf9241645, 32'shf9561237, 32'shf9881245, 
               32'shf9ba1651, 32'shf9ec1e3b, 32'shfa1e29e5, 32'shfa503930, 32'shfa824bfd, 32'shfab4622d, 32'shfae67ba2, 32'shfb18983b, 
               32'shfb4ab7db, 32'shfb7cda63, 32'shfbaeffb3, 32'shfbe127ac, 32'shfc135231, 32'shfc457f21, 32'shfc77ae5e, 32'shfca9dfc8, 
               32'shfcdc1342, 32'shfd0e48ab, 32'shfd407fe6, 32'shfd72b8d2, 32'shfda4f351, 32'shfdd72f45, 32'shfe096c8d, 32'shfe3bab0b, 
               32'shfe6deaa1, 32'shfea02b2e, 32'shfed26c94, 32'shff04aeb5, 32'shff36f170, 32'shff6934a8, 32'shff9b783c, 32'shffcdbc0f
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 12)
         begin
            reg signed [31:0] W_Re_table[2048] = '{
               32'sh40000000, 32'sh3ffffb11, 32'sh3fffec43, 32'sh3fffd396, 32'sh3fffb10b, 32'sh3fff84a1, 32'sh3fff4e59, 32'sh3fff0e32, 
               32'sh3ffec42d, 32'sh3ffe704a, 32'sh3ffe1288, 32'sh3ffdaae7, 32'sh3ffd3969, 32'sh3ffcbe0c, 32'sh3ffc38d1, 32'sh3ffba9b8, 
               32'sh3ffb10c1, 32'sh3ffa6dec, 32'sh3ff9c13a, 32'sh3ff90aaa, 32'sh3ff84a3c, 32'sh3ff77ff1, 32'sh3ff6abc8, 32'sh3ff5cdc3, 
               32'sh3ff4e5e0, 32'sh3ff3f420, 32'sh3ff2f884, 32'sh3ff1f30b, 32'sh3ff0e3b6, 32'sh3fefca84, 32'sh3feea776, 32'sh3fed7a8c, 
               32'sh3fec43c7, 32'sh3feb0326, 32'sh3fe9b8a9, 32'sh3fe86452, 32'sh3fe7061f, 32'sh3fe59e12, 32'sh3fe42c2a, 32'sh3fe2b067, 
               32'sh3fe12acb, 32'sh3fdf9b55, 32'sh3fde0205, 32'sh3fdc5edc, 32'sh3fdab1d9, 32'sh3fd8fafe, 32'sh3fd73a4a, 32'sh3fd56fbe, 
               32'sh3fd39b5a, 32'sh3fd1bd1e, 32'sh3fcfd50b, 32'sh3fcde320, 32'sh3fcbe75e, 32'sh3fc9e1c6, 32'sh3fc7d258, 32'sh3fc5b913, 
               32'sh3fc395f9, 32'sh3fc1690a, 32'sh3fbf3246, 32'sh3fbcf1ad, 32'sh3fbaa740, 32'sh3fb852ff, 32'sh3fb5f4ea, 32'sh3fb38d02, 
               32'sh3fb11b48, 32'sh3fae9fbb, 32'sh3fac1a5b, 32'sh3fa98b2a, 32'sh3fa6f228, 32'sh3fa44f55, 32'sh3fa1a2b2, 32'sh3f9eec3e, 
               32'sh3f9c2bfb, 32'sh3f9961e8, 32'sh3f968e07, 32'sh3f93b058, 32'sh3f90c8da, 32'sh3f8dd78f, 32'sh3f8adc77, 32'sh3f87d792, 
               32'sh3f84c8e2, 32'sh3f81b065, 32'sh3f7e8e1e, 32'sh3f7b620c, 32'sh3f782c30, 32'sh3f74ec8a, 32'sh3f71a31b, 32'sh3f6e4fe3, 
               32'sh3f6af2e3, 32'sh3f678c1c, 32'sh3f641b8d, 32'sh3f60a138, 32'sh3f5d1d1d, 32'sh3f598f3c, 32'sh3f55f796, 32'sh3f52562c, 
               32'sh3f4eaafe, 32'sh3f4af60d, 32'sh3f473759, 32'sh3f436ee3, 32'sh3f3f9cab, 32'sh3f3bc0b3, 32'sh3f37dafa, 32'sh3f33eb81, 
               32'sh3f2ff24a, 32'sh3f2bef53, 32'sh3f27e29f, 32'sh3f23cc2e, 32'sh3f1fabff, 32'sh3f1b8215, 32'sh3f174e70, 32'sh3f13110f, 
               32'sh3f0ec9f5, 32'sh3f0a7921, 32'sh3f061e95, 32'sh3f01ba50, 32'sh3efd4c54, 32'sh3ef8d4a1, 32'sh3ef45338, 32'sh3eefc81a, 
               32'sh3eeb3347, 32'sh3ee694c1, 32'sh3ee1ec87, 32'sh3edd3a9a, 32'sh3ed87efc, 32'sh3ed3b9ad, 32'sh3eceeaad, 32'sh3eca11fe, 
               32'sh3ec52fa0, 32'sh3ec04394, 32'sh3ebb4ddb, 32'sh3eb64e75, 32'sh3eb14563, 32'sh3eac32a6, 32'sh3ea7163f, 32'sh3ea1f02f, 
               32'sh3e9cc076, 32'sh3e978715, 32'sh3e92440d, 32'sh3e8cf75f, 32'sh3e87a10c, 32'sh3e824114, 32'sh3e7cd778, 32'sh3e77643a, 
               32'sh3e71e759, 32'sh3e6c60d7, 32'sh3e66d0b4, 32'sh3e6136f3, 32'sh3e5b9392, 32'sh3e55e694, 32'sh3e502ff9, 32'sh3e4a6fc1, 
               32'sh3e44a5ef, 32'sh3e3ed282, 32'sh3e38f57c, 32'sh3e330ede, 32'sh3e2d1ea8, 32'sh3e2724db, 32'sh3e212179, 32'sh3e1b1482, 
               32'sh3e14fdf7, 32'sh3e0eddd9, 32'sh3e08b42a, 32'sh3e0280e9, 32'sh3dfc4418, 32'sh3df5fdb8, 32'sh3defadca, 32'sh3de9544f, 
               32'sh3de2f148, 32'sh3ddc84b5, 32'sh3dd60e99, 32'sh3dcf8ef3, 32'sh3dc905c5, 32'sh3dc2730f, 32'sh3dbbd6d4, 32'sh3db53113, 
               32'sh3dae81cf, 32'sh3da7c907, 32'sh3da106bd, 32'sh3d9a3af2, 32'sh3d9365a8, 32'sh3d8c86de, 32'sh3d859e96, 32'sh3d7eacd2, 
               32'sh3d77b192, 32'sh3d70acd7, 32'sh3d699ea3, 32'sh3d6286f6, 32'sh3d5b65d2, 32'sh3d543b37, 32'sh3d4d0728, 32'sh3d45c9a4, 
               32'sh3d3e82ae, 32'sh3d373245, 32'sh3d2fd86c, 32'sh3d287523, 32'sh3d21086c, 32'sh3d199248, 32'sh3d1212b7, 32'sh3d0a89bc, 
               32'sh3d02f757, 32'sh3cfb5b89, 32'sh3cf3b653, 32'sh3cec07b8, 32'sh3ce44fb7, 32'sh3cdc8e52, 32'sh3cd4c38b, 32'sh3cccef62, 
               32'sh3cc511d9, 32'sh3cbd2af0, 32'sh3cb53aaa, 32'sh3cad4107, 32'sh3ca53e09, 32'sh3c9d31b0, 32'sh3c951bff, 32'sh3c8cfcf6, 
               32'sh3c84d496, 32'sh3c7ca2e2, 32'sh3c7467d9, 32'sh3c6c237e, 32'sh3c63d5d1, 32'sh3c5b7ed4, 32'sh3c531e88, 32'sh3c4ab4ef, 
               32'sh3c42420a, 32'sh3c39c5da, 32'sh3c314060, 32'sh3c28b19e, 32'sh3c201994, 32'sh3c177845, 32'sh3c0ecdb2, 32'sh3c0619dc, 
               32'sh3bfd5cc4, 32'sh3bf4966c, 32'sh3bebc6d5, 32'sh3be2ee01, 32'sh3bda0bf0, 32'sh3bd120a4, 32'sh3bc82c1f, 32'sh3bbf2e62, 
               32'sh3bb6276e, 32'sh3bad1744, 32'sh3ba3fde7, 32'sh3b9adb57, 32'sh3b91af97, 32'sh3b887aa6, 32'sh3b7f3c87, 32'sh3b75f53c, 
               32'sh3b6ca4c4, 32'sh3b634b23, 32'sh3b59e85a, 32'sh3b507c69, 32'sh3b470753, 32'sh3b3d8918, 32'sh3b3401bb, 32'sh3b2a713d, 
               32'sh3b20d79e, 32'sh3b1734e2, 32'sh3b0d8909, 32'sh3b03d414, 32'sh3afa1605, 32'sh3af04edf, 32'sh3ae67ea1, 32'sh3adca54e, 
               32'sh3ad2c2e8, 32'sh3ac8d76f, 32'sh3abee2e5, 32'sh3ab4e54c, 32'sh3aaadea6, 32'sh3aa0cef3, 32'sh3a96b636, 32'sh3a8c9470, 
               32'sh3a8269a3, 32'sh3a7835cf, 32'sh3a6df8f8, 32'sh3a63b31d, 32'sh3a596442, 32'sh3a4f0c67, 32'sh3a44ab8e, 32'sh3a3a41b9, 
               32'sh3a2fcee8, 32'sh3a25531f, 32'sh3a1ace5f, 32'sh3a1040a8, 32'sh3a05a9fd, 32'sh39fb0a60, 32'sh39f061d2, 32'sh39e5b054, 
               32'sh39daf5e8, 32'sh39d03291, 32'sh39c5664f, 32'sh39ba9125, 32'sh39afb313, 32'sh39a4cc1c, 32'sh3999dc42, 32'sh398ee385, 
               32'sh3983e1e8, 32'sh3978d76c, 32'sh396dc414, 32'sh3962a7e0, 32'sh395782d3, 32'sh394c54ee, 32'sh39411e33, 32'sh3935dea4, 
               32'sh392a9642, 32'sh391f4510, 32'sh3913eb0e, 32'sh3908883f, 32'sh38fd1ca4, 32'sh38f1a840, 32'sh38e62b13, 32'sh38daa520, 
               32'sh38cf1669, 32'sh38c37eef, 32'sh38b7deb4, 32'sh38ac35ba, 32'sh38a08402, 32'sh3894c98f, 32'sh38890663, 32'sh387d3a7e, 
               32'sh387165e3, 32'sh38658894, 32'sh3859a292, 32'sh384db3e0, 32'sh3841bc7f, 32'sh3835bc71, 32'sh3829b3b9, 32'sh381da256, 
               32'sh3811884d, 32'sh3805659e, 32'sh37f93a4b, 32'sh37ed0657, 32'sh37e0c9c3, 32'sh37d48490, 32'sh37c836c2, 32'sh37bbe05a, 
               32'sh37af8159, 32'sh37a319c2, 32'sh3796a996, 32'sh378a30d8, 32'sh377daf89, 32'sh377125ac, 32'sh37649341, 32'sh3757f84c, 
               32'sh374b54ce, 32'sh373ea8ca, 32'sh3731f440, 32'sh37253733, 32'sh371871a5, 32'sh370ba398, 32'sh36fecd0e, 32'sh36f1ee09, 
               32'sh36e5068a, 32'sh36d81695, 32'sh36cb1e2a, 32'sh36be1d4c, 32'sh36b113fd, 32'sh36a4023f, 32'sh3696e814, 32'sh3689c57d, 
               32'sh367c9a7e, 32'sh366f6717, 32'sh36622b4c, 32'sh3654e71d, 32'sh36479a8e, 32'sh363a45a0, 32'sh362ce855, 32'sh361f82af, 
               32'sh361214b0, 32'sh36049e5b, 32'sh35f71fb1, 32'sh35e998b5, 32'sh35dc0968, 32'sh35ce71ce, 32'sh35c0d1e7, 32'sh35b329b5, 
               32'sh35a5793c, 32'sh3597c07d, 32'sh3589ff7a, 32'sh357c3636, 32'sh356e64b2, 32'sh35608af1, 32'sh3552a8f4, 32'sh3544bebf, 
               32'sh3536cc52, 32'sh3528d1b1, 32'sh351acedd, 32'sh350cc3d8, 32'sh34feb0a5, 32'sh34f09546, 32'sh34e271bd, 32'sh34d4460c, 
               32'sh34c61236, 32'sh34b7d63c, 32'sh34a99221, 32'sh349b45e7, 32'sh348cf190, 32'sh347e951f, 32'sh34703095, 32'sh3461c3f5, 
               32'sh34534f41, 32'sh3444d27b, 32'sh34364da6, 32'sh3427c0c3, 32'sh34192bd5, 32'sh340a8edf, 32'sh33fbe9e2, 32'sh33ed3ce1, 
               32'sh33de87de, 32'sh33cfcadc, 32'sh33c105db, 32'sh33b238e0, 32'sh33a363ec, 32'sh33948701, 32'sh3385a222, 32'sh3376b551, 
               32'sh3367c090, 32'sh3358c3e2, 32'sh3349bf48, 32'sh333ab2c6, 32'sh332b9e5e, 32'sh331c8211, 32'sh330d5de3, 32'sh32fe31d5, 
               32'sh32eefdea, 32'sh32dfc224, 32'sh32d07e85, 32'sh32c13311, 32'sh32b1dfc9, 32'sh32a284b0, 32'sh329321c7, 32'sh3283b712, 
               32'sh32744493, 32'sh3264ca4c, 32'sh32554840, 32'sh3245be70, 32'sh32362ce0, 32'sh32269391, 32'sh3216f287, 32'sh320749c3, 
               32'sh31f79948, 32'sh31e7e118, 32'sh31d82137, 32'sh31c859a5, 32'sh31b88a66, 32'sh31a8b37c, 32'sh3198d4ea, 32'sh3188eeb2, 
               32'sh317900d6, 32'sh31690b59, 32'sh31590e3e, 32'sh31490986, 32'sh3138fd35, 32'sh3128e94c, 32'sh3118cdcf, 32'sh3108aabf, 
               32'sh30f8801f, 32'sh30e84df3, 32'sh30d8143b, 32'sh30c7d2fb, 32'sh30b78a36, 32'sh30a739ed, 32'sh3096e223, 32'sh308682dc, 
               32'sh30761c18, 32'sh3065addb, 32'sh30553828, 32'sh3044bb00, 32'sh30343667, 32'sh3023aa5f, 32'sh301316eb, 32'sh30027c0c, 
               32'sh2ff1d9c7, 32'sh2fe1301c, 32'sh2fd07f0f, 32'sh2fbfc6a3, 32'sh2faf06da, 32'sh2f9e3fb6, 32'sh2f8d713a, 32'sh2f7c9b69, 
               32'sh2f6bbe45, 32'sh2f5ad9d1, 32'sh2f49ee0f, 32'sh2f38fb03, 32'sh2f2800af, 32'sh2f16ff14, 32'sh2f05f637, 32'sh2ef4e619, 
               32'sh2ee3cebe, 32'sh2ed2b027, 32'sh2ec18a58, 32'sh2eb05d53, 32'sh2e9f291b, 32'sh2e8dedb3, 32'sh2e7cab1c, 32'sh2e6b615a, 
               32'sh2e5a1070, 32'sh2e48b860, 32'sh2e37592c, 32'sh2e25f2d8, 32'sh2e148566, 32'sh2e0310d9, 32'sh2df19534, 32'sh2de01278, 
               32'sh2dce88aa, 32'sh2dbcf7cb, 32'sh2dab5fdf, 32'sh2d99c0e7, 32'sh2d881ae8, 32'sh2d766de2, 32'sh2d64b9da, 32'sh2d52fed2, 
               32'sh2d413ccd, 32'sh2d2f73cd, 32'sh2d1da3d5, 32'sh2d0bcce8, 32'sh2cf9ef09, 32'sh2ce80a3a, 32'sh2cd61e7f, 32'sh2cc42bd9, 
               32'sh2cb2324c, 32'sh2ca031da, 32'sh2c8e2a87, 32'sh2c7c1c55, 32'sh2c6a0746, 32'sh2c57eb5e, 32'sh2c45c8a0, 32'sh2c339f0e, 
               32'sh2c216eaa, 32'sh2c0f3779, 32'sh2bfcf97c, 32'sh2beab4b6, 32'sh2bd8692b, 32'sh2bc616dd, 32'sh2bb3bdce, 32'sh2ba15e03, 
               32'sh2b8ef77d, 32'sh2b7c8a3f, 32'sh2b6a164d, 32'sh2b579ba8, 32'sh2b451a55, 32'sh2b329255, 32'sh2b2003ac, 32'sh2b0d6e5c, 
               32'sh2afad269, 32'sh2ae82fd5, 32'sh2ad586a3, 32'sh2ac2d6d6, 32'sh2ab02071, 32'sh2a9d6377, 32'sh2a8a9fea, 32'sh2a77d5ce, 
               32'sh2a650525, 32'sh2a522df3, 32'sh2a3f503a, 32'sh2a2c6bfd, 32'sh2a19813f, 32'sh2a069003, 32'sh29f3984c, 32'sh29e09a1c, 
               32'sh29cd9578, 32'sh29ba8a61, 32'sh29a778db, 32'sh299460e8, 32'sh2981428c, 32'sh296e1dc9, 32'sh295af2a3, 32'sh2947c11c, 
               32'sh29348937, 32'sh29214af8, 32'sh290e0661, 32'sh28fabb75, 32'sh28e76a37, 32'sh28d412ab, 32'sh28c0b4d2, 32'sh28ad50b1, 
               32'sh2899e64a, 32'sh288675a0, 32'sh2872feb6, 32'sh285f8190, 32'sh284bfe2f, 32'sh28387498, 32'sh2824e4cc, 32'sh28114ed0, 
               32'sh27fdb2a7, 32'sh27ea1052, 32'sh27d667d5, 32'sh27c2b934, 32'sh27af0472, 32'sh279b4990, 32'sh27878893, 32'sh2773c17d, 
               32'sh275ff452, 32'sh274c2115, 32'sh273847c8, 32'sh2724686e, 32'sh2710830c, 32'sh26fc97a3, 32'sh26e8a637, 32'sh26d4aecb, 
               32'sh26c0b162, 32'sh26acadff, 32'sh2698a4a6, 32'sh26849558, 32'sh2670801a, 32'sh265c64ef, 32'sh264843d9, 32'sh26341cdb, 
               32'sh261feffa, 32'sh260bbd37, 32'sh25f78497, 32'sh25e3461b, 32'sh25cf01c8, 32'sh25bab7a0, 32'sh25a667a7, 32'sh259211df, 
               32'sh257db64c, 32'sh256954f1, 32'sh2554edd1, 32'sh254080ef, 32'sh252c0e4f, 32'sh251795f3, 32'sh250317df, 32'sh24ee9415, 
               32'sh24da0a9a, 32'sh24c57b6f, 32'sh24b0e699, 32'sh249c4c1b, 32'sh2487abf7, 32'sh24730631, 32'sh245e5acc, 32'sh2449a9cc, 
               32'sh2434f332, 32'sh24203704, 32'sh240b7543, 32'sh23f6adf3, 32'sh23e1e117, 32'sh23cd0eb3, 32'sh23b836ca, 32'sh23a3595e, 
               32'sh238e7673, 32'sh23798e0d, 32'sh2364a02e, 32'sh234facda, 32'sh233ab414, 32'sh2325b5df, 32'sh2310b23e, 32'sh22fba936, 
               32'sh22e69ac8, 32'sh22d186f8, 32'sh22bc6dca, 32'sh22a74f40, 32'sh22922b5e, 32'sh227d0228, 32'sh2267d3a0, 32'sh22529fca, 
               32'sh223d66a8, 32'sh2228283f, 32'sh2212e492, 32'sh21fd9ba3, 32'sh21e84d76, 32'sh21d2fa0f, 32'sh21bda171, 32'sh21a8439e, 
               32'sh2192e09b, 32'sh217d786a, 32'sh21680b0f, 32'sh2152988d, 32'sh213d20e8, 32'sh2127a423, 32'sh21122240, 32'sh20fc9b44, 
               32'sh20e70f32, 32'sh20d17e0d, 32'sh20bbe7d8, 32'sh20a64c97, 32'sh2090ac4d, 32'sh207b06fe, 32'sh20655cac, 32'sh204fad5b, 
               32'sh2039f90f, 32'sh20243fca, 32'sh200e8190, 32'sh1ff8be65, 32'sh1fe2f64c, 32'sh1fcd2948, 32'sh1fb7575c, 32'sh1fa1808c, 
               32'sh1f8ba4dc, 32'sh1f75c44e, 32'sh1f5fdee6, 32'sh1f49f4a8, 32'sh1f340596, 32'sh1f1e11b5, 32'sh1f081907, 32'sh1ef21b90, 
               32'sh1edc1953, 32'sh1ec61254, 32'sh1eb00696, 32'sh1e99f61d, 32'sh1e83e0eb, 32'sh1e6dc705, 32'sh1e57a86d, 32'sh1e418528, 
               32'sh1e2b5d38, 32'sh1e1530a1, 32'sh1dfeff67, 32'sh1de8c98c, 32'sh1dd28f15, 32'sh1dbc5004, 32'sh1da60c5d, 32'sh1d8fc424, 
               32'sh1d79775c, 32'sh1d632608, 32'sh1d4cd02c, 32'sh1d3675cb, 32'sh1d2016e9, 32'sh1d09b389, 32'sh1cf34baf, 32'sh1cdcdf5e, 
               32'sh1cc66e99, 32'sh1caff965, 32'sh1c997fc4, 32'sh1c8301b9, 32'sh1c6c7f4a, 32'sh1c55f878, 32'sh1c3f6d47, 32'sh1c28ddbb, 
               32'sh1c1249d8, 32'sh1bfbb1a0, 32'sh1be51518, 32'sh1bce7442, 32'sh1bb7cf23, 32'sh1ba125bd, 32'sh1b8a7815, 32'sh1b73c62d, 
               32'sh1b5d100a, 32'sh1b4655ae, 32'sh1b2f971e, 32'sh1b18d45c, 32'sh1b020d6c, 32'sh1aeb4253, 32'sh1ad47312, 32'sh1abd9faf, 
               32'sh1aa6c82b, 32'sh1a8fec8c, 32'sh1a790cd4, 32'sh1a622907, 32'sh1a4b4128, 32'sh1a34553b, 32'sh1a1d6544, 32'sh1a067145, 
               32'sh19ef7944, 32'sh19d87d42, 32'sh19c17d44, 32'sh19aa794d, 32'sh19937161, 32'sh197c6584, 32'sh196555b8, 32'sh194e4201, 
               32'sh19372a64, 32'sh19200ee3, 32'sh1908ef82, 32'sh18f1cc45, 32'sh18daa52f, 32'sh18c37a44, 32'sh18ac4b87, 32'sh189518fc, 
               32'sh187de2a7, 32'sh1866a88a, 32'sh184f6aab, 32'sh1838290c, 32'sh1820e3b0, 32'sh18099a9c, 32'sh17f24dd3, 32'sh17dafd59, 
               32'sh17c3a931, 32'sh17ac515f, 32'sh1794f5e6, 32'sh177d96ca, 32'sh1766340f, 32'sh174ecdb8, 32'sh173763c9, 32'sh171ff646, 
               32'sh17088531, 32'sh16f1108f, 32'sh16d99864, 32'sh16c21cb2, 32'sh16aa9d7e, 32'sh16931acb, 32'sh167b949d, 32'sh16640af7, 
               32'sh164c7ddd, 32'sh1634ed53, 32'sh161d595d, 32'sh1605c1fd, 32'sh15ee2738, 32'sh15d68911, 32'sh15bee78c, 32'sh15a742ac, 
               32'sh158f9a76, 32'sh1577eeec, 32'sh15604013, 32'sh15488dee, 32'sh1530d881, 32'sh15191fcf, 32'sh150163dc, 32'sh14e9a4ac, 
               32'sh14d1e242, 32'sh14ba1ca3, 32'sh14a253d1, 32'sh148a87d1, 32'sh1472b8a5, 32'sh145ae653, 32'sh144310dd, 32'sh142b3846, 
               32'sh14135c94, 32'sh13fb7dc9, 32'sh13e39be9, 32'sh13cbb6f8, 32'sh13b3cefa, 32'sh139be3f2, 32'sh1383f5e3, 32'sh136c04d2, 
               32'sh135410c3, 32'sh133c19b8, 32'sh13241fb6, 32'sh130c22c1, 32'sh12f422db, 32'sh12dc2009, 32'sh12c41a4f, 32'sh12ac11af, 
               32'sh1294062f, 32'sh127bf7d1, 32'sh1263e699, 32'sh124bd28c, 32'sh1233bbac, 32'sh121ba1fd, 32'sh12038584, 32'sh11eb6643, 
               32'sh11d3443f, 32'sh11bb1f7c, 32'sh11a2f7fc, 32'sh118acdc4, 32'sh1172a0d7, 32'sh115a713a, 32'sh11423ef0, 32'sh112a09fc, 
               32'sh1111d263, 32'sh10f99827, 32'sh10e15b4e, 32'sh10c91bda, 32'sh10b0d9d0, 32'sh10989532, 32'sh10804e06, 32'sh1068044e, 
               32'sh104fb80e, 32'sh1037694b, 32'sh101f1807, 32'sh1006c446, 32'sh0fee6e0d, 32'sh0fd6155f, 32'sh0fbdba40, 32'sh0fa55cb4, 
               32'sh0f8cfcbe, 32'sh0f749a61, 32'sh0f5c35a3, 32'sh0f43ce86, 32'sh0f2b650f, 32'sh0f12f941, 32'sh0efa8b20, 32'sh0ee21aaf, 
               32'sh0ec9a7f3, 32'sh0eb132ef, 32'sh0e98bba7, 32'sh0e80421e, 32'sh0e67c65a, 32'sh0e4f485c, 32'sh0e36c82a, 32'sh0e1e45c6, 
               32'sh0e05c135, 32'sh0ded3a7b, 32'sh0dd4b19a, 32'sh0dbc2698, 32'sh0da39978, 32'sh0d8b0a3d, 32'sh0d7278eb, 32'sh0d59e586, 
               32'sh0d415013, 32'sh0d28b894, 32'sh0d101f0e, 32'sh0cf78383, 32'sh0cdee5f9, 32'sh0cc64673, 32'sh0cada4f5, 32'sh0c950182, 
               32'sh0c7c5c1e, 32'sh0c63b4ce, 32'sh0c4b0b94, 32'sh0c326075, 32'sh0c19b374, 32'sh0c010496, 32'sh0be853de, 32'sh0bcfa150, 
               32'sh0bb6ecef, 32'sh0b9e36c0, 32'sh0b857ec7, 32'sh0b6cc506, 32'sh0b540982, 32'sh0b3b4c40, 32'sh0b228d42, 32'sh0b09cc8c, 
               32'sh0af10a22, 32'sh0ad84609, 32'sh0abf8043, 32'sh0aa6b8d5, 32'sh0a8defc3, 32'sh0a752510, 32'sh0a5c58c0, 32'sh0a438ad7, 
               32'sh0a2abb59, 32'sh0a11ea49, 32'sh09f917ac, 32'sh09e04385, 32'sh09c76dd8, 32'sh09ae96aa, 32'sh0995bdfd, 32'sh097ce3d5, 
               32'sh09640837, 32'sh094b2b27, 32'sh09324ca7, 32'sh09196cbc, 32'sh09008b6a, 32'sh08e7a8b5, 32'sh08cec4a0, 32'sh08b5df30, 
               32'sh089cf867, 32'sh0884104b, 32'sh086b26de, 32'sh08523c25, 32'sh08395024, 32'sh082062de, 32'sh08077457, 32'sh07ee8493, 
               32'sh07d59396, 32'sh07bca163, 32'sh07a3adff, 32'sh078ab96e, 32'sh0771c3b3, 32'sh0758ccd2, 32'sh073fd4cf, 32'sh0726dbae, 
               32'sh070de172, 32'sh06f4e620, 32'sh06dbe9bb, 32'sh06c2ec48, 32'sh06a9edc9, 32'sh0690ee44, 32'sh0677edbb, 32'sh065eec33, 
               32'sh0645e9af, 32'sh062ce634, 32'sh0613e1c5, 32'sh05fadc66, 32'sh05e1d61b, 32'sh05c8cee7, 32'sh05afc6d0, 32'sh0596bdd7, 
               32'sh057db403, 32'sh0564a955, 32'sh054b9dd3, 32'sh0532917f, 32'sh0519845e, 32'sh05007674, 32'sh04e767c5, 32'sh04ce5854, 
               32'sh04b54825, 32'sh049c373c, 32'sh0483259d, 32'sh046a134c, 32'sh0451004d, 32'sh0437eca4, 32'sh041ed854, 32'sh0405c361, 
               32'sh03ecadcf, 32'sh03d397a3, 32'sh03ba80df, 32'sh03a16988, 32'sh038851a2, 32'sh036f3931, 32'sh03562038, 32'sh033d06bb, 
               32'sh0323ecbe, 32'sh030ad245, 32'sh02f1b755, 32'sh02d89bf0, 32'sh02bf801a, 32'sh02a663d8, 32'sh028d472e, 32'sh02742a1f, 
               32'sh025b0caf, 32'sh0241eee2, 32'sh0228d0bb, 32'sh020fb240, 32'sh01f69373, 32'sh01dd7459, 32'sh01c454f5, 32'sh01ab354b, 
               32'sh0192155f, 32'sh0178f536, 32'sh015fd4d2, 32'sh0146b438, 32'sh012d936c, 32'sh01147271, 32'sh00fb514b, 32'sh00e22fff, 
               32'sh00c90e90, 32'sh00afed02, 32'sh0096cb58, 32'sh007da998, 32'sh006487c4, 32'sh004b65e1, 32'sh003243f1, 32'sh001921fb, 
               32'sh00000000, 32'shffe6de05, 32'shffcdbc0f, 32'shffb49a1f, 32'shff9b783c, 32'shff825668, 32'shff6934a8, 32'shff5012fe, 
               32'shff36f170, 32'shff1dd001, 32'shff04aeb5, 32'shfeeb8d8f, 32'shfed26c94, 32'shfeb94bc8, 32'shfea02b2e, 32'shfe870aca, 
               32'shfe6deaa1, 32'shfe54cab5, 32'shfe3bab0b, 32'shfe228ba7, 32'shfe096c8d, 32'shfdf04dc0, 32'shfdd72f45, 32'shfdbe111e, 
               32'shfda4f351, 32'shfd8bd5e1, 32'shfd72b8d2, 32'shfd599c28, 32'shfd407fe6, 32'shfd276410, 32'shfd0e48ab, 32'shfcf52dbb, 
               32'shfcdc1342, 32'shfcc2f945, 32'shfca9dfc8, 32'shfc90c6cf, 32'shfc77ae5e, 32'shfc5e9678, 32'shfc457f21, 32'shfc2c685d, 
               32'shfc135231, 32'shfbfa3c9f, 32'shfbe127ac, 32'shfbc8135c, 32'shfbaeffb3, 32'shfb95ecb4, 32'shfb7cda63, 32'shfb63c8c4, 
               32'shfb4ab7db, 32'shfb31a7ac, 32'shfb18983b, 32'shfaff898c, 32'shfae67ba2, 32'shfacd6e81, 32'shfab4622d, 32'shfa9b56ab, 
               32'shfa824bfd, 32'shfa694229, 32'shfa503930, 32'shfa373119, 32'shfa1e29e5, 32'shfa05239a, 32'shf9ec1e3b, 32'shf9d319cc, 
               32'shf9ba1651, 32'shf9a113cd, 32'shf9881245, 32'shf96f11bc, 32'shf9561237, 32'shf93d13b8, 32'shf9241645, 32'shf90b19e0, 
               32'shf8f21e8e, 32'shf8d92452, 32'shf8c02b31, 32'shf8a7332e, 32'shf88e3c4d, 32'shf8754692, 32'shf85c5201, 32'shf8435e9d, 
               32'shf82a6c6a, 32'shf8117b6d, 32'shf7f88ba9, 32'shf7df9d22, 32'shf7c6afdc, 32'shf7adc3db, 32'shf794d922, 32'shf77befb5, 
               32'shf7630799, 32'shf74a20d0, 32'shf7313b60, 32'shf718574b, 32'shf6ff7496, 32'shf6e69344, 32'shf6cdb359, 32'shf6b4d4d9, 
               32'shf69bf7c9, 32'shf6831c2b, 32'shf66a4203, 32'shf6516956, 32'shf6389228, 32'shf61fbc7b, 32'shf606e854, 32'shf5ee15b7, 
               32'shf5d544a7, 32'shf5bc7529, 32'shf5a3a740, 32'shf58adaf0, 32'shf572103d, 32'shf559472b, 32'shf5407fbd, 32'shf527b9f7, 
               32'shf50ef5de, 32'shf4f63374, 32'shf4dd72be, 32'shf4c4b3c0, 32'shf4abf67e, 32'shf4933afa, 32'shf47a8139, 32'shf461c940, 
               32'shf4491311, 32'shf4305eb0, 32'shf417ac22, 32'shf3fefb6a, 32'shf3e64c8c, 32'shf3cd9f8b, 32'shf3b4f46c, 32'shf39c4b32, 
               32'shf383a3e2, 32'shf36afe7e, 32'shf3525b0b, 32'shf339b98d, 32'shf3211a07, 32'shf3087c7d, 32'shf2efe0f2, 32'shf2d7476c, 
               32'shf2beafed, 32'shf2a61a7a, 32'shf28d8715, 32'shf274f5c3, 32'shf25c6688, 32'shf243d968, 32'shf22b4e66, 32'shf212c585, 
               32'shf1fa3ecb, 32'shf1e1ba3a, 32'shf1c937d6, 32'shf1b0b7a4, 32'shf19839a6, 32'shf17fbde2, 32'shf1674459, 32'shf14ecd11, 
               32'shf136580d, 32'shf11de551, 32'shf10574e0, 32'shf0ed06bf, 32'shf0d49af1, 32'shf0bc317a, 32'shf0a3ca5d, 32'shf08b659f, 
               32'shf0730342, 32'shf05aa34c, 32'shf04245c0, 32'shf029eaa1, 32'shf01191f3, 32'sheff93bba, 32'shefe0e7f9, 32'shefc896b5, 
               32'shefb047f2, 32'shef97fbb2, 32'shef7fb1fa, 32'shef676ace, 32'shef4f2630, 32'shef36e426, 32'shef1ea4b2, 32'shef0667d9, 
               32'sheeee2d9d, 32'sheed5f604, 32'sheebdc110, 32'sheea58ec6, 32'shee8d5f29, 32'shee75323c, 32'shee5d0804, 32'shee44e084, 
               32'shee2cbbc1, 32'shee1499bd, 32'shedfc7a7c, 32'shede45e03, 32'shedcc4454, 32'shedb42d74, 32'shed9c1967, 32'shed84082f, 
               32'shed6bf9d1, 32'shed53ee51, 32'shed3be5b1, 32'shed23dff7, 32'shed0bdd25, 32'shecf3dd3f, 32'shecdbe04a, 32'shecc3e648, 
               32'shecabef3d, 32'shec93fb2e, 32'shec7c0a1d, 32'shec641c0e, 32'shec4c3106, 32'shec344908, 32'shec1c6417, 32'shec048237, 
               32'shebeca36c, 32'shebd4c7ba, 32'shebbcef23, 32'sheba519ad, 32'sheb8d475b, 32'sheb75782f, 32'sheb5dac2f, 32'sheb45e35d, 
               32'sheb2e1dbe, 32'sheb165b54, 32'sheafe9c24, 32'sheae6e031, 32'sheacf277f, 32'sheab77212, 32'shea9fbfed, 32'shea881114, 
               32'shea70658a, 32'shea58bd54, 32'shea411874, 32'shea2976ef, 32'shea11d8c8, 32'she9fa3e03, 32'she9e2a6a3, 32'she9cb12ad, 
               32'she9b38223, 32'she99bf509, 32'she9846b63, 32'she96ce535, 32'she9556282, 32'she93de34e, 32'she926679c, 32'she90eef71, 
               32'she8f77acf, 32'she8e009ba, 32'she8c89c37, 32'she8b13248, 32'she899cbf1, 32'she8826936, 32'she86b0a1a, 32'she853aea1, 
               32'she83c56cf, 32'she82502a7, 32'she80db22d, 32'she7f66564, 32'she7df1c50, 32'she7c7d6f4, 32'she7b09555, 32'she7995776, 
               32'she7821d59, 32'she76ae704, 32'she753b479, 32'she73c85bc, 32'she7255ad1, 32'she70e33bb, 32'she6f7107e, 32'she6dff11d, 
               32'she6c8d59c, 32'she6b1bdff, 32'she69aaa48, 32'she6839a7c, 32'she66c8e9f, 32'she65586b3, 32'she63e82bc, 32'she62782be, 
               32'she61086bc, 32'she5f98ebb, 32'she5e29abc, 32'she5cbaac5, 32'she5b4bed8, 32'she59dd6f9, 32'she586f32c, 32'she5701374, 
               32'she55937d5, 32'she5426051, 32'she52b8cee, 32'she514bdad, 32'she4fdf294, 32'she4e72ba4, 32'she4d068e2, 32'she4b9aa52, 
               32'she4a2eff6, 32'she48c39d3, 32'she47587eb, 32'she45eda43, 32'she44830dd, 32'she4318bbe, 32'she41aeae8, 32'she4044e60, 
               32'she3edb628, 32'she3d72245, 32'she3c092b9, 32'she3aa0788, 32'she39380b6, 32'she37cfe47, 32'she366803c, 32'she350069b, 
               32'she3399167, 32'she32320a2, 32'she30cb451, 32'she2f64c77, 32'she2dfe917, 32'she2c98a35, 32'she2b32fd4, 32'she29cd9f8, 
               32'she28688a4, 32'she2703bdc, 32'she259f3a3, 32'she243affc, 32'she22d70eb, 32'she2173674, 32'she2010099, 32'she1eacf5f, 
               32'she1d4a2c8, 32'she1be7ad8, 32'she1a85793, 32'she19238fb, 32'she17c1f15, 32'she16609e3, 32'she14ff96a, 32'she139edac, 
               32'she123e6ad, 32'she10de470, 32'she0f7e6f9, 32'she0e1ee4b, 32'she0cbfa6a, 32'she0b60b58, 32'she0a0211a, 32'she08a3bb2, 
               32'she0745b24, 32'she05e7f74, 32'she048a8a4, 32'she032d6b8, 32'she01d09b4, 32'she007419b, 32'shdff17e70, 32'shdfdbc036, 
               32'shdfc606f1, 32'shdfb052a5, 32'shdf9aa354, 32'shdf84f902, 32'shdf6f53b3, 32'shdf59b369, 32'shdf441828, 32'shdf2e81f3, 
               32'shdf18f0ce, 32'shdf0364bc, 32'shdeedddc0, 32'shded85bdd, 32'shdec2df18, 32'shdead6773, 32'shde97f4f1, 32'shde828796, 
               32'shde6d1f65, 32'shde57bc62, 32'shde425e8f, 32'shde2d05f1, 32'shde17b28a, 32'shde02645d, 32'shdded1b6e, 32'shddd7d7c1, 
               32'shddc29958, 32'shddad6036, 32'shdd982c60, 32'shdd82fdd8, 32'shdd6dd4a2, 32'shdd58b0c0, 32'shdd439236, 32'shdd2e7908, 
               32'shdd196538, 32'shdd0456ca, 32'shdcef4dc2, 32'shdcda4a21, 32'shdcc54bec, 32'shdcb05326, 32'shdc9b5fd2, 32'shdc8671f3, 
               32'shdc71898d, 32'shdc5ca6a2, 32'shdc47c936, 32'shdc32f14d, 32'shdc1e1ee9, 32'shdc09520d, 32'shdbf48abd, 32'shdbdfc8fc, 
               32'shdbcb0cce, 32'shdbb65634, 32'shdba1a534, 32'shdb8cf9cf, 32'shdb785409, 32'shdb63b3e5, 32'shdb4f1967, 32'shdb3a8491, 
               32'shdb25f566, 32'shdb116beb, 32'shdafce821, 32'shdae86a0d, 32'shdad3f1b1, 32'shdabf7f11, 32'shdaab122f, 32'shda96ab0f, 
               32'shda8249b4, 32'shda6dee21, 32'shda599859, 32'shda454860, 32'shda30fe38, 32'shda1cb9e5, 32'shda087b69, 32'shd9f442c9, 
               32'shd9e01006, 32'shd9cbe325, 32'shd9b7bc27, 32'shd9a39b11, 32'shd98f7fe6, 32'shd97b6aa8, 32'shd9675b5a, 32'shd9535201, 
               32'shd93f4e9e, 32'shd92b5135, 32'shd91759c9, 32'shd903685d, 32'shd8ef7cf4, 32'shd8db9792, 32'shd8c7b838, 32'shd8b3deeb, 
               32'shd8a00bae, 32'shd88c3e83, 32'shd878776d, 32'shd864b670, 32'shd850fb8e, 32'shd83d46cc, 32'shd829982b, 32'shd815efae, 
               32'shd8024d59, 32'shd7eeb130, 32'shd7db1b34, 32'shd7c78b68, 32'shd7b401d1, 32'shd7a07e70, 32'shd78d014a, 32'shd7798a60, 
               32'shd76619b6, 32'shd752af4f, 32'shd73f4b2e, 32'shd72bed55, 32'shd71895c9, 32'shd705448b, 32'shd6f1f99f, 32'shd6deb508, 
               32'shd6cb76c9, 32'shd6b83ee4, 32'shd6a50d5d, 32'shd691e237, 32'shd67ebd74, 32'shd66b9f18, 32'shd6588725, 32'shd645759f, 
               32'shd6326a88, 32'shd61f65e4, 32'shd60c67b4, 32'shd5f96ffd, 32'shd5e67ec1, 32'shd5d39403, 32'shd5c0afc6, 32'shd5add20d, 
               32'shd59afadb, 32'shd5882a32, 32'shd5756016, 32'shd5629c89, 32'shd54fdf8f, 32'shd53d292a, 32'shd52a795d, 32'shd517d02b, 
               32'shd5052d97, 32'shd4f291a4, 32'shd4dffc54, 32'shd4cd6dab, 32'shd4bae5ab, 32'shd4a86458, 32'shd495e9b3, 32'shd48375c1, 
               32'shd4710883, 32'shd45ea1fd, 32'shd44c4232, 32'shd439e923, 32'shd42796d5, 32'shd4154b4a, 32'shd4030684, 32'shd3f0c887, 
               32'shd3de9156, 32'shd3cc60f2, 32'shd3ba3760, 32'shd3a814a2, 32'shd395f8ba, 32'shd383e3ab, 32'shd371d579, 32'shd35fce26, 
               32'shd34dcdb4, 32'shd33bd427, 32'shd329e181, 32'shd317f5c6, 32'shd30610f7, 32'shd2f43318, 32'shd2e25c2b, 32'shd2d08c33, 
               32'shd2bec333, 32'shd2ad012e, 32'shd29b4626, 32'shd289921e, 32'shd277e518, 32'shd2663f19, 32'shd254a021, 32'shd2430835, 
               32'shd2317756, 32'shd21fed88, 32'shd20e6acc, 32'shd1fcef27, 32'shd1eb7a9a, 32'shd1da0d28, 32'shd1c8a6d4, 32'shd1b747a0, 
               32'shd1a5ef90, 32'shd1949ea6, 32'shd18354e4, 32'shd172124d, 32'shd160d6e5, 32'shd14fa2ad, 32'shd13e75a8, 32'shd12d4fd9, 
               32'shd11c3142, 32'shd10b19e7, 32'shd0fa09c9, 32'shd0e900ec, 32'shd0d7ff51, 32'shd0c704fd, 32'shd0b611f1, 32'shd0a5262f, 
               32'shd09441bb, 32'shd0836497, 32'shd0728ec6, 32'shd061c04a, 32'shd050f926, 32'shd040395d, 32'shd02f80f1, 32'shd01ecfe4, 
               32'shd00e2639, 32'shcffd83f4, 32'shcfece915, 32'shcfdc55a1, 32'shcfcbc999, 32'shcfbb4500, 32'shcfaac7d8, 32'shcf9a5225, 
               32'shcf89e3e8, 32'shcf797d24, 32'shcf691ddd, 32'shcf58c613, 32'shcf4875ca, 32'shcf382d05, 32'shcf27ebc5, 32'shcf17b20d, 
               32'shcf077fe1, 32'shcef75541, 32'shcee73231, 32'shced716b4, 32'shcec702cb, 32'shceb6f67a, 32'shcea6f1c2, 32'shce96f4a7, 
               32'shce86ff2a, 32'shce77114e, 32'shce672b16, 32'shce574c84, 32'shce47759a, 32'shce37a65b, 32'shce27dec9, 32'shce181ee8, 
               32'shce0866b8, 32'shcdf8b63d, 32'shcde90d79, 32'shcdd96c6f, 32'shcdc9d320, 32'shcdba4190, 32'shcdaab7c0, 32'shcd9b35b4, 
               32'shcd8bbb6d, 32'shcd7c48ee, 32'shcd6cde39, 32'shcd5d7b50, 32'shcd4e2037, 32'shcd3eccef, 32'shcd2f817b, 32'shcd203ddc, 
               32'shcd110216, 32'shcd01ce2b, 32'shccf2a21d, 32'shcce37def, 32'shccd461a2, 32'shccc54d3a, 32'shccb640b8, 32'shcca73c1e, 
               32'shcc983f70, 32'shcc894aaf, 32'shcc7a5dde, 32'shcc6b78ff, 32'shcc5c9c14, 32'shcc4dc720, 32'shcc3efa25, 32'shcc303524, 
               32'shcc217822, 32'shcc12c31f, 32'shcc04161e, 32'shcbf57121, 32'shcbe6d42b, 32'shcbd83f3d, 32'shcbc9b25a, 32'shcbbb2d85, 
               32'shcbacb0bf, 32'shcb9e3c0b, 32'shcb8fcf6b, 32'shcb816ae1, 32'shcb730e70, 32'shcb64ba19, 32'shcb566ddf, 32'shcb4829c4, 
               32'shcb39edca, 32'shcb2bb9f4, 32'shcb1d8e43, 32'shcb0f6aba, 32'shcb014f5b, 32'shcaf33c28, 32'shcae53123, 32'shcad72e4f, 
               32'shcac933ae, 32'shcabb4141, 32'shcaad570c, 32'shca9f750f, 32'shca919b4e, 32'shca83c9ca, 32'shca760086, 32'shca683f83, 
               32'shca5a86c4, 32'shca4cd64b, 32'shca3f2e19, 32'shca318e32, 32'shca23f698, 32'shca16674b, 32'shca08e04f, 32'shc9fb61a5, 
               32'shc9edeb50, 32'shc9e07d51, 32'shc9d317ab, 32'shc9c5ba60, 32'shc9b86572, 32'shc9ab18e3, 32'shc99dd4b4, 32'shc99098e9, 
               32'shc9836582, 32'shc9763a83, 32'shc96917ec, 32'shc95bfdc1, 32'shc94eec03, 32'shc941e2b4, 32'shc934e1d6, 32'shc927e96b, 
               32'shc91af976, 32'shc90e11f7, 32'shc90132f2, 32'shc8f45c68, 32'shc8e78e5b, 32'shc8dac8cd, 32'shc8ce0bc0, 32'shc8c15736, 
               32'shc8b4ab32, 32'shc8a807b4, 32'shc89b6cbf, 32'shc88eda54, 32'shc8825077, 32'shc875cf28, 32'shc869566a, 32'shc85ce63e, 
               32'shc8507ea7, 32'shc8441fa6, 32'shc837c93e, 32'shc82b7b70, 32'shc81f363d, 32'shc812f9a9, 32'shc806c5b5, 32'shc7fa9a62, 
               32'shc7ee77b3, 32'shc7e25daa, 32'shc7d64c47, 32'shc7ca438f, 32'shc7be4381, 32'shc7b24c20, 32'shc7a65d6e, 32'shc79a776c, 
               32'shc78e9a1d, 32'shc782c582, 32'shc776f99d, 32'shc76b3671, 32'shc75f7bfe, 32'shc753ca46, 32'shc748214c, 32'shc73c8111, 
               32'shc730e997, 32'shc7255ae0, 32'shc719d4ed, 32'shc70e57c0, 32'shc702e35c, 32'shc6f777c1, 32'shc6ec14f2, 32'shc6e0baf0, 
               32'shc6d569be, 32'shc6ca215c, 32'shc6bee1cd, 32'shc6b3ab12, 32'shc6a87d2d, 32'shc69d5820, 32'shc6923bec, 32'shc6872894, 
               32'shc67c1e18, 32'shc6711c7b, 32'shc66623be, 32'shc65b33e4, 32'shc6504ced, 32'shc6456edb, 32'shc63a99b1, 32'shc62fcd6f, 
               32'shc6250a18, 32'shc61a4fac, 32'shc60f9e2e, 32'shc604f5a0, 32'shc5fa5603, 32'shc5efbf58, 32'shc5e531a1, 32'shc5daace1, 
               32'shc5d03118, 32'shc5c5be47, 32'shc5bb5472, 32'shc5b0f399, 32'shc5a69bbe, 32'shc59c4ce3, 32'shc5920708, 32'shc587ca31, 
               32'shc57d965d, 32'shc5736b90, 32'shc56949ca, 32'shc55f310d, 32'shc555215a, 32'shc54b1ab4, 32'shc5411d1b, 32'shc5372891, 
               32'shc52d3d18, 32'shc5235ab2, 32'shc519815f, 32'shc50fb121, 32'shc505e9fb, 32'shc4fc2bec, 32'shc4f276f7, 32'shc4e8cb1e, 
               32'shc4df2862, 32'shc4d58ec3, 32'shc4cbfe45, 32'shc4c276e8, 32'shc4b8f8ad, 32'shc4af8397, 32'shc4a617a6, 32'shc49cb4dd, 
               32'shc4935b3c, 32'shc48a0ac4, 32'shc480c379, 32'shc477855a, 32'shc46e5069, 32'shc46524a9, 32'shc45c0219, 32'shc452e8bc, 
               32'shc449d892, 32'shc440d19e, 32'shc437d3e1, 32'shc42edf5c, 32'shc425f410, 32'shc41d11ff, 32'shc414392b, 32'shc40b6994, 
               32'shc402a33c, 32'shc3f9e624, 32'shc3f1324e, 32'shc3e887bb, 32'shc3dfe66c, 32'shc3d74e62, 32'shc3cebfa0, 32'shc3c63a26, 
               32'shc3bdbdf6, 32'shc3b54b11, 32'shc3ace178, 32'shc3a4812c, 32'shc39c2a2f, 32'shc393dc82, 32'shc38b9827, 32'shc3835d1e, 
               32'shc37b2b6a, 32'shc373030a, 32'shc36ae401, 32'shc362ce50, 32'shc35ac1f7, 32'shc352bef9, 32'shc34ac556, 32'shc342d510, 
               32'shc33aee27, 32'shc333109e, 32'shc32b3c75, 32'shc32371ae, 32'shc31bb049, 32'shc313f848, 32'shc30c49ad, 32'shc304a477, 
               32'shc2fd08a9, 32'shc2f57644, 32'shc2eded49, 32'shc2e66db8, 32'shc2def794, 32'shc2d78add, 32'shc2d02794, 32'shc2c8cdbb, 
               32'shc2c17d52, 32'shc2ba365c, 32'shc2b2f8d8, 32'shc2abc4c9, 32'shc2a49a2e, 32'shc29d790a, 32'shc296615d, 32'shc28f5329, 
               32'shc2884e6e, 32'shc281532e, 32'shc27a616a, 32'shc2737922, 32'shc26c9a58, 32'shc265c50e, 32'shc25ef943, 32'shc25836f9, 
               32'shc2517e31, 32'shc24aceed, 32'shc244292c, 32'shc23d8cf1, 32'shc236fa3b, 32'shc230710d, 32'shc229f167, 32'shc2237b4b, 
               32'shc21d0eb8, 32'shc216abb1, 32'shc2105236, 32'shc20a0248, 32'shc203bbe8, 32'shc1fd7f17, 32'shc1f74bd6, 32'shc1f12227, 
               32'shc1eb0209, 32'shc1e4eb7e, 32'shc1dede87, 32'shc1d8db25, 32'shc1d2e158, 32'shc1ccf122, 32'shc1c70a84, 32'shc1c12d7e, 
               32'shc1bb5a11, 32'shc1b5903f, 32'shc1afd007, 32'shc1aa196c, 32'shc1a46c6e, 32'shc19ec90d, 32'shc1992f4c, 32'shc1939f29, 
               32'shc18e18a7, 32'shc1889bc6, 32'shc1832888, 32'shc17dbeec, 32'shc1785ef4, 32'shc17308a1, 32'shc16dbbf3, 32'shc16878eb, 
               32'shc1633f8a, 32'shc15e0fd1, 32'shc158e9c1, 32'shc153cd5a, 32'shc14eba9d, 32'shc149b18b, 32'shc144b225, 32'shc13fbc6c, 
               32'shc13ad060, 32'shc135ee02, 32'shc1311553, 32'shc12c4653, 32'shc1278104, 32'shc122c566, 32'shc11e1379, 32'shc1196b3f, 
               32'shc114ccb9, 32'shc11037e6, 32'shc10bacc8, 32'shc1072b5f, 32'shc102b3ac, 32'shc0fe45b0, 32'shc0f9e16b, 32'shc0f586df, 
               32'shc0f1360b, 32'shc0eceef1, 32'shc0e8b190, 32'shc0e47deb, 32'shc0e05401, 32'shc0dc33d2, 32'shc0d81d61, 32'shc0d410ad, 
               32'shc0d00db6, 32'shc0cc147f, 32'shc0c82506, 32'shc0c43f4d, 32'shc0c06355, 32'shc0bc911d, 32'shc0b8c8a7, 32'shc0b509f3, 
               32'shc0b15502, 32'shc0ada9d4, 32'shc0aa086a, 32'shc0a670c4, 32'shc0a2e2e3, 32'shc09f5ec8, 32'shc09be473, 32'shc09873e4, 
               32'shc0950d1d, 32'shc091b01d, 32'shc08e5ce5, 32'shc08b1376, 32'shc087d3d0, 32'shc0849df4, 32'shc08171e2, 32'shc07e4f9b, 
               32'shc07b371e, 32'shc078286e, 32'shc0752389, 32'shc0722871, 32'shc06f3726, 32'shc06c4fa8, 32'shc06971f9, 32'shc0669e18, 
               32'shc063d405, 32'shc06113c2, 32'shc05e5d4e, 32'shc05bb0ab, 32'shc0590dd8, 32'shc05674d6, 32'shc053e5a5, 32'shc0516045, 
               32'shc04ee4b8, 32'shc04c72fe, 32'shc04a0b16, 32'shc047ad01, 32'shc04558c0, 32'shc0430e53, 32'shc040cdba, 32'shc03e96f6, 
               32'shc03c6a07, 32'shc03a46ed, 32'shc0382da8, 32'shc0361e3a, 32'shc03418a2, 32'shc0321ce0, 32'shc0302af5, 32'shc02e42e2, 
               32'shc02c64a6, 32'shc02a9042, 32'shc028c5b6, 32'shc0270502, 32'shc0254e27, 32'shc023a124, 32'shc021fdfb, 32'shc02064ab, 
               32'shc01ed535, 32'shc01d4f99, 32'shc01bd3d6, 32'shc01a61ee, 32'shc018f9e1, 32'shc0179bae, 32'shc0164757, 32'shc014fcda, 
               32'shc013bc39, 32'shc0128574, 32'shc011588a, 32'shc010357c, 32'shc00f1c4a, 32'shc00e0cf5, 32'shc00d077c, 32'shc00c0be0, 
               32'shc00b1a20, 32'shc00a323d, 32'shc0095438, 32'shc008800f, 32'shc007b5c4, 32'shc006f556, 32'shc0063ec6, 32'shc0059214, 
               32'shc004ef3f, 32'shc0045648, 32'shc003c72f, 32'shc00341f4, 32'shc002c697, 32'shc0025519, 32'shc001ed78, 32'shc0018fb6, 
               32'shc0013bd3, 32'shc000f1ce, 32'shc000b1a7, 32'shc0007b5f, 32'shc0004ef5, 32'shc0002c6a, 32'shc00013bd, 32'shc00004ef
            };

            reg signed [31:0] W_Im_table[2048] = '{
               32'sh00000000, 32'shffe6de05, 32'shffcdbc0f, 32'shffb49a1f, 32'shff9b783c, 32'shff825668, 32'shff6934a8, 32'shff5012fe, 
               32'shff36f170, 32'shff1dd001, 32'shff04aeb5, 32'shfeeb8d8f, 32'shfed26c94, 32'shfeb94bc8, 32'shfea02b2e, 32'shfe870aca, 
               32'shfe6deaa1, 32'shfe54cab5, 32'shfe3bab0b, 32'shfe228ba7, 32'shfe096c8d, 32'shfdf04dc0, 32'shfdd72f45, 32'shfdbe111e, 
               32'shfda4f351, 32'shfd8bd5e1, 32'shfd72b8d2, 32'shfd599c28, 32'shfd407fe6, 32'shfd276410, 32'shfd0e48ab, 32'shfcf52dbb, 
               32'shfcdc1342, 32'shfcc2f945, 32'shfca9dfc8, 32'shfc90c6cf, 32'shfc77ae5e, 32'shfc5e9678, 32'shfc457f21, 32'shfc2c685d, 
               32'shfc135231, 32'shfbfa3c9f, 32'shfbe127ac, 32'shfbc8135c, 32'shfbaeffb3, 32'shfb95ecb4, 32'shfb7cda63, 32'shfb63c8c4, 
               32'shfb4ab7db, 32'shfb31a7ac, 32'shfb18983b, 32'shfaff898c, 32'shfae67ba2, 32'shfacd6e81, 32'shfab4622d, 32'shfa9b56ab, 
               32'shfa824bfd, 32'shfa694229, 32'shfa503930, 32'shfa373119, 32'shfa1e29e5, 32'shfa05239a, 32'shf9ec1e3b, 32'shf9d319cc, 
               32'shf9ba1651, 32'shf9a113cd, 32'shf9881245, 32'shf96f11bc, 32'shf9561237, 32'shf93d13b8, 32'shf9241645, 32'shf90b19e0, 
               32'shf8f21e8e, 32'shf8d92452, 32'shf8c02b31, 32'shf8a7332e, 32'shf88e3c4d, 32'shf8754692, 32'shf85c5201, 32'shf8435e9d, 
               32'shf82a6c6a, 32'shf8117b6d, 32'shf7f88ba9, 32'shf7df9d22, 32'shf7c6afdc, 32'shf7adc3db, 32'shf794d922, 32'shf77befb5, 
               32'shf7630799, 32'shf74a20d0, 32'shf7313b60, 32'shf718574b, 32'shf6ff7496, 32'shf6e69344, 32'shf6cdb359, 32'shf6b4d4d9, 
               32'shf69bf7c9, 32'shf6831c2b, 32'shf66a4203, 32'shf6516956, 32'shf6389228, 32'shf61fbc7b, 32'shf606e854, 32'shf5ee15b7, 
               32'shf5d544a7, 32'shf5bc7529, 32'shf5a3a740, 32'shf58adaf0, 32'shf572103d, 32'shf559472b, 32'shf5407fbd, 32'shf527b9f7, 
               32'shf50ef5de, 32'shf4f63374, 32'shf4dd72be, 32'shf4c4b3c0, 32'shf4abf67e, 32'shf4933afa, 32'shf47a8139, 32'shf461c940, 
               32'shf4491311, 32'shf4305eb0, 32'shf417ac22, 32'shf3fefb6a, 32'shf3e64c8c, 32'shf3cd9f8b, 32'shf3b4f46c, 32'shf39c4b32, 
               32'shf383a3e2, 32'shf36afe7e, 32'shf3525b0b, 32'shf339b98d, 32'shf3211a07, 32'shf3087c7d, 32'shf2efe0f2, 32'shf2d7476c, 
               32'shf2beafed, 32'shf2a61a7a, 32'shf28d8715, 32'shf274f5c3, 32'shf25c6688, 32'shf243d968, 32'shf22b4e66, 32'shf212c585, 
               32'shf1fa3ecb, 32'shf1e1ba3a, 32'shf1c937d6, 32'shf1b0b7a4, 32'shf19839a6, 32'shf17fbde2, 32'shf1674459, 32'shf14ecd11, 
               32'shf136580d, 32'shf11de551, 32'shf10574e0, 32'shf0ed06bf, 32'shf0d49af1, 32'shf0bc317a, 32'shf0a3ca5d, 32'shf08b659f, 
               32'shf0730342, 32'shf05aa34c, 32'shf04245c0, 32'shf029eaa1, 32'shf01191f3, 32'sheff93bba, 32'shefe0e7f9, 32'shefc896b5, 
               32'shefb047f2, 32'shef97fbb2, 32'shef7fb1fa, 32'shef676ace, 32'shef4f2630, 32'shef36e426, 32'shef1ea4b2, 32'shef0667d9, 
               32'sheeee2d9d, 32'sheed5f604, 32'sheebdc110, 32'sheea58ec6, 32'shee8d5f29, 32'shee75323c, 32'shee5d0804, 32'shee44e084, 
               32'shee2cbbc1, 32'shee1499bd, 32'shedfc7a7c, 32'shede45e03, 32'shedcc4454, 32'shedb42d74, 32'shed9c1967, 32'shed84082f, 
               32'shed6bf9d1, 32'shed53ee51, 32'shed3be5b1, 32'shed23dff7, 32'shed0bdd25, 32'shecf3dd3f, 32'shecdbe04a, 32'shecc3e648, 
               32'shecabef3d, 32'shec93fb2e, 32'shec7c0a1d, 32'shec641c0e, 32'shec4c3106, 32'shec344908, 32'shec1c6417, 32'shec048237, 
               32'shebeca36c, 32'shebd4c7ba, 32'shebbcef23, 32'sheba519ad, 32'sheb8d475b, 32'sheb75782f, 32'sheb5dac2f, 32'sheb45e35d, 
               32'sheb2e1dbe, 32'sheb165b54, 32'sheafe9c24, 32'sheae6e031, 32'sheacf277f, 32'sheab77212, 32'shea9fbfed, 32'shea881114, 
               32'shea70658a, 32'shea58bd54, 32'shea411874, 32'shea2976ef, 32'shea11d8c8, 32'she9fa3e03, 32'she9e2a6a3, 32'she9cb12ad, 
               32'she9b38223, 32'she99bf509, 32'she9846b63, 32'she96ce535, 32'she9556282, 32'she93de34e, 32'she926679c, 32'she90eef71, 
               32'she8f77acf, 32'she8e009ba, 32'she8c89c37, 32'she8b13248, 32'she899cbf1, 32'she8826936, 32'she86b0a1a, 32'she853aea1, 
               32'she83c56cf, 32'she82502a7, 32'she80db22d, 32'she7f66564, 32'she7df1c50, 32'she7c7d6f4, 32'she7b09555, 32'she7995776, 
               32'she7821d59, 32'she76ae704, 32'she753b479, 32'she73c85bc, 32'she7255ad1, 32'she70e33bb, 32'she6f7107e, 32'she6dff11d, 
               32'she6c8d59c, 32'she6b1bdff, 32'she69aaa48, 32'she6839a7c, 32'she66c8e9f, 32'she65586b3, 32'she63e82bc, 32'she62782be, 
               32'she61086bc, 32'she5f98ebb, 32'she5e29abc, 32'she5cbaac5, 32'she5b4bed8, 32'she59dd6f9, 32'she586f32c, 32'she5701374, 
               32'she55937d5, 32'she5426051, 32'she52b8cee, 32'she514bdad, 32'she4fdf294, 32'she4e72ba4, 32'she4d068e2, 32'she4b9aa52, 
               32'she4a2eff6, 32'she48c39d3, 32'she47587eb, 32'she45eda43, 32'she44830dd, 32'she4318bbe, 32'she41aeae8, 32'she4044e60, 
               32'she3edb628, 32'she3d72245, 32'she3c092b9, 32'she3aa0788, 32'she39380b6, 32'she37cfe47, 32'she366803c, 32'she350069b, 
               32'she3399167, 32'she32320a2, 32'she30cb451, 32'she2f64c77, 32'she2dfe917, 32'she2c98a35, 32'she2b32fd4, 32'she29cd9f8, 
               32'she28688a4, 32'she2703bdc, 32'she259f3a3, 32'she243affc, 32'she22d70eb, 32'she2173674, 32'she2010099, 32'she1eacf5f, 
               32'she1d4a2c8, 32'she1be7ad8, 32'she1a85793, 32'she19238fb, 32'she17c1f15, 32'she16609e3, 32'she14ff96a, 32'she139edac, 
               32'she123e6ad, 32'she10de470, 32'she0f7e6f9, 32'she0e1ee4b, 32'she0cbfa6a, 32'she0b60b58, 32'she0a0211a, 32'she08a3bb2, 
               32'she0745b24, 32'she05e7f74, 32'she048a8a4, 32'she032d6b8, 32'she01d09b4, 32'she007419b, 32'shdff17e70, 32'shdfdbc036, 
               32'shdfc606f1, 32'shdfb052a5, 32'shdf9aa354, 32'shdf84f902, 32'shdf6f53b3, 32'shdf59b369, 32'shdf441828, 32'shdf2e81f3, 
               32'shdf18f0ce, 32'shdf0364bc, 32'shdeedddc0, 32'shded85bdd, 32'shdec2df18, 32'shdead6773, 32'shde97f4f1, 32'shde828796, 
               32'shde6d1f65, 32'shde57bc62, 32'shde425e8f, 32'shde2d05f1, 32'shde17b28a, 32'shde02645d, 32'shdded1b6e, 32'shddd7d7c1, 
               32'shddc29958, 32'shddad6036, 32'shdd982c60, 32'shdd82fdd8, 32'shdd6dd4a2, 32'shdd58b0c0, 32'shdd439236, 32'shdd2e7908, 
               32'shdd196538, 32'shdd0456ca, 32'shdcef4dc2, 32'shdcda4a21, 32'shdcc54bec, 32'shdcb05326, 32'shdc9b5fd2, 32'shdc8671f3, 
               32'shdc71898d, 32'shdc5ca6a2, 32'shdc47c936, 32'shdc32f14d, 32'shdc1e1ee9, 32'shdc09520d, 32'shdbf48abd, 32'shdbdfc8fc, 
               32'shdbcb0cce, 32'shdbb65634, 32'shdba1a534, 32'shdb8cf9cf, 32'shdb785409, 32'shdb63b3e5, 32'shdb4f1967, 32'shdb3a8491, 
               32'shdb25f566, 32'shdb116beb, 32'shdafce821, 32'shdae86a0d, 32'shdad3f1b1, 32'shdabf7f11, 32'shdaab122f, 32'shda96ab0f, 
               32'shda8249b4, 32'shda6dee21, 32'shda599859, 32'shda454860, 32'shda30fe38, 32'shda1cb9e5, 32'shda087b69, 32'shd9f442c9, 
               32'shd9e01006, 32'shd9cbe325, 32'shd9b7bc27, 32'shd9a39b11, 32'shd98f7fe6, 32'shd97b6aa8, 32'shd9675b5a, 32'shd9535201, 
               32'shd93f4e9e, 32'shd92b5135, 32'shd91759c9, 32'shd903685d, 32'shd8ef7cf4, 32'shd8db9792, 32'shd8c7b838, 32'shd8b3deeb, 
               32'shd8a00bae, 32'shd88c3e83, 32'shd878776d, 32'shd864b670, 32'shd850fb8e, 32'shd83d46cc, 32'shd829982b, 32'shd815efae, 
               32'shd8024d59, 32'shd7eeb130, 32'shd7db1b34, 32'shd7c78b68, 32'shd7b401d1, 32'shd7a07e70, 32'shd78d014a, 32'shd7798a60, 
               32'shd76619b6, 32'shd752af4f, 32'shd73f4b2e, 32'shd72bed55, 32'shd71895c9, 32'shd705448b, 32'shd6f1f99f, 32'shd6deb508, 
               32'shd6cb76c9, 32'shd6b83ee4, 32'shd6a50d5d, 32'shd691e237, 32'shd67ebd74, 32'shd66b9f18, 32'shd6588725, 32'shd645759f, 
               32'shd6326a88, 32'shd61f65e4, 32'shd60c67b4, 32'shd5f96ffd, 32'shd5e67ec1, 32'shd5d39403, 32'shd5c0afc6, 32'shd5add20d, 
               32'shd59afadb, 32'shd5882a32, 32'shd5756016, 32'shd5629c89, 32'shd54fdf8f, 32'shd53d292a, 32'shd52a795d, 32'shd517d02b, 
               32'shd5052d97, 32'shd4f291a4, 32'shd4dffc54, 32'shd4cd6dab, 32'shd4bae5ab, 32'shd4a86458, 32'shd495e9b3, 32'shd48375c1, 
               32'shd4710883, 32'shd45ea1fd, 32'shd44c4232, 32'shd439e923, 32'shd42796d5, 32'shd4154b4a, 32'shd4030684, 32'shd3f0c887, 
               32'shd3de9156, 32'shd3cc60f2, 32'shd3ba3760, 32'shd3a814a2, 32'shd395f8ba, 32'shd383e3ab, 32'shd371d579, 32'shd35fce26, 
               32'shd34dcdb4, 32'shd33bd427, 32'shd329e181, 32'shd317f5c6, 32'shd30610f7, 32'shd2f43318, 32'shd2e25c2b, 32'shd2d08c33, 
               32'shd2bec333, 32'shd2ad012e, 32'shd29b4626, 32'shd289921e, 32'shd277e518, 32'shd2663f19, 32'shd254a021, 32'shd2430835, 
               32'shd2317756, 32'shd21fed88, 32'shd20e6acc, 32'shd1fcef27, 32'shd1eb7a9a, 32'shd1da0d28, 32'shd1c8a6d4, 32'shd1b747a0, 
               32'shd1a5ef90, 32'shd1949ea6, 32'shd18354e4, 32'shd172124d, 32'shd160d6e5, 32'shd14fa2ad, 32'shd13e75a8, 32'shd12d4fd9, 
               32'shd11c3142, 32'shd10b19e7, 32'shd0fa09c9, 32'shd0e900ec, 32'shd0d7ff51, 32'shd0c704fd, 32'shd0b611f1, 32'shd0a5262f, 
               32'shd09441bb, 32'shd0836497, 32'shd0728ec6, 32'shd061c04a, 32'shd050f926, 32'shd040395d, 32'shd02f80f1, 32'shd01ecfe4, 
               32'shd00e2639, 32'shcffd83f4, 32'shcfece915, 32'shcfdc55a1, 32'shcfcbc999, 32'shcfbb4500, 32'shcfaac7d8, 32'shcf9a5225, 
               32'shcf89e3e8, 32'shcf797d24, 32'shcf691ddd, 32'shcf58c613, 32'shcf4875ca, 32'shcf382d05, 32'shcf27ebc5, 32'shcf17b20d, 
               32'shcf077fe1, 32'shcef75541, 32'shcee73231, 32'shced716b4, 32'shcec702cb, 32'shceb6f67a, 32'shcea6f1c2, 32'shce96f4a7, 
               32'shce86ff2a, 32'shce77114e, 32'shce672b16, 32'shce574c84, 32'shce47759a, 32'shce37a65b, 32'shce27dec9, 32'shce181ee8, 
               32'shce0866b8, 32'shcdf8b63d, 32'shcde90d79, 32'shcdd96c6f, 32'shcdc9d320, 32'shcdba4190, 32'shcdaab7c0, 32'shcd9b35b4, 
               32'shcd8bbb6d, 32'shcd7c48ee, 32'shcd6cde39, 32'shcd5d7b50, 32'shcd4e2037, 32'shcd3eccef, 32'shcd2f817b, 32'shcd203ddc, 
               32'shcd110216, 32'shcd01ce2b, 32'shccf2a21d, 32'shcce37def, 32'shccd461a2, 32'shccc54d3a, 32'shccb640b8, 32'shcca73c1e, 
               32'shcc983f70, 32'shcc894aaf, 32'shcc7a5dde, 32'shcc6b78ff, 32'shcc5c9c14, 32'shcc4dc720, 32'shcc3efa25, 32'shcc303524, 
               32'shcc217822, 32'shcc12c31f, 32'shcc04161e, 32'shcbf57121, 32'shcbe6d42b, 32'shcbd83f3d, 32'shcbc9b25a, 32'shcbbb2d85, 
               32'shcbacb0bf, 32'shcb9e3c0b, 32'shcb8fcf6b, 32'shcb816ae1, 32'shcb730e70, 32'shcb64ba19, 32'shcb566ddf, 32'shcb4829c4, 
               32'shcb39edca, 32'shcb2bb9f4, 32'shcb1d8e43, 32'shcb0f6aba, 32'shcb014f5b, 32'shcaf33c28, 32'shcae53123, 32'shcad72e4f, 
               32'shcac933ae, 32'shcabb4141, 32'shcaad570c, 32'shca9f750f, 32'shca919b4e, 32'shca83c9ca, 32'shca760086, 32'shca683f83, 
               32'shca5a86c4, 32'shca4cd64b, 32'shca3f2e19, 32'shca318e32, 32'shca23f698, 32'shca16674b, 32'shca08e04f, 32'shc9fb61a5, 
               32'shc9edeb50, 32'shc9e07d51, 32'shc9d317ab, 32'shc9c5ba60, 32'shc9b86572, 32'shc9ab18e3, 32'shc99dd4b4, 32'shc99098e9, 
               32'shc9836582, 32'shc9763a83, 32'shc96917ec, 32'shc95bfdc1, 32'shc94eec03, 32'shc941e2b4, 32'shc934e1d6, 32'shc927e96b, 
               32'shc91af976, 32'shc90e11f7, 32'shc90132f2, 32'shc8f45c68, 32'shc8e78e5b, 32'shc8dac8cd, 32'shc8ce0bc0, 32'shc8c15736, 
               32'shc8b4ab32, 32'shc8a807b4, 32'shc89b6cbf, 32'shc88eda54, 32'shc8825077, 32'shc875cf28, 32'shc869566a, 32'shc85ce63e, 
               32'shc8507ea7, 32'shc8441fa6, 32'shc837c93e, 32'shc82b7b70, 32'shc81f363d, 32'shc812f9a9, 32'shc806c5b5, 32'shc7fa9a62, 
               32'shc7ee77b3, 32'shc7e25daa, 32'shc7d64c47, 32'shc7ca438f, 32'shc7be4381, 32'shc7b24c20, 32'shc7a65d6e, 32'shc79a776c, 
               32'shc78e9a1d, 32'shc782c582, 32'shc776f99d, 32'shc76b3671, 32'shc75f7bfe, 32'shc753ca46, 32'shc748214c, 32'shc73c8111, 
               32'shc730e997, 32'shc7255ae0, 32'shc719d4ed, 32'shc70e57c0, 32'shc702e35c, 32'shc6f777c1, 32'shc6ec14f2, 32'shc6e0baf0, 
               32'shc6d569be, 32'shc6ca215c, 32'shc6bee1cd, 32'shc6b3ab12, 32'shc6a87d2d, 32'shc69d5820, 32'shc6923bec, 32'shc6872894, 
               32'shc67c1e18, 32'shc6711c7b, 32'shc66623be, 32'shc65b33e4, 32'shc6504ced, 32'shc6456edb, 32'shc63a99b1, 32'shc62fcd6f, 
               32'shc6250a18, 32'shc61a4fac, 32'shc60f9e2e, 32'shc604f5a0, 32'shc5fa5603, 32'shc5efbf58, 32'shc5e531a1, 32'shc5daace1, 
               32'shc5d03118, 32'shc5c5be47, 32'shc5bb5472, 32'shc5b0f399, 32'shc5a69bbe, 32'shc59c4ce3, 32'shc5920708, 32'shc587ca31, 
               32'shc57d965d, 32'shc5736b90, 32'shc56949ca, 32'shc55f310d, 32'shc555215a, 32'shc54b1ab4, 32'shc5411d1b, 32'shc5372891, 
               32'shc52d3d18, 32'shc5235ab2, 32'shc519815f, 32'shc50fb121, 32'shc505e9fb, 32'shc4fc2bec, 32'shc4f276f7, 32'shc4e8cb1e, 
               32'shc4df2862, 32'shc4d58ec3, 32'shc4cbfe45, 32'shc4c276e8, 32'shc4b8f8ad, 32'shc4af8397, 32'shc4a617a6, 32'shc49cb4dd, 
               32'shc4935b3c, 32'shc48a0ac4, 32'shc480c379, 32'shc477855a, 32'shc46e5069, 32'shc46524a9, 32'shc45c0219, 32'shc452e8bc, 
               32'shc449d892, 32'shc440d19e, 32'shc437d3e1, 32'shc42edf5c, 32'shc425f410, 32'shc41d11ff, 32'shc414392b, 32'shc40b6994, 
               32'shc402a33c, 32'shc3f9e624, 32'shc3f1324e, 32'shc3e887bb, 32'shc3dfe66c, 32'shc3d74e62, 32'shc3cebfa0, 32'shc3c63a26, 
               32'shc3bdbdf6, 32'shc3b54b11, 32'shc3ace178, 32'shc3a4812c, 32'shc39c2a2f, 32'shc393dc82, 32'shc38b9827, 32'shc3835d1e, 
               32'shc37b2b6a, 32'shc373030a, 32'shc36ae401, 32'shc362ce50, 32'shc35ac1f7, 32'shc352bef9, 32'shc34ac556, 32'shc342d510, 
               32'shc33aee27, 32'shc333109e, 32'shc32b3c75, 32'shc32371ae, 32'shc31bb049, 32'shc313f848, 32'shc30c49ad, 32'shc304a477, 
               32'shc2fd08a9, 32'shc2f57644, 32'shc2eded49, 32'shc2e66db8, 32'shc2def794, 32'shc2d78add, 32'shc2d02794, 32'shc2c8cdbb, 
               32'shc2c17d52, 32'shc2ba365c, 32'shc2b2f8d8, 32'shc2abc4c9, 32'shc2a49a2e, 32'shc29d790a, 32'shc296615d, 32'shc28f5329, 
               32'shc2884e6e, 32'shc281532e, 32'shc27a616a, 32'shc2737922, 32'shc26c9a58, 32'shc265c50e, 32'shc25ef943, 32'shc25836f9, 
               32'shc2517e31, 32'shc24aceed, 32'shc244292c, 32'shc23d8cf1, 32'shc236fa3b, 32'shc230710d, 32'shc229f167, 32'shc2237b4b, 
               32'shc21d0eb8, 32'shc216abb1, 32'shc2105236, 32'shc20a0248, 32'shc203bbe8, 32'shc1fd7f17, 32'shc1f74bd6, 32'shc1f12227, 
               32'shc1eb0209, 32'shc1e4eb7e, 32'shc1dede87, 32'shc1d8db25, 32'shc1d2e158, 32'shc1ccf122, 32'shc1c70a84, 32'shc1c12d7e, 
               32'shc1bb5a11, 32'shc1b5903f, 32'shc1afd007, 32'shc1aa196c, 32'shc1a46c6e, 32'shc19ec90d, 32'shc1992f4c, 32'shc1939f29, 
               32'shc18e18a7, 32'shc1889bc6, 32'shc1832888, 32'shc17dbeec, 32'shc1785ef4, 32'shc17308a1, 32'shc16dbbf3, 32'shc16878eb, 
               32'shc1633f8a, 32'shc15e0fd1, 32'shc158e9c1, 32'shc153cd5a, 32'shc14eba9d, 32'shc149b18b, 32'shc144b225, 32'shc13fbc6c, 
               32'shc13ad060, 32'shc135ee02, 32'shc1311553, 32'shc12c4653, 32'shc1278104, 32'shc122c566, 32'shc11e1379, 32'shc1196b3f, 
               32'shc114ccb9, 32'shc11037e6, 32'shc10bacc8, 32'shc1072b5f, 32'shc102b3ac, 32'shc0fe45b0, 32'shc0f9e16b, 32'shc0f586df, 
               32'shc0f1360b, 32'shc0eceef1, 32'shc0e8b190, 32'shc0e47deb, 32'shc0e05401, 32'shc0dc33d2, 32'shc0d81d61, 32'shc0d410ad, 
               32'shc0d00db6, 32'shc0cc147f, 32'shc0c82506, 32'shc0c43f4d, 32'shc0c06355, 32'shc0bc911d, 32'shc0b8c8a7, 32'shc0b509f3, 
               32'shc0b15502, 32'shc0ada9d4, 32'shc0aa086a, 32'shc0a670c4, 32'shc0a2e2e3, 32'shc09f5ec8, 32'shc09be473, 32'shc09873e4, 
               32'shc0950d1d, 32'shc091b01d, 32'shc08e5ce5, 32'shc08b1376, 32'shc087d3d0, 32'shc0849df4, 32'shc08171e2, 32'shc07e4f9b, 
               32'shc07b371e, 32'shc078286e, 32'shc0752389, 32'shc0722871, 32'shc06f3726, 32'shc06c4fa8, 32'shc06971f9, 32'shc0669e18, 
               32'shc063d405, 32'shc06113c2, 32'shc05e5d4e, 32'shc05bb0ab, 32'shc0590dd8, 32'shc05674d6, 32'shc053e5a5, 32'shc0516045, 
               32'shc04ee4b8, 32'shc04c72fe, 32'shc04a0b16, 32'shc047ad01, 32'shc04558c0, 32'shc0430e53, 32'shc040cdba, 32'shc03e96f6, 
               32'shc03c6a07, 32'shc03a46ed, 32'shc0382da8, 32'shc0361e3a, 32'shc03418a2, 32'shc0321ce0, 32'shc0302af5, 32'shc02e42e2, 
               32'shc02c64a6, 32'shc02a9042, 32'shc028c5b6, 32'shc0270502, 32'shc0254e27, 32'shc023a124, 32'shc021fdfb, 32'shc02064ab, 
               32'shc01ed535, 32'shc01d4f99, 32'shc01bd3d6, 32'shc01a61ee, 32'shc018f9e1, 32'shc0179bae, 32'shc0164757, 32'shc014fcda, 
               32'shc013bc39, 32'shc0128574, 32'shc011588a, 32'shc010357c, 32'shc00f1c4a, 32'shc00e0cf5, 32'shc00d077c, 32'shc00c0be0, 
               32'shc00b1a20, 32'shc00a323d, 32'shc0095438, 32'shc008800f, 32'shc007b5c4, 32'shc006f556, 32'shc0063ec6, 32'shc0059214, 
               32'shc004ef3f, 32'shc0045648, 32'shc003c72f, 32'shc00341f4, 32'shc002c697, 32'shc0025519, 32'shc001ed78, 32'shc0018fb6, 
               32'shc0013bd3, 32'shc000f1ce, 32'shc000b1a7, 32'shc0007b5f, 32'shc0004ef5, 32'shc0002c6a, 32'shc00013bd, 32'shc00004ef, 
               32'shc0000000, 32'shc00004ef, 32'shc00013bd, 32'shc0002c6a, 32'shc0004ef5, 32'shc0007b5f, 32'shc000b1a7, 32'shc000f1ce, 
               32'shc0013bd3, 32'shc0018fb6, 32'shc001ed78, 32'shc0025519, 32'shc002c697, 32'shc00341f4, 32'shc003c72f, 32'shc0045648, 
               32'shc004ef3f, 32'shc0059214, 32'shc0063ec6, 32'shc006f556, 32'shc007b5c4, 32'shc008800f, 32'shc0095438, 32'shc00a323d, 
               32'shc00b1a20, 32'shc00c0be0, 32'shc00d077c, 32'shc00e0cf5, 32'shc00f1c4a, 32'shc010357c, 32'shc011588a, 32'shc0128574, 
               32'shc013bc39, 32'shc014fcda, 32'shc0164757, 32'shc0179bae, 32'shc018f9e1, 32'shc01a61ee, 32'shc01bd3d6, 32'shc01d4f99, 
               32'shc01ed535, 32'shc02064ab, 32'shc021fdfb, 32'shc023a124, 32'shc0254e27, 32'shc0270502, 32'shc028c5b6, 32'shc02a9042, 
               32'shc02c64a6, 32'shc02e42e2, 32'shc0302af5, 32'shc0321ce0, 32'shc03418a2, 32'shc0361e3a, 32'shc0382da8, 32'shc03a46ed, 
               32'shc03c6a07, 32'shc03e96f6, 32'shc040cdba, 32'shc0430e53, 32'shc04558c0, 32'shc047ad01, 32'shc04a0b16, 32'shc04c72fe, 
               32'shc04ee4b8, 32'shc0516045, 32'shc053e5a5, 32'shc05674d6, 32'shc0590dd8, 32'shc05bb0ab, 32'shc05e5d4e, 32'shc06113c2, 
               32'shc063d405, 32'shc0669e18, 32'shc06971f9, 32'shc06c4fa8, 32'shc06f3726, 32'shc0722871, 32'shc0752389, 32'shc078286e, 
               32'shc07b371e, 32'shc07e4f9b, 32'shc08171e2, 32'shc0849df4, 32'shc087d3d0, 32'shc08b1376, 32'shc08e5ce5, 32'shc091b01d, 
               32'shc0950d1d, 32'shc09873e4, 32'shc09be473, 32'shc09f5ec8, 32'shc0a2e2e3, 32'shc0a670c4, 32'shc0aa086a, 32'shc0ada9d4, 
               32'shc0b15502, 32'shc0b509f3, 32'shc0b8c8a7, 32'shc0bc911d, 32'shc0c06355, 32'shc0c43f4d, 32'shc0c82506, 32'shc0cc147f, 
               32'shc0d00db6, 32'shc0d410ad, 32'shc0d81d61, 32'shc0dc33d2, 32'shc0e05401, 32'shc0e47deb, 32'shc0e8b190, 32'shc0eceef1, 
               32'shc0f1360b, 32'shc0f586df, 32'shc0f9e16b, 32'shc0fe45b0, 32'shc102b3ac, 32'shc1072b5f, 32'shc10bacc8, 32'shc11037e6, 
               32'shc114ccb9, 32'shc1196b3f, 32'shc11e1379, 32'shc122c566, 32'shc1278104, 32'shc12c4653, 32'shc1311553, 32'shc135ee02, 
               32'shc13ad060, 32'shc13fbc6c, 32'shc144b225, 32'shc149b18b, 32'shc14eba9d, 32'shc153cd5a, 32'shc158e9c1, 32'shc15e0fd1, 
               32'shc1633f8a, 32'shc16878eb, 32'shc16dbbf3, 32'shc17308a1, 32'shc1785ef4, 32'shc17dbeec, 32'shc1832888, 32'shc1889bc6, 
               32'shc18e18a7, 32'shc1939f29, 32'shc1992f4c, 32'shc19ec90d, 32'shc1a46c6e, 32'shc1aa196c, 32'shc1afd007, 32'shc1b5903f, 
               32'shc1bb5a11, 32'shc1c12d7e, 32'shc1c70a84, 32'shc1ccf122, 32'shc1d2e158, 32'shc1d8db25, 32'shc1dede87, 32'shc1e4eb7e, 
               32'shc1eb0209, 32'shc1f12227, 32'shc1f74bd6, 32'shc1fd7f17, 32'shc203bbe8, 32'shc20a0248, 32'shc2105236, 32'shc216abb1, 
               32'shc21d0eb8, 32'shc2237b4b, 32'shc229f167, 32'shc230710d, 32'shc236fa3b, 32'shc23d8cf1, 32'shc244292c, 32'shc24aceed, 
               32'shc2517e31, 32'shc25836f9, 32'shc25ef943, 32'shc265c50e, 32'shc26c9a58, 32'shc2737922, 32'shc27a616a, 32'shc281532e, 
               32'shc2884e6e, 32'shc28f5329, 32'shc296615d, 32'shc29d790a, 32'shc2a49a2e, 32'shc2abc4c9, 32'shc2b2f8d8, 32'shc2ba365c, 
               32'shc2c17d52, 32'shc2c8cdbb, 32'shc2d02794, 32'shc2d78add, 32'shc2def794, 32'shc2e66db8, 32'shc2eded49, 32'shc2f57644, 
               32'shc2fd08a9, 32'shc304a477, 32'shc30c49ad, 32'shc313f848, 32'shc31bb049, 32'shc32371ae, 32'shc32b3c75, 32'shc333109e, 
               32'shc33aee27, 32'shc342d510, 32'shc34ac556, 32'shc352bef9, 32'shc35ac1f7, 32'shc362ce50, 32'shc36ae401, 32'shc373030a, 
               32'shc37b2b6a, 32'shc3835d1e, 32'shc38b9827, 32'shc393dc82, 32'shc39c2a2f, 32'shc3a4812c, 32'shc3ace178, 32'shc3b54b11, 
               32'shc3bdbdf6, 32'shc3c63a26, 32'shc3cebfa0, 32'shc3d74e62, 32'shc3dfe66c, 32'shc3e887bb, 32'shc3f1324e, 32'shc3f9e624, 
               32'shc402a33c, 32'shc40b6994, 32'shc414392b, 32'shc41d11ff, 32'shc425f410, 32'shc42edf5c, 32'shc437d3e1, 32'shc440d19e, 
               32'shc449d892, 32'shc452e8bc, 32'shc45c0219, 32'shc46524a9, 32'shc46e5069, 32'shc477855a, 32'shc480c379, 32'shc48a0ac4, 
               32'shc4935b3c, 32'shc49cb4dd, 32'shc4a617a6, 32'shc4af8397, 32'shc4b8f8ad, 32'shc4c276e8, 32'shc4cbfe45, 32'shc4d58ec3, 
               32'shc4df2862, 32'shc4e8cb1e, 32'shc4f276f7, 32'shc4fc2bec, 32'shc505e9fb, 32'shc50fb121, 32'shc519815f, 32'shc5235ab2, 
               32'shc52d3d18, 32'shc5372891, 32'shc5411d1b, 32'shc54b1ab4, 32'shc555215a, 32'shc55f310d, 32'shc56949ca, 32'shc5736b90, 
               32'shc57d965d, 32'shc587ca31, 32'shc5920708, 32'shc59c4ce3, 32'shc5a69bbe, 32'shc5b0f399, 32'shc5bb5472, 32'shc5c5be47, 
               32'shc5d03118, 32'shc5daace1, 32'shc5e531a1, 32'shc5efbf58, 32'shc5fa5603, 32'shc604f5a0, 32'shc60f9e2e, 32'shc61a4fac, 
               32'shc6250a18, 32'shc62fcd6f, 32'shc63a99b1, 32'shc6456edb, 32'shc6504ced, 32'shc65b33e4, 32'shc66623be, 32'shc6711c7b, 
               32'shc67c1e18, 32'shc6872894, 32'shc6923bec, 32'shc69d5820, 32'shc6a87d2d, 32'shc6b3ab12, 32'shc6bee1cd, 32'shc6ca215c, 
               32'shc6d569be, 32'shc6e0baf0, 32'shc6ec14f2, 32'shc6f777c1, 32'shc702e35c, 32'shc70e57c0, 32'shc719d4ed, 32'shc7255ae0, 
               32'shc730e997, 32'shc73c8111, 32'shc748214c, 32'shc753ca46, 32'shc75f7bfe, 32'shc76b3671, 32'shc776f99d, 32'shc782c582, 
               32'shc78e9a1d, 32'shc79a776c, 32'shc7a65d6e, 32'shc7b24c20, 32'shc7be4381, 32'shc7ca438f, 32'shc7d64c47, 32'shc7e25daa, 
               32'shc7ee77b3, 32'shc7fa9a62, 32'shc806c5b5, 32'shc812f9a9, 32'shc81f363d, 32'shc82b7b70, 32'shc837c93e, 32'shc8441fa6, 
               32'shc8507ea7, 32'shc85ce63e, 32'shc869566a, 32'shc875cf28, 32'shc8825077, 32'shc88eda54, 32'shc89b6cbf, 32'shc8a807b4, 
               32'shc8b4ab32, 32'shc8c15736, 32'shc8ce0bc0, 32'shc8dac8cd, 32'shc8e78e5b, 32'shc8f45c68, 32'shc90132f2, 32'shc90e11f7, 
               32'shc91af976, 32'shc927e96b, 32'shc934e1d6, 32'shc941e2b4, 32'shc94eec03, 32'shc95bfdc1, 32'shc96917ec, 32'shc9763a83, 
               32'shc9836582, 32'shc99098e9, 32'shc99dd4b4, 32'shc9ab18e3, 32'shc9b86572, 32'shc9c5ba60, 32'shc9d317ab, 32'shc9e07d51, 
               32'shc9edeb50, 32'shc9fb61a5, 32'shca08e04f, 32'shca16674b, 32'shca23f698, 32'shca318e32, 32'shca3f2e19, 32'shca4cd64b, 
               32'shca5a86c4, 32'shca683f83, 32'shca760086, 32'shca83c9ca, 32'shca919b4e, 32'shca9f750f, 32'shcaad570c, 32'shcabb4141, 
               32'shcac933ae, 32'shcad72e4f, 32'shcae53123, 32'shcaf33c28, 32'shcb014f5b, 32'shcb0f6aba, 32'shcb1d8e43, 32'shcb2bb9f4, 
               32'shcb39edca, 32'shcb4829c4, 32'shcb566ddf, 32'shcb64ba19, 32'shcb730e70, 32'shcb816ae1, 32'shcb8fcf6b, 32'shcb9e3c0b, 
               32'shcbacb0bf, 32'shcbbb2d85, 32'shcbc9b25a, 32'shcbd83f3d, 32'shcbe6d42b, 32'shcbf57121, 32'shcc04161e, 32'shcc12c31f, 
               32'shcc217822, 32'shcc303524, 32'shcc3efa25, 32'shcc4dc720, 32'shcc5c9c14, 32'shcc6b78ff, 32'shcc7a5dde, 32'shcc894aaf, 
               32'shcc983f70, 32'shcca73c1e, 32'shccb640b8, 32'shccc54d3a, 32'shccd461a2, 32'shcce37def, 32'shccf2a21d, 32'shcd01ce2b, 
               32'shcd110216, 32'shcd203ddc, 32'shcd2f817b, 32'shcd3eccef, 32'shcd4e2037, 32'shcd5d7b50, 32'shcd6cde39, 32'shcd7c48ee, 
               32'shcd8bbb6d, 32'shcd9b35b4, 32'shcdaab7c0, 32'shcdba4190, 32'shcdc9d320, 32'shcdd96c6f, 32'shcde90d79, 32'shcdf8b63d, 
               32'shce0866b8, 32'shce181ee8, 32'shce27dec9, 32'shce37a65b, 32'shce47759a, 32'shce574c84, 32'shce672b16, 32'shce77114e, 
               32'shce86ff2a, 32'shce96f4a7, 32'shcea6f1c2, 32'shceb6f67a, 32'shcec702cb, 32'shced716b4, 32'shcee73231, 32'shcef75541, 
               32'shcf077fe1, 32'shcf17b20d, 32'shcf27ebc5, 32'shcf382d05, 32'shcf4875ca, 32'shcf58c613, 32'shcf691ddd, 32'shcf797d24, 
               32'shcf89e3e8, 32'shcf9a5225, 32'shcfaac7d8, 32'shcfbb4500, 32'shcfcbc999, 32'shcfdc55a1, 32'shcfece915, 32'shcffd83f4, 
               32'shd00e2639, 32'shd01ecfe4, 32'shd02f80f1, 32'shd040395d, 32'shd050f926, 32'shd061c04a, 32'shd0728ec6, 32'shd0836497, 
               32'shd09441bb, 32'shd0a5262f, 32'shd0b611f1, 32'shd0c704fd, 32'shd0d7ff51, 32'shd0e900ec, 32'shd0fa09c9, 32'shd10b19e7, 
               32'shd11c3142, 32'shd12d4fd9, 32'shd13e75a8, 32'shd14fa2ad, 32'shd160d6e5, 32'shd172124d, 32'shd18354e4, 32'shd1949ea6, 
               32'shd1a5ef90, 32'shd1b747a0, 32'shd1c8a6d4, 32'shd1da0d28, 32'shd1eb7a9a, 32'shd1fcef27, 32'shd20e6acc, 32'shd21fed88, 
               32'shd2317756, 32'shd2430835, 32'shd254a021, 32'shd2663f19, 32'shd277e518, 32'shd289921e, 32'shd29b4626, 32'shd2ad012e, 
               32'shd2bec333, 32'shd2d08c33, 32'shd2e25c2b, 32'shd2f43318, 32'shd30610f7, 32'shd317f5c6, 32'shd329e181, 32'shd33bd427, 
               32'shd34dcdb4, 32'shd35fce26, 32'shd371d579, 32'shd383e3ab, 32'shd395f8ba, 32'shd3a814a2, 32'shd3ba3760, 32'shd3cc60f2, 
               32'shd3de9156, 32'shd3f0c887, 32'shd4030684, 32'shd4154b4a, 32'shd42796d5, 32'shd439e923, 32'shd44c4232, 32'shd45ea1fd, 
               32'shd4710883, 32'shd48375c1, 32'shd495e9b3, 32'shd4a86458, 32'shd4bae5ab, 32'shd4cd6dab, 32'shd4dffc54, 32'shd4f291a4, 
               32'shd5052d97, 32'shd517d02b, 32'shd52a795d, 32'shd53d292a, 32'shd54fdf8f, 32'shd5629c89, 32'shd5756016, 32'shd5882a32, 
               32'shd59afadb, 32'shd5add20d, 32'shd5c0afc6, 32'shd5d39403, 32'shd5e67ec1, 32'shd5f96ffd, 32'shd60c67b4, 32'shd61f65e4, 
               32'shd6326a88, 32'shd645759f, 32'shd6588725, 32'shd66b9f18, 32'shd67ebd74, 32'shd691e237, 32'shd6a50d5d, 32'shd6b83ee4, 
               32'shd6cb76c9, 32'shd6deb508, 32'shd6f1f99f, 32'shd705448b, 32'shd71895c9, 32'shd72bed55, 32'shd73f4b2e, 32'shd752af4f, 
               32'shd76619b6, 32'shd7798a60, 32'shd78d014a, 32'shd7a07e70, 32'shd7b401d1, 32'shd7c78b68, 32'shd7db1b34, 32'shd7eeb130, 
               32'shd8024d59, 32'shd815efae, 32'shd829982b, 32'shd83d46cc, 32'shd850fb8e, 32'shd864b670, 32'shd878776d, 32'shd88c3e83, 
               32'shd8a00bae, 32'shd8b3deeb, 32'shd8c7b838, 32'shd8db9792, 32'shd8ef7cf4, 32'shd903685d, 32'shd91759c9, 32'shd92b5135, 
               32'shd93f4e9e, 32'shd9535201, 32'shd9675b5a, 32'shd97b6aa8, 32'shd98f7fe6, 32'shd9a39b11, 32'shd9b7bc27, 32'shd9cbe325, 
               32'shd9e01006, 32'shd9f442c9, 32'shda087b69, 32'shda1cb9e5, 32'shda30fe38, 32'shda454860, 32'shda599859, 32'shda6dee21, 
               32'shda8249b4, 32'shda96ab0f, 32'shdaab122f, 32'shdabf7f11, 32'shdad3f1b1, 32'shdae86a0d, 32'shdafce821, 32'shdb116beb, 
               32'shdb25f566, 32'shdb3a8491, 32'shdb4f1967, 32'shdb63b3e5, 32'shdb785409, 32'shdb8cf9cf, 32'shdba1a534, 32'shdbb65634, 
               32'shdbcb0cce, 32'shdbdfc8fc, 32'shdbf48abd, 32'shdc09520d, 32'shdc1e1ee9, 32'shdc32f14d, 32'shdc47c936, 32'shdc5ca6a2, 
               32'shdc71898d, 32'shdc8671f3, 32'shdc9b5fd2, 32'shdcb05326, 32'shdcc54bec, 32'shdcda4a21, 32'shdcef4dc2, 32'shdd0456ca, 
               32'shdd196538, 32'shdd2e7908, 32'shdd439236, 32'shdd58b0c0, 32'shdd6dd4a2, 32'shdd82fdd8, 32'shdd982c60, 32'shddad6036, 
               32'shddc29958, 32'shddd7d7c1, 32'shdded1b6e, 32'shde02645d, 32'shde17b28a, 32'shde2d05f1, 32'shde425e8f, 32'shde57bc62, 
               32'shde6d1f65, 32'shde828796, 32'shde97f4f1, 32'shdead6773, 32'shdec2df18, 32'shded85bdd, 32'shdeedddc0, 32'shdf0364bc, 
               32'shdf18f0ce, 32'shdf2e81f3, 32'shdf441828, 32'shdf59b369, 32'shdf6f53b3, 32'shdf84f902, 32'shdf9aa354, 32'shdfb052a5, 
               32'shdfc606f1, 32'shdfdbc036, 32'shdff17e70, 32'she007419b, 32'she01d09b4, 32'she032d6b8, 32'she048a8a4, 32'she05e7f74, 
               32'she0745b24, 32'she08a3bb2, 32'she0a0211a, 32'she0b60b58, 32'she0cbfa6a, 32'she0e1ee4b, 32'she0f7e6f9, 32'she10de470, 
               32'she123e6ad, 32'she139edac, 32'she14ff96a, 32'she16609e3, 32'she17c1f15, 32'she19238fb, 32'she1a85793, 32'she1be7ad8, 
               32'she1d4a2c8, 32'she1eacf5f, 32'she2010099, 32'she2173674, 32'she22d70eb, 32'she243affc, 32'she259f3a3, 32'she2703bdc, 
               32'she28688a4, 32'she29cd9f8, 32'she2b32fd4, 32'she2c98a35, 32'she2dfe917, 32'she2f64c77, 32'she30cb451, 32'she32320a2, 
               32'she3399167, 32'she350069b, 32'she366803c, 32'she37cfe47, 32'she39380b6, 32'she3aa0788, 32'she3c092b9, 32'she3d72245, 
               32'she3edb628, 32'she4044e60, 32'she41aeae8, 32'she4318bbe, 32'she44830dd, 32'she45eda43, 32'she47587eb, 32'she48c39d3, 
               32'she4a2eff6, 32'she4b9aa52, 32'she4d068e2, 32'she4e72ba4, 32'she4fdf294, 32'she514bdad, 32'she52b8cee, 32'she5426051, 
               32'she55937d5, 32'she5701374, 32'she586f32c, 32'she59dd6f9, 32'she5b4bed8, 32'she5cbaac5, 32'she5e29abc, 32'she5f98ebb, 
               32'she61086bc, 32'she62782be, 32'she63e82bc, 32'she65586b3, 32'she66c8e9f, 32'she6839a7c, 32'she69aaa48, 32'she6b1bdff, 
               32'she6c8d59c, 32'she6dff11d, 32'she6f7107e, 32'she70e33bb, 32'she7255ad1, 32'she73c85bc, 32'she753b479, 32'she76ae704, 
               32'she7821d59, 32'she7995776, 32'she7b09555, 32'she7c7d6f4, 32'she7df1c50, 32'she7f66564, 32'she80db22d, 32'she82502a7, 
               32'she83c56cf, 32'she853aea1, 32'she86b0a1a, 32'she8826936, 32'she899cbf1, 32'she8b13248, 32'she8c89c37, 32'she8e009ba, 
               32'she8f77acf, 32'she90eef71, 32'she926679c, 32'she93de34e, 32'she9556282, 32'she96ce535, 32'she9846b63, 32'she99bf509, 
               32'she9b38223, 32'she9cb12ad, 32'she9e2a6a3, 32'she9fa3e03, 32'shea11d8c8, 32'shea2976ef, 32'shea411874, 32'shea58bd54, 
               32'shea70658a, 32'shea881114, 32'shea9fbfed, 32'sheab77212, 32'sheacf277f, 32'sheae6e031, 32'sheafe9c24, 32'sheb165b54, 
               32'sheb2e1dbe, 32'sheb45e35d, 32'sheb5dac2f, 32'sheb75782f, 32'sheb8d475b, 32'sheba519ad, 32'shebbcef23, 32'shebd4c7ba, 
               32'shebeca36c, 32'shec048237, 32'shec1c6417, 32'shec344908, 32'shec4c3106, 32'shec641c0e, 32'shec7c0a1d, 32'shec93fb2e, 
               32'shecabef3d, 32'shecc3e648, 32'shecdbe04a, 32'shecf3dd3f, 32'shed0bdd25, 32'shed23dff7, 32'shed3be5b1, 32'shed53ee51, 
               32'shed6bf9d1, 32'shed84082f, 32'shed9c1967, 32'shedb42d74, 32'shedcc4454, 32'shede45e03, 32'shedfc7a7c, 32'shee1499bd, 
               32'shee2cbbc1, 32'shee44e084, 32'shee5d0804, 32'shee75323c, 32'shee8d5f29, 32'sheea58ec6, 32'sheebdc110, 32'sheed5f604, 
               32'sheeee2d9d, 32'shef0667d9, 32'shef1ea4b2, 32'shef36e426, 32'shef4f2630, 32'shef676ace, 32'shef7fb1fa, 32'shef97fbb2, 
               32'shefb047f2, 32'shefc896b5, 32'shefe0e7f9, 32'sheff93bba, 32'shf01191f3, 32'shf029eaa1, 32'shf04245c0, 32'shf05aa34c, 
               32'shf0730342, 32'shf08b659f, 32'shf0a3ca5d, 32'shf0bc317a, 32'shf0d49af1, 32'shf0ed06bf, 32'shf10574e0, 32'shf11de551, 
               32'shf136580d, 32'shf14ecd11, 32'shf1674459, 32'shf17fbde2, 32'shf19839a6, 32'shf1b0b7a4, 32'shf1c937d6, 32'shf1e1ba3a, 
               32'shf1fa3ecb, 32'shf212c585, 32'shf22b4e66, 32'shf243d968, 32'shf25c6688, 32'shf274f5c3, 32'shf28d8715, 32'shf2a61a7a, 
               32'shf2beafed, 32'shf2d7476c, 32'shf2efe0f2, 32'shf3087c7d, 32'shf3211a07, 32'shf339b98d, 32'shf3525b0b, 32'shf36afe7e, 
               32'shf383a3e2, 32'shf39c4b32, 32'shf3b4f46c, 32'shf3cd9f8b, 32'shf3e64c8c, 32'shf3fefb6a, 32'shf417ac22, 32'shf4305eb0, 
               32'shf4491311, 32'shf461c940, 32'shf47a8139, 32'shf4933afa, 32'shf4abf67e, 32'shf4c4b3c0, 32'shf4dd72be, 32'shf4f63374, 
               32'shf50ef5de, 32'shf527b9f7, 32'shf5407fbd, 32'shf559472b, 32'shf572103d, 32'shf58adaf0, 32'shf5a3a740, 32'shf5bc7529, 
               32'shf5d544a7, 32'shf5ee15b7, 32'shf606e854, 32'shf61fbc7b, 32'shf6389228, 32'shf6516956, 32'shf66a4203, 32'shf6831c2b, 
               32'shf69bf7c9, 32'shf6b4d4d9, 32'shf6cdb359, 32'shf6e69344, 32'shf6ff7496, 32'shf718574b, 32'shf7313b60, 32'shf74a20d0, 
               32'shf7630799, 32'shf77befb5, 32'shf794d922, 32'shf7adc3db, 32'shf7c6afdc, 32'shf7df9d22, 32'shf7f88ba9, 32'shf8117b6d, 
               32'shf82a6c6a, 32'shf8435e9d, 32'shf85c5201, 32'shf8754692, 32'shf88e3c4d, 32'shf8a7332e, 32'shf8c02b31, 32'shf8d92452, 
               32'shf8f21e8e, 32'shf90b19e0, 32'shf9241645, 32'shf93d13b8, 32'shf9561237, 32'shf96f11bc, 32'shf9881245, 32'shf9a113cd, 
               32'shf9ba1651, 32'shf9d319cc, 32'shf9ec1e3b, 32'shfa05239a, 32'shfa1e29e5, 32'shfa373119, 32'shfa503930, 32'shfa694229, 
               32'shfa824bfd, 32'shfa9b56ab, 32'shfab4622d, 32'shfacd6e81, 32'shfae67ba2, 32'shfaff898c, 32'shfb18983b, 32'shfb31a7ac, 
               32'shfb4ab7db, 32'shfb63c8c4, 32'shfb7cda63, 32'shfb95ecb4, 32'shfbaeffb3, 32'shfbc8135c, 32'shfbe127ac, 32'shfbfa3c9f, 
               32'shfc135231, 32'shfc2c685d, 32'shfc457f21, 32'shfc5e9678, 32'shfc77ae5e, 32'shfc90c6cf, 32'shfca9dfc8, 32'shfcc2f945, 
               32'shfcdc1342, 32'shfcf52dbb, 32'shfd0e48ab, 32'shfd276410, 32'shfd407fe6, 32'shfd599c28, 32'shfd72b8d2, 32'shfd8bd5e1, 
               32'shfda4f351, 32'shfdbe111e, 32'shfdd72f45, 32'shfdf04dc0, 32'shfe096c8d, 32'shfe228ba7, 32'shfe3bab0b, 32'shfe54cab5, 
               32'shfe6deaa1, 32'shfe870aca, 32'shfea02b2e, 32'shfeb94bc8, 32'shfed26c94, 32'shfeeb8d8f, 32'shff04aeb5, 32'shff1dd001, 
               32'shff36f170, 32'shff5012fe, 32'shff6934a8, 32'shff825668, 32'shff9b783c, 32'shffb49a1f, 32'shffcdbc0f, 32'shffe6de05
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 13)
         begin
            reg signed [31:0] W_Re_table[4096] = '{
               32'sh40000000, 32'sh3ffffec4, 32'sh3ffffb11, 32'sh3ffff4e6, 32'sh3fffec43, 32'sh3fffe128, 32'sh3fffd396, 32'sh3fffc38c, 
               32'sh3fffb10b, 32'sh3fff9c12, 32'sh3fff84a1, 32'sh3fff6ab9, 32'sh3fff4e59, 32'sh3fff2f82, 32'sh3fff0e32, 32'sh3ffeea6c, 
               32'sh3ffec42d, 32'sh3ffe9b77, 32'sh3ffe704a, 32'sh3ffe42a4, 32'sh3ffe1288, 32'sh3ffddff3, 32'sh3ffdaae7, 32'sh3ffd7364, 
               32'sh3ffd3969, 32'sh3ffcfcf6, 32'sh3ffcbe0c, 32'sh3ffc7caa, 32'sh3ffc38d1, 32'sh3ffbf280, 32'sh3ffba9b8, 32'sh3ffb5e78, 
               32'sh3ffb10c1, 32'sh3ffac092, 32'sh3ffa6dec, 32'sh3ffa18cf, 32'sh3ff9c13a, 32'sh3ff9672d, 32'sh3ff90aaa, 32'sh3ff8abae, 
               32'sh3ff84a3c, 32'sh3ff7e652, 32'sh3ff77ff1, 32'sh3ff71718, 32'sh3ff6abc8, 32'sh3ff63e01, 32'sh3ff5cdc3, 32'sh3ff55b0d, 
               32'sh3ff4e5e0, 32'sh3ff46e3c, 32'sh3ff3f420, 32'sh3ff3778e, 32'sh3ff2f884, 32'sh3ff27703, 32'sh3ff1f30b, 32'sh3ff16c9c, 
               32'sh3ff0e3b6, 32'sh3ff05858, 32'sh3fefca84, 32'sh3fef3a39, 32'sh3feea776, 32'sh3fee123d, 32'sh3fed7a8c, 32'sh3fece065, 
               32'sh3fec43c7, 32'sh3feba4b2, 32'sh3feb0326, 32'sh3fea5f23, 32'sh3fe9b8a9, 32'sh3fe90fb9, 32'sh3fe86452, 32'sh3fe7b674, 
               32'sh3fe7061f, 32'sh3fe65354, 32'sh3fe59e12, 32'sh3fe4e659, 32'sh3fe42c2a, 32'sh3fe36f84, 32'sh3fe2b067, 32'sh3fe1eed5, 
               32'sh3fe12acb, 32'sh3fe0644b, 32'sh3fdf9b55, 32'sh3fdecfe8, 32'sh3fde0205, 32'sh3fdd31ac, 32'sh3fdc5edc, 32'sh3fdb8996, 
               32'sh3fdab1d9, 32'sh3fd9d7a7, 32'sh3fd8fafe, 32'sh3fd81bdf, 32'sh3fd73a4a, 32'sh3fd6563f, 32'sh3fd56fbe, 32'sh3fd486c7, 
               32'sh3fd39b5a, 32'sh3fd2ad77, 32'sh3fd1bd1e, 32'sh3fd0ca4f, 32'sh3fcfd50b, 32'sh3fcedd50, 32'sh3fcde320, 32'sh3fcce67a, 
               32'sh3fcbe75e, 32'sh3fcae5cd, 32'sh3fc9e1c6, 32'sh3fc8db4a, 32'sh3fc7d258, 32'sh3fc6c6f0, 32'sh3fc5b913, 32'sh3fc4a8c1, 
               32'sh3fc395f9, 32'sh3fc280bc, 32'sh3fc1690a, 32'sh3fc04ee3, 32'sh3fbf3246, 32'sh3fbe1334, 32'sh3fbcf1ad, 32'sh3fbbcdb1, 
               32'sh3fbaa740, 32'sh3fb97e5a, 32'sh3fb852ff, 32'sh3fb7252f, 32'sh3fb5f4ea, 32'sh3fb4c231, 32'sh3fb38d02, 32'sh3fb2555f, 
               32'sh3fb11b48, 32'sh3fafdebb, 32'sh3fae9fbb, 32'sh3fad5e45, 32'sh3fac1a5b, 32'sh3faad3fd, 32'sh3fa98b2a, 32'sh3fa83fe3, 
               32'sh3fa6f228, 32'sh3fa5a1f9, 32'sh3fa44f55, 32'sh3fa2fa3d, 32'sh3fa1a2b2, 32'sh3fa048b2, 32'sh3f9eec3e, 32'sh3f9d8d56, 
               32'sh3f9c2bfb, 32'sh3f9ac82c, 32'sh3f9961e8, 32'sh3f97f932, 32'sh3f968e07, 32'sh3f952069, 32'sh3f93b058, 32'sh3f923dd2, 
               32'sh3f90c8da, 32'sh3f8f516e, 32'sh3f8dd78f, 32'sh3f8c5b3d, 32'sh3f8adc77, 32'sh3f895b3e, 32'sh3f87d792, 32'sh3f865174, 
               32'sh3f84c8e2, 32'sh3f833ddd, 32'sh3f81b065, 32'sh3f80207b, 32'sh3f7e8e1e, 32'sh3f7cf94e, 32'sh3f7b620c, 32'sh3f79c857, 
               32'sh3f782c30, 32'sh3f768d96, 32'sh3f74ec8a, 32'sh3f73490b, 32'sh3f71a31b, 32'sh3f6ffab8, 32'sh3f6e4fe3, 32'sh3f6ca29c, 
               32'sh3f6af2e3, 32'sh3f6940b8, 32'sh3f678c1c, 32'sh3f65d50d, 32'sh3f641b8d, 32'sh3f625f9b, 32'sh3f60a138, 32'sh3f5ee063, 
               32'sh3f5d1d1d, 32'sh3f5b5765, 32'sh3f598f3c, 32'sh3f57c4a2, 32'sh3f55f796, 32'sh3f54281a, 32'sh3f52562c, 32'sh3f5081cd, 
               32'sh3f4eaafe, 32'sh3f4cd1be, 32'sh3f4af60d, 32'sh3f4917eb, 32'sh3f473759, 32'sh3f455456, 32'sh3f436ee3, 32'sh3f4186ff, 
               32'sh3f3f9cab, 32'sh3f3dafe7, 32'sh3f3bc0b3, 32'sh3f39cf0e, 32'sh3f37dafa, 32'sh3f35e476, 32'sh3f33eb81, 32'sh3f31f01d, 
               32'sh3f2ff24a, 32'sh3f2df206, 32'sh3f2bef53, 32'sh3f29ea31, 32'sh3f27e29f, 32'sh3f25d89e, 32'sh3f23cc2e, 32'sh3f21bd4e, 
               32'sh3f1fabff, 32'sh3f1d9842, 32'sh3f1b8215, 32'sh3f19697a, 32'sh3f174e70, 32'sh3f1530f7, 32'sh3f13110f, 32'sh3f10eeb9, 
               32'sh3f0ec9f5, 32'sh3f0ca2c2, 32'sh3f0a7921, 32'sh3f084d12, 32'sh3f061e95, 32'sh3f03eda9, 32'sh3f01ba50, 32'sh3eff8489, 
               32'sh3efd4c54, 32'sh3efb11b1, 32'sh3ef8d4a1, 32'sh3ef69523, 32'sh3ef45338, 32'sh3ef20ee0, 32'sh3eefc81a, 32'sh3eed7ee7, 
               32'sh3eeb3347, 32'sh3ee8e53a, 32'sh3ee694c1, 32'sh3ee441da, 32'sh3ee1ec87, 32'sh3edf94c7, 32'sh3edd3a9a, 32'sh3edade01, 
               32'sh3ed87efc, 32'sh3ed61d8a, 32'sh3ed3b9ad, 32'sh3ed15363, 32'sh3eceeaad, 32'sh3ecc7f8b, 32'sh3eca11fe, 32'sh3ec7a205, 
               32'sh3ec52fa0, 32'sh3ec2bad0, 32'sh3ec04394, 32'sh3ebdc9ed, 32'sh3ebb4ddb, 32'sh3eb8cf5d, 32'sh3eb64e75, 32'sh3eb3cb21, 
               32'sh3eb14563, 32'sh3eaebd3a, 32'sh3eac32a6, 32'sh3ea9a5a8, 32'sh3ea7163f, 32'sh3ea4846c, 32'sh3ea1f02f, 32'sh3e9f5988, 
               32'sh3e9cc076, 32'sh3e9a24fb, 32'sh3e978715, 32'sh3e94e6c6, 32'sh3e92440d, 32'sh3e8f9eeb, 32'sh3e8cf75f, 32'sh3e8a4d6a, 
               32'sh3e87a10c, 32'sh3e84f245, 32'sh3e824114, 32'sh3e7f8d7b, 32'sh3e7cd778, 32'sh3e7a1f0d, 32'sh3e77643a, 32'sh3e74a6fd, 
               32'sh3e71e759, 32'sh3e6f254c, 32'sh3e6c60d7, 32'sh3e6999fa, 32'sh3e66d0b4, 32'sh3e640507, 32'sh3e6136f3, 32'sh3e5e6676, 
               32'sh3e5b9392, 32'sh3e58be47, 32'sh3e55e694, 32'sh3e530c7a, 32'sh3e502ff9, 32'sh3e4d5110, 32'sh3e4a6fc1, 32'sh3e478c0b, 
               32'sh3e44a5ef, 32'sh3e41bd6c, 32'sh3e3ed282, 32'sh3e3be532, 32'sh3e38f57c, 32'sh3e360360, 32'sh3e330ede, 32'sh3e3017f6, 
               32'sh3e2d1ea8, 32'sh3e2a22f4, 32'sh3e2724db, 32'sh3e24245d, 32'sh3e212179, 32'sh3e1e1c30, 32'sh3e1b1482, 32'sh3e180a6f, 
               32'sh3e14fdf7, 32'sh3e11ef1b, 32'sh3e0eddd9, 32'sh3e0bca34, 32'sh3e08b42a, 32'sh3e059bbb, 32'sh3e0280e9, 32'sh3dff63b2, 
               32'sh3dfc4418, 32'sh3df9221a, 32'sh3df5fdb8, 32'sh3df2d6f3, 32'sh3defadca, 32'sh3dec823e, 32'sh3de9544f, 32'sh3de623fd, 
               32'sh3de2f148, 32'sh3ddfbc30, 32'sh3ddc84b5, 32'sh3dd94ad8, 32'sh3dd60e99, 32'sh3dd2cff7, 32'sh3dcf8ef3, 32'sh3dcc4b8d, 
               32'sh3dc905c5, 32'sh3dc5bd9b, 32'sh3dc2730f, 32'sh3dbf2622, 32'sh3dbbd6d4, 32'sh3db88524, 32'sh3db53113, 32'sh3db1daa2, 
               32'sh3dae81cf, 32'sh3dab269b, 32'sh3da7c907, 32'sh3da46912, 32'sh3da106bd, 32'sh3d9da208, 32'sh3d9a3af2, 32'sh3d96d17d, 
               32'sh3d9365a8, 32'sh3d8ff772, 32'sh3d8c86de, 32'sh3d8913ea, 32'sh3d859e96, 32'sh3d8226e4, 32'sh3d7eacd2, 32'sh3d7b3061, 
               32'sh3d77b192, 32'sh3d743064, 32'sh3d70acd7, 32'sh3d6d26ec, 32'sh3d699ea3, 32'sh3d6613fb, 32'sh3d6286f6, 32'sh3d5ef793, 
               32'sh3d5b65d2, 32'sh3d57d1b3, 32'sh3d543b37, 32'sh3d50a25e, 32'sh3d4d0728, 32'sh3d496994, 32'sh3d45c9a4, 32'sh3d422757, 
               32'sh3d3e82ae, 32'sh3d3adba7, 32'sh3d373245, 32'sh3d338687, 32'sh3d2fd86c, 32'sh3d2c27f6, 32'sh3d287523, 32'sh3d24bff6, 
               32'sh3d21086c, 32'sh3d1d4e88, 32'sh3d199248, 32'sh3d15d3ad, 32'sh3d1212b7, 32'sh3d0e4f67, 32'sh3d0a89bc, 32'sh3d06c1b6, 
               32'sh3d02f757, 32'sh3cff2a9d, 32'sh3cfb5b89, 32'sh3cf78a1b, 32'sh3cf3b653, 32'sh3cefe032, 32'sh3cec07b8, 32'sh3ce82ce4, 
               32'sh3ce44fb7, 32'sh3ce07031, 32'sh3cdc8e52, 32'sh3cd8aa1b, 32'sh3cd4c38b, 32'sh3cd0daa2, 32'sh3cccef62, 32'sh3cc901c9, 
               32'sh3cc511d9, 32'sh3cc11f90, 32'sh3cbd2af0, 32'sh3cb933f9, 32'sh3cb53aaa, 32'sh3cb13f04, 32'sh3cad4107, 32'sh3ca940b3, 
               32'sh3ca53e09, 32'sh3ca13908, 32'sh3c9d31b0, 32'sh3c992803, 32'sh3c951bff, 32'sh3c910da5, 32'sh3c8cfcf6, 32'sh3c88e9f1, 
               32'sh3c84d496, 32'sh3c80bce7, 32'sh3c7ca2e2, 32'sh3c788688, 32'sh3c7467d9, 32'sh3c7046d6, 32'sh3c6c237e, 32'sh3c67fdd1, 
               32'sh3c63d5d1, 32'sh3c5fab7c, 32'sh3c5b7ed4, 32'sh3c574fd8, 32'sh3c531e88, 32'sh3c4eeae5, 32'sh3c4ab4ef, 32'sh3c467ca6, 
               32'sh3c42420a, 32'sh3c3e051b, 32'sh3c39c5da, 32'sh3c358446, 32'sh3c314060, 32'sh3c2cfa28, 32'sh3c28b19e, 32'sh3c2466c2, 
               32'sh3c201994, 32'sh3c1bca16, 32'sh3c177845, 32'sh3c132424, 32'sh3c0ecdb2, 32'sh3c0a74f0, 32'sh3c0619dc, 32'sh3c01bc78, 
               32'sh3bfd5cc4, 32'sh3bf8fac0, 32'sh3bf4966c, 32'sh3bf02fc9, 32'sh3bebc6d5, 32'sh3be75b93, 32'sh3be2ee01, 32'sh3bde7e20, 
               32'sh3bda0bf0, 32'sh3bd59771, 32'sh3bd120a4, 32'sh3bcca789, 32'sh3bc82c1f, 32'sh3bc3ae67, 32'sh3bbf2e62, 32'sh3bbaac0e, 
               32'sh3bb6276e, 32'sh3bb1a080, 32'sh3bad1744, 32'sh3ba88bbc, 32'sh3ba3fde7, 32'sh3b9f6dc5, 32'sh3b9adb57, 32'sh3b96469d, 
               32'sh3b91af97, 32'sh3b8d1644, 32'sh3b887aa6, 32'sh3b83dcbc, 32'sh3b7f3c87, 32'sh3b7a9a07, 32'sh3b75f53c, 32'sh3b714e25, 
               32'sh3b6ca4c4, 32'sh3b67f919, 32'sh3b634b23, 32'sh3b5e9ae4, 32'sh3b59e85a, 32'sh3b553386, 32'sh3b507c69, 32'sh3b4bc303, 
               32'sh3b470753, 32'sh3b42495a, 32'sh3b3d8918, 32'sh3b38c68e, 32'sh3b3401bb, 32'sh3b2f3aa0, 32'sh3b2a713d, 32'sh3b25a591, 
               32'sh3b20d79e, 32'sh3b1c0764, 32'sh3b1734e2, 32'sh3b126019, 32'sh3b0d8909, 32'sh3b08afb2, 32'sh3b03d414, 32'sh3afef630, 
               32'sh3afa1605, 32'sh3af53395, 32'sh3af04edf, 32'sh3aeb67e3, 32'sh3ae67ea1, 32'sh3ae1931a, 32'sh3adca54e, 32'sh3ad7b53d, 
               32'sh3ad2c2e8, 32'sh3acdce4d, 32'sh3ac8d76f, 32'sh3ac3de4c, 32'sh3abee2e5, 32'sh3ab9e53a, 32'sh3ab4e54c, 32'sh3aafe31b, 
               32'sh3aaadea6, 32'sh3aa5d7ee, 32'sh3aa0cef3, 32'sh3a9bc3b6, 32'sh3a96b636, 32'sh3a91a674, 32'sh3a8c9470, 32'sh3a87802a, 
               32'sh3a8269a3, 32'sh3a7d50da, 32'sh3a7835cf, 32'sh3a731884, 32'sh3a6df8f8, 32'sh3a68d72b, 32'sh3a63b31d, 32'sh3a5e8cd0, 
               32'sh3a596442, 32'sh3a543974, 32'sh3a4f0c67, 32'sh3a49dd1a, 32'sh3a44ab8e, 32'sh3a3f77c3, 32'sh3a3a41b9, 32'sh3a350970, 
               32'sh3a2fcee8, 32'sh3a2a9223, 32'sh3a25531f, 32'sh3a2011de, 32'sh3a1ace5f, 32'sh3a1588a2, 32'sh3a1040a8, 32'sh3a0af671, 
               32'sh3a05a9fd, 32'sh3a005b4d, 32'sh39fb0a60, 32'sh39f5b737, 32'sh39f061d2, 32'sh39eb0a31, 32'sh39e5b054, 32'sh39e0543c, 
               32'sh39daf5e8, 32'sh39d5955a, 32'sh39d03291, 32'sh39cacd8d, 32'sh39c5664f, 32'sh39bffcd7, 32'sh39ba9125, 32'sh39b52339, 
               32'sh39afb313, 32'sh39aa40b4, 32'sh39a4cc1c, 32'sh399f554b, 32'sh3999dc42, 32'sh399460ff, 32'sh398ee385, 32'sh398963d2, 
               32'sh3983e1e8, 32'sh397e5dc6, 32'sh3978d76c, 32'sh39734edc, 32'sh396dc414, 32'sh39683715, 32'sh3962a7e0, 32'sh395d1675, 
               32'sh395782d3, 32'sh3951ecfc, 32'sh394c54ee, 32'sh3946baac, 32'sh39411e33, 32'sh393b7f86, 32'sh3935dea4, 32'sh39303b8e, 
               32'sh392a9642, 32'sh3924eec3, 32'sh391f4510, 32'sh39199929, 32'sh3913eb0e, 32'sh390e3ac0, 32'sh3908883f, 32'sh3902d38b, 
               32'sh38fd1ca4, 32'sh38f7638b, 32'sh38f1a840, 32'sh38ebeac2, 32'sh38e62b13, 32'sh38e06932, 32'sh38daa520, 32'sh38d4dedd, 
               32'sh38cf1669, 32'sh38c94bc4, 32'sh38c37eef, 32'sh38bdafea, 32'sh38b7deb4, 32'sh38b20b4f, 32'sh38ac35ba, 32'sh38a65df6, 
               32'sh38a08402, 32'sh389aa7e0, 32'sh3894c98f, 32'sh388ee910, 32'sh38890663, 32'sh38832187, 32'sh387d3a7e, 32'sh38775147, 
               32'sh387165e3, 32'sh386b7852, 32'sh38658894, 32'sh385f96a9, 32'sh3859a292, 32'sh3853ac4f, 32'sh384db3e0, 32'sh3847b946, 
               32'sh3841bc7f, 32'sh383bbd8e, 32'sh3835bc71, 32'sh382fb92a, 32'sh3829b3b9, 32'sh3823ac1d, 32'sh381da256, 32'sh38179666, 
               32'sh3811884d, 32'sh380b780a, 32'sh3805659e, 32'sh37ff5109, 32'sh37f93a4b, 32'sh37f32165, 32'sh37ed0657, 32'sh37e6e921, 
               32'sh37e0c9c3, 32'sh37daa83d, 32'sh37d48490, 32'sh37ce5ebd, 32'sh37c836c2, 32'sh37c20ca1, 32'sh37bbe05a, 32'sh37b5b1ec, 
               32'sh37af8159, 32'sh37a94ea0, 32'sh37a319c2, 32'sh379ce2be, 32'sh3796a996, 32'sh37906e49, 32'sh378a30d8, 32'sh3783f143, 
               32'sh377daf89, 32'sh37776bac, 32'sh377125ac, 32'sh376add88, 32'sh37649341, 32'sh375e46d8, 32'sh3757f84c, 32'sh3751a79e, 
               32'sh374b54ce, 32'sh3744ffdd, 32'sh373ea8ca, 32'sh37384f95, 32'sh3731f440, 32'sh372b96ca, 32'sh37253733, 32'sh371ed57c, 
               32'sh371871a5, 32'sh37120bae, 32'sh370ba398, 32'sh37053962, 32'sh36fecd0e, 32'sh36f85e9a, 32'sh36f1ee09, 32'sh36eb7b58, 
               32'sh36e5068a, 32'sh36de8f9e, 32'sh36d81695, 32'sh36d19b6e, 32'sh36cb1e2a, 32'sh36c49ec9, 32'sh36be1d4c, 32'sh36b799b3, 
               32'sh36b113fd, 32'sh36aa8c2c, 32'sh36a4023f, 32'sh369d7637, 32'sh3696e814, 32'sh369057d6, 32'sh3689c57d, 32'sh3683310b, 
               32'sh367c9a7e, 32'sh367601d7, 32'sh366f6717, 32'sh3668ca3e, 32'sh36622b4c, 32'sh365b8a41, 32'sh3654e71d, 32'sh364e41e2, 
               32'sh36479a8e, 32'sh3640f123, 32'sh363a45a0, 32'sh36339806, 32'sh362ce855, 32'sh3626368d, 32'sh361f82af, 32'sh3618ccba, 
               32'sh361214b0, 32'sh360b5a90, 32'sh36049e5b, 32'sh35fde011, 32'sh35f71fb1, 32'sh35f05d3d, 32'sh35e998b5, 32'sh35e2d219, 
               32'sh35dc0968, 32'sh35d53ea5, 32'sh35ce71ce, 32'sh35c7a2e3, 32'sh35c0d1e7, 32'sh35b9fed7, 32'sh35b329b5, 32'sh35ac5282, 
               32'sh35a5793c, 32'sh359e9de5, 32'sh3597c07d, 32'sh3590e104, 32'sh3589ff7a, 32'sh35831be0, 32'sh357c3636, 32'sh35754e7c, 
               32'sh356e64b2, 32'sh356778d9, 32'sh35608af1, 32'sh35599afa, 32'sh3552a8f4, 32'sh354bb4e1, 32'sh3544bebf, 32'sh353dc68f, 
               32'sh3536cc52, 32'sh352fd008, 32'sh3528d1b1, 32'sh3521d14d, 32'sh351acedd, 32'sh3513ca60, 32'sh350cc3d8, 32'sh3505bb44, 
               32'sh34feb0a5, 32'sh34f7a3fb, 32'sh34f09546, 32'sh34e98487, 32'sh34e271bd, 32'sh34db5cea, 32'sh34d4460c, 32'sh34cd2d26, 
               32'sh34c61236, 32'sh34bef53d, 32'sh34b7d63c, 32'sh34b0b533, 32'sh34a99221, 32'sh34a26d08, 32'sh349b45e7, 32'sh34941cbf, 
               32'sh348cf190, 32'sh3485c45b, 32'sh347e951f, 32'sh347763dd, 32'sh34703095, 32'sh3468fb47, 32'sh3461c3f5, 32'sh345a8a9d, 
               32'sh34534f41, 32'sh344c11e0, 32'sh3444d27b, 32'sh343d9112, 32'sh34364da6, 32'sh342f0836, 32'sh3427c0c3, 32'sh3420774d, 
               32'sh34192bd5, 32'sh3411de5b, 32'sh340a8edf, 32'sh34033d61, 32'sh33fbe9e2, 32'sh33f49462, 32'sh33ed3ce1, 32'sh33e5e360, 
               32'sh33de87de, 32'sh33d72a5d, 32'sh33cfcadc, 32'sh33c8695b, 32'sh33c105db, 32'sh33b9a05d, 32'sh33b238e0, 32'sh33aacf65, 
               32'sh33a363ec, 32'sh339bf675, 32'sh33948701, 32'sh338d1590, 32'sh3385a222, 32'sh337e2cb7, 32'sh3376b551, 32'sh336f3bee, 
               32'sh3367c090, 32'sh33604336, 32'sh3358c3e2, 32'sh33514292, 32'sh3349bf48, 32'sh33423a04, 32'sh333ab2c6, 32'sh3333298f, 
               32'sh332b9e5e, 32'sh33241134, 32'sh331c8211, 32'sh3314f0f6, 32'sh330d5de3, 32'sh3305c8d7, 32'sh32fe31d5, 32'sh32f698db, 
               32'sh32eefdea, 32'sh32e76102, 32'sh32dfc224, 32'sh32d82150, 32'sh32d07e85, 32'sh32c8d9c6, 32'sh32c13311, 32'sh32b98a67, 
               32'sh32b1dfc9, 32'sh32aa3336, 32'sh32a284b0, 32'sh329ad435, 32'sh329321c7, 32'sh328b6d66, 32'sh3283b712, 32'sh327bfecc, 
               32'sh32744493, 32'sh326c8868, 32'sh3264ca4c, 32'sh325d0a3e, 32'sh32554840, 32'sh324d8450, 32'sh3245be70, 32'sh323df6a0, 
               32'sh32362ce0, 32'sh322e6130, 32'sh32269391, 32'sh321ec403, 32'sh3216f287, 32'sh320f1f1c, 32'sh320749c3, 32'sh31ff727c, 
               32'sh31f79948, 32'sh31efbe27, 32'sh31e7e118, 32'sh31e0021e, 32'sh31d82137, 32'sh31d03e64, 32'sh31c859a5, 32'sh31c072fb, 
               32'sh31b88a66, 32'sh31b09fe7, 32'sh31a8b37c, 32'sh31a0c528, 32'sh3198d4ea, 32'sh3190e2c3, 32'sh3188eeb2, 32'sh3180f8b8, 
               32'sh317900d6, 32'sh3171070c, 32'sh31690b59, 32'sh31610dbf, 32'sh31590e3e, 32'sh31510cd5, 32'sh31490986, 32'sh31410450, 
               32'sh3138fd35, 32'sh3130f433, 32'sh3128e94c, 32'sh3120dc80, 32'sh3118cdcf, 32'sh3110bd39, 32'sh3108aabf, 32'sh31009661, 
               32'sh30f8801f, 32'sh30f067fb, 32'sh30e84df3, 32'sh30e03208, 32'sh30d8143b, 32'sh30cff48c, 32'sh30c7d2fb, 32'sh30bfaf89, 
               32'sh30b78a36, 32'sh30af6302, 32'sh30a739ed, 32'sh309f0ef8, 32'sh3096e223, 32'sh308eb36f, 32'sh308682dc, 32'sh307e5069, 
               32'sh30761c18, 32'sh306de5e9, 32'sh3065addb, 32'sh305d73f0, 32'sh30553828, 32'sh304cfa83, 32'sh3044bb00, 32'sh303c79a2, 
               32'sh30343667, 32'sh302bf151, 32'sh3023aa5f, 32'sh301b6193, 32'sh301316eb, 32'sh300aca69, 32'sh30027c0c, 32'sh2ffa2bd6, 
               32'sh2ff1d9c7, 32'sh2fe985de, 32'sh2fe1301c, 32'sh2fd8d882, 32'sh2fd07f0f, 32'sh2fc823c5, 32'sh2fbfc6a3, 32'sh2fb767aa, 
               32'sh2faf06da, 32'sh2fa6a433, 32'sh2f9e3fb6, 32'sh2f95d963, 32'sh2f8d713a, 32'sh2f85073c, 32'sh2f7c9b69, 32'sh2f742dc1, 
               32'sh2f6bbe45, 32'sh2f634cf5, 32'sh2f5ad9d1, 32'sh2f5264da, 32'sh2f49ee0f, 32'sh2f417573, 32'sh2f38fb03, 32'sh2f307ec2, 
               32'sh2f2800af, 32'sh2f1f80ca, 32'sh2f16ff14, 32'sh2f0e7b8e, 32'sh2f05f637, 32'sh2efd6f10, 32'sh2ef4e619, 32'sh2eec5b53, 
               32'sh2ee3cebe, 32'sh2edb405a, 32'sh2ed2b027, 32'sh2eca1e27, 32'sh2ec18a58, 32'sh2eb8f4bc, 32'sh2eb05d53, 32'sh2ea7c41e, 
               32'sh2e9f291b, 32'sh2e968c4d, 32'sh2e8dedb3, 32'sh2e854d4d, 32'sh2e7cab1c, 32'sh2e740720, 32'sh2e6b615a, 32'sh2e62b9ca, 
               32'sh2e5a1070, 32'sh2e51654c, 32'sh2e48b860, 32'sh2e4009aa, 32'sh2e37592c, 32'sh2e2ea6e6, 32'sh2e25f2d8, 32'sh2e1d3d03, 
               32'sh2e148566, 32'sh2e0bcc03, 32'sh2e0310d9, 32'sh2dfa53e9, 32'sh2df19534, 32'sh2de8d4b8, 32'sh2de01278, 32'sh2dd74e73, 
               32'sh2dce88aa, 32'sh2dc5c11c, 32'sh2dbcf7cb, 32'sh2db42cb6, 32'sh2dab5fdf, 32'sh2da29144, 32'sh2d99c0e7, 32'sh2d90eec8, 
               32'sh2d881ae8, 32'sh2d7f4545, 32'sh2d766de2, 32'sh2d6d94bf, 32'sh2d64b9da, 32'sh2d5bdd36, 32'sh2d52fed2, 32'sh2d4a1eaf, 
               32'sh2d413ccd, 32'sh2d38592c, 32'sh2d2f73cd, 32'sh2d268cb0, 32'sh2d1da3d5, 32'sh2d14b93d, 32'sh2d0bcce8, 32'sh2d02ded7, 
               32'sh2cf9ef09, 32'sh2cf0fd80, 32'sh2ce80a3a, 32'sh2cdf153a, 32'sh2cd61e7f, 32'sh2ccd2609, 32'sh2cc42bd9, 32'sh2cbb2fef, 
               32'sh2cb2324c, 32'sh2ca932ef, 32'sh2ca031da, 32'sh2c972f0d, 32'sh2c8e2a87, 32'sh2c85244a, 32'sh2c7c1c55, 32'sh2c7312a9, 
               32'sh2c6a0746, 32'sh2c60fa2d, 32'sh2c57eb5e, 32'sh2c4edada, 32'sh2c45c8a0, 32'sh2c3cb4b1, 32'sh2c339f0e, 32'sh2c2a87b6, 
               32'sh2c216eaa, 32'sh2c1853eb, 32'sh2c0f3779, 32'sh2c061953, 32'sh2bfcf97c, 32'sh2bf3d7f2, 32'sh2beab4b6, 32'sh2be18fc9, 
               32'sh2bd8692b, 32'sh2bcf40dc, 32'sh2bc616dd, 32'sh2bbceb2d, 32'sh2bb3bdce, 32'sh2baa8ec0, 32'sh2ba15e03, 32'sh2b982b97, 
               32'sh2b8ef77d, 32'sh2b85c1b5, 32'sh2b7c8a3f, 32'sh2b73511c, 32'sh2b6a164d, 32'sh2b60d9d0, 32'sh2b579ba8, 32'sh2b4e5bd4, 
               32'sh2b451a55, 32'sh2b3bd72a, 32'sh2b329255, 32'sh2b294bd5, 32'sh2b2003ac, 32'sh2b16b9d9, 32'sh2b0d6e5c, 32'sh2b042137, 
               32'sh2afad269, 32'sh2af181f3, 32'sh2ae82fd5, 32'sh2adedc10, 32'sh2ad586a3, 32'sh2acc2f90, 32'sh2ac2d6d6, 32'sh2ab97c77, 
               32'sh2ab02071, 32'sh2aa6c2c6, 32'sh2a9d6377, 32'sh2a940283, 32'sh2a8a9fea, 32'sh2a813bae, 32'sh2a77d5ce, 32'sh2a6e6e4b, 
               32'sh2a650525, 32'sh2a5b9a5d, 32'sh2a522df3, 32'sh2a48bfe7, 32'sh2a3f503a, 32'sh2a35deeb, 32'sh2a2c6bfd, 32'sh2a22f76e, 
               32'sh2a19813f, 32'sh2a100970, 32'sh2a069003, 32'sh29fd14f6, 32'sh29f3984c, 32'sh29ea1a03, 32'sh29e09a1c, 32'sh29d71899, 
               32'sh29cd9578, 32'sh29c410ba, 32'sh29ba8a61, 32'sh29b1026c, 32'sh29a778db, 32'sh299dedaf, 32'sh299460e8, 32'sh298ad287, 
               32'sh2981428c, 32'sh2977b0f7, 32'sh296e1dc9, 32'sh29648902, 32'sh295af2a3, 32'sh29515aab, 32'sh2947c11c, 32'sh293e25f5, 
               32'sh29348937, 32'sh292aeae3, 32'sh29214af8, 32'sh2917a977, 32'sh290e0661, 32'sh290461b5, 32'sh28fabb75, 32'sh28f113a0, 
               32'sh28e76a37, 32'sh28ddbf3b, 32'sh28d412ab, 32'sh28ca6488, 32'sh28c0b4d2, 32'sh28b7038b, 32'sh28ad50b1, 32'sh28a39c46, 
               32'sh2899e64a, 32'sh28902ebd, 32'sh288675a0, 32'sh287cbaf3, 32'sh2872feb6, 32'sh286940ea, 32'sh285f8190, 32'sh2855c0a6, 
               32'sh284bfe2f, 32'sh28423a2a, 32'sh28387498, 32'sh282ead78, 32'sh2824e4cc, 32'sh281b1a94, 32'sh28114ed0, 32'sh28078181, 
               32'sh27fdb2a7, 32'sh27f3e241, 32'sh27ea1052, 32'sh27e03cd8, 32'sh27d667d5, 32'sh27cc9149, 32'sh27c2b934, 32'sh27b8df97, 
               32'sh27af0472, 32'sh27a527c4, 32'sh279b4990, 32'sh279169d5, 32'sh27878893, 32'sh277da5cb, 32'sh2773c17d, 32'sh2769dbaa, 
               32'sh275ff452, 32'sh27560b76, 32'sh274c2115, 32'sh27423530, 32'sh273847c8, 32'sh272e58dc, 32'sh2724686e, 32'sh271a767e, 
               32'sh2710830c, 32'sh27068e18, 32'sh26fc97a3, 32'sh26f29fad, 32'sh26e8a637, 32'sh26deab41, 32'sh26d4aecb, 32'sh26cab0d6, 
               32'sh26c0b162, 32'sh26b6b070, 32'sh26acadff, 32'sh26a2aa11, 32'sh2698a4a6, 32'sh268e9dbd, 32'sh26849558, 32'sh267a8b77, 
               32'sh2670801a, 32'sh26667342, 32'sh265c64ef, 32'sh26525521, 32'sh264843d9, 32'sh263e3117, 32'sh26341cdb, 32'sh262a0727, 
               32'sh261feffa, 32'sh2615d754, 32'sh260bbd37, 32'sh2601a1a2, 32'sh25f78497, 32'sh25ed6614, 32'sh25e3461b, 32'sh25d924ac, 
               32'sh25cf01c8, 32'sh25c4dd6e, 32'sh25bab7a0, 32'sh25b0905d, 32'sh25a667a7, 32'sh259c3d7c, 32'sh259211df, 32'sh2587e4cf, 
               32'sh257db64c, 32'sh25738657, 32'sh256954f1, 32'sh255f2219, 32'sh2554edd1, 32'sh254ab818, 32'sh254080ef, 32'sh25364857, 
               32'sh252c0e4f, 32'sh2521d2d8, 32'sh251795f3, 32'sh250d57a0, 32'sh250317df, 32'sh24f8d6b0, 32'sh24ee9415, 32'sh24e4500e, 
               32'sh24da0a9a, 32'sh24cfc3ba, 32'sh24c57b6f, 32'sh24bb31ba, 32'sh24b0e699, 32'sh24a69a0f, 32'sh249c4c1b, 32'sh2491fcbe, 
               32'sh2487abf7, 32'sh247d59c8, 32'sh24730631, 32'sh2468b132, 32'sh245e5acc, 32'sh245402ff, 32'sh2449a9cc, 32'sh243f4f32, 
               32'sh2434f332, 32'sh242a95ce, 32'sh24203704, 32'sh2415d6d5, 32'sh240b7543, 32'sh2401124d, 32'sh23f6adf3, 32'sh23ec4837, 
               32'sh23e1e117, 32'sh23d77896, 32'sh23cd0eb3, 32'sh23c2a36f, 32'sh23b836ca, 32'sh23adc8c4, 32'sh23a3595e, 32'sh2398e898, 
               32'sh238e7673, 32'sh238402ef, 32'sh23798e0d, 32'sh236f17cc, 32'sh2364a02e, 32'sh235a2733, 32'sh234facda, 32'sh23453125, 
               32'sh233ab414, 32'sh233035a7, 32'sh2325b5df, 32'sh231b34bc, 32'sh2310b23e, 32'sh23062e67, 32'sh22fba936, 32'sh22f122ab, 
               32'sh22e69ac8, 32'sh22dc118c, 32'sh22d186f8, 32'sh22c6fb0c, 32'sh22bc6dca, 32'sh22b1df30, 32'sh22a74f40, 32'sh229cbdfa, 
               32'sh22922b5e, 32'sh2287976e, 32'sh227d0228, 32'sh22726b8e, 32'sh2267d3a0, 32'sh225d3a5e, 32'sh22529fca, 32'sh224803e2, 
               32'sh223d66a8, 32'sh2232c81c, 32'sh2228283f, 32'sh221d8711, 32'sh2212e492, 32'sh220840c2, 32'sh21fd9ba3, 32'sh21f2f534, 
               32'sh21e84d76, 32'sh21dda46a, 32'sh21d2fa0f, 32'sh21c84e67, 32'sh21bda171, 32'sh21b2f32e, 32'sh21a8439e, 32'sh219d92c2, 
               32'sh2192e09b, 32'sh21882d28, 32'sh217d786a, 32'sh2172c262, 32'sh21680b0f, 32'sh215d5273, 32'sh2152988d, 32'sh2147dd5f, 
               32'sh213d20e8, 32'sh21326329, 32'sh2127a423, 32'sh211ce3d5, 32'sh21122240, 32'sh21075f65, 32'sh20fc9b44, 32'sh20f1d5de, 
               32'sh20e70f32, 32'sh20dc4742, 32'sh20d17e0d, 32'sh20c6b395, 32'sh20bbe7d8, 32'sh20b11ad9, 32'sh20a64c97, 32'sh209b7d13, 
               32'sh2090ac4d, 32'sh2085da46, 32'sh207b06fe, 32'sh20703275, 32'sh20655cac, 32'sh205a85a3, 32'sh204fad5b, 32'sh2044d3d4, 
               32'sh2039f90f, 32'sh202f1d0b, 32'sh20243fca, 32'sh2019614c, 32'sh200e8190, 32'sh2003a099, 32'sh1ff8be65, 32'sh1feddaf6, 
               32'sh1fe2f64c, 32'sh1fd81067, 32'sh1fcd2948, 32'sh1fc240ef, 32'sh1fb7575c, 32'sh1fac6c91, 32'sh1fa1808c, 32'sh1f969350, 
               32'sh1f8ba4dc, 32'sh1f80b531, 32'sh1f75c44e, 32'sh1f6ad235, 32'sh1f5fdee6, 32'sh1f54ea62, 32'sh1f49f4a8, 32'sh1f3efdb9, 
               32'sh1f340596, 32'sh1f290c3f, 32'sh1f1e11b5, 32'sh1f1315f7, 32'sh1f081907, 32'sh1efd1ae4, 32'sh1ef21b90, 32'sh1ee71b0a, 
               32'sh1edc1953, 32'sh1ed1166b, 32'sh1ec61254, 32'sh1ebb0d0d, 32'sh1eb00696, 32'sh1ea4fef0, 32'sh1e99f61d, 32'sh1e8eec1b, 
               32'sh1e83e0eb, 32'sh1e78d48e, 32'sh1e6dc705, 32'sh1e62b84f, 32'sh1e57a86d, 32'sh1e4c9760, 32'sh1e418528, 32'sh1e3671c5, 
               32'sh1e2b5d38, 32'sh1e204781, 32'sh1e1530a1, 32'sh1e0a1898, 32'sh1dfeff67, 32'sh1df3e50d, 32'sh1de8c98c, 32'sh1dddace4, 
               32'sh1dd28f15, 32'sh1dc7701f, 32'sh1dbc5004, 32'sh1db12ec3, 32'sh1da60c5d, 32'sh1d9ae8d2, 32'sh1d8fc424, 32'sh1d849e51, 
               32'sh1d79775c, 32'sh1d6e4f43, 32'sh1d632608, 32'sh1d57fbaa, 32'sh1d4cd02c, 32'sh1d41a38c, 32'sh1d3675cb, 32'sh1d2b46ea, 
               32'sh1d2016e9, 32'sh1d14e5c9, 32'sh1d09b389, 32'sh1cfe802b, 32'sh1cf34baf, 32'sh1ce81615, 32'sh1cdcdf5e, 32'sh1cd1a78a, 
               32'sh1cc66e99, 32'sh1cbb348d, 32'sh1caff965, 32'sh1ca4bd21, 32'sh1c997fc4, 32'sh1c8e414b, 32'sh1c8301b9, 32'sh1c77c10e, 
               32'sh1c6c7f4a, 32'sh1c613c6d, 32'sh1c55f878, 32'sh1c4ab36b, 32'sh1c3f6d47, 32'sh1c34260c, 32'sh1c28ddbb, 32'sh1c1d9454, 
               32'sh1c1249d8, 32'sh1c06fe46, 32'sh1bfbb1a0, 32'sh1bf063e6, 32'sh1be51518, 32'sh1bd9c537, 32'sh1bce7442, 32'sh1bc3223c, 
               32'sh1bb7cf23, 32'sh1bac7af9, 32'sh1ba125bd, 32'sh1b95cf71, 32'sh1b8a7815, 32'sh1b7f1fa9, 32'sh1b73c62d, 32'sh1b686ba3, 
               32'sh1b5d100a, 32'sh1b51b363, 32'sh1b4655ae, 32'sh1b3af6ec, 32'sh1b2f971e, 32'sh1b243643, 32'sh1b18d45c, 32'sh1b0d716a, 
               32'sh1b020d6c, 32'sh1af6a865, 32'sh1aeb4253, 32'sh1adfdb37, 32'sh1ad47312, 32'sh1ac909e5, 32'sh1abd9faf, 32'sh1ab23471, 
               32'sh1aa6c82b, 32'sh1a9b5adf, 32'sh1a8fec8c, 32'sh1a847d33, 32'sh1a790cd4, 32'sh1a6d9b70, 32'sh1a622907, 32'sh1a56b599, 
               32'sh1a4b4128, 32'sh1a3fcbb3, 32'sh1a34553b, 32'sh1a28ddc0, 32'sh1a1d6544, 32'sh1a11ebc5, 32'sh1a067145, 32'sh19faf5c5, 
               32'sh19ef7944, 32'sh19e3fbc3, 32'sh19d87d42, 32'sh19ccfdc2, 32'sh19c17d44, 32'sh19b5fbc8, 32'sh19aa794d, 32'sh199ef5d6, 
               32'sh19937161, 32'sh1987ebf0, 32'sh197c6584, 32'sh1970de1b, 32'sh196555b8, 32'sh1959cc5a, 32'sh194e4201, 32'sh1942b6af, 
               32'sh19372a64, 32'sh192b9d1f, 32'sh19200ee3, 32'sh19147fae, 32'sh1908ef82, 32'sh18fd5e5f, 32'sh18f1cc45, 32'sh18e63935, 
               32'sh18daa52f, 32'sh18cf1034, 32'sh18c37a44, 32'sh18b7e35f, 32'sh18ac4b87, 32'sh18a0b2bb, 32'sh189518fc, 32'sh18897e4a, 
               32'sh187de2a7, 32'sh18724611, 32'sh1866a88a, 32'sh185b0a13, 32'sh184f6aab, 32'sh1843ca53, 32'sh1838290c, 32'sh182c86d5, 
               32'sh1820e3b0, 32'sh18153f9d, 32'sh18099a9c, 32'sh17fdf4ae, 32'sh17f24dd3, 32'sh17e6a60c, 32'sh17dafd59, 32'sh17cf53bb, 
               32'sh17c3a931, 32'sh17b7fdbd, 32'sh17ac515f, 32'sh17a0a417, 32'sh1794f5e6, 32'sh178946cc, 32'sh177d96ca, 32'sh1771e5e0, 
               32'sh1766340f, 32'sh175a8157, 32'sh174ecdb8, 32'sh17431933, 32'sh173763c9, 32'sh172bad7a, 32'sh171ff646, 32'sh17143e2d, 
               32'sh17088531, 32'sh16fccb51, 32'sh16f1108f, 32'sh16e554ea, 32'sh16d99864, 32'sh16cddafb, 32'sh16c21cb2, 32'sh16b65d88, 
               32'sh16aa9d7e, 32'sh169edc94, 32'sh16931acb, 32'sh16875823, 32'sh167b949d, 32'sh166fd039, 32'sh16640af7, 32'sh165844d8, 
               32'sh164c7ddd, 32'sh1640b606, 32'sh1634ed53, 32'sh162923c5, 32'sh161d595d, 32'sh16118e1a, 32'sh1605c1fd, 32'sh15f9f507, 
               32'sh15ee2738, 32'sh15e25890, 32'sh15d68911, 32'sh15cab8ba, 32'sh15bee78c, 32'sh15b31587, 32'sh15a742ac, 32'sh159b6efb, 
               32'sh158f9a76, 32'sh1583c51b, 32'sh1577eeec, 32'sh156c17e9, 32'sh15604013, 32'sh1554676a, 32'sh15488dee, 32'sh153cb3a0, 
               32'sh1530d881, 32'sh1524fc90, 32'sh15191fcf, 32'sh150d423d, 32'sh150163dc, 32'sh14f584ac, 32'sh14e9a4ac, 32'sh14ddc3de, 
               32'sh14d1e242, 32'sh14c5ffd9, 32'sh14ba1ca3, 32'sh14ae38a0, 32'sh14a253d1, 32'sh14966e36, 32'sh148a87d1, 32'sh147ea0a0, 
               32'sh1472b8a5, 32'sh1466cfe1, 32'sh145ae653, 32'sh144efbfc, 32'sh144310dd, 32'sh143724f5, 32'sh142b3846, 32'sh141f4ad1, 
               32'sh14135c94, 32'sh14076d91, 32'sh13fb7dc9, 32'sh13ef8d3c, 32'sh13e39be9, 32'sh13d7a9d3, 32'sh13cbb6f8, 32'sh13bfc35b, 
               32'sh13b3cefa, 32'sh13a7d9d7, 32'sh139be3f2, 32'sh138fed4b, 32'sh1383f5e3, 32'sh1377fdbb, 32'sh136c04d2, 32'sh13600b2a, 
               32'sh135410c3, 32'sh1348159d, 32'sh133c19b8, 32'sh13301d16, 32'sh13241fb6, 32'sh1318219a, 32'sh130c22c1, 32'sh1300232c, 
               32'sh12f422db, 32'sh12e821cf, 32'sh12dc2009, 32'sh12d01d89, 32'sh12c41a4f, 32'sh12b8165b, 32'sh12ac11af, 32'sh12a00c4b, 
               32'sh1294062f, 32'sh1287ff5b, 32'sh127bf7d1, 32'sh126fef90, 32'sh1263e699, 32'sh1257dced, 32'sh124bd28c, 32'sh123fc776, 
               32'sh1233bbac, 32'sh1227af2e, 32'sh121ba1fd, 32'sh120f941a, 32'sh12038584, 32'sh11f7763c, 32'sh11eb6643, 32'sh11df5599, 
               32'sh11d3443f, 32'sh11c73235, 32'sh11bb1f7c, 32'sh11af0c13, 32'sh11a2f7fc, 32'sh1196e337, 32'sh118acdc4, 32'sh117eb7a4, 
               32'sh1172a0d7, 32'sh1166895f, 32'sh115a713a, 32'sh114e586a, 32'sh11423ef0, 32'sh113624cb, 32'sh112a09fc, 32'sh111dee84, 
               32'sh1111d263, 32'sh1105b599, 32'sh10f99827, 32'sh10ed7a0e, 32'sh10e15b4e, 32'sh10d53be7, 32'sh10c91bda, 32'sh10bcfb28, 
               32'sh10b0d9d0, 32'sh10a4b7d3, 32'sh10989532, 32'sh108c71ee, 32'sh10804e06, 32'sh1074297b, 32'sh1068044e, 32'sh105bde7f, 
               32'sh104fb80e, 32'sh104390fd, 32'sh1037694b, 32'sh102b40f8, 32'sh101f1807, 32'sh1012ee76, 32'sh1006c446, 32'sh0ffa9979, 
               32'sh0fee6e0d, 32'sh0fe24205, 32'sh0fd6155f, 32'sh0fc9e81e, 32'sh0fbdba40, 32'sh0fb18bc8, 32'sh0fa55cb4, 32'sh0f992d06, 
               32'sh0f8cfcbe, 32'sh0f80cbdc, 32'sh0f749a61, 32'sh0f68684e, 32'sh0f5c35a3, 32'sh0f500260, 32'sh0f43ce86, 32'sh0f379a16, 
               32'sh0f2b650f, 32'sh0f1f2f73, 32'sh0f12f941, 32'sh0f06c27a, 32'sh0efa8b20, 32'sh0eee5331, 32'sh0ee21aaf, 32'sh0ed5e19a, 
               32'sh0ec9a7f3, 32'sh0ebd6db9, 32'sh0eb132ef, 32'sh0ea4f793, 32'sh0e98bba7, 32'sh0e8c7f2a, 32'sh0e80421e, 32'sh0e740483, 
               32'sh0e67c65a, 32'sh0e5b87a2, 32'sh0e4f485c, 32'sh0e430889, 32'sh0e36c82a, 32'sh0e2a873e, 32'sh0e1e45c6, 32'sh0e1203c3, 
               32'sh0e05c135, 32'sh0df97e1d, 32'sh0ded3a7b, 32'sh0de0f64f, 32'sh0dd4b19a, 32'sh0dc86c5d, 32'sh0dbc2698, 32'sh0dafe04b, 
               32'sh0da39978, 32'sh0d97521d, 32'sh0d8b0a3d, 32'sh0d7ec1d6, 32'sh0d7278eb, 32'sh0d662f7b, 32'sh0d59e586, 32'sh0d4d9b0e, 
               32'sh0d415013, 32'sh0d350495, 32'sh0d28b894, 32'sh0d1c6c11, 32'sh0d101f0e, 32'sh0d03d189, 32'sh0cf78383, 32'sh0ceb34fe, 
               32'sh0cdee5f9, 32'sh0cd29676, 32'sh0cc64673, 32'sh0cb9f5f3, 32'sh0cada4f5, 32'sh0ca1537a, 32'sh0c950182, 32'sh0c88af0e, 
               32'sh0c7c5c1e, 32'sh0c7008b3, 32'sh0c63b4ce, 32'sh0c57606e, 32'sh0c4b0b94, 32'sh0c3eb641, 32'sh0c326075, 32'sh0c260a31, 
               32'sh0c19b374, 32'sh0c0d5c41, 32'sh0c010496, 32'sh0bf4ac75, 32'sh0be853de, 32'sh0bdbfad1, 32'sh0bcfa150, 32'sh0bc34759, 
               32'sh0bb6ecef, 32'sh0baa9211, 32'sh0b9e36c0, 32'sh0b91dafc, 32'sh0b857ec7, 32'sh0b79221f, 32'sh0b6cc506, 32'sh0b60677c, 
               32'sh0b540982, 32'sh0b47ab19, 32'sh0b3b4c40, 32'sh0b2eecf8, 32'sh0b228d42, 32'sh0b162d1d, 32'sh0b09cc8c, 32'sh0afd6b8d, 
               32'sh0af10a22, 32'sh0ae4a84b, 32'sh0ad84609, 32'sh0acbe35b, 32'sh0abf8043, 32'sh0ab31cc1, 32'sh0aa6b8d5, 32'sh0a9a5480, 
               32'sh0a8defc3, 32'sh0a818a9d, 32'sh0a752510, 32'sh0a68bf1b, 32'sh0a5c58c0, 32'sh0a4ff1fe, 32'sh0a438ad7, 32'sh0a37234a, 
               32'sh0a2abb59, 32'sh0a1e5303, 32'sh0a11ea49, 32'sh0a05812c, 32'sh09f917ac, 32'sh09ecadc9, 32'sh09e04385, 32'sh09d3d8df, 
               32'sh09c76dd8, 32'sh09bb0271, 32'sh09ae96aa, 32'sh09a22a83, 32'sh0995bdfd, 32'sh09895118, 32'sh097ce3d5, 32'sh09707635, 
               32'sh09640837, 32'sh095799dd, 32'sh094b2b27, 32'sh093ebc14, 32'sh09324ca7, 32'sh0925dcdf, 32'sh09196cbc, 32'sh090cfc40, 
               32'sh09008b6a, 32'sh08f41a3c, 32'sh08e7a8b5, 32'sh08db36d6, 32'sh08cec4a0, 32'sh08c25213, 32'sh08b5df30, 32'sh08a96bf6, 
               32'sh089cf867, 32'sh08908483, 32'sh0884104b, 32'sh08779bbe, 32'sh086b26de, 32'sh085eb1ab, 32'sh08523c25, 32'sh0845c64d, 
               32'sh08395024, 32'sh082cd9a9, 32'sh082062de, 32'sh0813ebc2, 32'sh08077457, 32'sh07fafc9c, 32'sh07ee8493, 32'sh07e20c3b, 
               32'sh07d59396, 32'sh07c91aa3, 32'sh07bca163, 32'sh07b027d7, 32'sh07a3adff, 32'sh079733dc, 32'sh078ab96e, 32'sh077e3eb5, 
               32'sh0771c3b3, 32'sh07654867, 32'sh0758ccd2, 32'sh074c50f4, 32'sh073fd4cf, 32'sh07335862, 32'sh0726dbae, 32'sh071a5eb3, 
               32'sh070de172, 32'sh070163eb, 32'sh06f4e620, 32'sh06e86810, 32'sh06dbe9bb, 32'sh06cf6b23, 32'sh06c2ec48, 32'sh06b66d29, 
               32'sh06a9edc9, 32'sh069d6e27, 32'sh0690ee44, 32'sh06846e1f, 32'sh0677edbb, 32'sh066b6d16, 32'sh065eec33, 32'sh06526b10, 
               32'sh0645e9af, 32'sh06396810, 32'sh062ce634, 32'sh0620641a, 32'sh0613e1c5, 32'sh06075f33, 32'sh05fadc66, 32'sh05ee595d, 
               32'sh05e1d61b, 32'sh05d5529e, 32'sh05c8cee7, 32'sh05bc4af8, 32'sh05afc6d0, 32'sh05a3426f, 32'sh0596bdd7, 32'sh058a3908, 
               32'sh057db403, 32'sh05712ec7, 32'sh0564a955, 32'sh055823ae, 32'sh054b9dd3, 32'sh053f17c3, 32'sh0532917f, 32'sh05260b08, 
               32'sh0519845e, 32'sh050cfd82, 32'sh05007674, 32'sh04f3ef35, 32'sh04e767c5, 32'sh04dae024, 32'sh04ce5854, 32'sh04c1d054, 
               32'sh04b54825, 32'sh04a8bfc7, 32'sh049c373c, 32'sh048fae83, 32'sh0483259d, 32'sh04769c8b, 32'sh046a134c, 32'sh045d89e2, 
               32'sh0451004d, 32'sh0444768d, 32'sh0437eca4, 32'sh042b6290, 32'sh041ed854, 32'sh04124dee, 32'sh0405c361, 32'sh03f938ac, 
               32'sh03ecadcf, 32'sh03e022cc, 32'sh03d397a3, 32'sh03c70c54, 32'sh03ba80df, 32'sh03adf546, 32'sh03a16988, 32'sh0394dda7, 
               32'sh038851a2, 32'sh037bc57b, 32'sh036f3931, 32'sh0362acc5, 32'sh03562038, 32'sh03499389, 32'sh033d06bb, 32'sh033079cc, 
               32'sh0323ecbe, 32'sh03175f91, 32'sh030ad245, 32'sh02fe44dc, 32'sh02f1b755, 32'sh02e529b0, 32'sh02d89bf0, 32'sh02cc0e13, 
               32'sh02bf801a, 32'sh02b2f207, 32'sh02a663d8, 32'sh0299d590, 32'sh028d472e, 32'sh0280b8b3, 32'sh02742a1f, 32'sh02679b73, 
               32'sh025b0caf, 32'sh024e7dd4, 32'sh0241eee2, 32'sh02355fd9, 32'sh0228d0bb, 32'sh021c4188, 32'sh020fb240, 32'sh020322e3, 
               32'sh01f69373, 32'sh01ea03ef, 32'sh01dd7459, 32'sh01d0e4b0, 32'sh01c454f5, 32'sh01b7c528, 32'sh01ab354b, 32'sh019ea55d, 
               32'sh0192155f, 32'sh01858552, 32'sh0178f536, 32'sh016c650b, 32'sh015fd4d2, 32'sh0153448c, 32'sh0146b438, 32'sh013a23d8, 
               32'sh012d936c, 32'sh012102f4, 32'sh01147271, 32'sh0107e1e3, 32'sh00fb514b, 32'sh00eec0aa, 32'sh00e22fff, 32'sh00d59f4c, 
               32'sh00c90e90, 32'sh00bc7dcc, 32'sh00afed02, 32'sh00a35c30, 32'sh0096cb58, 32'sh008a3a7b, 32'sh007da998, 32'sh007118b0, 
               32'sh006487c4, 32'sh0057f6d4, 32'sh004b65e1, 32'sh003ed4ea, 32'sh003243f1, 32'sh0025b2f7, 32'sh001921fb, 32'sh000c90fe, 
               32'sh00000000, 32'shfff36f02, 32'shffe6de05, 32'shffda4d09, 32'shffcdbc0f, 32'shffc12b16, 32'shffb49a1f, 32'shffa8092c, 
               32'shff9b783c, 32'shff8ee750, 32'shff825668, 32'shff75c585, 32'shff6934a8, 32'shff5ca3d0, 32'shff5012fe, 32'shff438234, 
               32'shff36f170, 32'shff2a60b4, 32'shff1dd001, 32'shff113f56, 32'shff04aeb5, 32'shfef81e1d, 32'shfeeb8d8f, 32'shfedefd0c, 
               32'shfed26c94, 32'shfec5dc28, 32'shfeb94bc8, 32'shfeacbb74, 32'shfea02b2e, 32'shfe939af5, 32'shfe870aca, 32'shfe7a7aae, 
               32'shfe6deaa1, 32'shfe615aa3, 32'shfe54cab5, 32'shfe483ad8, 32'shfe3bab0b, 32'shfe2f1b50, 32'shfe228ba7, 32'shfe15fc11, 
               32'shfe096c8d, 32'shfdfcdd1d, 32'shfdf04dc0, 32'shfde3be78, 32'shfdd72f45, 32'shfdcaa027, 32'shfdbe111e, 32'shfdb1822c, 
               32'shfda4f351, 32'shfd98648d, 32'shfd8bd5e1, 32'shfd7f474d, 32'shfd72b8d2, 32'shfd662a70, 32'shfd599c28, 32'shfd4d0df9, 
               32'shfd407fe6, 32'shfd33f1ed, 32'shfd276410, 32'shfd1ad650, 32'shfd0e48ab, 32'shfd01bb24, 32'shfcf52dbb, 32'shfce8a06f, 
               32'shfcdc1342, 32'shfccf8634, 32'shfcc2f945, 32'shfcb66c77, 32'shfca9dfc8, 32'shfc9d533b, 32'shfc90c6cf, 32'shfc843a85, 
               32'shfc77ae5e, 32'shfc6b2259, 32'shfc5e9678, 32'shfc520aba, 32'shfc457f21, 32'shfc38f3ac, 32'shfc2c685d, 32'shfc1fdd34, 
               32'shfc135231, 32'shfc06c754, 32'shfbfa3c9f, 32'shfbedb212, 32'shfbe127ac, 32'shfbd49d70, 32'shfbc8135c, 32'shfbbb8973, 
               32'shfbaeffb3, 32'shfba2761e, 32'shfb95ecb4, 32'shfb896375, 32'shfb7cda63, 32'shfb70517d, 32'shfb63c8c4, 32'shfb574039, 
               32'shfb4ab7db, 32'shfb3e2fac, 32'shfb31a7ac, 32'shfb251fdc, 32'shfb18983b, 32'shfb0c10cb, 32'shfaff898c, 32'shfaf3027e, 
               32'shfae67ba2, 32'shfad9f4f8, 32'shfacd6e81, 32'shfac0e83d, 32'shfab4622d, 32'shfaa7dc52, 32'shfa9b56ab, 32'shfa8ed139, 
               32'shfa824bfd, 32'shfa75c6f8, 32'shfa694229, 32'shfa5cbd91, 32'shfa503930, 32'shfa43b508, 32'shfa373119, 32'shfa2aad62, 
               32'shfa1e29e5, 32'shfa11a6a3, 32'shfa05239a, 32'shf9f8a0cd, 32'shf9ec1e3b, 32'shf9df9be6, 32'shf9d319cc, 32'shf9c697f0, 
               32'shf9ba1651, 32'shf9ad94f0, 32'shf9a113cd, 32'shf99492ea, 32'shf9881245, 32'shf97b91e1, 32'shf96f11bc, 32'shf96291d9, 
               32'shf9561237, 32'shf94992d7, 32'shf93d13b8, 32'shf93094dd, 32'shf9241645, 32'shf91797f0, 32'shf90b19e0, 32'shf8fe9c15, 
               32'shf8f21e8e, 32'shf8e5a14d, 32'shf8d92452, 32'shf8cca79e, 32'shf8c02b31, 32'shf8b3af0c, 32'shf8a7332e, 32'shf89ab799, 
               32'shf88e3c4d, 32'shf881c14b, 32'shf8754692, 32'shf868cc24, 32'shf85c5201, 32'shf84fd829, 32'shf8435e9d, 32'shf836e55d, 
               32'shf82a6c6a, 32'shf81df3c5, 32'shf8117b6d, 32'shf8050364, 32'shf7f88ba9, 32'shf7ec143e, 32'shf7df9d22, 32'shf7d32657, 
               32'shf7c6afdc, 32'shf7ba39b3, 32'shf7adc3db, 32'shf7a14e55, 32'shf794d922, 32'shf7886442, 32'shf77befb5, 32'shf76f7b7d, 
               32'shf7630799, 32'shf756940a, 32'shf74a20d0, 32'shf73daded, 32'shf7313b60, 32'shf724c92a, 32'shf718574b, 32'shf70be5c4, 
               32'shf6ff7496, 32'shf6f303c0, 32'shf6e69344, 32'shf6da2321, 32'shf6cdb359, 32'shf6c143ec, 32'shf6b4d4d9, 32'shf6a86623, 
               32'shf69bf7c9, 32'shf68f89cb, 32'shf6831c2b, 32'shf676aee8, 32'shf66a4203, 32'shf65dd57d, 32'shf6516956, 32'shf644fd8f, 
               32'shf6389228, 32'shf62c2721, 32'shf61fbc7b, 32'shf6135237, 32'shf606e854, 32'shf5fa7ed4, 32'shf5ee15b7, 32'shf5e1acfd, 
               32'shf5d544a7, 32'shf5c8dcb6, 32'shf5bc7529, 32'shf5b00e02, 32'shf5a3a740, 32'shf59740e5, 32'shf58adaf0, 32'shf57e7563, 
               32'shf572103d, 32'shf565ab80, 32'shf559472b, 32'shf54ce33f, 32'shf5407fbd, 32'shf5341ca5, 32'shf527b9f7, 32'shf51b57b5, 
               32'shf50ef5de, 32'shf5029473, 32'shf4f63374, 32'shf4e9d2e3, 32'shf4dd72be, 32'shf4d11308, 32'shf4c4b3c0, 32'shf4b854e7, 
               32'shf4abf67e, 32'shf49f9884, 32'shf4933afa, 32'shf486dde1, 32'shf47a8139, 32'shf46e2504, 32'shf461c940, 32'shf4556def, 
               32'shf4491311, 32'shf43cb8a7, 32'shf4305eb0, 32'shf424052f, 32'shf417ac22, 32'shf40b538b, 32'shf3fefb6a, 32'shf3f2a3bf, 
               32'shf3e64c8c, 32'shf3d9f5cf, 32'shf3cd9f8b, 32'shf3c149bf, 32'shf3b4f46c, 32'shf3a89f92, 32'shf39c4b32, 32'shf38ff74d, 
               32'shf383a3e2, 32'shf37750f2, 32'shf36afe7e, 32'shf35eac86, 32'shf3525b0b, 32'shf3460a0d, 32'shf339b98d, 32'shf32d698a, 
               32'shf3211a07, 32'shf314cb02, 32'shf3087c7d, 32'shf2fc2e77, 32'shf2efe0f2, 32'shf2e393ef, 32'shf2d7476c, 32'shf2cafb6b, 
               32'shf2beafed, 32'shf2b264f2, 32'shf2a61a7a, 32'shf299d085, 32'shf28d8715, 32'shf2813e2a, 32'shf274f5c3, 32'shf268ade3, 
               32'shf25c6688, 32'shf2501fb5, 32'shf243d968, 32'shf23793a3, 32'shf22b4e66, 32'shf21f09b1, 32'shf212c585, 32'shf20681e3, 
               32'shf1fa3ecb, 32'shf1edfc3d, 32'shf1e1ba3a, 32'shf1d578c2, 32'shf1c937d6, 32'shf1bcf777, 32'shf1b0b7a4, 32'shf1a4785e, 
               32'shf19839a6, 32'shf18bfb7d, 32'shf17fbde2, 32'shf17380d6, 32'shf1674459, 32'shf15b086d, 32'shf14ecd11, 32'shf1429247, 
               32'shf136580d, 32'shf12a1e66, 32'shf11de551, 32'shf111accf, 32'shf10574e0, 32'shf0f93d86, 32'shf0ed06bf, 32'shf0e0d08d, 
               32'shf0d49af1, 32'shf0c865ea, 32'shf0bc317a, 32'shf0affda0, 32'shf0a3ca5d, 32'shf09797b2, 32'shf08b659f, 32'shf07f3424, 
               32'shf0730342, 32'shf066d2fa, 32'shf05aa34c, 32'shf04e7438, 32'shf04245c0, 32'shf03617e2, 32'shf029eaa1, 32'shf01dbdfb, 
               32'shf01191f3, 32'shf0056687, 32'sheff93bba, 32'shefed118a, 32'shefe0e7f9, 32'shefd4bf08, 32'shefc896b5, 32'shefbc6f03, 
               32'shefb047f2, 32'shefa42181, 32'shef97fbb2, 32'shef8bd685, 32'shef7fb1fa, 32'shef738e12, 32'shef676ace, 32'shef5b482d, 
               32'shef4f2630, 32'shef4304d8, 32'shef36e426, 32'shef2ac419, 32'shef1ea4b2, 32'shef1285f2, 32'shef0667d9, 32'sheefa4a67, 
               32'sheeee2d9d, 32'sheee2117c, 32'sheed5f604, 32'sheec9db35, 32'sheebdc110, 32'sheeb1a796, 32'sheea58ec6, 32'shee9976a1, 
               32'shee8d5f29, 32'shee81485c, 32'shee75323c, 32'shee691cc9, 32'shee5d0804, 32'shee50f3ed, 32'shee44e084, 32'shee38cdcb, 
               32'shee2cbbc1, 32'shee20aa67, 32'shee1499bd, 32'shee0889c4, 32'shedfc7a7c, 32'shedf06be6, 32'shede45e03, 32'shedd850d2, 
               32'shedcc4454, 32'shedc0388a, 32'shedb42d74, 32'sheda82313, 32'shed9c1967, 32'shed901070, 32'shed84082f, 32'shed7800a5, 
               32'shed6bf9d1, 32'shed5ff3b5, 32'shed53ee51, 32'shed47e9a5, 32'shed3be5b1, 32'shed2fe277, 32'shed23dff7, 32'shed17de31, 
               32'shed0bdd25, 32'shecffdcd4, 32'shecf3dd3f, 32'shece7de66, 32'shecdbe04a, 32'sheccfe2ea, 32'shecc3e648, 32'shecb7ea63, 
               32'shecabef3d, 32'shec9ff4d6, 32'shec93fb2e, 32'shec880245, 32'shec7c0a1d, 32'shec7012b5, 32'shec641c0e, 32'shec582629, 
               32'shec4c3106, 32'shec403ca5, 32'shec344908, 32'shec28562d, 32'shec1c6417, 32'shec1072c4, 32'shec048237, 32'shebf8926f, 
               32'shebeca36c, 32'shebe0b52f, 32'shebd4c7ba, 32'shebc8db0b, 32'shebbcef23, 32'shebb10404, 32'sheba519ad, 32'sheb99301f, 
               32'sheb8d475b, 32'sheb815f60, 32'sheb75782f, 32'sheb6991ca, 32'sheb5dac2f, 32'sheb51c760, 32'sheb45e35d, 32'sheb3a0027, 
               32'sheb2e1dbe, 32'sheb223c22, 32'sheb165b54, 32'sheb0a7b54, 32'sheafe9c24, 32'sheaf2bdc3, 32'sheae6e031, 32'sheadb0370, 
               32'sheacf277f, 32'sheac34c60, 32'sheab77212, 32'sheaab9896, 32'shea9fbfed, 32'shea93e817, 32'shea881114, 32'shea7c3ae5, 
               32'shea70658a, 32'shea649105, 32'shea58bd54, 32'shea4cea79, 32'shea411874, 32'shea354746, 32'shea2976ef, 32'shea1da770, 
               32'shea11d8c8, 32'shea060af9, 32'she9fa3e03, 32'she9ee71e6, 32'she9e2a6a3, 32'she9d6dc3b, 32'she9cb12ad, 32'she9bf49fa, 
               32'she9b38223, 32'she9a7bb28, 32'she99bf509, 32'she9902fc7, 32'she9846b63, 32'she978a7dd, 32'she96ce535, 32'she961236c, 
               32'she9556282, 32'she949a278, 32'she93de34e, 32'she9322505, 32'she926679c, 32'she91aab16, 32'she90eef71, 32'she90334af, 
               32'she8f77acf, 32'she8ebc1d3, 32'she8e009ba, 32'she8d45286, 32'she8c89c37, 32'she8bce6cd, 32'she8b13248, 32'she8a57ea9, 
               32'she899cbf1, 32'she88e1a20, 32'she8826936, 32'she876b934, 32'she86b0a1a, 32'she85f5be9, 32'she853aea1, 32'she8480243, 
               32'she83c56cf, 32'she830ac45, 32'she82502a7, 32'she81959f4, 32'she80db22d, 32'she8020b52, 32'she7f66564, 32'she7eac063, 
               32'she7df1c50, 32'she7d3792b, 32'she7c7d6f4, 32'she7bc35ad, 32'she7b09555, 32'she7a4f5ed, 32'she7995776, 32'she78db9ef, 
               32'she7821d59, 32'she77681b6, 32'she76ae704, 32'she75f4d45, 32'she753b479, 32'she7481ca1, 32'she73c85bc, 32'she730efcc, 
               32'she7255ad1, 32'she719c6cb, 32'she70e33bb, 32'she702a1a1, 32'she6f7107e, 32'she6eb8052, 32'she6dff11d, 32'she6d462e1, 
               32'she6c8d59c, 32'she6bd4951, 32'she6b1bdff, 32'she6a633a6, 32'she69aaa48, 32'she68f21e5, 32'she6839a7c, 32'she6781410, 
               32'she66c8e9f, 32'she6610a2a, 32'she65586b3, 32'she64a0438, 32'she63e82bc, 32'she633023e, 32'she62782be, 32'she61c043d, 
               32'she61086bc, 32'she6050a3b, 32'she5f98ebb, 32'she5ee143b, 32'she5e29abc, 32'she5d72240, 32'she5cbaac5, 32'she5c0344d, 
               32'she5b4bed8, 32'she5a94a67, 32'she59dd6f9, 32'she5926490, 32'she586f32c, 32'she57b82cd, 32'she5701374, 32'she564a521, 
               32'she55937d5, 32'she54dcb8f, 32'she5426051, 32'she536f61b, 32'she52b8cee, 32'she52024c9, 32'she514bdad, 32'she509579b, 
               32'she4fdf294, 32'she4f28e96, 32'she4e72ba4, 32'she4dbc9bd, 32'she4d068e2, 32'she4c50914, 32'she4b9aa52, 32'she4ae4c9d, 
               32'she4a2eff6, 32'she497945d, 32'she48c39d3, 32'she480e057, 32'she47587eb, 32'she46a308f, 32'she45eda43, 32'she4538507, 
               32'she44830dd, 32'she43cddc4, 32'she4318bbe, 32'she4263ac9, 32'she41aeae8, 32'she40f9c1a, 32'she4044e60, 32'she3f901ba, 
               32'she3edb628, 32'she3e26bac, 32'she3d72245, 32'she3cbd9f4, 32'she3c092b9, 32'she3b54c95, 32'she3aa0788, 32'she39ec393, 
               32'she39380b6, 32'she3883ef2, 32'she37cfe47, 32'she371beb5, 32'she366803c, 32'she35b42df, 32'she350069b, 32'she344cb73, 
               32'she3399167, 32'she32e5876, 32'she32320a2, 32'she317e9eb, 32'she30cb451, 32'she3017fd5, 32'she2f64c77, 32'she2eb1a37, 
               32'she2dfe917, 32'she2d4b916, 32'she2c98a35, 32'she2be5c74, 32'she2b32fd4, 32'she2a80456, 32'she29cd9f8, 32'she291b0bd, 
               32'she28688a4, 32'she27b61af, 32'she2703bdc, 32'she265172e, 32'she259f3a3, 32'she24ed13d, 32'she243affc, 32'she2388fe1, 
               32'she22d70eb, 32'she222531c, 32'she2173674, 32'she20c1af3, 32'she2010099, 32'she1f5e768, 32'she1eacf5f, 32'she1dfb87f, 
               32'she1d4a2c8, 32'she1c98e3b, 32'she1be7ad8, 32'she1b368a0, 32'she1a85793, 32'she19d47b1, 32'she19238fb, 32'she1872b72, 
               32'she17c1f15, 32'she17113e5, 32'she16609e3, 32'she15b0110, 32'she14ff96a, 32'she144f2f3, 32'she139edac, 32'she12ee995, 
               32'she123e6ad, 32'she118e4f6, 32'she10de470, 32'she102e51c, 32'she0f7e6f9, 32'she0ecea09, 32'she0e1ee4b, 32'she0d6f3c1, 
               32'she0cbfa6a, 32'she0c10247, 32'she0b60b58, 32'she0ab159e, 32'she0a0211a, 32'she0952dcb, 32'she08a3bb2, 32'she07f4acf, 
               32'she0745b24, 32'she0696cb0, 32'she05e7f74, 32'she053936f, 32'she048a8a4, 32'she03dbf11, 32'she032d6b8, 32'she027ef99, 
               32'she01d09b4, 32'she012250a, 32'she007419b, 32'shdffc5f67, 32'shdff17e70, 32'shdfe69eb4, 32'shdfdbc036, 32'shdfd0e2f5, 
               32'shdfc606f1, 32'shdfbb2c2c, 32'shdfb052a5, 32'shdfa57a5d, 32'shdf9aa354, 32'shdf8fcd8b, 32'shdf84f902, 32'shdf7a25ba, 
               32'shdf6f53b3, 32'shdf6482ed, 32'shdf59b369, 32'shdf4ee527, 32'shdf441828, 32'shdf394c6b, 32'shdf2e81f3, 32'shdf23b8be, 
               32'shdf18f0ce, 32'shdf0e2a22, 32'shdf0364bc, 32'shdef8a09b, 32'shdeedddc0, 32'shdee31c2b, 32'shded85bdd, 32'shdecd9cd7, 
               32'shdec2df18, 32'shdeb822a1, 32'shdead6773, 32'shdea2ad8d, 32'shde97f4f1, 32'shde8d3d9e, 32'shde828796, 32'shde77d2d8, 
               32'shde6d1f65, 32'shde626d3e, 32'shde57bc62, 32'shde4d0cd2, 32'shde425e8f, 32'shde37b199, 32'shde2d05f1, 32'shde225b96, 
               32'shde17b28a, 32'shde0d0acc, 32'shde02645d, 32'shddf7bf3e, 32'shdded1b6e, 32'shdde278ef, 32'shddd7d7c1, 32'shddcd37e4, 
               32'shddc29958, 32'shddb7fc1e, 32'shddad6036, 32'shdda2c5a2, 32'shdd982c60, 32'shdd8d9472, 32'shdd82fdd8, 32'shdd786892, 
               32'shdd6dd4a2, 32'shdd634206, 32'shdd58b0c0, 32'shdd4e20d0, 32'shdd439236, 32'shdd3904f4, 32'shdd2e7908, 32'shdd23ee74, 
               32'shdd196538, 32'shdd0edd55, 32'shdd0456ca, 32'shdcf9d199, 32'shdcef4dc2, 32'shdce4cb44, 32'shdcda4a21, 32'shdccfca59, 
               32'shdcc54bec, 32'shdcbacedb, 32'shdcb05326, 32'shdca5d8cd, 32'shdc9b5fd2, 32'shdc90e834, 32'shdc8671f3, 32'shdc7bfd11, 
               32'shdc71898d, 32'shdc671768, 32'shdc5ca6a2, 32'shdc52373c, 32'shdc47c936, 32'shdc3d5c91, 32'shdc32f14d, 32'shdc28876a, 
               32'shdc1e1ee9, 32'shdc13b7c9, 32'shdc09520d, 32'shdbfeedb3, 32'shdbf48abd, 32'shdbea292b, 32'shdbdfc8fc, 32'shdbd56a32, 
               32'shdbcb0cce, 32'shdbc0b0ce, 32'shdbb65634, 32'shdbabfd01, 32'shdba1a534, 32'shdb974ece, 32'shdb8cf9cf, 32'shdb82a638, 
               32'shdb785409, 32'shdb6e0342, 32'shdb63b3e5, 32'shdb5965f1, 32'shdb4f1967, 32'shdb44ce46, 32'shdb3a8491, 32'shdb303c46, 
               32'shdb25f566, 32'shdb1baff2, 32'shdb116beb, 32'shdb072950, 32'shdafce821, 32'shdaf2a860, 32'shdae86a0d, 32'shdade2d28, 
               32'shdad3f1b1, 32'shdac9b7a9, 32'shdabf7f11, 32'shdab547e8, 32'shdaab122f, 32'shdaa0dde7, 32'shda96ab0f, 32'shda8c79a9, 
               32'shda8249b4, 32'shda781b31, 32'shda6dee21, 32'shda63c284, 32'shda599859, 32'shda4f6fa3, 32'shda454860, 32'shda3b2292, 
               32'shda30fe38, 32'shda26db54, 32'shda1cb9e5, 32'shda1299ec, 32'shda087b69, 32'shd9fe5e5e, 32'shd9f442c9, 32'shd9ea28ac, 
               32'shd9e01006, 32'shd9d5f8d9, 32'shd9cbe325, 32'shd9c1cee9, 32'shd9b7bc27, 32'shd9adaadf, 32'shd9a39b11, 32'shd9998cbe, 
               32'shd98f7fe6, 32'shd9857489, 32'shd97b6aa8, 32'shd9716243, 32'shd9675b5a, 32'shd95d55ef, 32'shd9535201, 32'shd9494f90, 
               32'shd93f4e9e, 32'shd9354f2a, 32'shd92b5135, 32'shd92154bf, 32'shd91759c9, 32'shd90d6053, 32'shd903685d, 32'shd8f971e8, 
               32'shd8ef7cf4, 32'shd8e58982, 32'shd8db9792, 32'shd8d1a724, 32'shd8c7b838, 32'shd8bdcad0, 32'shd8b3deeb, 32'shd8a9f48a, 
               32'shd8a00bae, 32'shd8962456, 32'shd88c3e83, 32'shd8825a35, 32'shd878776d, 32'shd86e962b, 32'shd864b670, 32'shd85ad83c, 
               32'shd850fb8e, 32'shd8472069, 32'shd83d46cc, 32'shd8336eb7, 32'shd829982b, 32'shd81fc328, 32'shd815efae, 32'shd80c1dbf, 
               32'shd8024d59, 32'shd7f87e7f, 32'shd7eeb130, 32'shd7e4e56c, 32'shd7db1b34, 32'shd7d15288, 32'shd7c78b68, 32'shd7bdc5d6, 
               32'shd7b401d1, 32'shd7aa3f5a, 32'shd7a07e70, 32'shd796bf16, 32'shd78d014a, 32'shd783450d, 32'shd7798a60, 32'shd76fd143, 
               32'shd76619b6, 32'shd75c63ba, 32'shd752af4f, 32'shd748fc75, 32'shd73f4b2e, 32'shd7359b78, 32'shd72bed55, 32'shd72240c5, 
               32'shd71895c9, 32'shd70eec60, 32'shd705448b, 32'shd6fb9e4b, 32'shd6f1f99f, 32'shd6e85689, 32'shd6deb508, 32'shd6d5151d, 
               32'shd6cb76c9, 32'shd6c1da0b, 32'shd6b83ee4, 32'shd6aea555, 32'shd6a50d5d, 32'shd69b76fe, 32'shd691e237, 32'shd6884f09, 
               32'shd67ebd74, 32'shd6752d79, 32'shd66b9f18, 32'shd6621251, 32'shd6588725, 32'shd64efd94, 32'shd645759f, 32'shd63bef46, 
               32'shd6326a88, 32'shd628e767, 32'shd61f65e4, 32'shd615e5fd, 32'shd60c67b4, 32'shd602eb0a, 32'shd5f96ffd, 32'shd5eff690, 
               32'shd5e67ec1, 32'shd5dd0892, 32'shd5d39403, 32'shd5ca2115, 32'shd5c0afc6, 32'shd5b74019, 32'shd5add20d, 32'shd5a465a3, 
               32'shd59afadb, 32'shd59191b5, 32'shd5882a32, 32'shd57ec452, 32'shd5756016, 32'shd56bfd7d, 32'shd5629c89, 32'shd5593d3a, 
               32'shd54fdf8f, 32'shd5468389, 32'shd53d292a, 32'shd533d070, 32'shd52a795d, 32'shd52123f0, 32'shd517d02b, 32'shd50e7e0d, 
               32'shd5052d97, 32'shd4fbdec9, 32'shd4f291a4, 32'shd4e94627, 32'shd4dffc54, 32'shd4d6b42b, 32'shd4cd6dab, 32'shd4c428d6, 
               32'shd4bae5ab, 32'shd4b1a42c, 32'shd4a86458, 32'shd49f2630, 32'shd495e9b3, 32'shd48caee4, 32'shd48375c1, 32'shd47a3e4b, 
               32'shd4710883, 32'shd467d469, 32'shd45ea1fd, 32'shd4557140, 32'shd44c4232, 32'shd44314d3, 32'shd439e923, 32'shd430bf24, 
               32'shd42796d5, 32'shd41e7037, 32'shd4154b4a, 32'shd40c280e, 32'shd4030684, 32'shd3f9e6ad, 32'shd3f0c887, 32'shd3e7ac15, 
               32'shd3de9156, 32'shd3d5784a, 32'shd3cc60f2, 32'shd3c34b4f, 32'shd3ba3760, 32'shd3b12526, 32'shd3a814a2, 32'shd39f05d3, 
               32'shd395f8ba, 32'shd38ced57, 32'shd383e3ab, 32'shd37adbb6, 32'shd371d579, 32'shd368d0f3, 32'shd35fce26, 32'shd356cd11, 
               32'shd34dcdb4, 32'shd344d011, 32'shd33bd427, 32'shd332d9f7, 32'shd329e181, 32'shd320eac6, 32'shd317f5c6, 32'shd30f0280, 
               32'shd30610f7, 32'shd2fd2129, 32'shd2f43318, 32'shd2eb46c3, 32'shd2e25c2b, 32'shd2d97350, 32'shd2d08c33, 32'shd2c7a6d4, 
               32'shd2bec333, 32'shd2b5e151, 32'shd2ad012e, 32'shd2a422ca, 32'shd29b4626, 32'shd2926b41, 32'shd289921e, 32'shd280babb, 
               32'shd277e518, 32'shd26f1138, 32'shd2663f19, 32'shd25d6ebc, 32'shd254a021, 32'shd24bd34a, 32'shd2430835, 32'shd23a3ee4, 
               32'shd2317756, 32'shd228b18d, 32'shd21fed88, 32'shd2172b48, 32'shd20e6acc, 32'shd205ac17, 32'shd1fcef27, 32'shd1f433fd, 
               32'shd1eb7a9a, 32'shd1e2c2fd, 32'shd1da0d28, 32'shd1d1591a, 32'shd1c8a6d4, 32'shd1bff656, 32'shd1b747a0, 32'shd1ae9ab4, 
               32'shd1a5ef90, 32'shd19d4636, 32'shd1949ea6, 32'shd18bf8e0, 32'shd18354e4, 32'shd17ab2b3, 32'shd172124d, 32'shd16973b3, 
               32'shd160d6e5, 32'shd1583be2, 32'shd14fa2ad, 32'shd1470b44, 32'shd13e75a8, 32'shd135e1d9, 32'shd12d4fd9, 32'shd124bfa6, 
               32'shd11c3142, 32'shd113a4ad, 32'shd10b19e7, 32'shd10290f0, 32'shd0fa09c9, 32'shd0f18472, 32'shd0e900ec, 32'shd0e07f36, 
               32'shd0d7ff51, 32'shd0cf813e, 32'shd0c704fd, 32'shd0be8a8d, 32'shd0b611f1, 32'shd0ad9b26, 32'shd0a5262f, 32'shd09cb30b, 
               32'shd09441bb, 32'shd08bd23f, 32'shd0836497, 32'shd07af8c4, 32'shd0728ec6, 32'shd06a269d, 32'shd061c04a, 32'shd0595bcd, 
               32'shd050f926, 32'shd0489856, 32'shd040395d, 32'shd037dc3b, 32'shd02f80f1, 32'shd027277e, 32'shd01ecfe4, 32'shd0167a22, 
               32'shd00e2639, 32'shd005d42a, 32'shcffd83f4, 32'shcff53597, 32'shcfece915, 32'shcfe49e6d, 32'shcfdc55a1, 32'shcfd40eaf, 
               32'shcfcbc999, 32'shcfc3865e, 32'shcfbb4500, 32'shcfb3057d, 32'shcfaac7d8, 32'shcfa28c10, 32'shcf9a5225, 32'shcf921a17, 
               32'shcf89e3e8, 32'shcf81af97, 32'shcf797d24, 32'shcf714c91, 32'shcf691ddd, 32'shcf60f108, 32'shcf58c613, 32'shcf509cfe, 
               32'shcf4875ca, 32'shcf405077, 32'shcf382d05, 32'shcf300b74, 32'shcf27ebc5, 32'shcf1fcdf8, 32'shcf17b20d, 32'shcf0f9805, 
               32'shcf077fe1, 32'shceff699f, 32'shcef75541, 32'shceef42c7, 32'shcee73231, 32'shcedf2380, 32'shced716b4, 32'shcecf0bcd, 
               32'shcec702cb, 32'shcebefbb0, 32'shceb6f67a, 32'shceaef32b, 32'shcea6f1c2, 32'shce9ef241, 32'shce96f4a7, 32'shce8ef8f4, 
               32'shce86ff2a, 32'shce7f0748, 32'shce77114e, 32'shce6f1d3d, 32'shce672b16, 32'shce5f3ad8, 32'shce574c84, 32'shce4f6019, 
               32'shce47759a, 32'shce3f8d05, 32'shce37a65b, 32'shce2fc19c, 32'shce27dec9, 32'shce1ffde2, 32'shce181ee8, 32'shce1041d9, 
               32'shce0866b8, 32'shce008d84, 32'shcdf8b63d, 32'shcdf0e0e4, 32'shcde90d79, 32'shcde13bfd, 32'shcdd96c6f, 32'shcdd19ed0, 
               32'shcdc9d320, 32'shcdc20960, 32'shcdba4190, 32'shcdb27bb0, 32'shcdaab7c0, 32'shcda2f5c2, 32'shcd9b35b4, 32'shcd937798, 
               32'shcd8bbb6d, 32'shcd840134, 32'shcd7c48ee, 32'shcd74929a, 32'shcd6cde39, 32'shcd652bcb, 32'shcd5d7b50, 32'shcd55ccca, 
               32'shcd4e2037, 32'shcd467599, 32'shcd3eccef, 32'shcd37263a, 32'shcd2f817b, 32'shcd27deb0, 32'shcd203ddc, 32'shcd189efe, 
               32'shcd110216, 32'shcd096725, 32'shcd01ce2b, 32'shccfa3729, 32'shccf2a21d, 32'shcceb0f0a, 32'shcce37def, 32'shccdbeecc, 
               32'shccd461a2, 32'shccccd671, 32'shccc54d3a, 32'shccbdc5fc, 32'shccb640b8, 32'shccaebd6e, 32'shcca73c1e, 32'shcc9fbcca, 
               32'shcc983f70, 32'shcc90c412, 32'shcc894aaf, 32'shcc81d349, 32'shcc7a5dde, 32'shcc72ea70, 32'shcc6b78ff, 32'shcc64098b, 
               32'shcc5c9c14, 32'shcc55309b, 32'shcc4dc720, 32'shcc465fa3, 32'shcc3efa25, 32'shcc3796a5, 32'shcc303524, 32'shcc28d5a3, 
               32'shcc217822, 32'shcc1a1ca0, 32'shcc12c31f, 32'shcc0b6b9e, 32'shcc04161e, 32'shcbfcc29f, 32'shcbf57121, 32'shcbee21a5, 
               32'shcbe6d42b, 32'shcbdf88b3, 32'shcbd83f3d, 32'shcbd0f7ca, 32'shcbc9b25a, 32'shcbc26eee, 32'shcbbb2d85, 32'shcbb3ee20, 
               32'shcbacb0bf, 32'shcba57563, 32'shcb9e3c0b, 32'shcb9704b9, 32'shcb8fcf6b, 32'shcb889c23, 32'shcb816ae1, 32'shcb7a3ba5, 
               32'shcb730e70, 32'shcb6be341, 32'shcb64ba19, 32'shcb5d92f8, 32'shcb566ddf, 32'shcb4f4acd, 32'shcb4829c4, 32'shcb410ac3, 
               32'shcb39edca, 32'shcb32d2da, 32'shcb2bb9f4, 32'shcb24a316, 32'shcb1d8e43, 32'shcb167b79, 32'shcb0f6aba, 32'shcb085c05, 
               32'shcb014f5b, 32'shcafa44bc, 32'shcaf33c28, 32'shcaec35a0, 32'shcae53123, 32'shcade2eb3, 32'shcad72e4f, 32'shcad02ff8, 
               32'shcac933ae, 32'shcac23971, 32'shcabb4141, 32'shcab44b1f, 32'shcaad570c, 32'shcaa66506, 32'shca9f750f, 32'shca988727, 
               32'shca919b4e, 32'shca8ab184, 32'shca83c9ca, 32'shca7ce420, 32'shca760086, 32'shca6f1efc, 32'shca683f83, 32'shca61621b, 
               32'shca5a86c4, 32'shca53ad7e, 32'shca4cd64b, 32'shca460129, 32'shca3f2e19, 32'shca385d1d, 32'shca318e32, 32'shca2ac15b, 
               32'shca23f698, 32'shca1d2de7, 32'shca16674b, 32'shca0fa2c3, 32'shca08e04f, 32'shca021fef, 32'shc9fb61a5, 32'shc9f4a570, 
               32'shc9edeb50, 32'shc9e73346, 32'shc9e07d51, 32'shc9d9c973, 32'shc9d317ab, 32'shc9cc67fa, 32'shc9c5ba60, 32'shc9bf0edd, 
               32'shc9b86572, 32'shc9b1be1e, 32'shc9ab18e3, 32'shc9a475bf, 32'shc99dd4b4, 32'shc99735c2, 32'shc99098e9, 32'shc989fe29, 
               32'shc9836582, 32'shc97ccef5, 32'shc9763a83, 32'shc96fa82a, 32'shc96917ec, 32'shc96289c9, 32'shc95bfdc1, 32'shc95573d4, 
               32'shc94eec03, 32'shc948664d, 32'shc941e2b4, 32'shc93b6137, 32'shc934e1d6, 32'shc92e6492, 32'shc927e96b, 32'shc9217062, 
               32'shc91af976, 32'shc91484a8, 32'shc90e11f7, 32'shc907a166, 32'shc90132f2, 32'shc8fac69e, 32'shc8f45c68, 32'shc8edf452, 
               32'shc8e78e5b, 32'shc8e12a84, 32'shc8dac8cd, 32'shc8d46936, 32'shc8ce0bc0, 32'shc8c7b06b, 32'shc8c15736, 32'shc8bb0023, 
               32'shc8b4ab32, 32'shc8ae5862, 32'shc8a807b4, 32'shc8a1b928, 32'shc89b6cbf, 32'shc8952278, 32'shc88eda54, 32'shc8889454, 
               32'shc8825077, 32'shc87c0ebd, 32'shc875cf28, 32'shc86f91b7, 32'shc869566a, 32'shc8631d42, 32'shc85ce63e, 32'shc856b160, 
               32'shc8507ea7, 32'shc84a4e14, 32'shc8441fa6, 32'shc83df35f, 32'shc837c93e, 32'shc831a143, 32'shc82b7b70, 32'shc82557c3, 
               32'shc81f363d, 32'shc81916df, 32'shc812f9a9, 32'shc80cde9b, 32'shc806c5b5, 32'shc800aef7, 32'shc7fa9a62, 32'shc7f487f6, 
               32'shc7ee77b3, 32'shc7e8699a, 32'shc7e25daa, 32'shc7dc53e3, 32'shc7d64c47, 32'shc7d046d6, 32'shc7ca438f, 32'shc7c44272, 
               32'shc7be4381, 32'shc7b846ba, 32'shc7b24c20, 32'shc7ac53b1, 32'shc7a65d6e, 32'shc7a06957, 32'shc79a776c, 32'shc79487ae, 
               32'shc78e9a1d, 32'shc788aeb9, 32'shc782c582, 32'shc77cde79, 32'shc776f99d, 32'shc77116f0, 32'shc76b3671, 32'shc7655820, 
               32'shc75f7bfe, 32'shc759a20a, 32'shc753ca46, 32'shc74df4b1, 32'shc748214c, 32'shc7425016, 32'shc73c8111, 32'shc736b43c, 
               32'shc730e997, 32'shc72b2123, 32'shc7255ae0, 32'shc71f96ce, 32'shc719d4ed, 32'shc714153e, 32'shc70e57c0, 32'shc7089c75, 
               32'shc702e35c, 32'shc6fd2c75, 32'shc6f777c1, 32'shc6f1c540, 32'shc6ec14f2, 32'shc6e666d7, 32'shc6e0baf0, 32'shc6db113d, 
               32'shc6d569be, 32'shc6cfc472, 32'shc6ca215c, 32'shc6c4807a, 32'shc6bee1cd, 32'shc6b94554, 32'shc6b3ab12, 32'shc6ae1304, 
               32'shc6a87d2d, 32'shc6a2e98b, 32'shc69d5820, 32'shc697c8eb, 32'shc6923bec, 32'shc68cb124, 32'shc6872894, 32'shc681a23a, 
               32'shc67c1e18, 32'shc6769c2e, 32'shc6711c7b, 32'shc66b9f01, 32'shc66623be, 32'shc660aab5, 32'shc65b33e4, 32'shc655bf4c, 
               32'shc6504ced, 32'shc64adcc7, 32'shc6456edb, 32'shc6400329, 32'shc63a99b1, 32'shc6353273, 32'shc62fcd6f, 32'shc62a6aa6, 
               32'shc6250a18, 32'shc61fabc4, 32'shc61a4fac, 32'shc614f5cf, 32'shc60f9e2e, 32'shc60a48c9, 32'shc604f5a0, 32'shc5ffa4b3, 
               32'shc5fa5603, 32'shc5f5098f, 32'shc5efbf58, 32'shc5ea775e, 32'shc5e531a1, 32'shc5dfee22, 32'shc5daace1, 32'shc5d56ddd, 
               32'shc5d03118, 32'shc5caf690, 32'shc5c5be47, 32'shc5c0883d, 32'shc5bb5472, 32'shc5b622e6, 32'shc5b0f399, 32'shc5abc68c, 
               32'shc5a69bbe, 32'shc5a17330, 32'shc59c4ce3, 32'shc59728d5, 32'shc5920708, 32'shc58ce77c, 32'shc587ca31, 32'shc582af26, 
               32'shc57d965d, 32'shc5787fd6, 32'shc5736b90, 32'shc56e598c, 32'shc56949ca, 32'shc5643c4a, 32'shc55f310d, 32'shc55a2812, 
               32'shc555215a, 32'shc5501ce5, 32'shc54b1ab4, 32'shc5461ac6, 32'shc5411d1b, 32'shc53c21b4, 32'shc5372891, 32'shc53231b3, 
               32'shc52d3d18, 32'shc5284ac3, 32'shc5235ab2, 32'shc51e6ce6, 32'shc519815f, 32'shc514981d, 32'shc50fb121, 32'shc50acc6b, 
               32'shc505e9fb, 32'shc50109d0, 32'shc4fc2bec, 32'shc4f7504e, 32'shc4f276f7, 32'shc4ed9fe7, 32'shc4e8cb1e, 32'shc4e3f89c, 
               32'shc4df2862, 32'shc4da5a6f, 32'shc4d58ec3, 32'shc4d0c560, 32'shc4cbfe45, 32'shc4c73972, 32'shc4c276e8, 32'shc4bdb6a6, 
               32'shc4b8f8ad, 32'shc4b43cfd, 32'shc4af8397, 32'shc4aacc7a, 32'shc4a617a6, 32'shc4a1651c, 32'shc49cb4dd, 32'shc49806e7, 
               32'shc4935b3c, 32'shc48eb1db, 32'shc48a0ac4, 32'shc48565f9, 32'shc480c379, 32'shc47c2344, 32'shc477855a, 32'shc472e9bc, 
               32'shc46e5069, 32'shc469b963, 32'shc46524a9, 32'shc460923b, 32'shc45c0219, 32'shc4577444, 32'shc452e8bc, 32'shc44e5f80, 
               32'shc449d892, 32'shc44553f2, 32'shc440d19e, 32'shc43c5199, 32'shc437d3e1, 32'shc4335877, 32'shc42edf5c, 32'shc42a688f, 
               32'shc425f410, 32'shc42181e0, 32'shc41d11ff, 32'shc418a46d, 32'shc414392b, 32'shc40fd037, 32'shc40b6994, 32'shc4070540, 
               32'shc402a33c, 32'shc3fe4388, 32'shc3f9e624, 32'shc3f58b10, 32'shc3f1324e, 32'shc3ecdbdc, 32'shc3e887bb, 32'shc3e435ea, 
               32'shc3dfe66c, 32'shc3db993e, 32'shc3d74e62, 32'shc3d305d8, 32'shc3cebfa0, 32'shc3ca7bba, 32'shc3c63a26, 32'shc3c1fae5, 
               32'shc3bdbdf6, 32'shc3b9835a, 32'shc3b54b11, 32'shc3b1151b, 32'shc3ace178, 32'shc3a8b028, 32'shc3a4812c, 32'shc3a05484, 
               32'shc39c2a2f, 32'shc398022f, 32'shc393dc82, 32'shc38fb92a, 32'shc38b9827, 32'shc3877978, 32'shc3835d1e, 32'shc37f4319, 
               32'shc37b2b6a, 32'shc377160f, 32'shc373030a, 32'shc36ef25b, 32'shc36ae401, 32'shc366d7fd, 32'shc362ce50, 32'shc35ec6f8, 
               32'shc35ac1f7, 32'shc356bf4d, 32'shc352bef9, 32'shc34ec0fc, 32'shc34ac556, 32'shc346cc07, 32'shc342d510, 32'shc33ee070, 
               32'shc33aee27, 32'shc336fe37, 32'shc333109e, 32'shc32f255e, 32'shc32b3c75, 32'shc32755e5, 32'shc32371ae, 32'shc31f8fcf, 
               32'shc31bb049, 32'shc317d31c, 32'shc313f848, 32'shc3101fce, 32'shc30c49ad, 32'shc30875e5, 32'shc304a477, 32'shc300d563, 
               32'shc2fd08a9, 32'shc2f93e4a, 32'shc2f57644, 32'shc2f1b099, 32'shc2eded49, 32'shc2ea2c53, 32'shc2e66db8, 32'shc2e2b178, 
               32'shc2def794, 32'shc2db400a, 32'shc2d78add, 32'shc2d3d80a, 32'shc2d02794, 32'shc2cc7979, 32'shc2c8cdbb, 32'shc2c52459, 
               32'shc2c17d52, 32'shc2bdd8a9, 32'shc2ba365c, 32'shc2b6966c, 32'shc2b2f8d8, 32'shc2af5da2, 32'shc2abc4c9, 32'shc2a82e4d, 
               32'shc2a49a2e, 32'shc2a1086d, 32'shc29d790a, 32'shc299ec05, 32'shc296615d, 32'shc292d914, 32'shc28f5329, 32'shc28bcf9c, 
               32'shc2884e6e, 32'shc284cf9f, 32'shc281532e, 32'shc27dd91c, 32'shc27a616a, 32'shc276ec16, 32'shc2737922, 32'shc270088e, 
               32'shc26c9a58, 32'shc2692e83, 32'shc265c50e, 32'shc2625df8, 32'shc25ef943, 32'shc25b96ee, 32'shc25836f9, 32'shc254d965, 
               32'shc2517e31, 32'shc24e255e, 32'shc24aceed, 32'shc2477adc, 32'shc244292c, 32'shc240d9de, 32'shc23d8cf1, 32'shc23a4265, 
               32'shc236fa3b, 32'shc233b473, 32'shc230710d, 32'shc22d3009, 32'shc229f167, 32'shc226b528, 32'shc2237b4b, 32'shc22043d0, 
               32'shc21d0eb8, 32'shc219dc03, 32'shc216abb1, 32'shc2137dc2, 32'shc2105236, 32'shc20d290d, 32'shc20a0248, 32'shc206dde6, 
               32'shc203bbe8, 32'shc2009c4e, 32'shc1fd7f17, 32'shc1fa6445, 32'shc1f74bd6, 32'shc1f435cc, 32'shc1f12227, 32'shc1ee10e5, 
               32'shc1eb0209, 32'shc1e7f591, 32'shc1e4eb7e, 32'shc1e1e3d0, 32'shc1dede87, 32'shc1dbdba3, 32'shc1d8db25, 32'shc1d5dd0c, 
               32'shc1d2e158, 32'shc1cfe80a, 32'shc1ccf122, 32'shc1c9fca0, 32'shc1c70a84, 32'shc1c41ace, 32'shc1c12d7e, 32'shc1be4294, 
               32'shc1bb5a11, 32'shc1b873f5, 32'shc1b5903f, 32'shc1b2aef0, 32'shc1afd007, 32'shc1acf386, 32'shc1aa196c, 32'shc1a741b9, 
               32'shc1a46c6e, 32'shc1a1998a, 32'shc19ec90d, 32'shc19bfaf9, 32'shc1992f4c, 32'shc1966606, 32'shc1939f29, 32'shc190dab4, 
               32'shc18e18a7, 32'shc18b5903, 32'shc1889bc6, 32'shc185e0f3, 32'shc1832888, 32'shc1807285, 32'shc17dbeec, 32'shc17b0dbb, 
               32'shc1785ef4, 32'shc175b296, 32'shc17308a1, 32'shc1706115, 32'shc16dbbf3, 32'shc16b193a, 32'shc16878eb, 32'shc165db05, 
               32'shc1633f8a, 32'shc160a678, 32'shc15e0fd1, 32'shc15b7b94, 32'shc158e9c1, 32'shc1565a58, 32'shc153cd5a, 32'shc15142c6, 
               32'shc14eba9d, 32'shc14c34df, 32'shc149b18b, 32'shc14730a3, 32'shc144b225, 32'shc1423613, 32'shc13fbc6c, 32'shc13d4530, 
               32'shc13ad060, 32'shc1385dfb, 32'shc135ee02, 32'shc1338075, 32'shc1311553, 32'shc12eac9d, 32'shc12c4653, 32'shc129e276, 
               32'shc1278104, 32'shc12521ff, 32'shc122c566, 32'shc1206b39, 32'shc11e1379, 32'shc11bbe26, 32'shc1196b3f, 32'shc1171ac6, 
               32'shc114ccb9, 32'shc1128119, 32'shc11037e6, 32'shc10df120, 32'shc10bacc8, 32'shc1096add, 32'shc1072b5f, 32'shc104ee4f, 
               32'shc102b3ac, 32'shc1007b77, 32'shc0fe45b0, 32'shc0fc1257, 32'shc0f9e16b, 32'shc0f7b2ee, 32'shc0f586df, 32'shc0f35d3e, 
               32'shc0f1360b, 32'shc0ef1147, 32'shc0eceef1, 32'shc0eacf09, 32'shc0e8b190, 32'shc0e69686, 32'shc0e47deb, 32'shc0e267be, 
               32'shc0e05401, 32'shc0de42b2, 32'shc0dc33d2, 32'shc0da2762, 32'shc0d81d61, 32'shc0d615cf, 32'shc0d410ad, 32'shc0d20dfa, 
               32'shc0d00db6, 32'shc0ce0fe3, 32'shc0cc147f, 32'shc0ca1b8a, 32'shc0c82506, 32'shc0c630f2, 32'shc0c43f4d, 32'shc0c25019, 
               32'shc0c06355, 32'shc0be7901, 32'shc0bc911d, 32'shc0baabaa, 32'shc0b8c8a7, 32'shc0b6e815, 32'shc0b509f3, 32'shc0b32e42, 
               32'shc0b15502, 32'shc0af7e33, 32'shc0ada9d4, 32'shc0abd7e6, 32'shc0aa086a, 32'shc0a83b5e, 32'shc0a670c4, 32'shc0a4a89b, 
               32'shc0a2e2e3, 32'shc0a11f9d, 32'shc09f5ec8, 32'shc09da065, 32'shc09be473, 32'shc09a2af3, 32'shc09873e4, 32'shc096bf48, 
               32'shc0950d1d, 32'shc0935d64, 32'shc091b01d, 32'shc0900548, 32'shc08e5ce5, 32'shc08cb6f5, 32'shc08b1376, 32'shc089726a, 
               32'shc087d3d0, 32'shc08637a9, 32'shc0849df4, 32'shc08306b2, 32'shc08171e2, 32'shc07fdf85, 32'shc07e4f9b, 32'shc07cc223, 
               32'shc07b371e, 32'shc079ae8c, 32'shc078286e, 32'shc076a4c2, 32'shc0752389, 32'shc073a4c3, 32'shc0722871, 32'shc070ae92, 
               32'shc06f3726, 32'shc06dc22e, 32'shc06c4fa8, 32'shc06adf97, 32'shc06971f9, 32'shc06806ce, 32'shc0669e18, 32'shc06537d4, 
               32'shc063d405, 32'shc06272aa, 32'shc06113c2, 32'shc05fb74e, 32'shc05e5d4e, 32'shc05d05c3, 32'shc05bb0ab, 32'shc05a5e07, 
               32'shc0590dd8, 32'shc057c01d, 32'shc05674d6, 32'shc0552c03, 32'shc053e5a5, 32'shc052a1bb, 32'shc0516045, 32'shc0502145, 
               32'shc04ee4b8, 32'shc04daaa1, 32'shc04c72fe, 32'shc04b3dcf, 32'shc04a0b16, 32'shc048dad1, 32'shc047ad01, 32'shc04681a6, 
               32'shc04558c0, 32'shc044324f, 32'shc0430e53, 32'shc041eccc, 32'shc040cdba, 32'shc03fb11d, 32'shc03e96f6, 32'shc03d7f44, 
               32'shc03c6a07, 32'shc03b573f, 32'shc03a46ed, 32'shc0393910, 32'shc0382da8, 32'shc03724b6, 32'shc0361e3a, 32'shc0351a33, 
               32'shc03418a2, 32'shc0331986, 32'shc0321ce0, 32'shc03122b0, 32'shc0302af5, 32'shc02f35b1, 32'shc02e42e2, 32'shc02d5289, 
               32'shc02c64a6, 32'shc02b7939, 32'shc02a9042, 32'shc029a9c1, 32'shc028c5b6, 32'shc027e421, 32'shc0270502, 32'shc0262859, 
               32'shc0254e27, 32'shc024766a, 32'shc023a124, 32'shc022ce54, 32'shc021fdfb, 32'shc0213018, 32'shc02064ab, 32'shc01f9bb5, 
               32'shc01ed535, 32'shc01e112b, 32'shc01d4f99, 32'shc01c907c, 32'shc01bd3d6, 32'shc01b19a7, 32'shc01a61ee, 32'shc019acac, 
               32'shc018f9e1, 32'shc018498c, 32'shc0179bae, 32'shc016f047, 32'shc0164757, 32'shc015a0dd, 32'shc014fcda, 32'shc0145b4e, 
               32'shc013bc39, 32'shc0131f9b, 32'shc0128574, 32'shc011edc3, 32'shc011588a, 32'shc010c5c7, 32'shc010357c, 32'shc00fa7a8, 
               32'shc00f1c4a, 32'shc00e9364, 32'shc00e0cf5, 32'shc00d88fd, 32'shc00d077c, 32'shc00c8872, 32'shc00c0be0, 32'shc00b91c4, 
               32'shc00b1a20, 32'shc00aa4f3, 32'shc00a323d, 32'shc009c1ff, 32'shc0095438, 32'shc008e8e8, 32'shc008800f, 32'shc00819ae, 
               32'shc007b5c4, 32'shc0075452, 32'shc006f556, 32'shc00698d3, 32'shc0063ec6, 32'shc005e731, 32'shc0059214, 32'shc0053f6e, 
               32'shc004ef3f, 32'shc004a188, 32'shc0045648, 32'shc0040d80, 32'shc003c72f, 32'shc0038356, 32'shc00341f4, 32'shc003030a, 
               32'shc002c697, 32'shc0028c9c, 32'shc0025519, 32'shc002200d, 32'shc001ed78, 32'shc001bd5c, 32'shc0018fb6, 32'shc0016489, 
               32'shc0013bd3, 32'shc0011594, 32'shc000f1ce, 32'shc000d07e, 32'shc000b1a7, 32'shc0009547, 32'shc0007b5f, 32'shc00063ee, 
               32'shc0004ef5, 32'shc0003c74, 32'shc0002c6a, 32'shc0001ed8, 32'shc00013bd, 32'shc0000b1a, 32'shc00004ef, 32'shc000013c
            };

            reg signed [31:0] W_Im_table[4096] = '{
               32'sh00000000, 32'shfff36f02, 32'shffe6de05, 32'shffda4d09, 32'shffcdbc0f, 32'shffc12b16, 32'shffb49a1f, 32'shffa8092c, 
               32'shff9b783c, 32'shff8ee750, 32'shff825668, 32'shff75c585, 32'shff6934a8, 32'shff5ca3d0, 32'shff5012fe, 32'shff438234, 
               32'shff36f170, 32'shff2a60b4, 32'shff1dd001, 32'shff113f56, 32'shff04aeb5, 32'shfef81e1d, 32'shfeeb8d8f, 32'shfedefd0c, 
               32'shfed26c94, 32'shfec5dc28, 32'shfeb94bc8, 32'shfeacbb74, 32'shfea02b2e, 32'shfe939af5, 32'shfe870aca, 32'shfe7a7aae, 
               32'shfe6deaa1, 32'shfe615aa3, 32'shfe54cab5, 32'shfe483ad8, 32'shfe3bab0b, 32'shfe2f1b50, 32'shfe228ba7, 32'shfe15fc11, 
               32'shfe096c8d, 32'shfdfcdd1d, 32'shfdf04dc0, 32'shfde3be78, 32'shfdd72f45, 32'shfdcaa027, 32'shfdbe111e, 32'shfdb1822c, 
               32'shfda4f351, 32'shfd98648d, 32'shfd8bd5e1, 32'shfd7f474d, 32'shfd72b8d2, 32'shfd662a70, 32'shfd599c28, 32'shfd4d0df9, 
               32'shfd407fe6, 32'shfd33f1ed, 32'shfd276410, 32'shfd1ad650, 32'shfd0e48ab, 32'shfd01bb24, 32'shfcf52dbb, 32'shfce8a06f, 
               32'shfcdc1342, 32'shfccf8634, 32'shfcc2f945, 32'shfcb66c77, 32'shfca9dfc8, 32'shfc9d533b, 32'shfc90c6cf, 32'shfc843a85, 
               32'shfc77ae5e, 32'shfc6b2259, 32'shfc5e9678, 32'shfc520aba, 32'shfc457f21, 32'shfc38f3ac, 32'shfc2c685d, 32'shfc1fdd34, 
               32'shfc135231, 32'shfc06c754, 32'shfbfa3c9f, 32'shfbedb212, 32'shfbe127ac, 32'shfbd49d70, 32'shfbc8135c, 32'shfbbb8973, 
               32'shfbaeffb3, 32'shfba2761e, 32'shfb95ecb4, 32'shfb896375, 32'shfb7cda63, 32'shfb70517d, 32'shfb63c8c4, 32'shfb574039, 
               32'shfb4ab7db, 32'shfb3e2fac, 32'shfb31a7ac, 32'shfb251fdc, 32'shfb18983b, 32'shfb0c10cb, 32'shfaff898c, 32'shfaf3027e, 
               32'shfae67ba2, 32'shfad9f4f8, 32'shfacd6e81, 32'shfac0e83d, 32'shfab4622d, 32'shfaa7dc52, 32'shfa9b56ab, 32'shfa8ed139, 
               32'shfa824bfd, 32'shfa75c6f8, 32'shfa694229, 32'shfa5cbd91, 32'shfa503930, 32'shfa43b508, 32'shfa373119, 32'shfa2aad62, 
               32'shfa1e29e5, 32'shfa11a6a3, 32'shfa05239a, 32'shf9f8a0cd, 32'shf9ec1e3b, 32'shf9df9be6, 32'shf9d319cc, 32'shf9c697f0, 
               32'shf9ba1651, 32'shf9ad94f0, 32'shf9a113cd, 32'shf99492ea, 32'shf9881245, 32'shf97b91e1, 32'shf96f11bc, 32'shf96291d9, 
               32'shf9561237, 32'shf94992d7, 32'shf93d13b8, 32'shf93094dd, 32'shf9241645, 32'shf91797f0, 32'shf90b19e0, 32'shf8fe9c15, 
               32'shf8f21e8e, 32'shf8e5a14d, 32'shf8d92452, 32'shf8cca79e, 32'shf8c02b31, 32'shf8b3af0c, 32'shf8a7332e, 32'shf89ab799, 
               32'shf88e3c4d, 32'shf881c14b, 32'shf8754692, 32'shf868cc24, 32'shf85c5201, 32'shf84fd829, 32'shf8435e9d, 32'shf836e55d, 
               32'shf82a6c6a, 32'shf81df3c5, 32'shf8117b6d, 32'shf8050364, 32'shf7f88ba9, 32'shf7ec143e, 32'shf7df9d22, 32'shf7d32657, 
               32'shf7c6afdc, 32'shf7ba39b3, 32'shf7adc3db, 32'shf7a14e55, 32'shf794d922, 32'shf7886442, 32'shf77befb5, 32'shf76f7b7d, 
               32'shf7630799, 32'shf756940a, 32'shf74a20d0, 32'shf73daded, 32'shf7313b60, 32'shf724c92a, 32'shf718574b, 32'shf70be5c4, 
               32'shf6ff7496, 32'shf6f303c0, 32'shf6e69344, 32'shf6da2321, 32'shf6cdb359, 32'shf6c143ec, 32'shf6b4d4d9, 32'shf6a86623, 
               32'shf69bf7c9, 32'shf68f89cb, 32'shf6831c2b, 32'shf676aee8, 32'shf66a4203, 32'shf65dd57d, 32'shf6516956, 32'shf644fd8f, 
               32'shf6389228, 32'shf62c2721, 32'shf61fbc7b, 32'shf6135237, 32'shf606e854, 32'shf5fa7ed4, 32'shf5ee15b7, 32'shf5e1acfd, 
               32'shf5d544a7, 32'shf5c8dcb6, 32'shf5bc7529, 32'shf5b00e02, 32'shf5a3a740, 32'shf59740e5, 32'shf58adaf0, 32'shf57e7563, 
               32'shf572103d, 32'shf565ab80, 32'shf559472b, 32'shf54ce33f, 32'shf5407fbd, 32'shf5341ca5, 32'shf527b9f7, 32'shf51b57b5, 
               32'shf50ef5de, 32'shf5029473, 32'shf4f63374, 32'shf4e9d2e3, 32'shf4dd72be, 32'shf4d11308, 32'shf4c4b3c0, 32'shf4b854e7, 
               32'shf4abf67e, 32'shf49f9884, 32'shf4933afa, 32'shf486dde1, 32'shf47a8139, 32'shf46e2504, 32'shf461c940, 32'shf4556def, 
               32'shf4491311, 32'shf43cb8a7, 32'shf4305eb0, 32'shf424052f, 32'shf417ac22, 32'shf40b538b, 32'shf3fefb6a, 32'shf3f2a3bf, 
               32'shf3e64c8c, 32'shf3d9f5cf, 32'shf3cd9f8b, 32'shf3c149bf, 32'shf3b4f46c, 32'shf3a89f92, 32'shf39c4b32, 32'shf38ff74d, 
               32'shf383a3e2, 32'shf37750f2, 32'shf36afe7e, 32'shf35eac86, 32'shf3525b0b, 32'shf3460a0d, 32'shf339b98d, 32'shf32d698a, 
               32'shf3211a07, 32'shf314cb02, 32'shf3087c7d, 32'shf2fc2e77, 32'shf2efe0f2, 32'shf2e393ef, 32'shf2d7476c, 32'shf2cafb6b, 
               32'shf2beafed, 32'shf2b264f2, 32'shf2a61a7a, 32'shf299d085, 32'shf28d8715, 32'shf2813e2a, 32'shf274f5c3, 32'shf268ade3, 
               32'shf25c6688, 32'shf2501fb5, 32'shf243d968, 32'shf23793a3, 32'shf22b4e66, 32'shf21f09b1, 32'shf212c585, 32'shf20681e3, 
               32'shf1fa3ecb, 32'shf1edfc3d, 32'shf1e1ba3a, 32'shf1d578c2, 32'shf1c937d6, 32'shf1bcf777, 32'shf1b0b7a4, 32'shf1a4785e, 
               32'shf19839a6, 32'shf18bfb7d, 32'shf17fbde2, 32'shf17380d6, 32'shf1674459, 32'shf15b086d, 32'shf14ecd11, 32'shf1429247, 
               32'shf136580d, 32'shf12a1e66, 32'shf11de551, 32'shf111accf, 32'shf10574e0, 32'shf0f93d86, 32'shf0ed06bf, 32'shf0e0d08d, 
               32'shf0d49af1, 32'shf0c865ea, 32'shf0bc317a, 32'shf0affda0, 32'shf0a3ca5d, 32'shf09797b2, 32'shf08b659f, 32'shf07f3424, 
               32'shf0730342, 32'shf066d2fa, 32'shf05aa34c, 32'shf04e7438, 32'shf04245c0, 32'shf03617e2, 32'shf029eaa1, 32'shf01dbdfb, 
               32'shf01191f3, 32'shf0056687, 32'sheff93bba, 32'shefed118a, 32'shefe0e7f9, 32'shefd4bf08, 32'shefc896b5, 32'shefbc6f03, 
               32'shefb047f2, 32'shefa42181, 32'shef97fbb2, 32'shef8bd685, 32'shef7fb1fa, 32'shef738e12, 32'shef676ace, 32'shef5b482d, 
               32'shef4f2630, 32'shef4304d8, 32'shef36e426, 32'shef2ac419, 32'shef1ea4b2, 32'shef1285f2, 32'shef0667d9, 32'sheefa4a67, 
               32'sheeee2d9d, 32'sheee2117c, 32'sheed5f604, 32'sheec9db35, 32'sheebdc110, 32'sheeb1a796, 32'sheea58ec6, 32'shee9976a1, 
               32'shee8d5f29, 32'shee81485c, 32'shee75323c, 32'shee691cc9, 32'shee5d0804, 32'shee50f3ed, 32'shee44e084, 32'shee38cdcb, 
               32'shee2cbbc1, 32'shee20aa67, 32'shee1499bd, 32'shee0889c4, 32'shedfc7a7c, 32'shedf06be6, 32'shede45e03, 32'shedd850d2, 
               32'shedcc4454, 32'shedc0388a, 32'shedb42d74, 32'sheda82313, 32'shed9c1967, 32'shed901070, 32'shed84082f, 32'shed7800a5, 
               32'shed6bf9d1, 32'shed5ff3b5, 32'shed53ee51, 32'shed47e9a5, 32'shed3be5b1, 32'shed2fe277, 32'shed23dff7, 32'shed17de31, 
               32'shed0bdd25, 32'shecffdcd4, 32'shecf3dd3f, 32'shece7de66, 32'shecdbe04a, 32'sheccfe2ea, 32'shecc3e648, 32'shecb7ea63, 
               32'shecabef3d, 32'shec9ff4d6, 32'shec93fb2e, 32'shec880245, 32'shec7c0a1d, 32'shec7012b5, 32'shec641c0e, 32'shec582629, 
               32'shec4c3106, 32'shec403ca5, 32'shec344908, 32'shec28562d, 32'shec1c6417, 32'shec1072c4, 32'shec048237, 32'shebf8926f, 
               32'shebeca36c, 32'shebe0b52f, 32'shebd4c7ba, 32'shebc8db0b, 32'shebbcef23, 32'shebb10404, 32'sheba519ad, 32'sheb99301f, 
               32'sheb8d475b, 32'sheb815f60, 32'sheb75782f, 32'sheb6991ca, 32'sheb5dac2f, 32'sheb51c760, 32'sheb45e35d, 32'sheb3a0027, 
               32'sheb2e1dbe, 32'sheb223c22, 32'sheb165b54, 32'sheb0a7b54, 32'sheafe9c24, 32'sheaf2bdc3, 32'sheae6e031, 32'sheadb0370, 
               32'sheacf277f, 32'sheac34c60, 32'sheab77212, 32'sheaab9896, 32'shea9fbfed, 32'shea93e817, 32'shea881114, 32'shea7c3ae5, 
               32'shea70658a, 32'shea649105, 32'shea58bd54, 32'shea4cea79, 32'shea411874, 32'shea354746, 32'shea2976ef, 32'shea1da770, 
               32'shea11d8c8, 32'shea060af9, 32'she9fa3e03, 32'she9ee71e6, 32'she9e2a6a3, 32'she9d6dc3b, 32'she9cb12ad, 32'she9bf49fa, 
               32'she9b38223, 32'she9a7bb28, 32'she99bf509, 32'she9902fc7, 32'she9846b63, 32'she978a7dd, 32'she96ce535, 32'she961236c, 
               32'she9556282, 32'she949a278, 32'she93de34e, 32'she9322505, 32'she926679c, 32'she91aab16, 32'she90eef71, 32'she90334af, 
               32'she8f77acf, 32'she8ebc1d3, 32'she8e009ba, 32'she8d45286, 32'she8c89c37, 32'she8bce6cd, 32'she8b13248, 32'she8a57ea9, 
               32'she899cbf1, 32'she88e1a20, 32'she8826936, 32'she876b934, 32'she86b0a1a, 32'she85f5be9, 32'she853aea1, 32'she8480243, 
               32'she83c56cf, 32'she830ac45, 32'she82502a7, 32'she81959f4, 32'she80db22d, 32'she8020b52, 32'she7f66564, 32'she7eac063, 
               32'she7df1c50, 32'she7d3792b, 32'she7c7d6f4, 32'she7bc35ad, 32'she7b09555, 32'she7a4f5ed, 32'she7995776, 32'she78db9ef, 
               32'she7821d59, 32'she77681b6, 32'she76ae704, 32'she75f4d45, 32'she753b479, 32'she7481ca1, 32'she73c85bc, 32'she730efcc, 
               32'she7255ad1, 32'she719c6cb, 32'she70e33bb, 32'she702a1a1, 32'she6f7107e, 32'she6eb8052, 32'she6dff11d, 32'she6d462e1, 
               32'she6c8d59c, 32'she6bd4951, 32'she6b1bdff, 32'she6a633a6, 32'she69aaa48, 32'she68f21e5, 32'she6839a7c, 32'she6781410, 
               32'she66c8e9f, 32'she6610a2a, 32'she65586b3, 32'she64a0438, 32'she63e82bc, 32'she633023e, 32'she62782be, 32'she61c043d, 
               32'she61086bc, 32'she6050a3b, 32'she5f98ebb, 32'she5ee143b, 32'she5e29abc, 32'she5d72240, 32'she5cbaac5, 32'she5c0344d, 
               32'she5b4bed8, 32'she5a94a67, 32'she59dd6f9, 32'she5926490, 32'she586f32c, 32'she57b82cd, 32'she5701374, 32'she564a521, 
               32'she55937d5, 32'she54dcb8f, 32'she5426051, 32'she536f61b, 32'she52b8cee, 32'she52024c9, 32'she514bdad, 32'she509579b, 
               32'she4fdf294, 32'she4f28e96, 32'she4e72ba4, 32'she4dbc9bd, 32'she4d068e2, 32'she4c50914, 32'she4b9aa52, 32'she4ae4c9d, 
               32'she4a2eff6, 32'she497945d, 32'she48c39d3, 32'she480e057, 32'she47587eb, 32'she46a308f, 32'she45eda43, 32'she4538507, 
               32'she44830dd, 32'she43cddc4, 32'she4318bbe, 32'she4263ac9, 32'she41aeae8, 32'she40f9c1a, 32'she4044e60, 32'she3f901ba, 
               32'she3edb628, 32'she3e26bac, 32'she3d72245, 32'she3cbd9f4, 32'she3c092b9, 32'she3b54c95, 32'she3aa0788, 32'she39ec393, 
               32'she39380b6, 32'she3883ef2, 32'she37cfe47, 32'she371beb5, 32'she366803c, 32'she35b42df, 32'she350069b, 32'she344cb73, 
               32'she3399167, 32'she32e5876, 32'she32320a2, 32'she317e9eb, 32'she30cb451, 32'she3017fd5, 32'she2f64c77, 32'she2eb1a37, 
               32'she2dfe917, 32'she2d4b916, 32'she2c98a35, 32'she2be5c74, 32'she2b32fd4, 32'she2a80456, 32'she29cd9f8, 32'she291b0bd, 
               32'she28688a4, 32'she27b61af, 32'she2703bdc, 32'she265172e, 32'she259f3a3, 32'she24ed13d, 32'she243affc, 32'she2388fe1, 
               32'she22d70eb, 32'she222531c, 32'she2173674, 32'she20c1af3, 32'she2010099, 32'she1f5e768, 32'she1eacf5f, 32'she1dfb87f, 
               32'she1d4a2c8, 32'she1c98e3b, 32'she1be7ad8, 32'she1b368a0, 32'she1a85793, 32'she19d47b1, 32'she19238fb, 32'she1872b72, 
               32'she17c1f15, 32'she17113e5, 32'she16609e3, 32'she15b0110, 32'she14ff96a, 32'she144f2f3, 32'she139edac, 32'she12ee995, 
               32'she123e6ad, 32'she118e4f6, 32'she10de470, 32'she102e51c, 32'she0f7e6f9, 32'she0ecea09, 32'she0e1ee4b, 32'she0d6f3c1, 
               32'she0cbfa6a, 32'she0c10247, 32'she0b60b58, 32'she0ab159e, 32'she0a0211a, 32'she0952dcb, 32'she08a3bb2, 32'she07f4acf, 
               32'she0745b24, 32'she0696cb0, 32'she05e7f74, 32'she053936f, 32'she048a8a4, 32'she03dbf11, 32'she032d6b8, 32'she027ef99, 
               32'she01d09b4, 32'she012250a, 32'she007419b, 32'shdffc5f67, 32'shdff17e70, 32'shdfe69eb4, 32'shdfdbc036, 32'shdfd0e2f5, 
               32'shdfc606f1, 32'shdfbb2c2c, 32'shdfb052a5, 32'shdfa57a5d, 32'shdf9aa354, 32'shdf8fcd8b, 32'shdf84f902, 32'shdf7a25ba, 
               32'shdf6f53b3, 32'shdf6482ed, 32'shdf59b369, 32'shdf4ee527, 32'shdf441828, 32'shdf394c6b, 32'shdf2e81f3, 32'shdf23b8be, 
               32'shdf18f0ce, 32'shdf0e2a22, 32'shdf0364bc, 32'shdef8a09b, 32'shdeedddc0, 32'shdee31c2b, 32'shded85bdd, 32'shdecd9cd7, 
               32'shdec2df18, 32'shdeb822a1, 32'shdead6773, 32'shdea2ad8d, 32'shde97f4f1, 32'shde8d3d9e, 32'shde828796, 32'shde77d2d8, 
               32'shde6d1f65, 32'shde626d3e, 32'shde57bc62, 32'shde4d0cd2, 32'shde425e8f, 32'shde37b199, 32'shde2d05f1, 32'shde225b96, 
               32'shde17b28a, 32'shde0d0acc, 32'shde02645d, 32'shddf7bf3e, 32'shdded1b6e, 32'shdde278ef, 32'shddd7d7c1, 32'shddcd37e4, 
               32'shddc29958, 32'shddb7fc1e, 32'shddad6036, 32'shdda2c5a2, 32'shdd982c60, 32'shdd8d9472, 32'shdd82fdd8, 32'shdd786892, 
               32'shdd6dd4a2, 32'shdd634206, 32'shdd58b0c0, 32'shdd4e20d0, 32'shdd439236, 32'shdd3904f4, 32'shdd2e7908, 32'shdd23ee74, 
               32'shdd196538, 32'shdd0edd55, 32'shdd0456ca, 32'shdcf9d199, 32'shdcef4dc2, 32'shdce4cb44, 32'shdcda4a21, 32'shdccfca59, 
               32'shdcc54bec, 32'shdcbacedb, 32'shdcb05326, 32'shdca5d8cd, 32'shdc9b5fd2, 32'shdc90e834, 32'shdc8671f3, 32'shdc7bfd11, 
               32'shdc71898d, 32'shdc671768, 32'shdc5ca6a2, 32'shdc52373c, 32'shdc47c936, 32'shdc3d5c91, 32'shdc32f14d, 32'shdc28876a, 
               32'shdc1e1ee9, 32'shdc13b7c9, 32'shdc09520d, 32'shdbfeedb3, 32'shdbf48abd, 32'shdbea292b, 32'shdbdfc8fc, 32'shdbd56a32, 
               32'shdbcb0cce, 32'shdbc0b0ce, 32'shdbb65634, 32'shdbabfd01, 32'shdba1a534, 32'shdb974ece, 32'shdb8cf9cf, 32'shdb82a638, 
               32'shdb785409, 32'shdb6e0342, 32'shdb63b3e5, 32'shdb5965f1, 32'shdb4f1967, 32'shdb44ce46, 32'shdb3a8491, 32'shdb303c46, 
               32'shdb25f566, 32'shdb1baff2, 32'shdb116beb, 32'shdb072950, 32'shdafce821, 32'shdaf2a860, 32'shdae86a0d, 32'shdade2d28, 
               32'shdad3f1b1, 32'shdac9b7a9, 32'shdabf7f11, 32'shdab547e8, 32'shdaab122f, 32'shdaa0dde7, 32'shda96ab0f, 32'shda8c79a9, 
               32'shda8249b4, 32'shda781b31, 32'shda6dee21, 32'shda63c284, 32'shda599859, 32'shda4f6fa3, 32'shda454860, 32'shda3b2292, 
               32'shda30fe38, 32'shda26db54, 32'shda1cb9e5, 32'shda1299ec, 32'shda087b69, 32'shd9fe5e5e, 32'shd9f442c9, 32'shd9ea28ac, 
               32'shd9e01006, 32'shd9d5f8d9, 32'shd9cbe325, 32'shd9c1cee9, 32'shd9b7bc27, 32'shd9adaadf, 32'shd9a39b11, 32'shd9998cbe, 
               32'shd98f7fe6, 32'shd9857489, 32'shd97b6aa8, 32'shd9716243, 32'shd9675b5a, 32'shd95d55ef, 32'shd9535201, 32'shd9494f90, 
               32'shd93f4e9e, 32'shd9354f2a, 32'shd92b5135, 32'shd92154bf, 32'shd91759c9, 32'shd90d6053, 32'shd903685d, 32'shd8f971e8, 
               32'shd8ef7cf4, 32'shd8e58982, 32'shd8db9792, 32'shd8d1a724, 32'shd8c7b838, 32'shd8bdcad0, 32'shd8b3deeb, 32'shd8a9f48a, 
               32'shd8a00bae, 32'shd8962456, 32'shd88c3e83, 32'shd8825a35, 32'shd878776d, 32'shd86e962b, 32'shd864b670, 32'shd85ad83c, 
               32'shd850fb8e, 32'shd8472069, 32'shd83d46cc, 32'shd8336eb7, 32'shd829982b, 32'shd81fc328, 32'shd815efae, 32'shd80c1dbf, 
               32'shd8024d59, 32'shd7f87e7f, 32'shd7eeb130, 32'shd7e4e56c, 32'shd7db1b34, 32'shd7d15288, 32'shd7c78b68, 32'shd7bdc5d6, 
               32'shd7b401d1, 32'shd7aa3f5a, 32'shd7a07e70, 32'shd796bf16, 32'shd78d014a, 32'shd783450d, 32'shd7798a60, 32'shd76fd143, 
               32'shd76619b6, 32'shd75c63ba, 32'shd752af4f, 32'shd748fc75, 32'shd73f4b2e, 32'shd7359b78, 32'shd72bed55, 32'shd72240c5, 
               32'shd71895c9, 32'shd70eec60, 32'shd705448b, 32'shd6fb9e4b, 32'shd6f1f99f, 32'shd6e85689, 32'shd6deb508, 32'shd6d5151d, 
               32'shd6cb76c9, 32'shd6c1da0b, 32'shd6b83ee4, 32'shd6aea555, 32'shd6a50d5d, 32'shd69b76fe, 32'shd691e237, 32'shd6884f09, 
               32'shd67ebd74, 32'shd6752d79, 32'shd66b9f18, 32'shd6621251, 32'shd6588725, 32'shd64efd94, 32'shd645759f, 32'shd63bef46, 
               32'shd6326a88, 32'shd628e767, 32'shd61f65e4, 32'shd615e5fd, 32'shd60c67b4, 32'shd602eb0a, 32'shd5f96ffd, 32'shd5eff690, 
               32'shd5e67ec1, 32'shd5dd0892, 32'shd5d39403, 32'shd5ca2115, 32'shd5c0afc6, 32'shd5b74019, 32'shd5add20d, 32'shd5a465a3, 
               32'shd59afadb, 32'shd59191b5, 32'shd5882a32, 32'shd57ec452, 32'shd5756016, 32'shd56bfd7d, 32'shd5629c89, 32'shd5593d3a, 
               32'shd54fdf8f, 32'shd5468389, 32'shd53d292a, 32'shd533d070, 32'shd52a795d, 32'shd52123f0, 32'shd517d02b, 32'shd50e7e0d, 
               32'shd5052d97, 32'shd4fbdec9, 32'shd4f291a4, 32'shd4e94627, 32'shd4dffc54, 32'shd4d6b42b, 32'shd4cd6dab, 32'shd4c428d6, 
               32'shd4bae5ab, 32'shd4b1a42c, 32'shd4a86458, 32'shd49f2630, 32'shd495e9b3, 32'shd48caee4, 32'shd48375c1, 32'shd47a3e4b, 
               32'shd4710883, 32'shd467d469, 32'shd45ea1fd, 32'shd4557140, 32'shd44c4232, 32'shd44314d3, 32'shd439e923, 32'shd430bf24, 
               32'shd42796d5, 32'shd41e7037, 32'shd4154b4a, 32'shd40c280e, 32'shd4030684, 32'shd3f9e6ad, 32'shd3f0c887, 32'shd3e7ac15, 
               32'shd3de9156, 32'shd3d5784a, 32'shd3cc60f2, 32'shd3c34b4f, 32'shd3ba3760, 32'shd3b12526, 32'shd3a814a2, 32'shd39f05d3, 
               32'shd395f8ba, 32'shd38ced57, 32'shd383e3ab, 32'shd37adbb6, 32'shd371d579, 32'shd368d0f3, 32'shd35fce26, 32'shd356cd11, 
               32'shd34dcdb4, 32'shd344d011, 32'shd33bd427, 32'shd332d9f7, 32'shd329e181, 32'shd320eac6, 32'shd317f5c6, 32'shd30f0280, 
               32'shd30610f7, 32'shd2fd2129, 32'shd2f43318, 32'shd2eb46c3, 32'shd2e25c2b, 32'shd2d97350, 32'shd2d08c33, 32'shd2c7a6d4, 
               32'shd2bec333, 32'shd2b5e151, 32'shd2ad012e, 32'shd2a422ca, 32'shd29b4626, 32'shd2926b41, 32'shd289921e, 32'shd280babb, 
               32'shd277e518, 32'shd26f1138, 32'shd2663f19, 32'shd25d6ebc, 32'shd254a021, 32'shd24bd34a, 32'shd2430835, 32'shd23a3ee4, 
               32'shd2317756, 32'shd228b18d, 32'shd21fed88, 32'shd2172b48, 32'shd20e6acc, 32'shd205ac17, 32'shd1fcef27, 32'shd1f433fd, 
               32'shd1eb7a9a, 32'shd1e2c2fd, 32'shd1da0d28, 32'shd1d1591a, 32'shd1c8a6d4, 32'shd1bff656, 32'shd1b747a0, 32'shd1ae9ab4, 
               32'shd1a5ef90, 32'shd19d4636, 32'shd1949ea6, 32'shd18bf8e0, 32'shd18354e4, 32'shd17ab2b3, 32'shd172124d, 32'shd16973b3, 
               32'shd160d6e5, 32'shd1583be2, 32'shd14fa2ad, 32'shd1470b44, 32'shd13e75a8, 32'shd135e1d9, 32'shd12d4fd9, 32'shd124bfa6, 
               32'shd11c3142, 32'shd113a4ad, 32'shd10b19e7, 32'shd10290f0, 32'shd0fa09c9, 32'shd0f18472, 32'shd0e900ec, 32'shd0e07f36, 
               32'shd0d7ff51, 32'shd0cf813e, 32'shd0c704fd, 32'shd0be8a8d, 32'shd0b611f1, 32'shd0ad9b26, 32'shd0a5262f, 32'shd09cb30b, 
               32'shd09441bb, 32'shd08bd23f, 32'shd0836497, 32'shd07af8c4, 32'shd0728ec6, 32'shd06a269d, 32'shd061c04a, 32'shd0595bcd, 
               32'shd050f926, 32'shd0489856, 32'shd040395d, 32'shd037dc3b, 32'shd02f80f1, 32'shd027277e, 32'shd01ecfe4, 32'shd0167a22, 
               32'shd00e2639, 32'shd005d42a, 32'shcffd83f4, 32'shcff53597, 32'shcfece915, 32'shcfe49e6d, 32'shcfdc55a1, 32'shcfd40eaf, 
               32'shcfcbc999, 32'shcfc3865e, 32'shcfbb4500, 32'shcfb3057d, 32'shcfaac7d8, 32'shcfa28c10, 32'shcf9a5225, 32'shcf921a17, 
               32'shcf89e3e8, 32'shcf81af97, 32'shcf797d24, 32'shcf714c91, 32'shcf691ddd, 32'shcf60f108, 32'shcf58c613, 32'shcf509cfe, 
               32'shcf4875ca, 32'shcf405077, 32'shcf382d05, 32'shcf300b74, 32'shcf27ebc5, 32'shcf1fcdf8, 32'shcf17b20d, 32'shcf0f9805, 
               32'shcf077fe1, 32'shceff699f, 32'shcef75541, 32'shceef42c7, 32'shcee73231, 32'shcedf2380, 32'shced716b4, 32'shcecf0bcd, 
               32'shcec702cb, 32'shcebefbb0, 32'shceb6f67a, 32'shceaef32b, 32'shcea6f1c2, 32'shce9ef241, 32'shce96f4a7, 32'shce8ef8f4, 
               32'shce86ff2a, 32'shce7f0748, 32'shce77114e, 32'shce6f1d3d, 32'shce672b16, 32'shce5f3ad8, 32'shce574c84, 32'shce4f6019, 
               32'shce47759a, 32'shce3f8d05, 32'shce37a65b, 32'shce2fc19c, 32'shce27dec9, 32'shce1ffde2, 32'shce181ee8, 32'shce1041d9, 
               32'shce0866b8, 32'shce008d84, 32'shcdf8b63d, 32'shcdf0e0e4, 32'shcde90d79, 32'shcde13bfd, 32'shcdd96c6f, 32'shcdd19ed0, 
               32'shcdc9d320, 32'shcdc20960, 32'shcdba4190, 32'shcdb27bb0, 32'shcdaab7c0, 32'shcda2f5c2, 32'shcd9b35b4, 32'shcd937798, 
               32'shcd8bbb6d, 32'shcd840134, 32'shcd7c48ee, 32'shcd74929a, 32'shcd6cde39, 32'shcd652bcb, 32'shcd5d7b50, 32'shcd55ccca, 
               32'shcd4e2037, 32'shcd467599, 32'shcd3eccef, 32'shcd37263a, 32'shcd2f817b, 32'shcd27deb0, 32'shcd203ddc, 32'shcd189efe, 
               32'shcd110216, 32'shcd096725, 32'shcd01ce2b, 32'shccfa3729, 32'shccf2a21d, 32'shcceb0f0a, 32'shcce37def, 32'shccdbeecc, 
               32'shccd461a2, 32'shccccd671, 32'shccc54d3a, 32'shccbdc5fc, 32'shccb640b8, 32'shccaebd6e, 32'shcca73c1e, 32'shcc9fbcca, 
               32'shcc983f70, 32'shcc90c412, 32'shcc894aaf, 32'shcc81d349, 32'shcc7a5dde, 32'shcc72ea70, 32'shcc6b78ff, 32'shcc64098b, 
               32'shcc5c9c14, 32'shcc55309b, 32'shcc4dc720, 32'shcc465fa3, 32'shcc3efa25, 32'shcc3796a5, 32'shcc303524, 32'shcc28d5a3, 
               32'shcc217822, 32'shcc1a1ca0, 32'shcc12c31f, 32'shcc0b6b9e, 32'shcc04161e, 32'shcbfcc29f, 32'shcbf57121, 32'shcbee21a5, 
               32'shcbe6d42b, 32'shcbdf88b3, 32'shcbd83f3d, 32'shcbd0f7ca, 32'shcbc9b25a, 32'shcbc26eee, 32'shcbbb2d85, 32'shcbb3ee20, 
               32'shcbacb0bf, 32'shcba57563, 32'shcb9e3c0b, 32'shcb9704b9, 32'shcb8fcf6b, 32'shcb889c23, 32'shcb816ae1, 32'shcb7a3ba5, 
               32'shcb730e70, 32'shcb6be341, 32'shcb64ba19, 32'shcb5d92f8, 32'shcb566ddf, 32'shcb4f4acd, 32'shcb4829c4, 32'shcb410ac3, 
               32'shcb39edca, 32'shcb32d2da, 32'shcb2bb9f4, 32'shcb24a316, 32'shcb1d8e43, 32'shcb167b79, 32'shcb0f6aba, 32'shcb085c05, 
               32'shcb014f5b, 32'shcafa44bc, 32'shcaf33c28, 32'shcaec35a0, 32'shcae53123, 32'shcade2eb3, 32'shcad72e4f, 32'shcad02ff8, 
               32'shcac933ae, 32'shcac23971, 32'shcabb4141, 32'shcab44b1f, 32'shcaad570c, 32'shcaa66506, 32'shca9f750f, 32'shca988727, 
               32'shca919b4e, 32'shca8ab184, 32'shca83c9ca, 32'shca7ce420, 32'shca760086, 32'shca6f1efc, 32'shca683f83, 32'shca61621b, 
               32'shca5a86c4, 32'shca53ad7e, 32'shca4cd64b, 32'shca460129, 32'shca3f2e19, 32'shca385d1d, 32'shca318e32, 32'shca2ac15b, 
               32'shca23f698, 32'shca1d2de7, 32'shca16674b, 32'shca0fa2c3, 32'shca08e04f, 32'shca021fef, 32'shc9fb61a5, 32'shc9f4a570, 
               32'shc9edeb50, 32'shc9e73346, 32'shc9e07d51, 32'shc9d9c973, 32'shc9d317ab, 32'shc9cc67fa, 32'shc9c5ba60, 32'shc9bf0edd, 
               32'shc9b86572, 32'shc9b1be1e, 32'shc9ab18e3, 32'shc9a475bf, 32'shc99dd4b4, 32'shc99735c2, 32'shc99098e9, 32'shc989fe29, 
               32'shc9836582, 32'shc97ccef5, 32'shc9763a83, 32'shc96fa82a, 32'shc96917ec, 32'shc96289c9, 32'shc95bfdc1, 32'shc95573d4, 
               32'shc94eec03, 32'shc948664d, 32'shc941e2b4, 32'shc93b6137, 32'shc934e1d6, 32'shc92e6492, 32'shc927e96b, 32'shc9217062, 
               32'shc91af976, 32'shc91484a8, 32'shc90e11f7, 32'shc907a166, 32'shc90132f2, 32'shc8fac69e, 32'shc8f45c68, 32'shc8edf452, 
               32'shc8e78e5b, 32'shc8e12a84, 32'shc8dac8cd, 32'shc8d46936, 32'shc8ce0bc0, 32'shc8c7b06b, 32'shc8c15736, 32'shc8bb0023, 
               32'shc8b4ab32, 32'shc8ae5862, 32'shc8a807b4, 32'shc8a1b928, 32'shc89b6cbf, 32'shc8952278, 32'shc88eda54, 32'shc8889454, 
               32'shc8825077, 32'shc87c0ebd, 32'shc875cf28, 32'shc86f91b7, 32'shc869566a, 32'shc8631d42, 32'shc85ce63e, 32'shc856b160, 
               32'shc8507ea7, 32'shc84a4e14, 32'shc8441fa6, 32'shc83df35f, 32'shc837c93e, 32'shc831a143, 32'shc82b7b70, 32'shc82557c3, 
               32'shc81f363d, 32'shc81916df, 32'shc812f9a9, 32'shc80cde9b, 32'shc806c5b5, 32'shc800aef7, 32'shc7fa9a62, 32'shc7f487f6, 
               32'shc7ee77b3, 32'shc7e8699a, 32'shc7e25daa, 32'shc7dc53e3, 32'shc7d64c47, 32'shc7d046d6, 32'shc7ca438f, 32'shc7c44272, 
               32'shc7be4381, 32'shc7b846ba, 32'shc7b24c20, 32'shc7ac53b1, 32'shc7a65d6e, 32'shc7a06957, 32'shc79a776c, 32'shc79487ae, 
               32'shc78e9a1d, 32'shc788aeb9, 32'shc782c582, 32'shc77cde79, 32'shc776f99d, 32'shc77116f0, 32'shc76b3671, 32'shc7655820, 
               32'shc75f7bfe, 32'shc759a20a, 32'shc753ca46, 32'shc74df4b1, 32'shc748214c, 32'shc7425016, 32'shc73c8111, 32'shc736b43c, 
               32'shc730e997, 32'shc72b2123, 32'shc7255ae0, 32'shc71f96ce, 32'shc719d4ed, 32'shc714153e, 32'shc70e57c0, 32'shc7089c75, 
               32'shc702e35c, 32'shc6fd2c75, 32'shc6f777c1, 32'shc6f1c540, 32'shc6ec14f2, 32'shc6e666d7, 32'shc6e0baf0, 32'shc6db113d, 
               32'shc6d569be, 32'shc6cfc472, 32'shc6ca215c, 32'shc6c4807a, 32'shc6bee1cd, 32'shc6b94554, 32'shc6b3ab12, 32'shc6ae1304, 
               32'shc6a87d2d, 32'shc6a2e98b, 32'shc69d5820, 32'shc697c8eb, 32'shc6923bec, 32'shc68cb124, 32'shc6872894, 32'shc681a23a, 
               32'shc67c1e18, 32'shc6769c2e, 32'shc6711c7b, 32'shc66b9f01, 32'shc66623be, 32'shc660aab5, 32'shc65b33e4, 32'shc655bf4c, 
               32'shc6504ced, 32'shc64adcc7, 32'shc6456edb, 32'shc6400329, 32'shc63a99b1, 32'shc6353273, 32'shc62fcd6f, 32'shc62a6aa6, 
               32'shc6250a18, 32'shc61fabc4, 32'shc61a4fac, 32'shc614f5cf, 32'shc60f9e2e, 32'shc60a48c9, 32'shc604f5a0, 32'shc5ffa4b3, 
               32'shc5fa5603, 32'shc5f5098f, 32'shc5efbf58, 32'shc5ea775e, 32'shc5e531a1, 32'shc5dfee22, 32'shc5daace1, 32'shc5d56ddd, 
               32'shc5d03118, 32'shc5caf690, 32'shc5c5be47, 32'shc5c0883d, 32'shc5bb5472, 32'shc5b622e6, 32'shc5b0f399, 32'shc5abc68c, 
               32'shc5a69bbe, 32'shc5a17330, 32'shc59c4ce3, 32'shc59728d5, 32'shc5920708, 32'shc58ce77c, 32'shc587ca31, 32'shc582af26, 
               32'shc57d965d, 32'shc5787fd6, 32'shc5736b90, 32'shc56e598c, 32'shc56949ca, 32'shc5643c4a, 32'shc55f310d, 32'shc55a2812, 
               32'shc555215a, 32'shc5501ce5, 32'shc54b1ab4, 32'shc5461ac6, 32'shc5411d1b, 32'shc53c21b4, 32'shc5372891, 32'shc53231b3, 
               32'shc52d3d18, 32'shc5284ac3, 32'shc5235ab2, 32'shc51e6ce6, 32'shc519815f, 32'shc514981d, 32'shc50fb121, 32'shc50acc6b, 
               32'shc505e9fb, 32'shc50109d0, 32'shc4fc2bec, 32'shc4f7504e, 32'shc4f276f7, 32'shc4ed9fe7, 32'shc4e8cb1e, 32'shc4e3f89c, 
               32'shc4df2862, 32'shc4da5a6f, 32'shc4d58ec3, 32'shc4d0c560, 32'shc4cbfe45, 32'shc4c73972, 32'shc4c276e8, 32'shc4bdb6a6, 
               32'shc4b8f8ad, 32'shc4b43cfd, 32'shc4af8397, 32'shc4aacc7a, 32'shc4a617a6, 32'shc4a1651c, 32'shc49cb4dd, 32'shc49806e7, 
               32'shc4935b3c, 32'shc48eb1db, 32'shc48a0ac4, 32'shc48565f9, 32'shc480c379, 32'shc47c2344, 32'shc477855a, 32'shc472e9bc, 
               32'shc46e5069, 32'shc469b963, 32'shc46524a9, 32'shc460923b, 32'shc45c0219, 32'shc4577444, 32'shc452e8bc, 32'shc44e5f80, 
               32'shc449d892, 32'shc44553f2, 32'shc440d19e, 32'shc43c5199, 32'shc437d3e1, 32'shc4335877, 32'shc42edf5c, 32'shc42a688f, 
               32'shc425f410, 32'shc42181e0, 32'shc41d11ff, 32'shc418a46d, 32'shc414392b, 32'shc40fd037, 32'shc40b6994, 32'shc4070540, 
               32'shc402a33c, 32'shc3fe4388, 32'shc3f9e624, 32'shc3f58b10, 32'shc3f1324e, 32'shc3ecdbdc, 32'shc3e887bb, 32'shc3e435ea, 
               32'shc3dfe66c, 32'shc3db993e, 32'shc3d74e62, 32'shc3d305d8, 32'shc3cebfa0, 32'shc3ca7bba, 32'shc3c63a26, 32'shc3c1fae5, 
               32'shc3bdbdf6, 32'shc3b9835a, 32'shc3b54b11, 32'shc3b1151b, 32'shc3ace178, 32'shc3a8b028, 32'shc3a4812c, 32'shc3a05484, 
               32'shc39c2a2f, 32'shc398022f, 32'shc393dc82, 32'shc38fb92a, 32'shc38b9827, 32'shc3877978, 32'shc3835d1e, 32'shc37f4319, 
               32'shc37b2b6a, 32'shc377160f, 32'shc373030a, 32'shc36ef25b, 32'shc36ae401, 32'shc366d7fd, 32'shc362ce50, 32'shc35ec6f8, 
               32'shc35ac1f7, 32'shc356bf4d, 32'shc352bef9, 32'shc34ec0fc, 32'shc34ac556, 32'shc346cc07, 32'shc342d510, 32'shc33ee070, 
               32'shc33aee27, 32'shc336fe37, 32'shc333109e, 32'shc32f255e, 32'shc32b3c75, 32'shc32755e5, 32'shc32371ae, 32'shc31f8fcf, 
               32'shc31bb049, 32'shc317d31c, 32'shc313f848, 32'shc3101fce, 32'shc30c49ad, 32'shc30875e5, 32'shc304a477, 32'shc300d563, 
               32'shc2fd08a9, 32'shc2f93e4a, 32'shc2f57644, 32'shc2f1b099, 32'shc2eded49, 32'shc2ea2c53, 32'shc2e66db8, 32'shc2e2b178, 
               32'shc2def794, 32'shc2db400a, 32'shc2d78add, 32'shc2d3d80a, 32'shc2d02794, 32'shc2cc7979, 32'shc2c8cdbb, 32'shc2c52459, 
               32'shc2c17d52, 32'shc2bdd8a9, 32'shc2ba365c, 32'shc2b6966c, 32'shc2b2f8d8, 32'shc2af5da2, 32'shc2abc4c9, 32'shc2a82e4d, 
               32'shc2a49a2e, 32'shc2a1086d, 32'shc29d790a, 32'shc299ec05, 32'shc296615d, 32'shc292d914, 32'shc28f5329, 32'shc28bcf9c, 
               32'shc2884e6e, 32'shc284cf9f, 32'shc281532e, 32'shc27dd91c, 32'shc27a616a, 32'shc276ec16, 32'shc2737922, 32'shc270088e, 
               32'shc26c9a58, 32'shc2692e83, 32'shc265c50e, 32'shc2625df8, 32'shc25ef943, 32'shc25b96ee, 32'shc25836f9, 32'shc254d965, 
               32'shc2517e31, 32'shc24e255e, 32'shc24aceed, 32'shc2477adc, 32'shc244292c, 32'shc240d9de, 32'shc23d8cf1, 32'shc23a4265, 
               32'shc236fa3b, 32'shc233b473, 32'shc230710d, 32'shc22d3009, 32'shc229f167, 32'shc226b528, 32'shc2237b4b, 32'shc22043d0, 
               32'shc21d0eb8, 32'shc219dc03, 32'shc216abb1, 32'shc2137dc2, 32'shc2105236, 32'shc20d290d, 32'shc20a0248, 32'shc206dde6, 
               32'shc203bbe8, 32'shc2009c4e, 32'shc1fd7f17, 32'shc1fa6445, 32'shc1f74bd6, 32'shc1f435cc, 32'shc1f12227, 32'shc1ee10e5, 
               32'shc1eb0209, 32'shc1e7f591, 32'shc1e4eb7e, 32'shc1e1e3d0, 32'shc1dede87, 32'shc1dbdba3, 32'shc1d8db25, 32'shc1d5dd0c, 
               32'shc1d2e158, 32'shc1cfe80a, 32'shc1ccf122, 32'shc1c9fca0, 32'shc1c70a84, 32'shc1c41ace, 32'shc1c12d7e, 32'shc1be4294, 
               32'shc1bb5a11, 32'shc1b873f5, 32'shc1b5903f, 32'shc1b2aef0, 32'shc1afd007, 32'shc1acf386, 32'shc1aa196c, 32'shc1a741b9, 
               32'shc1a46c6e, 32'shc1a1998a, 32'shc19ec90d, 32'shc19bfaf9, 32'shc1992f4c, 32'shc1966606, 32'shc1939f29, 32'shc190dab4, 
               32'shc18e18a7, 32'shc18b5903, 32'shc1889bc6, 32'shc185e0f3, 32'shc1832888, 32'shc1807285, 32'shc17dbeec, 32'shc17b0dbb, 
               32'shc1785ef4, 32'shc175b296, 32'shc17308a1, 32'shc1706115, 32'shc16dbbf3, 32'shc16b193a, 32'shc16878eb, 32'shc165db05, 
               32'shc1633f8a, 32'shc160a678, 32'shc15e0fd1, 32'shc15b7b94, 32'shc158e9c1, 32'shc1565a58, 32'shc153cd5a, 32'shc15142c6, 
               32'shc14eba9d, 32'shc14c34df, 32'shc149b18b, 32'shc14730a3, 32'shc144b225, 32'shc1423613, 32'shc13fbc6c, 32'shc13d4530, 
               32'shc13ad060, 32'shc1385dfb, 32'shc135ee02, 32'shc1338075, 32'shc1311553, 32'shc12eac9d, 32'shc12c4653, 32'shc129e276, 
               32'shc1278104, 32'shc12521ff, 32'shc122c566, 32'shc1206b39, 32'shc11e1379, 32'shc11bbe26, 32'shc1196b3f, 32'shc1171ac6, 
               32'shc114ccb9, 32'shc1128119, 32'shc11037e6, 32'shc10df120, 32'shc10bacc8, 32'shc1096add, 32'shc1072b5f, 32'shc104ee4f, 
               32'shc102b3ac, 32'shc1007b77, 32'shc0fe45b0, 32'shc0fc1257, 32'shc0f9e16b, 32'shc0f7b2ee, 32'shc0f586df, 32'shc0f35d3e, 
               32'shc0f1360b, 32'shc0ef1147, 32'shc0eceef1, 32'shc0eacf09, 32'shc0e8b190, 32'shc0e69686, 32'shc0e47deb, 32'shc0e267be, 
               32'shc0e05401, 32'shc0de42b2, 32'shc0dc33d2, 32'shc0da2762, 32'shc0d81d61, 32'shc0d615cf, 32'shc0d410ad, 32'shc0d20dfa, 
               32'shc0d00db6, 32'shc0ce0fe3, 32'shc0cc147f, 32'shc0ca1b8a, 32'shc0c82506, 32'shc0c630f2, 32'shc0c43f4d, 32'shc0c25019, 
               32'shc0c06355, 32'shc0be7901, 32'shc0bc911d, 32'shc0baabaa, 32'shc0b8c8a7, 32'shc0b6e815, 32'shc0b509f3, 32'shc0b32e42, 
               32'shc0b15502, 32'shc0af7e33, 32'shc0ada9d4, 32'shc0abd7e6, 32'shc0aa086a, 32'shc0a83b5e, 32'shc0a670c4, 32'shc0a4a89b, 
               32'shc0a2e2e3, 32'shc0a11f9d, 32'shc09f5ec8, 32'shc09da065, 32'shc09be473, 32'shc09a2af3, 32'shc09873e4, 32'shc096bf48, 
               32'shc0950d1d, 32'shc0935d64, 32'shc091b01d, 32'shc0900548, 32'shc08e5ce5, 32'shc08cb6f5, 32'shc08b1376, 32'shc089726a, 
               32'shc087d3d0, 32'shc08637a9, 32'shc0849df4, 32'shc08306b2, 32'shc08171e2, 32'shc07fdf85, 32'shc07e4f9b, 32'shc07cc223, 
               32'shc07b371e, 32'shc079ae8c, 32'shc078286e, 32'shc076a4c2, 32'shc0752389, 32'shc073a4c3, 32'shc0722871, 32'shc070ae92, 
               32'shc06f3726, 32'shc06dc22e, 32'shc06c4fa8, 32'shc06adf97, 32'shc06971f9, 32'shc06806ce, 32'shc0669e18, 32'shc06537d4, 
               32'shc063d405, 32'shc06272aa, 32'shc06113c2, 32'shc05fb74e, 32'shc05e5d4e, 32'shc05d05c3, 32'shc05bb0ab, 32'shc05a5e07, 
               32'shc0590dd8, 32'shc057c01d, 32'shc05674d6, 32'shc0552c03, 32'shc053e5a5, 32'shc052a1bb, 32'shc0516045, 32'shc0502145, 
               32'shc04ee4b8, 32'shc04daaa1, 32'shc04c72fe, 32'shc04b3dcf, 32'shc04a0b16, 32'shc048dad1, 32'shc047ad01, 32'shc04681a6, 
               32'shc04558c0, 32'shc044324f, 32'shc0430e53, 32'shc041eccc, 32'shc040cdba, 32'shc03fb11d, 32'shc03e96f6, 32'shc03d7f44, 
               32'shc03c6a07, 32'shc03b573f, 32'shc03a46ed, 32'shc0393910, 32'shc0382da8, 32'shc03724b6, 32'shc0361e3a, 32'shc0351a33, 
               32'shc03418a2, 32'shc0331986, 32'shc0321ce0, 32'shc03122b0, 32'shc0302af5, 32'shc02f35b1, 32'shc02e42e2, 32'shc02d5289, 
               32'shc02c64a6, 32'shc02b7939, 32'shc02a9042, 32'shc029a9c1, 32'shc028c5b6, 32'shc027e421, 32'shc0270502, 32'shc0262859, 
               32'shc0254e27, 32'shc024766a, 32'shc023a124, 32'shc022ce54, 32'shc021fdfb, 32'shc0213018, 32'shc02064ab, 32'shc01f9bb5, 
               32'shc01ed535, 32'shc01e112b, 32'shc01d4f99, 32'shc01c907c, 32'shc01bd3d6, 32'shc01b19a7, 32'shc01a61ee, 32'shc019acac, 
               32'shc018f9e1, 32'shc018498c, 32'shc0179bae, 32'shc016f047, 32'shc0164757, 32'shc015a0dd, 32'shc014fcda, 32'shc0145b4e, 
               32'shc013bc39, 32'shc0131f9b, 32'shc0128574, 32'shc011edc3, 32'shc011588a, 32'shc010c5c7, 32'shc010357c, 32'shc00fa7a8, 
               32'shc00f1c4a, 32'shc00e9364, 32'shc00e0cf5, 32'shc00d88fd, 32'shc00d077c, 32'shc00c8872, 32'shc00c0be0, 32'shc00b91c4, 
               32'shc00b1a20, 32'shc00aa4f3, 32'shc00a323d, 32'shc009c1ff, 32'shc0095438, 32'shc008e8e8, 32'shc008800f, 32'shc00819ae, 
               32'shc007b5c4, 32'shc0075452, 32'shc006f556, 32'shc00698d3, 32'shc0063ec6, 32'shc005e731, 32'shc0059214, 32'shc0053f6e, 
               32'shc004ef3f, 32'shc004a188, 32'shc0045648, 32'shc0040d80, 32'shc003c72f, 32'shc0038356, 32'shc00341f4, 32'shc003030a, 
               32'shc002c697, 32'shc0028c9c, 32'shc0025519, 32'shc002200d, 32'shc001ed78, 32'shc001bd5c, 32'shc0018fb6, 32'shc0016489, 
               32'shc0013bd3, 32'shc0011594, 32'shc000f1ce, 32'shc000d07e, 32'shc000b1a7, 32'shc0009547, 32'shc0007b5f, 32'shc00063ee, 
               32'shc0004ef5, 32'shc0003c74, 32'shc0002c6a, 32'shc0001ed8, 32'shc00013bd, 32'shc0000b1a, 32'shc00004ef, 32'shc000013c, 
               32'shc0000000, 32'shc000013c, 32'shc00004ef, 32'shc0000b1a, 32'shc00013bd, 32'shc0001ed8, 32'shc0002c6a, 32'shc0003c74, 
               32'shc0004ef5, 32'shc00063ee, 32'shc0007b5f, 32'shc0009547, 32'shc000b1a7, 32'shc000d07e, 32'shc000f1ce, 32'shc0011594, 
               32'shc0013bd3, 32'shc0016489, 32'shc0018fb6, 32'shc001bd5c, 32'shc001ed78, 32'shc002200d, 32'shc0025519, 32'shc0028c9c, 
               32'shc002c697, 32'shc003030a, 32'shc00341f4, 32'shc0038356, 32'shc003c72f, 32'shc0040d80, 32'shc0045648, 32'shc004a188, 
               32'shc004ef3f, 32'shc0053f6e, 32'shc0059214, 32'shc005e731, 32'shc0063ec6, 32'shc00698d3, 32'shc006f556, 32'shc0075452, 
               32'shc007b5c4, 32'shc00819ae, 32'shc008800f, 32'shc008e8e8, 32'shc0095438, 32'shc009c1ff, 32'shc00a323d, 32'shc00aa4f3, 
               32'shc00b1a20, 32'shc00b91c4, 32'shc00c0be0, 32'shc00c8872, 32'shc00d077c, 32'shc00d88fd, 32'shc00e0cf5, 32'shc00e9364, 
               32'shc00f1c4a, 32'shc00fa7a8, 32'shc010357c, 32'shc010c5c7, 32'shc011588a, 32'shc011edc3, 32'shc0128574, 32'shc0131f9b, 
               32'shc013bc39, 32'shc0145b4e, 32'shc014fcda, 32'shc015a0dd, 32'shc0164757, 32'shc016f047, 32'shc0179bae, 32'shc018498c, 
               32'shc018f9e1, 32'shc019acac, 32'shc01a61ee, 32'shc01b19a7, 32'shc01bd3d6, 32'shc01c907c, 32'shc01d4f99, 32'shc01e112b, 
               32'shc01ed535, 32'shc01f9bb5, 32'shc02064ab, 32'shc0213018, 32'shc021fdfb, 32'shc022ce54, 32'shc023a124, 32'shc024766a, 
               32'shc0254e27, 32'shc0262859, 32'shc0270502, 32'shc027e421, 32'shc028c5b6, 32'shc029a9c1, 32'shc02a9042, 32'shc02b7939, 
               32'shc02c64a6, 32'shc02d5289, 32'shc02e42e2, 32'shc02f35b1, 32'shc0302af5, 32'shc03122b0, 32'shc0321ce0, 32'shc0331986, 
               32'shc03418a2, 32'shc0351a33, 32'shc0361e3a, 32'shc03724b6, 32'shc0382da8, 32'shc0393910, 32'shc03a46ed, 32'shc03b573f, 
               32'shc03c6a07, 32'shc03d7f44, 32'shc03e96f6, 32'shc03fb11d, 32'shc040cdba, 32'shc041eccc, 32'shc0430e53, 32'shc044324f, 
               32'shc04558c0, 32'shc04681a6, 32'shc047ad01, 32'shc048dad1, 32'shc04a0b16, 32'shc04b3dcf, 32'shc04c72fe, 32'shc04daaa1, 
               32'shc04ee4b8, 32'shc0502145, 32'shc0516045, 32'shc052a1bb, 32'shc053e5a5, 32'shc0552c03, 32'shc05674d6, 32'shc057c01d, 
               32'shc0590dd8, 32'shc05a5e07, 32'shc05bb0ab, 32'shc05d05c3, 32'shc05e5d4e, 32'shc05fb74e, 32'shc06113c2, 32'shc06272aa, 
               32'shc063d405, 32'shc06537d4, 32'shc0669e18, 32'shc06806ce, 32'shc06971f9, 32'shc06adf97, 32'shc06c4fa8, 32'shc06dc22e, 
               32'shc06f3726, 32'shc070ae92, 32'shc0722871, 32'shc073a4c3, 32'shc0752389, 32'shc076a4c2, 32'shc078286e, 32'shc079ae8c, 
               32'shc07b371e, 32'shc07cc223, 32'shc07e4f9b, 32'shc07fdf85, 32'shc08171e2, 32'shc08306b2, 32'shc0849df4, 32'shc08637a9, 
               32'shc087d3d0, 32'shc089726a, 32'shc08b1376, 32'shc08cb6f5, 32'shc08e5ce5, 32'shc0900548, 32'shc091b01d, 32'shc0935d64, 
               32'shc0950d1d, 32'shc096bf48, 32'shc09873e4, 32'shc09a2af3, 32'shc09be473, 32'shc09da065, 32'shc09f5ec8, 32'shc0a11f9d, 
               32'shc0a2e2e3, 32'shc0a4a89b, 32'shc0a670c4, 32'shc0a83b5e, 32'shc0aa086a, 32'shc0abd7e6, 32'shc0ada9d4, 32'shc0af7e33, 
               32'shc0b15502, 32'shc0b32e42, 32'shc0b509f3, 32'shc0b6e815, 32'shc0b8c8a7, 32'shc0baabaa, 32'shc0bc911d, 32'shc0be7901, 
               32'shc0c06355, 32'shc0c25019, 32'shc0c43f4d, 32'shc0c630f2, 32'shc0c82506, 32'shc0ca1b8a, 32'shc0cc147f, 32'shc0ce0fe3, 
               32'shc0d00db6, 32'shc0d20dfa, 32'shc0d410ad, 32'shc0d615cf, 32'shc0d81d61, 32'shc0da2762, 32'shc0dc33d2, 32'shc0de42b2, 
               32'shc0e05401, 32'shc0e267be, 32'shc0e47deb, 32'shc0e69686, 32'shc0e8b190, 32'shc0eacf09, 32'shc0eceef1, 32'shc0ef1147, 
               32'shc0f1360b, 32'shc0f35d3e, 32'shc0f586df, 32'shc0f7b2ee, 32'shc0f9e16b, 32'shc0fc1257, 32'shc0fe45b0, 32'shc1007b77, 
               32'shc102b3ac, 32'shc104ee4f, 32'shc1072b5f, 32'shc1096add, 32'shc10bacc8, 32'shc10df120, 32'shc11037e6, 32'shc1128119, 
               32'shc114ccb9, 32'shc1171ac6, 32'shc1196b3f, 32'shc11bbe26, 32'shc11e1379, 32'shc1206b39, 32'shc122c566, 32'shc12521ff, 
               32'shc1278104, 32'shc129e276, 32'shc12c4653, 32'shc12eac9d, 32'shc1311553, 32'shc1338075, 32'shc135ee02, 32'shc1385dfb, 
               32'shc13ad060, 32'shc13d4530, 32'shc13fbc6c, 32'shc1423613, 32'shc144b225, 32'shc14730a3, 32'shc149b18b, 32'shc14c34df, 
               32'shc14eba9d, 32'shc15142c6, 32'shc153cd5a, 32'shc1565a58, 32'shc158e9c1, 32'shc15b7b94, 32'shc15e0fd1, 32'shc160a678, 
               32'shc1633f8a, 32'shc165db05, 32'shc16878eb, 32'shc16b193a, 32'shc16dbbf3, 32'shc1706115, 32'shc17308a1, 32'shc175b296, 
               32'shc1785ef4, 32'shc17b0dbb, 32'shc17dbeec, 32'shc1807285, 32'shc1832888, 32'shc185e0f3, 32'shc1889bc6, 32'shc18b5903, 
               32'shc18e18a7, 32'shc190dab4, 32'shc1939f29, 32'shc1966606, 32'shc1992f4c, 32'shc19bfaf9, 32'shc19ec90d, 32'shc1a1998a, 
               32'shc1a46c6e, 32'shc1a741b9, 32'shc1aa196c, 32'shc1acf386, 32'shc1afd007, 32'shc1b2aef0, 32'shc1b5903f, 32'shc1b873f5, 
               32'shc1bb5a11, 32'shc1be4294, 32'shc1c12d7e, 32'shc1c41ace, 32'shc1c70a84, 32'shc1c9fca0, 32'shc1ccf122, 32'shc1cfe80a, 
               32'shc1d2e158, 32'shc1d5dd0c, 32'shc1d8db25, 32'shc1dbdba3, 32'shc1dede87, 32'shc1e1e3d0, 32'shc1e4eb7e, 32'shc1e7f591, 
               32'shc1eb0209, 32'shc1ee10e5, 32'shc1f12227, 32'shc1f435cc, 32'shc1f74bd6, 32'shc1fa6445, 32'shc1fd7f17, 32'shc2009c4e, 
               32'shc203bbe8, 32'shc206dde6, 32'shc20a0248, 32'shc20d290d, 32'shc2105236, 32'shc2137dc2, 32'shc216abb1, 32'shc219dc03, 
               32'shc21d0eb8, 32'shc22043d0, 32'shc2237b4b, 32'shc226b528, 32'shc229f167, 32'shc22d3009, 32'shc230710d, 32'shc233b473, 
               32'shc236fa3b, 32'shc23a4265, 32'shc23d8cf1, 32'shc240d9de, 32'shc244292c, 32'shc2477adc, 32'shc24aceed, 32'shc24e255e, 
               32'shc2517e31, 32'shc254d965, 32'shc25836f9, 32'shc25b96ee, 32'shc25ef943, 32'shc2625df8, 32'shc265c50e, 32'shc2692e83, 
               32'shc26c9a58, 32'shc270088e, 32'shc2737922, 32'shc276ec16, 32'shc27a616a, 32'shc27dd91c, 32'shc281532e, 32'shc284cf9f, 
               32'shc2884e6e, 32'shc28bcf9c, 32'shc28f5329, 32'shc292d914, 32'shc296615d, 32'shc299ec05, 32'shc29d790a, 32'shc2a1086d, 
               32'shc2a49a2e, 32'shc2a82e4d, 32'shc2abc4c9, 32'shc2af5da2, 32'shc2b2f8d8, 32'shc2b6966c, 32'shc2ba365c, 32'shc2bdd8a9, 
               32'shc2c17d52, 32'shc2c52459, 32'shc2c8cdbb, 32'shc2cc7979, 32'shc2d02794, 32'shc2d3d80a, 32'shc2d78add, 32'shc2db400a, 
               32'shc2def794, 32'shc2e2b178, 32'shc2e66db8, 32'shc2ea2c53, 32'shc2eded49, 32'shc2f1b099, 32'shc2f57644, 32'shc2f93e4a, 
               32'shc2fd08a9, 32'shc300d563, 32'shc304a477, 32'shc30875e5, 32'shc30c49ad, 32'shc3101fce, 32'shc313f848, 32'shc317d31c, 
               32'shc31bb049, 32'shc31f8fcf, 32'shc32371ae, 32'shc32755e5, 32'shc32b3c75, 32'shc32f255e, 32'shc333109e, 32'shc336fe37, 
               32'shc33aee27, 32'shc33ee070, 32'shc342d510, 32'shc346cc07, 32'shc34ac556, 32'shc34ec0fc, 32'shc352bef9, 32'shc356bf4d, 
               32'shc35ac1f7, 32'shc35ec6f8, 32'shc362ce50, 32'shc366d7fd, 32'shc36ae401, 32'shc36ef25b, 32'shc373030a, 32'shc377160f, 
               32'shc37b2b6a, 32'shc37f4319, 32'shc3835d1e, 32'shc3877978, 32'shc38b9827, 32'shc38fb92a, 32'shc393dc82, 32'shc398022f, 
               32'shc39c2a2f, 32'shc3a05484, 32'shc3a4812c, 32'shc3a8b028, 32'shc3ace178, 32'shc3b1151b, 32'shc3b54b11, 32'shc3b9835a, 
               32'shc3bdbdf6, 32'shc3c1fae5, 32'shc3c63a26, 32'shc3ca7bba, 32'shc3cebfa0, 32'shc3d305d8, 32'shc3d74e62, 32'shc3db993e, 
               32'shc3dfe66c, 32'shc3e435ea, 32'shc3e887bb, 32'shc3ecdbdc, 32'shc3f1324e, 32'shc3f58b10, 32'shc3f9e624, 32'shc3fe4388, 
               32'shc402a33c, 32'shc4070540, 32'shc40b6994, 32'shc40fd037, 32'shc414392b, 32'shc418a46d, 32'shc41d11ff, 32'shc42181e0, 
               32'shc425f410, 32'shc42a688f, 32'shc42edf5c, 32'shc4335877, 32'shc437d3e1, 32'shc43c5199, 32'shc440d19e, 32'shc44553f2, 
               32'shc449d892, 32'shc44e5f80, 32'shc452e8bc, 32'shc4577444, 32'shc45c0219, 32'shc460923b, 32'shc46524a9, 32'shc469b963, 
               32'shc46e5069, 32'shc472e9bc, 32'shc477855a, 32'shc47c2344, 32'shc480c379, 32'shc48565f9, 32'shc48a0ac4, 32'shc48eb1db, 
               32'shc4935b3c, 32'shc49806e7, 32'shc49cb4dd, 32'shc4a1651c, 32'shc4a617a6, 32'shc4aacc7a, 32'shc4af8397, 32'shc4b43cfd, 
               32'shc4b8f8ad, 32'shc4bdb6a6, 32'shc4c276e8, 32'shc4c73972, 32'shc4cbfe45, 32'shc4d0c560, 32'shc4d58ec3, 32'shc4da5a6f, 
               32'shc4df2862, 32'shc4e3f89c, 32'shc4e8cb1e, 32'shc4ed9fe7, 32'shc4f276f7, 32'shc4f7504e, 32'shc4fc2bec, 32'shc50109d0, 
               32'shc505e9fb, 32'shc50acc6b, 32'shc50fb121, 32'shc514981d, 32'shc519815f, 32'shc51e6ce6, 32'shc5235ab2, 32'shc5284ac3, 
               32'shc52d3d18, 32'shc53231b3, 32'shc5372891, 32'shc53c21b4, 32'shc5411d1b, 32'shc5461ac6, 32'shc54b1ab4, 32'shc5501ce5, 
               32'shc555215a, 32'shc55a2812, 32'shc55f310d, 32'shc5643c4a, 32'shc56949ca, 32'shc56e598c, 32'shc5736b90, 32'shc5787fd6, 
               32'shc57d965d, 32'shc582af26, 32'shc587ca31, 32'shc58ce77c, 32'shc5920708, 32'shc59728d5, 32'shc59c4ce3, 32'shc5a17330, 
               32'shc5a69bbe, 32'shc5abc68c, 32'shc5b0f399, 32'shc5b622e6, 32'shc5bb5472, 32'shc5c0883d, 32'shc5c5be47, 32'shc5caf690, 
               32'shc5d03118, 32'shc5d56ddd, 32'shc5daace1, 32'shc5dfee22, 32'shc5e531a1, 32'shc5ea775e, 32'shc5efbf58, 32'shc5f5098f, 
               32'shc5fa5603, 32'shc5ffa4b3, 32'shc604f5a0, 32'shc60a48c9, 32'shc60f9e2e, 32'shc614f5cf, 32'shc61a4fac, 32'shc61fabc4, 
               32'shc6250a18, 32'shc62a6aa6, 32'shc62fcd6f, 32'shc6353273, 32'shc63a99b1, 32'shc6400329, 32'shc6456edb, 32'shc64adcc7, 
               32'shc6504ced, 32'shc655bf4c, 32'shc65b33e4, 32'shc660aab5, 32'shc66623be, 32'shc66b9f01, 32'shc6711c7b, 32'shc6769c2e, 
               32'shc67c1e18, 32'shc681a23a, 32'shc6872894, 32'shc68cb124, 32'shc6923bec, 32'shc697c8eb, 32'shc69d5820, 32'shc6a2e98b, 
               32'shc6a87d2d, 32'shc6ae1304, 32'shc6b3ab12, 32'shc6b94554, 32'shc6bee1cd, 32'shc6c4807a, 32'shc6ca215c, 32'shc6cfc472, 
               32'shc6d569be, 32'shc6db113d, 32'shc6e0baf0, 32'shc6e666d7, 32'shc6ec14f2, 32'shc6f1c540, 32'shc6f777c1, 32'shc6fd2c75, 
               32'shc702e35c, 32'shc7089c75, 32'shc70e57c0, 32'shc714153e, 32'shc719d4ed, 32'shc71f96ce, 32'shc7255ae0, 32'shc72b2123, 
               32'shc730e997, 32'shc736b43c, 32'shc73c8111, 32'shc7425016, 32'shc748214c, 32'shc74df4b1, 32'shc753ca46, 32'shc759a20a, 
               32'shc75f7bfe, 32'shc7655820, 32'shc76b3671, 32'shc77116f0, 32'shc776f99d, 32'shc77cde79, 32'shc782c582, 32'shc788aeb9, 
               32'shc78e9a1d, 32'shc79487ae, 32'shc79a776c, 32'shc7a06957, 32'shc7a65d6e, 32'shc7ac53b1, 32'shc7b24c20, 32'shc7b846ba, 
               32'shc7be4381, 32'shc7c44272, 32'shc7ca438f, 32'shc7d046d6, 32'shc7d64c47, 32'shc7dc53e3, 32'shc7e25daa, 32'shc7e8699a, 
               32'shc7ee77b3, 32'shc7f487f6, 32'shc7fa9a62, 32'shc800aef7, 32'shc806c5b5, 32'shc80cde9b, 32'shc812f9a9, 32'shc81916df, 
               32'shc81f363d, 32'shc82557c3, 32'shc82b7b70, 32'shc831a143, 32'shc837c93e, 32'shc83df35f, 32'shc8441fa6, 32'shc84a4e14, 
               32'shc8507ea7, 32'shc856b160, 32'shc85ce63e, 32'shc8631d42, 32'shc869566a, 32'shc86f91b7, 32'shc875cf28, 32'shc87c0ebd, 
               32'shc8825077, 32'shc8889454, 32'shc88eda54, 32'shc8952278, 32'shc89b6cbf, 32'shc8a1b928, 32'shc8a807b4, 32'shc8ae5862, 
               32'shc8b4ab32, 32'shc8bb0023, 32'shc8c15736, 32'shc8c7b06b, 32'shc8ce0bc0, 32'shc8d46936, 32'shc8dac8cd, 32'shc8e12a84, 
               32'shc8e78e5b, 32'shc8edf452, 32'shc8f45c68, 32'shc8fac69e, 32'shc90132f2, 32'shc907a166, 32'shc90e11f7, 32'shc91484a8, 
               32'shc91af976, 32'shc9217062, 32'shc927e96b, 32'shc92e6492, 32'shc934e1d6, 32'shc93b6137, 32'shc941e2b4, 32'shc948664d, 
               32'shc94eec03, 32'shc95573d4, 32'shc95bfdc1, 32'shc96289c9, 32'shc96917ec, 32'shc96fa82a, 32'shc9763a83, 32'shc97ccef5, 
               32'shc9836582, 32'shc989fe29, 32'shc99098e9, 32'shc99735c2, 32'shc99dd4b4, 32'shc9a475bf, 32'shc9ab18e3, 32'shc9b1be1e, 
               32'shc9b86572, 32'shc9bf0edd, 32'shc9c5ba60, 32'shc9cc67fa, 32'shc9d317ab, 32'shc9d9c973, 32'shc9e07d51, 32'shc9e73346, 
               32'shc9edeb50, 32'shc9f4a570, 32'shc9fb61a5, 32'shca021fef, 32'shca08e04f, 32'shca0fa2c3, 32'shca16674b, 32'shca1d2de7, 
               32'shca23f698, 32'shca2ac15b, 32'shca318e32, 32'shca385d1d, 32'shca3f2e19, 32'shca460129, 32'shca4cd64b, 32'shca53ad7e, 
               32'shca5a86c4, 32'shca61621b, 32'shca683f83, 32'shca6f1efc, 32'shca760086, 32'shca7ce420, 32'shca83c9ca, 32'shca8ab184, 
               32'shca919b4e, 32'shca988727, 32'shca9f750f, 32'shcaa66506, 32'shcaad570c, 32'shcab44b1f, 32'shcabb4141, 32'shcac23971, 
               32'shcac933ae, 32'shcad02ff8, 32'shcad72e4f, 32'shcade2eb3, 32'shcae53123, 32'shcaec35a0, 32'shcaf33c28, 32'shcafa44bc, 
               32'shcb014f5b, 32'shcb085c05, 32'shcb0f6aba, 32'shcb167b79, 32'shcb1d8e43, 32'shcb24a316, 32'shcb2bb9f4, 32'shcb32d2da, 
               32'shcb39edca, 32'shcb410ac3, 32'shcb4829c4, 32'shcb4f4acd, 32'shcb566ddf, 32'shcb5d92f8, 32'shcb64ba19, 32'shcb6be341, 
               32'shcb730e70, 32'shcb7a3ba5, 32'shcb816ae1, 32'shcb889c23, 32'shcb8fcf6b, 32'shcb9704b9, 32'shcb9e3c0b, 32'shcba57563, 
               32'shcbacb0bf, 32'shcbb3ee20, 32'shcbbb2d85, 32'shcbc26eee, 32'shcbc9b25a, 32'shcbd0f7ca, 32'shcbd83f3d, 32'shcbdf88b3, 
               32'shcbe6d42b, 32'shcbee21a5, 32'shcbf57121, 32'shcbfcc29f, 32'shcc04161e, 32'shcc0b6b9e, 32'shcc12c31f, 32'shcc1a1ca0, 
               32'shcc217822, 32'shcc28d5a3, 32'shcc303524, 32'shcc3796a5, 32'shcc3efa25, 32'shcc465fa3, 32'shcc4dc720, 32'shcc55309b, 
               32'shcc5c9c14, 32'shcc64098b, 32'shcc6b78ff, 32'shcc72ea70, 32'shcc7a5dde, 32'shcc81d349, 32'shcc894aaf, 32'shcc90c412, 
               32'shcc983f70, 32'shcc9fbcca, 32'shcca73c1e, 32'shccaebd6e, 32'shccb640b8, 32'shccbdc5fc, 32'shccc54d3a, 32'shccccd671, 
               32'shccd461a2, 32'shccdbeecc, 32'shcce37def, 32'shcceb0f0a, 32'shccf2a21d, 32'shccfa3729, 32'shcd01ce2b, 32'shcd096725, 
               32'shcd110216, 32'shcd189efe, 32'shcd203ddc, 32'shcd27deb0, 32'shcd2f817b, 32'shcd37263a, 32'shcd3eccef, 32'shcd467599, 
               32'shcd4e2037, 32'shcd55ccca, 32'shcd5d7b50, 32'shcd652bcb, 32'shcd6cde39, 32'shcd74929a, 32'shcd7c48ee, 32'shcd840134, 
               32'shcd8bbb6d, 32'shcd937798, 32'shcd9b35b4, 32'shcda2f5c2, 32'shcdaab7c0, 32'shcdb27bb0, 32'shcdba4190, 32'shcdc20960, 
               32'shcdc9d320, 32'shcdd19ed0, 32'shcdd96c6f, 32'shcde13bfd, 32'shcde90d79, 32'shcdf0e0e4, 32'shcdf8b63d, 32'shce008d84, 
               32'shce0866b8, 32'shce1041d9, 32'shce181ee8, 32'shce1ffde2, 32'shce27dec9, 32'shce2fc19c, 32'shce37a65b, 32'shce3f8d05, 
               32'shce47759a, 32'shce4f6019, 32'shce574c84, 32'shce5f3ad8, 32'shce672b16, 32'shce6f1d3d, 32'shce77114e, 32'shce7f0748, 
               32'shce86ff2a, 32'shce8ef8f4, 32'shce96f4a7, 32'shce9ef241, 32'shcea6f1c2, 32'shceaef32b, 32'shceb6f67a, 32'shcebefbb0, 
               32'shcec702cb, 32'shcecf0bcd, 32'shced716b4, 32'shcedf2380, 32'shcee73231, 32'shceef42c7, 32'shcef75541, 32'shceff699f, 
               32'shcf077fe1, 32'shcf0f9805, 32'shcf17b20d, 32'shcf1fcdf8, 32'shcf27ebc5, 32'shcf300b74, 32'shcf382d05, 32'shcf405077, 
               32'shcf4875ca, 32'shcf509cfe, 32'shcf58c613, 32'shcf60f108, 32'shcf691ddd, 32'shcf714c91, 32'shcf797d24, 32'shcf81af97, 
               32'shcf89e3e8, 32'shcf921a17, 32'shcf9a5225, 32'shcfa28c10, 32'shcfaac7d8, 32'shcfb3057d, 32'shcfbb4500, 32'shcfc3865e, 
               32'shcfcbc999, 32'shcfd40eaf, 32'shcfdc55a1, 32'shcfe49e6d, 32'shcfece915, 32'shcff53597, 32'shcffd83f4, 32'shd005d42a, 
               32'shd00e2639, 32'shd0167a22, 32'shd01ecfe4, 32'shd027277e, 32'shd02f80f1, 32'shd037dc3b, 32'shd040395d, 32'shd0489856, 
               32'shd050f926, 32'shd0595bcd, 32'shd061c04a, 32'shd06a269d, 32'shd0728ec6, 32'shd07af8c4, 32'shd0836497, 32'shd08bd23f, 
               32'shd09441bb, 32'shd09cb30b, 32'shd0a5262f, 32'shd0ad9b26, 32'shd0b611f1, 32'shd0be8a8d, 32'shd0c704fd, 32'shd0cf813e, 
               32'shd0d7ff51, 32'shd0e07f36, 32'shd0e900ec, 32'shd0f18472, 32'shd0fa09c9, 32'shd10290f0, 32'shd10b19e7, 32'shd113a4ad, 
               32'shd11c3142, 32'shd124bfa6, 32'shd12d4fd9, 32'shd135e1d9, 32'shd13e75a8, 32'shd1470b44, 32'shd14fa2ad, 32'shd1583be2, 
               32'shd160d6e5, 32'shd16973b3, 32'shd172124d, 32'shd17ab2b3, 32'shd18354e4, 32'shd18bf8e0, 32'shd1949ea6, 32'shd19d4636, 
               32'shd1a5ef90, 32'shd1ae9ab4, 32'shd1b747a0, 32'shd1bff656, 32'shd1c8a6d4, 32'shd1d1591a, 32'shd1da0d28, 32'shd1e2c2fd, 
               32'shd1eb7a9a, 32'shd1f433fd, 32'shd1fcef27, 32'shd205ac17, 32'shd20e6acc, 32'shd2172b48, 32'shd21fed88, 32'shd228b18d, 
               32'shd2317756, 32'shd23a3ee4, 32'shd2430835, 32'shd24bd34a, 32'shd254a021, 32'shd25d6ebc, 32'shd2663f19, 32'shd26f1138, 
               32'shd277e518, 32'shd280babb, 32'shd289921e, 32'shd2926b41, 32'shd29b4626, 32'shd2a422ca, 32'shd2ad012e, 32'shd2b5e151, 
               32'shd2bec333, 32'shd2c7a6d4, 32'shd2d08c33, 32'shd2d97350, 32'shd2e25c2b, 32'shd2eb46c3, 32'shd2f43318, 32'shd2fd2129, 
               32'shd30610f7, 32'shd30f0280, 32'shd317f5c6, 32'shd320eac6, 32'shd329e181, 32'shd332d9f7, 32'shd33bd427, 32'shd344d011, 
               32'shd34dcdb4, 32'shd356cd11, 32'shd35fce26, 32'shd368d0f3, 32'shd371d579, 32'shd37adbb6, 32'shd383e3ab, 32'shd38ced57, 
               32'shd395f8ba, 32'shd39f05d3, 32'shd3a814a2, 32'shd3b12526, 32'shd3ba3760, 32'shd3c34b4f, 32'shd3cc60f2, 32'shd3d5784a, 
               32'shd3de9156, 32'shd3e7ac15, 32'shd3f0c887, 32'shd3f9e6ad, 32'shd4030684, 32'shd40c280e, 32'shd4154b4a, 32'shd41e7037, 
               32'shd42796d5, 32'shd430bf24, 32'shd439e923, 32'shd44314d3, 32'shd44c4232, 32'shd4557140, 32'shd45ea1fd, 32'shd467d469, 
               32'shd4710883, 32'shd47a3e4b, 32'shd48375c1, 32'shd48caee4, 32'shd495e9b3, 32'shd49f2630, 32'shd4a86458, 32'shd4b1a42c, 
               32'shd4bae5ab, 32'shd4c428d6, 32'shd4cd6dab, 32'shd4d6b42b, 32'shd4dffc54, 32'shd4e94627, 32'shd4f291a4, 32'shd4fbdec9, 
               32'shd5052d97, 32'shd50e7e0d, 32'shd517d02b, 32'shd52123f0, 32'shd52a795d, 32'shd533d070, 32'shd53d292a, 32'shd5468389, 
               32'shd54fdf8f, 32'shd5593d3a, 32'shd5629c89, 32'shd56bfd7d, 32'shd5756016, 32'shd57ec452, 32'shd5882a32, 32'shd59191b5, 
               32'shd59afadb, 32'shd5a465a3, 32'shd5add20d, 32'shd5b74019, 32'shd5c0afc6, 32'shd5ca2115, 32'shd5d39403, 32'shd5dd0892, 
               32'shd5e67ec1, 32'shd5eff690, 32'shd5f96ffd, 32'shd602eb0a, 32'shd60c67b4, 32'shd615e5fd, 32'shd61f65e4, 32'shd628e767, 
               32'shd6326a88, 32'shd63bef46, 32'shd645759f, 32'shd64efd94, 32'shd6588725, 32'shd6621251, 32'shd66b9f18, 32'shd6752d79, 
               32'shd67ebd74, 32'shd6884f09, 32'shd691e237, 32'shd69b76fe, 32'shd6a50d5d, 32'shd6aea555, 32'shd6b83ee4, 32'shd6c1da0b, 
               32'shd6cb76c9, 32'shd6d5151d, 32'shd6deb508, 32'shd6e85689, 32'shd6f1f99f, 32'shd6fb9e4b, 32'shd705448b, 32'shd70eec60, 
               32'shd71895c9, 32'shd72240c5, 32'shd72bed55, 32'shd7359b78, 32'shd73f4b2e, 32'shd748fc75, 32'shd752af4f, 32'shd75c63ba, 
               32'shd76619b6, 32'shd76fd143, 32'shd7798a60, 32'shd783450d, 32'shd78d014a, 32'shd796bf16, 32'shd7a07e70, 32'shd7aa3f5a, 
               32'shd7b401d1, 32'shd7bdc5d6, 32'shd7c78b68, 32'shd7d15288, 32'shd7db1b34, 32'shd7e4e56c, 32'shd7eeb130, 32'shd7f87e7f, 
               32'shd8024d59, 32'shd80c1dbf, 32'shd815efae, 32'shd81fc328, 32'shd829982b, 32'shd8336eb7, 32'shd83d46cc, 32'shd8472069, 
               32'shd850fb8e, 32'shd85ad83c, 32'shd864b670, 32'shd86e962b, 32'shd878776d, 32'shd8825a35, 32'shd88c3e83, 32'shd8962456, 
               32'shd8a00bae, 32'shd8a9f48a, 32'shd8b3deeb, 32'shd8bdcad0, 32'shd8c7b838, 32'shd8d1a724, 32'shd8db9792, 32'shd8e58982, 
               32'shd8ef7cf4, 32'shd8f971e8, 32'shd903685d, 32'shd90d6053, 32'shd91759c9, 32'shd92154bf, 32'shd92b5135, 32'shd9354f2a, 
               32'shd93f4e9e, 32'shd9494f90, 32'shd9535201, 32'shd95d55ef, 32'shd9675b5a, 32'shd9716243, 32'shd97b6aa8, 32'shd9857489, 
               32'shd98f7fe6, 32'shd9998cbe, 32'shd9a39b11, 32'shd9adaadf, 32'shd9b7bc27, 32'shd9c1cee9, 32'shd9cbe325, 32'shd9d5f8d9, 
               32'shd9e01006, 32'shd9ea28ac, 32'shd9f442c9, 32'shd9fe5e5e, 32'shda087b69, 32'shda1299ec, 32'shda1cb9e5, 32'shda26db54, 
               32'shda30fe38, 32'shda3b2292, 32'shda454860, 32'shda4f6fa3, 32'shda599859, 32'shda63c284, 32'shda6dee21, 32'shda781b31, 
               32'shda8249b4, 32'shda8c79a9, 32'shda96ab0f, 32'shdaa0dde7, 32'shdaab122f, 32'shdab547e8, 32'shdabf7f11, 32'shdac9b7a9, 
               32'shdad3f1b1, 32'shdade2d28, 32'shdae86a0d, 32'shdaf2a860, 32'shdafce821, 32'shdb072950, 32'shdb116beb, 32'shdb1baff2, 
               32'shdb25f566, 32'shdb303c46, 32'shdb3a8491, 32'shdb44ce46, 32'shdb4f1967, 32'shdb5965f1, 32'shdb63b3e5, 32'shdb6e0342, 
               32'shdb785409, 32'shdb82a638, 32'shdb8cf9cf, 32'shdb974ece, 32'shdba1a534, 32'shdbabfd01, 32'shdbb65634, 32'shdbc0b0ce, 
               32'shdbcb0cce, 32'shdbd56a32, 32'shdbdfc8fc, 32'shdbea292b, 32'shdbf48abd, 32'shdbfeedb3, 32'shdc09520d, 32'shdc13b7c9, 
               32'shdc1e1ee9, 32'shdc28876a, 32'shdc32f14d, 32'shdc3d5c91, 32'shdc47c936, 32'shdc52373c, 32'shdc5ca6a2, 32'shdc671768, 
               32'shdc71898d, 32'shdc7bfd11, 32'shdc8671f3, 32'shdc90e834, 32'shdc9b5fd2, 32'shdca5d8cd, 32'shdcb05326, 32'shdcbacedb, 
               32'shdcc54bec, 32'shdccfca59, 32'shdcda4a21, 32'shdce4cb44, 32'shdcef4dc2, 32'shdcf9d199, 32'shdd0456ca, 32'shdd0edd55, 
               32'shdd196538, 32'shdd23ee74, 32'shdd2e7908, 32'shdd3904f4, 32'shdd439236, 32'shdd4e20d0, 32'shdd58b0c0, 32'shdd634206, 
               32'shdd6dd4a2, 32'shdd786892, 32'shdd82fdd8, 32'shdd8d9472, 32'shdd982c60, 32'shdda2c5a2, 32'shddad6036, 32'shddb7fc1e, 
               32'shddc29958, 32'shddcd37e4, 32'shddd7d7c1, 32'shdde278ef, 32'shdded1b6e, 32'shddf7bf3e, 32'shde02645d, 32'shde0d0acc, 
               32'shde17b28a, 32'shde225b96, 32'shde2d05f1, 32'shde37b199, 32'shde425e8f, 32'shde4d0cd2, 32'shde57bc62, 32'shde626d3e, 
               32'shde6d1f65, 32'shde77d2d8, 32'shde828796, 32'shde8d3d9e, 32'shde97f4f1, 32'shdea2ad8d, 32'shdead6773, 32'shdeb822a1, 
               32'shdec2df18, 32'shdecd9cd7, 32'shded85bdd, 32'shdee31c2b, 32'shdeedddc0, 32'shdef8a09b, 32'shdf0364bc, 32'shdf0e2a22, 
               32'shdf18f0ce, 32'shdf23b8be, 32'shdf2e81f3, 32'shdf394c6b, 32'shdf441828, 32'shdf4ee527, 32'shdf59b369, 32'shdf6482ed, 
               32'shdf6f53b3, 32'shdf7a25ba, 32'shdf84f902, 32'shdf8fcd8b, 32'shdf9aa354, 32'shdfa57a5d, 32'shdfb052a5, 32'shdfbb2c2c, 
               32'shdfc606f1, 32'shdfd0e2f5, 32'shdfdbc036, 32'shdfe69eb4, 32'shdff17e70, 32'shdffc5f67, 32'she007419b, 32'she012250a, 
               32'she01d09b4, 32'she027ef99, 32'she032d6b8, 32'she03dbf11, 32'she048a8a4, 32'she053936f, 32'she05e7f74, 32'she0696cb0, 
               32'she0745b24, 32'she07f4acf, 32'she08a3bb2, 32'she0952dcb, 32'she0a0211a, 32'she0ab159e, 32'she0b60b58, 32'she0c10247, 
               32'she0cbfa6a, 32'she0d6f3c1, 32'she0e1ee4b, 32'she0ecea09, 32'she0f7e6f9, 32'she102e51c, 32'she10de470, 32'she118e4f6, 
               32'she123e6ad, 32'she12ee995, 32'she139edac, 32'she144f2f3, 32'she14ff96a, 32'she15b0110, 32'she16609e3, 32'she17113e5, 
               32'she17c1f15, 32'she1872b72, 32'she19238fb, 32'she19d47b1, 32'she1a85793, 32'she1b368a0, 32'she1be7ad8, 32'she1c98e3b, 
               32'she1d4a2c8, 32'she1dfb87f, 32'she1eacf5f, 32'she1f5e768, 32'she2010099, 32'she20c1af3, 32'she2173674, 32'she222531c, 
               32'she22d70eb, 32'she2388fe1, 32'she243affc, 32'she24ed13d, 32'she259f3a3, 32'she265172e, 32'she2703bdc, 32'she27b61af, 
               32'she28688a4, 32'she291b0bd, 32'she29cd9f8, 32'she2a80456, 32'she2b32fd4, 32'she2be5c74, 32'she2c98a35, 32'she2d4b916, 
               32'she2dfe917, 32'she2eb1a37, 32'she2f64c77, 32'she3017fd5, 32'she30cb451, 32'she317e9eb, 32'she32320a2, 32'she32e5876, 
               32'she3399167, 32'she344cb73, 32'she350069b, 32'she35b42df, 32'she366803c, 32'she371beb5, 32'she37cfe47, 32'she3883ef2, 
               32'she39380b6, 32'she39ec393, 32'she3aa0788, 32'she3b54c95, 32'she3c092b9, 32'she3cbd9f4, 32'she3d72245, 32'she3e26bac, 
               32'she3edb628, 32'she3f901ba, 32'she4044e60, 32'she40f9c1a, 32'she41aeae8, 32'she4263ac9, 32'she4318bbe, 32'she43cddc4, 
               32'she44830dd, 32'she4538507, 32'she45eda43, 32'she46a308f, 32'she47587eb, 32'she480e057, 32'she48c39d3, 32'she497945d, 
               32'she4a2eff6, 32'she4ae4c9d, 32'she4b9aa52, 32'she4c50914, 32'she4d068e2, 32'she4dbc9bd, 32'she4e72ba4, 32'she4f28e96, 
               32'she4fdf294, 32'she509579b, 32'she514bdad, 32'she52024c9, 32'she52b8cee, 32'she536f61b, 32'she5426051, 32'she54dcb8f, 
               32'she55937d5, 32'she564a521, 32'she5701374, 32'she57b82cd, 32'she586f32c, 32'she5926490, 32'she59dd6f9, 32'she5a94a67, 
               32'she5b4bed8, 32'she5c0344d, 32'she5cbaac5, 32'she5d72240, 32'she5e29abc, 32'she5ee143b, 32'she5f98ebb, 32'she6050a3b, 
               32'she61086bc, 32'she61c043d, 32'she62782be, 32'she633023e, 32'she63e82bc, 32'she64a0438, 32'she65586b3, 32'she6610a2a, 
               32'she66c8e9f, 32'she6781410, 32'she6839a7c, 32'she68f21e5, 32'she69aaa48, 32'she6a633a6, 32'she6b1bdff, 32'she6bd4951, 
               32'she6c8d59c, 32'she6d462e1, 32'she6dff11d, 32'she6eb8052, 32'she6f7107e, 32'she702a1a1, 32'she70e33bb, 32'she719c6cb, 
               32'she7255ad1, 32'she730efcc, 32'she73c85bc, 32'she7481ca1, 32'she753b479, 32'she75f4d45, 32'she76ae704, 32'she77681b6, 
               32'she7821d59, 32'she78db9ef, 32'she7995776, 32'she7a4f5ed, 32'she7b09555, 32'she7bc35ad, 32'she7c7d6f4, 32'she7d3792b, 
               32'she7df1c50, 32'she7eac063, 32'she7f66564, 32'she8020b52, 32'she80db22d, 32'she81959f4, 32'she82502a7, 32'she830ac45, 
               32'she83c56cf, 32'she8480243, 32'she853aea1, 32'she85f5be9, 32'she86b0a1a, 32'she876b934, 32'she8826936, 32'she88e1a20, 
               32'she899cbf1, 32'she8a57ea9, 32'she8b13248, 32'she8bce6cd, 32'she8c89c37, 32'she8d45286, 32'she8e009ba, 32'she8ebc1d3, 
               32'she8f77acf, 32'she90334af, 32'she90eef71, 32'she91aab16, 32'she926679c, 32'she9322505, 32'she93de34e, 32'she949a278, 
               32'she9556282, 32'she961236c, 32'she96ce535, 32'she978a7dd, 32'she9846b63, 32'she9902fc7, 32'she99bf509, 32'she9a7bb28, 
               32'she9b38223, 32'she9bf49fa, 32'she9cb12ad, 32'she9d6dc3b, 32'she9e2a6a3, 32'she9ee71e6, 32'she9fa3e03, 32'shea060af9, 
               32'shea11d8c8, 32'shea1da770, 32'shea2976ef, 32'shea354746, 32'shea411874, 32'shea4cea79, 32'shea58bd54, 32'shea649105, 
               32'shea70658a, 32'shea7c3ae5, 32'shea881114, 32'shea93e817, 32'shea9fbfed, 32'sheaab9896, 32'sheab77212, 32'sheac34c60, 
               32'sheacf277f, 32'sheadb0370, 32'sheae6e031, 32'sheaf2bdc3, 32'sheafe9c24, 32'sheb0a7b54, 32'sheb165b54, 32'sheb223c22, 
               32'sheb2e1dbe, 32'sheb3a0027, 32'sheb45e35d, 32'sheb51c760, 32'sheb5dac2f, 32'sheb6991ca, 32'sheb75782f, 32'sheb815f60, 
               32'sheb8d475b, 32'sheb99301f, 32'sheba519ad, 32'shebb10404, 32'shebbcef23, 32'shebc8db0b, 32'shebd4c7ba, 32'shebe0b52f, 
               32'shebeca36c, 32'shebf8926f, 32'shec048237, 32'shec1072c4, 32'shec1c6417, 32'shec28562d, 32'shec344908, 32'shec403ca5, 
               32'shec4c3106, 32'shec582629, 32'shec641c0e, 32'shec7012b5, 32'shec7c0a1d, 32'shec880245, 32'shec93fb2e, 32'shec9ff4d6, 
               32'shecabef3d, 32'shecb7ea63, 32'shecc3e648, 32'sheccfe2ea, 32'shecdbe04a, 32'shece7de66, 32'shecf3dd3f, 32'shecffdcd4, 
               32'shed0bdd25, 32'shed17de31, 32'shed23dff7, 32'shed2fe277, 32'shed3be5b1, 32'shed47e9a5, 32'shed53ee51, 32'shed5ff3b5, 
               32'shed6bf9d1, 32'shed7800a5, 32'shed84082f, 32'shed901070, 32'shed9c1967, 32'sheda82313, 32'shedb42d74, 32'shedc0388a, 
               32'shedcc4454, 32'shedd850d2, 32'shede45e03, 32'shedf06be6, 32'shedfc7a7c, 32'shee0889c4, 32'shee1499bd, 32'shee20aa67, 
               32'shee2cbbc1, 32'shee38cdcb, 32'shee44e084, 32'shee50f3ed, 32'shee5d0804, 32'shee691cc9, 32'shee75323c, 32'shee81485c, 
               32'shee8d5f29, 32'shee9976a1, 32'sheea58ec6, 32'sheeb1a796, 32'sheebdc110, 32'sheec9db35, 32'sheed5f604, 32'sheee2117c, 
               32'sheeee2d9d, 32'sheefa4a67, 32'shef0667d9, 32'shef1285f2, 32'shef1ea4b2, 32'shef2ac419, 32'shef36e426, 32'shef4304d8, 
               32'shef4f2630, 32'shef5b482d, 32'shef676ace, 32'shef738e12, 32'shef7fb1fa, 32'shef8bd685, 32'shef97fbb2, 32'shefa42181, 
               32'shefb047f2, 32'shefbc6f03, 32'shefc896b5, 32'shefd4bf08, 32'shefe0e7f9, 32'shefed118a, 32'sheff93bba, 32'shf0056687, 
               32'shf01191f3, 32'shf01dbdfb, 32'shf029eaa1, 32'shf03617e2, 32'shf04245c0, 32'shf04e7438, 32'shf05aa34c, 32'shf066d2fa, 
               32'shf0730342, 32'shf07f3424, 32'shf08b659f, 32'shf09797b2, 32'shf0a3ca5d, 32'shf0affda0, 32'shf0bc317a, 32'shf0c865ea, 
               32'shf0d49af1, 32'shf0e0d08d, 32'shf0ed06bf, 32'shf0f93d86, 32'shf10574e0, 32'shf111accf, 32'shf11de551, 32'shf12a1e66, 
               32'shf136580d, 32'shf1429247, 32'shf14ecd11, 32'shf15b086d, 32'shf1674459, 32'shf17380d6, 32'shf17fbde2, 32'shf18bfb7d, 
               32'shf19839a6, 32'shf1a4785e, 32'shf1b0b7a4, 32'shf1bcf777, 32'shf1c937d6, 32'shf1d578c2, 32'shf1e1ba3a, 32'shf1edfc3d, 
               32'shf1fa3ecb, 32'shf20681e3, 32'shf212c585, 32'shf21f09b1, 32'shf22b4e66, 32'shf23793a3, 32'shf243d968, 32'shf2501fb5, 
               32'shf25c6688, 32'shf268ade3, 32'shf274f5c3, 32'shf2813e2a, 32'shf28d8715, 32'shf299d085, 32'shf2a61a7a, 32'shf2b264f2, 
               32'shf2beafed, 32'shf2cafb6b, 32'shf2d7476c, 32'shf2e393ef, 32'shf2efe0f2, 32'shf2fc2e77, 32'shf3087c7d, 32'shf314cb02, 
               32'shf3211a07, 32'shf32d698a, 32'shf339b98d, 32'shf3460a0d, 32'shf3525b0b, 32'shf35eac86, 32'shf36afe7e, 32'shf37750f2, 
               32'shf383a3e2, 32'shf38ff74d, 32'shf39c4b32, 32'shf3a89f92, 32'shf3b4f46c, 32'shf3c149bf, 32'shf3cd9f8b, 32'shf3d9f5cf, 
               32'shf3e64c8c, 32'shf3f2a3bf, 32'shf3fefb6a, 32'shf40b538b, 32'shf417ac22, 32'shf424052f, 32'shf4305eb0, 32'shf43cb8a7, 
               32'shf4491311, 32'shf4556def, 32'shf461c940, 32'shf46e2504, 32'shf47a8139, 32'shf486dde1, 32'shf4933afa, 32'shf49f9884, 
               32'shf4abf67e, 32'shf4b854e7, 32'shf4c4b3c0, 32'shf4d11308, 32'shf4dd72be, 32'shf4e9d2e3, 32'shf4f63374, 32'shf5029473, 
               32'shf50ef5de, 32'shf51b57b5, 32'shf527b9f7, 32'shf5341ca5, 32'shf5407fbd, 32'shf54ce33f, 32'shf559472b, 32'shf565ab80, 
               32'shf572103d, 32'shf57e7563, 32'shf58adaf0, 32'shf59740e5, 32'shf5a3a740, 32'shf5b00e02, 32'shf5bc7529, 32'shf5c8dcb6, 
               32'shf5d544a7, 32'shf5e1acfd, 32'shf5ee15b7, 32'shf5fa7ed4, 32'shf606e854, 32'shf6135237, 32'shf61fbc7b, 32'shf62c2721, 
               32'shf6389228, 32'shf644fd8f, 32'shf6516956, 32'shf65dd57d, 32'shf66a4203, 32'shf676aee8, 32'shf6831c2b, 32'shf68f89cb, 
               32'shf69bf7c9, 32'shf6a86623, 32'shf6b4d4d9, 32'shf6c143ec, 32'shf6cdb359, 32'shf6da2321, 32'shf6e69344, 32'shf6f303c0, 
               32'shf6ff7496, 32'shf70be5c4, 32'shf718574b, 32'shf724c92a, 32'shf7313b60, 32'shf73daded, 32'shf74a20d0, 32'shf756940a, 
               32'shf7630799, 32'shf76f7b7d, 32'shf77befb5, 32'shf7886442, 32'shf794d922, 32'shf7a14e55, 32'shf7adc3db, 32'shf7ba39b3, 
               32'shf7c6afdc, 32'shf7d32657, 32'shf7df9d22, 32'shf7ec143e, 32'shf7f88ba9, 32'shf8050364, 32'shf8117b6d, 32'shf81df3c5, 
               32'shf82a6c6a, 32'shf836e55d, 32'shf8435e9d, 32'shf84fd829, 32'shf85c5201, 32'shf868cc24, 32'shf8754692, 32'shf881c14b, 
               32'shf88e3c4d, 32'shf89ab799, 32'shf8a7332e, 32'shf8b3af0c, 32'shf8c02b31, 32'shf8cca79e, 32'shf8d92452, 32'shf8e5a14d, 
               32'shf8f21e8e, 32'shf8fe9c15, 32'shf90b19e0, 32'shf91797f0, 32'shf9241645, 32'shf93094dd, 32'shf93d13b8, 32'shf94992d7, 
               32'shf9561237, 32'shf96291d9, 32'shf96f11bc, 32'shf97b91e1, 32'shf9881245, 32'shf99492ea, 32'shf9a113cd, 32'shf9ad94f0, 
               32'shf9ba1651, 32'shf9c697f0, 32'shf9d319cc, 32'shf9df9be6, 32'shf9ec1e3b, 32'shf9f8a0cd, 32'shfa05239a, 32'shfa11a6a3, 
               32'shfa1e29e5, 32'shfa2aad62, 32'shfa373119, 32'shfa43b508, 32'shfa503930, 32'shfa5cbd91, 32'shfa694229, 32'shfa75c6f8, 
               32'shfa824bfd, 32'shfa8ed139, 32'shfa9b56ab, 32'shfaa7dc52, 32'shfab4622d, 32'shfac0e83d, 32'shfacd6e81, 32'shfad9f4f8, 
               32'shfae67ba2, 32'shfaf3027e, 32'shfaff898c, 32'shfb0c10cb, 32'shfb18983b, 32'shfb251fdc, 32'shfb31a7ac, 32'shfb3e2fac, 
               32'shfb4ab7db, 32'shfb574039, 32'shfb63c8c4, 32'shfb70517d, 32'shfb7cda63, 32'shfb896375, 32'shfb95ecb4, 32'shfba2761e, 
               32'shfbaeffb3, 32'shfbbb8973, 32'shfbc8135c, 32'shfbd49d70, 32'shfbe127ac, 32'shfbedb212, 32'shfbfa3c9f, 32'shfc06c754, 
               32'shfc135231, 32'shfc1fdd34, 32'shfc2c685d, 32'shfc38f3ac, 32'shfc457f21, 32'shfc520aba, 32'shfc5e9678, 32'shfc6b2259, 
               32'shfc77ae5e, 32'shfc843a85, 32'shfc90c6cf, 32'shfc9d533b, 32'shfca9dfc8, 32'shfcb66c77, 32'shfcc2f945, 32'shfccf8634, 
               32'shfcdc1342, 32'shfce8a06f, 32'shfcf52dbb, 32'shfd01bb24, 32'shfd0e48ab, 32'shfd1ad650, 32'shfd276410, 32'shfd33f1ed, 
               32'shfd407fe6, 32'shfd4d0df9, 32'shfd599c28, 32'shfd662a70, 32'shfd72b8d2, 32'shfd7f474d, 32'shfd8bd5e1, 32'shfd98648d, 
               32'shfda4f351, 32'shfdb1822c, 32'shfdbe111e, 32'shfdcaa027, 32'shfdd72f45, 32'shfde3be78, 32'shfdf04dc0, 32'shfdfcdd1d, 
               32'shfe096c8d, 32'shfe15fc11, 32'shfe228ba7, 32'shfe2f1b50, 32'shfe3bab0b, 32'shfe483ad8, 32'shfe54cab5, 32'shfe615aa3, 
               32'shfe6deaa1, 32'shfe7a7aae, 32'shfe870aca, 32'shfe939af5, 32'shfea02b2e, 32'shfeacbb74, 32'shfeb94bc8, 32'shfec5dc28, 
               32'shfed26c94, 32'shfedefd0c, 32'shfeeb8d8f, 32'shfef81e1d, 32'shff04aeb5, 32'shff113f56, 32'shff1dd001, 32'shff2a60b4, 
               32'shff36f170, 32'shff438234, 32'shff5012fe, 32'shff5ca3d0, 32'shff6934a8, 32'shff75c585, 32'shff825668, 32'shff8ee750, 
               32'shff9b783c, 32'shffa8092c, 32'shffb49a1f, 32'shffc12b16, 32'shffcdbc0f, 32'shffda4d09, 32'shffe6de05, 32'shfff36f02
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 14)
         begin
            reg signed [31:0] W_Re_table[8192] = '{
               32'sh40000000, 32'sh3fffffb1, 32'sh3ffffec4, 32'sh3ffffd39, 32'sh3ffffb11, 32'sh3ffff84a, 32'sh3ffff4e6, 32'sh3ffff0e3, 
               32'sh3fffec43, 32'sh3fffe705, 32'sh3fffe128, 32'sh3fffdaae, 32'sh3fffd396, 32'sh3fffcbe0, 32'sh3fffc38c, 32'sh3fffba9b, 
               32'sh3fffb10b, 32'sh3fffa6de, 32'sh3fff9c12, 32'sh3fff90a9, 32'sh3fff84a1, 32'sh3fff77fc, 32'sh3fff6ab9, 32'sh3fff5cd8, 
               32'sh3fff4e59, 32'sh3fff3f3c, 32'sh3fff2f82, 32'sh3fff1f29, 32'sh3fff0e32, 32'sh3ffefc9e, 32'sh3ffeea6c, 32'sh3ffed79b, 
               32'sh3ffec42d, 32'sh3ffeb021, 32'sh3ffe9b77, 32'sh3ffe862f, 32'sh3ffe704a, 32'sh3ffe59c6, 32'sh3ffe42a4, 32'sh3ffe2ae5, 
               32'sh3ffe1288, 32'sh3ffdf98c, 32'sh3ffddff3, 32'sh3ffdc5bc, 32'sh3ffdaae7, 32'sh3ffd8f74, 32'sh3ffd7364, 32'sh3ffd56b5, 
               32'sh3ffd3969, 32'sh3ffd1b7e, 32'sh3ffcfcf6, 32'sh3ffcddd0, 32'sh3ffcbe0c, 32'sh3ffc9daa, 32'sh3ffc7caa, 32'sh3ffc5b0c, 
               32'sh3ffc38d1, 32'sh3ffc15f7, 32'sh3ffbf280, 32'sh3ffbce6b, 32'sh3ffba9b8, 32'sh3ffb8467, 32'sh3ffb5e78, 32'sh3ffb37ec, 
               32'sh3ffb10c1, 32'sh3ffae8f9, 32'sh3ffac092, 32'sh3ffa978e, 32'sh3ffa6dec, 32'sh3ffa43ac, 32'sh3ffa18cf, 32'sh3ff9ed53, 
               32'sh3ff9c13a, 32'sh3ff99483, 32'sh3ff9672d, 32'sh3ff9393a, 32'sh3ff90aaa, 32'sh3ff8db7b, 32'sh3ff8abae, 32'sh3ff87b44, 
               32'sh3ff84a3c, 32'sh3ff81896, 32'sh3ff7e652, 32'sh3ff7b370, 32'sh3ff77ff1, 32'sh3ff74bd3, 32'sh3ff71718, 32'sh3ff6e1bf, 
               32'sh3ff6abc8, 32'sh3ff67534, 32'sh3ff63e01, 32'sh3ff60631, 32'sh3ff5cdc3, 32'sh3ff594b7, 32'sh3ff55b0d, 32'sh3ff520c5, 
               32'sh3ff4e5e0, 32'sh3ff4aa5d, 32'sh3ff46e3c, 32'sh3ff4317d, 32'sh3ff3f420, 32'sh3ff3b626, 32'sh3ff3778e, 32'sh3ff33858, 
               32'sh3ff2f884, 32'sh3ff2b813, 32'sh3ff27703, 32'sh3ff23556, 32'sh3ff1f30b, 32'sh3ff1b022, 32'sh3ff16c9c, 32'sh3ff12878, 
               32'sh3ff0e3b6, 32'sh3ff09e56, 32'sh3ff05858, 32'sh3ff011bd, 32'sh3fefca84, 32'sh3fef82ad, 32'sh3fef3a39, 32'sh3feef126, 
               32'sh3feea776, 32'sh3fee5d28, 32'sh3fee123d, 32'sh3fedc6b4, 32'sh3fed7a8c, 32'sh3fed2dc8, 32'sh3fece065, 32'sh3fec9265, 
               32'sh3fec43c7, 32'sh3febf48b, 32'sh3feba4b2, 32'sh3feb543b, 32'sh3feb0326, 32'sh3feab173, 32'sh3fea5f23, 32'sh3fea0c35, 
               32'sh3fe9b8a9, 32'sh3fe96480, 32'sh3fe90fb9, 32'sh3fe8ba54, 32'sh3fe86452, 32'sh3fe80db2, 32'sh3fe7b674, 32'sh3fe75e98, 
               32'sh3fe7061f, 32'sh3fe6ad08, 32'sh3fe65354, 32'sh3fe5f902, 32'sh3fe59e12, 32'sh3fe54284, 32'sh3fe4e659, 32'sh3fe48990, 
               32'sh3fe42c2a, 32'sh3fe3ce26, 32'sh3fe36f84, 32'sh3fe31045, 32'sh3fe2b067, 32'sh3fe24fed, 32'sh3fe1eed5, 32'sh3fe18d1f, 
               32'sh3fe12acb, 32'sh3fe0c7da, 32'sh3fe0644b, 32'sh3fe0001f, 32'sh3fdf9b55, 32'sh3fdf35ed, 32'sh3fdecfe8, 32'sh3fde6945, 
               32'sh3fde0205, 32'sh3fdd9a27, 32'sh3fdd31ac, 32'sh3fdcc892, 32'sh3fdc5edc, 32'sh3fdbf488, 32'sh3fdb8996, 32'sh3fdb1e06, 
               32'sh3fdab1d9, 32'sh3fda450f, 32'sh3fd9d7a7, 32'sh3fd969a1, 32'sh3fd8fafe, 32'sh3fd88bbe, 32'sh3fd81bdf, 32'sh3fd7ab64, 
               32'sh3fd73a4a, 32'sh3fd6c894, 32'sh3fd6563f, 32'sh3fd5e34e, 32'sh3fd56fbe, 32'sh3fd4fb91, 32'sh3fd486c7, 32'sh3fd4115f, 
               32'sh3fd39b5a, 32'sh3fd324b7, 32'sh3fd2ad77, 32'sh3fd23599, 32'sh3fd1bd1e, 32'sh3fd14405, 32'sh3fd0ca4f, 32'sh3fd04ffc, 
               32'sh3fcfd50b, 32'sh3fcf597c, 32'sh3fcedd50, 32'sh3fce6087, 32'sh3fcde320, 32'sh3fcd651c, 32'sh3fcce67a, 32'sh3fcc673b, 
               32'sh3fcbe75e, 32'sh3fcb66e4, 32'sh3fcae5cd, 32'sh3fca6418, 32'sh3fc9e1c6, 32'sh3fc95ed7, 32'sh3fc8db4a, 32'sh3fc8571f, 
               32'sh3fc7d258, 32'sh3fc74cf3, 32'sh3fc6c6f0, 32'sh3fc64051, 32'sh3fc5b913, 32'sh3fc53139, 32'sh3fc4a8c1, 32'sh3fc41fac, 
               32'sh3fc395f9, 32'sh3fc30baa, 32'sh3fc280bc, 32'sh3fc1f532, 32'sh3fc1690a, 32'sh3fc0dc45, 32'sh3fc04ee3, 32'sh3fbfc0e3, 
               32'sh3fbf3246, 32'sh3fbea30c, 32'sh3fbe1334, 32'sh3fbd82bf, 32'sh3fbcf1ad, 32'sh3fbc5ffe, 32'sh3fbbcdb1, 32'sh3fbb3ac7, 
               32'sh3fbaa740, 32'sh3fba131b, 32'sh3fb97e5a, 32'sh3fb8e8fb, 32'sh3fb852ff, 32'sh3fb7bc65, 32'sh3fb7252f, 32'sh3fb68d5b, 
               32'sh3fb5f4ea, 32'sh3fb55bdc, 32'sh3fb4c231, 32'sh3fb427e8, 32'sh3fb38d02, 32'sh3fb2f17f, 32'sh3fb2555f, 32'sh3fb1b8a2, 
               32'sh3fb11b48, 32'sh3fb07d50, 32'sh3fafdebb, 32'sh3faf3f89, 32'sh3fae9fbb, 32'sh3fadff4e, 32'sh3fad5e45, 32'sh3facbc9f, 
               32'sh3fac1a5b, 32'sh3fab777b, 32'sh3faad3fd, 32'sh3faa2fe2, 32'sh3fa98b2a, 32'sh3fa8e5d5, 32'sh3fa83fe3, 32'sh3fa79954, 
               32'sh3fa6f228, 32'sh3fa64a5f, 32'sh3fa5a1f9, 32'sh3fa4f8f6, 32'sh3fa44f55, 32'sh3fa3a518, 32'sh3fa2fa3d, 32'sh3fa24ec6, 
               32'sh3fa1a2b2, 32'sh3fa0f600, 32'sh3fa048b2, 32'sh3f9f9ac6, 32'sh3f9eec3e, 32'sh3f9e3d19, 32'sh3f9d8d56, 32'sh3f9cdcf7, 
               32'sh3f9c2bfb, 32'sh3f9b7a62, 32'sh3f9ac82c, 32'sh3f9a1558, 32'sh3f9961e8, 32'sh3f98addb, 32'sh3f97f932, 32'sh3f9743eb, 
               32'sh3f968e07, 32'sh3f95d787, 32'sh3f952069, 32'sh3f9468af, 32'sh3f93b058, 32'sh3f92f763, 32'sh3f923dd2, 32'sh3f9183a5, 
               32'sh3f90c8da, 32'sh3f900d72, 32'sh3f8f516e, 32'sh3f8e94cd, 32'sh3f8dd78f, 32'sh3f8d19b4, 32'sh3f8c5b3d, 32'sh3f8b9c28, 
               32'sh3f8adc77, 32'sh3f8a1c29, 32'sh3f895b3e, 32'sh3f8899b7, 32'sh3f87d792, 32'sh3f8714d1, 32'sh3f865174, 32'sh3f858d79, 
               32'sh3f84c8e2, 32'sh3f8403ae, 32'sh3f833ddd, 32'sh3f827770, 32'sh3f81b065, 32'sh3f80e8bf, 32'sh3f80207b, 32'sh3f7f579b, 
               32'sh3f7e8e1e, 32'sh3f7dc405, 32'sh3f7cf94e, 32'sh3f7c2dfc, 32'sh3f7b620c, 32'sh3f7a9580, 32'sh3f79c857, 32'sh3f78fa92, 
               32'sh3f782c30, 32'sh3f775d31, 32'sh3f768d96, 32'sh3f75bd5e, 32'sh3f74ec8a, 32'sh3f741b19, 32'sh3f73490b, 32'sh3f727661, 
               32'sh3f71a31b, 32'sh3f70cf38, 32'sh3f6ffab8, 32'sh3f6f259c, 32'sh3f6e4fe3, 32'sh3f6d798e, 32'sh3f6ca29c, 32'sh3f6bcb0e, 
               32'sh3f6af2e3, 32'sh3f6a1a1c, 32'sh3f6940b8, 32'sh3f6866b8, 32'sh3f678c1c, 32'sh3f66b0e3, 32'sh3f65d50d, 32'sh3f64f89b, 
               32'sh3f641b8d, 32'sh3f633de2, 32'sh3f625f9b, 32'sh3f6180b8, 32'sh3f60a138, 32'sh3f5fc11c, 32'sh3f5ee063, 32'sh3f5dff0e, 
               32'sh3f5d1d1d, 32'sh3f5c3a8f, 32'sh3f5b5765, 32'sh3f5a739e, 32'sh3f598f3c, 32'sh3f58aa3d, 32'sh3f57c4a2, 32'sh3f56de6a, 
               32'sh3f55f796, 32'sh3f551026, 32'sh3f54281a, 32'sh3f533f71, 32'sh3f52562c, 32'sh3f516c4b, 32'sh3f5081cd, 32'sh3f4f96b4, 
               32'sh3f4eaafe, 32'sh3f4dbeac, 32'sh3f4cd1be, 32'sh3f4be433, 32'sh3f4af60d, 32'sh3f4a074a, 32'sh3f4917eb, 32'sh3f4827f0, 
               32'sh3f473759, 32'sh3f464626, 32'sh3f455456, 32'sh3f4461eb, 32'sh3f436ee3, 32'sh3f427b3f, 32'sh3f4186ff, 32'sh3f409223, 
               32'sh3f3f9cab, 32'sh3f3ea697, 32'sh3f3dafe7, 32'sh3f3cb89b, 32'sh3f3bc0b3, 32'sh3f3ac82f, 32'sh3f39cf0e, 32'sh3f38d552, 
               32'sh3f37dafa, 32'sh3f36e006, 32'sh3f35e476, 32'sh3f34e849, 32'sh3f33eb81, 32'sh3f32ee1d, 32'sh3f31f01d, 32'sh3f30f181, 
               32'sh3f2ff24a, 32'sh3f2ef276, 32'sh3f2df206, 32'sh3f2cf0fb, 32'sh3f2bef53, 32'sh3f2aed10, 32'sh3f29ea31, 32'sh3f28e6b6, 
               32'sh3f27e29f, 32'sh3f26ddec, 32'sh3f25d89e, 32'sh3f24d2b4, 32'sh3f23cc2e, 32'sh3f22c50c, 32'sh3f21bd4e, 32'sh3f20b4f5, 
               32'sh3f1fabff, 32'sh3f1ea26e, 32'sh3f1d9842, 32'sh3f1c8d79, 32'sh3f1b8215, 32'sh3f1a7615, 32'sh3f19697a, 32'sh3f185c43, 
               32'sh3f174e70, 32'sh3f164001, 32'sh3f1530f7, 32'sh3f142151, 32'sh3f13110f, 32'sh3f120032, 32'sh3f10eeb9, 32'sh3f0fdca5, 
               32'sh3f0ec9f5, 32'sh3f0db6a9, 32'sh3f0ca2c2, 32'sh3f0b8e3f, 32'sh3f0a7921, 32'sh3f096367, 32'sh3f084d12, 32'sh3f073621, 
               32'sh3f061e95, 32'sh3f05066d, 32'sh3f03eda9, 32'sh3f02d44a, 32'sh3f01ba50, 32'sh3f009fba, 32'sh3eff8489, 32'sh3efe68bc, 
               32'sh3efd4c54, 32'sh3efc2f50, 32'sh3efb11b1, 32'sh3ef9f377, 32'sh3ef8d4a1, 32'sh3ef7b530, 32'sh3ef69523, 32'sh3ef5747b, 
               32'sh3ef45338, 32'sh3ef3315a, 32'sh3ef20ee0, 32'sh3ef0ebcb, 32'sh3eefc81a, 32'sh3eeea3ce, 32'sh3eed7ee7, 32'sh3eec5965, 
               32'sh3eeb3347, 32'sh3eea0c8e, 32'sh3ee8e53a, 32'sh3ee7bd4b, 32'sh3ee694c1, 32'sh3ee56b9b, 32'sh3ee441da, 32'sh3ee3177e, 
               32'sh3ee1ec87, 32'sh3ee0c0f4, 32'sh3edf94c7, 32'sh3ede67fe, 32'sh3edd3a9a, 32'sh3edc0c9b, 32'sh3edade01, 32'sh3ed9aecc, 
               32'sh3ed87efc, 32'sh3ed74e91, 32'sh3ed61d8a, 32'sh3ed4ebe9, 32'sh3ed3b9ad, 32'sh3ed286d5, 32'sh3ed15363, 32'sh3ed01f55, 
               32'sh3eceeaad, 32'sh3ecdb56a, 32'sh3ecc7f8b, 32'sh3ecb4912, 32'sh3eca11fe, 32'sh3ec8da4f, 32'sh3ec7a205, 32'sh3ec66920, 
               32'sh3ec52fa0, 32'sh3ec3f585, 32'sh3ec2bad0, 32'sh3ec17f7f, 32'sh3ec04394, 32'sh3ebf070e, 32'sh3ebdc9ed, 32'sh3ebc8c31, 
               32'sh3ebb4ddb, 32'sh3eba0ee9, 32'sh3eb8cf5d, 32'sh3eb78f36, 32'sh3eb64e75, 32'sh3eb50d18, 32'sh3eb3cb21, 32'sh3eb2888f, 
               32'sh3eb14563, 32'sh3eb0019c, 32'sh3eaebd3a, 32'sh3ead783d, 32'sh3eac32a6, 32'sh3eaaec74, 32'sh3ea9a5a8, 32'sh3ea85e41, 
               32'sh3ea7163f, 32'sh3ea5cda3, 32'sh3ea4846c, 32'sh3ea33a9b, 32'sh3ea1f02f, 32'sh3ea0a529, 32'sh3e9f5988, 32'sh3e9e0d4c, 
               32'sh3e9cc076, 32'sh3e9b7306, 32'sh3e9a24fb, 32'sh3e98d655, 32'sh3e978715, 32'sh3e96373b, 32'sh3e94e6c6, 32'sh3e9395b7, 
               32'sh3e92440d, 32'sh3e90f1ca, 32'sh3e8f9eeb, 32'sh3e8e4b72, 32'sh3e8cf75f, 32'sh3e8ba2b2, 32'sh3e8a4d6a, 32'sh3e88f788, 
               32'sh3e87a10c, 32'sh3e8649f5, 32'sh3e84f245, 32'sh3e8399f9, 32'sh3e824114, 32'sh3e80e794, 32'sh3e7f8d7b, 32'sh3e7e32c6, 
               32'sh3e7cd778, 32'sh3e7b7b90, 32'sh3e7a1f0d, 32'sh3e78c1f0, 32'sh3e77643a, 32'sh3e7605e9, 32'sh3e74a6fd, 32'sh3e734778, 
               32'sh3e71e759, 32'sh3e70869f, 32'sh3e6f254c, 32'sh3e6dc35e, 32'sh3e6c60d7, 32'sh3e6afdb5, 32'sh3e6999fa, 32'sh3e6835a4, 
               32'sh3e66d0b4, 32'sh3e656b2b, 32'sh3e640507, 32'sh3e629e4a, 32'sh3e6136f3, 32'sh3e5fcf01, 32'sh3e5e6676, 32'sh3e5cfd51, 
               32'sh3e5b9392, 32'sh3e5a2939, 32'sh3e58be47, 32'sh3e5752ba, 32'sh3e55e694, 32'sh3e5479d4, 32'sh3e530c7a, 32'sh3e519e86, 
               32'sh3e502ff9, 32'sh3e4ec0d1, 32'sh3e4d5110, 32'sh3e4be0b6, 32'sh3e4a6fc1, 32'sh3e48fe33, 32'sh3e478c0b, 32'sh3e46194a, 
               32'sh3e44a5ef, 32'sh3e4331fa, 32'sh3e41bd6c, 32'sh3e404844, 32'sh3e3ed282, 32'sh3e3d5c27, 32'sh3e3be532, 32'sh3e3a6da4, 
               32'sh3e38f57c, 32'sh3e377cbb, 32'sh3e360360, 32'sh3e34896c, 32'sh3e330ede, 32'sh3e3193b7, 32'sh3e3017f6, 32'sh3e2e9b9c, 
               32'sh3e2d1ea8, 32'sh3e2ba11b, 32'sh3e2a22f4, 32'sh3e28a435, 32'sh3e2724db, 32'sh3e25a4e9, 32'sh3e24245d, 32'sh3e22a338, 
               32'sh3e212179, 32'sh3e1f9f21, 32'sh3e1e1c30, 32'sh3e1c98a6, 32'sh3e1b1482, 32'sh3e198fc5, 32'sh3e180a6f, 32'sh3e168480, 
               32'sh3e14fdf7, 32'sh3e1376d5, 32'sh3e11ef1b, 32'sh3e1066c7, 32'sh3e0eddd9, 32'sh3e0d5453, 32'sh3e0bca34, 32'sh3e0a3f7b, 
               32'sh3e08b42a, 32'sh3e07283f, 32'sh3e059bbb, 32'sh3e040e9f, 32'sh3e0280e9, 32'sh3e00f29a, 32'sh3dff63b2, 32'sh3dfdd432, 
               32'sh3dfc4418, 32'sh3dfab365, 32'sh3df9221a, 32'sh3df79036, 32'sh3df5fdb8, 32'sh3df46aa2, 32'sh3df2d6f3, 32'sh3df142ab, 
               32'sh3defadca, 32'sh3dee1851, 32'sh3dec823e, 32'sh3deaeb93, 32'sh3de9544f, 32'sh3de7bc72, 32'sh3de623fd, 32'sh3de48aef, 
               32'sh3de2f148, 32'sh3de15708, 32'sh3ddfbc30, 32'sh3dde20bf, 32'sh3ddc84b5, 32'sh3ddae813, 32'sh3dd94ad8, 32'sh3dd7ad05, 
               32'sh3dd60e99, 32'sh3dd46f94, 32'sh3dd2cff7, 32'sh3dd12fc1, 32'sh3dcf8ef3, 32'sh3dcded8c, 32'sh3dcc4b8d, 32'sh3dcaa8f5, 
               32'sh3dc905c5, 32'sh3dc761fc, 32'sh3dc5bd9b, 32'sh3dc418a1, 32'sh3dc2730f, 32'sh3dc0cce5, 32'sh3dbf2622, 32'sh3dbd7ec7, 
               32'sh3dbbd6d4, 32'sh3dba2e48, 32'sh3db88524, 32'sh3db6db68, 32'sh3db53113, 32'sh3db38627, 32'sh3db1daa2, 32'sh3db02e84, 
               32'sh3dae81cf, 32'sh3dacd481, 32'sh3dab269b, 32'sh3da9781d, 32'sh3da7c907, 32'sh3da61959, 32'sh3da46912, 32'sh3da2b834, 
               32'sh3da106bd, 32'sh3d9f54af, 32'sh3d9da208, 32'sh3d9beec9, 32'sh3d9a3af2, 32'sh3d988684, 32'sh3d96d17d, 32'sh3d951bde, 
               32'sh3d9365a8, 32'sh3d91aed9, 32'sh3d8ff772, 32'sh3d8e3f74, 32'sh3d8c86de, 32'sh3d8acdb0, 32'sh3d8913ea, 32'sh3d87598c, 
               32'sh3d859e96, 32'sh3d83e309, 32'sh3d8226e4, 32'sh3d806a27, 32'sh3d7eacd2, 32'sh3d7ceee5, 32'sh3d7b3061, 32'sh3d797145, 
               32'sh3d77b192, 32'sh3d75f147, 32'sh3d743064, 32'sh3d726ee9, 32'sh3d70acd7, 32'sh3d6eea2d, 32'sh3d6d26ec, 32'sh3d6b6313, 
               32'sh3d699ea3, 32'sh3d67d99b, 32'sh3d6613fb, 32'sh3d644dc4, 32'sh3d6286f6, 32'sh3d60bf90, 32'sh3d5ef793, 32'sh3d5d2efe, 
               32'sh3d5b65d2, 32'sh3d599c0e, 32'sh3d57d1b3, 32'sh3d5606c1, 32'sh3d543b37, 32'sh3d526f16, 32'sh3d50a25e, 32'sh3d4ed50f, 
               32'sh3d4d0728, 32'sh3d4b38aa, 32'sh3d496994, 32'sh3d4799e8, 32'sh3d45c9a4, 32'sh3d43f8c9, 32'sh3d422757, 32'sh3d40554e, 
               32'sh3d3e82ae, 32'sh3d3caf76, 32'sh3d3adba7, 32'sh3d390742, 32'sh3d373245, 32'sh3d355cb1, 32'sh3d338687, 32'sh3d31afc5, 
               32'sh3d2fd86c, 32'sh3d2e007c, 32'sh3d2c27f6, 32'sh3d2a4ed8, 32'sh3d287523, 32'sh3d269ad8, 32'sh3d24bff6, 32'sh3d22e47c, 
               32'sh3d21086c, 32'sh3d1f2bc5, 32'sh3d1d4e88, 32'sh3d1b70b3, 32'sh3d199248, 32'sh3d17b346, 32'sh3d15d3ad, 32'sh3d13f37e, 
               32'sh3d1212b7, 32'sh3d10315a, 32'sh3d0e4f67, 32'sh3d0c6cdd, 32'sh3d0a89bc, 32'sh3d08a604, 32'sh3d06c1b6, 32'sh3d04dcd2, 
               32'sh3d02f757, 32'sh3d011145, 32'sh3cff2a9d, 32'sh3cfd435e, 32'sh3cfb5b89, 32'sh3cf9731d, 32'sh3cf78a1b, 32'sh3cf5a082, 
               32'sh3cf3b653, 32'sh3cf1cb8e, 32'sh3cefe032, 32'sh3cedf440, 32'sh3cec07b8, 32'sh3cea1a99, 32'sh3ce82ce4, 32'sh3ce63e98, 
               32'sh3ce44fb7, 32'sh3ce2603f, 32'sh3ce07031, 32'sh3cde7f8d, 32'sh3cdc8e52, 32'sh3cda9c81, 32'sh3cd8aa1b, 32'sh3cd6b71e, 
               32'sh3cd4c38b, 32'sh3cd2cf62, 32'sh3cd0daa2, 32'sh3ccee54d, 32'sh3cccef62, 32'sh3ccaf8e0, 32'sh3cc901c9, 32'sh3cc70a1c, 
               32'sh3cc511d9, 32'sh3cc318ff, 32'sh3cc11f90, 32'sh3cbf258b, 32'sh3cbd2af0, 32'sh3cbb2fbf, 32'sh3cb933f9, 32'sh3cb7379c, 
               32'sh3cb53aaa, 32'sh3cb33d22, 32'sh3cb13f04, 32'sh3caf4051, 32'sh3cad4107, 32'sh3cab4128, 32'sh3ca940b3, 32'sh3ca73fa9, 
               32'sh3ca53e09, 32'sh3ca33bd3, 32'sh3ca13908, 32'sh3c9f35a7, 32'sh3c9d31b0, 32'sh3c9b2d24, 32'sh3c992803, 32'sh3c97224c, 
               32'sh3c951bff, 32'sh3c93151d, 32'sh3c910da5, 32'sh3c8f0598, 32'sh3c8cfcf6, 32'sh3c8af3be, 32'sh3c88e9f1, 32'sh3c86df8e, 
               32'sh3c84d496, 32'sh3c82c909, 32'sh3c80bce7, 32'sh3c7eb02f, 32'sh3c7ca2e2, 32'sh3c7a94ff, 32'sh3c788688, 32'sh3c76777b, 
               32'sh3c7467d9, 32'sh3c7257a2, 32'sh3c7046d6, 32'sh3c6e3574, 32'sh3c6c237e, 32'sh3c6a10f2, 32'sh3c67fdd1, 32'sh3c65ea1c, 
               32'sh3c63d5d1, 32'sh3c61c0f1, 32'sh3c5fab7c, 32'sh3c5d9573, 32'sh3c5b7ed4, 32'sh3c5967a1, 32'sh3c574fd8, 32'sh3c55377b, 
               32'sh3c531e88, 32'sh3c510501, 32'sh3c4eeae5, 32'sh3c4cd035, 32'sh3c4ab4ef, 32'sh3c489915, 32'sh3c467ca6, 32'sh3c445fa2, 
               32'sh3c42420a, 32'sh3c4023dd, 32'sh3c3e051b, 32'sh3c3be5c5, 32'sh3c39c5da, 32'sh3c37a55a, 32'sh3c358446, 32'sh3c33629d, 
               32'sh3c314060, 32'sh3c2f1d8e, 32'sh3c2cfa28, 32'sh3c2ad62d, 32'sh3c28b19e, 32'sh3c268c7a, 32'sh3c2466c2, 32'sh3c224075, 
               32'sh3c201994, 32'sh3c1df21f, 32'sh3c1bca16, 32'sh3c19a178, 32'sh3c177845, 32'sh3c154e7f, 32'sh3c132424, 32'sh3c10f935, 
               32'sh3c0ecdb2, 32'sh3c0ca19b, 32'sh3c0a74f0, 32'sh3c0847b0, 32'sh3c0619dc, 32'sh3c03eb74, 32'sh3c01bc78, 32'sh3bff8ce8, 
               32'sh3bfd5cc4, 32'sh3bfb2c0c, 32'sh3bf8fac0, 32'sh3bf6c8e0, 32'sh3bf4966c, 32'sh3bf26364, 32'sh3bf02fc9, 32'sh3bedfb99, 
               32'sh3bebc6d5, 32'sh3be9917e, 32'sh3be75b93, 32'sh3be52513, 32'sh3be2ee01, 32'sh3be0b65a, 32'sh3bde7e20, 32'sh3bdc4552, 
               32'sh3bda0bf0, 32'sh3bd7d1fa, 32'sh3bd59771, 32'sh3bd35c54, 32'sh3bd120a4, 32'sh3bcee460, 32'sh3bcca789, 32'sh3bca6a1d, 
               32'sh3bc82c1f, 32'sh3bc5ed8d, 32'sh3bc3ae67, 32'sh3bc16eae, 32'sh3bbf2e62, 32'sh3bbced82, 32'sh3bbaac0e, 32'sh3bb86a08, 
               32'sh3bb6276e, 32'sh3bb3e440, 32'sh3bb1a080, 32'sh3baf5c2c, 32'sh3bad1744, 32'sh3baad1ca, 32'sh3ba88bbc, 32'sh3ba6451b, 
               32'sh3ba3fde7, 32'sh3ba1b620, 32'sh3b9f6dc5, 32'sh3b9d24d8, 32'sh3b9adb57, 32'sh3b989144, 32'sh3b96469d, 32'sh3b93fb63, 
               32'sh3b91af97, 32'sh3b8f6337, 32'sh3b8d1644, 32'sh3b8ac8bf, 32'sh3b887aa6, 32'sh3b862bfb, 32'sh3b83dcbc, 32'sh3b818ceb, 
               32'sh3b7f3c87, 32'sh3b7ceb90, 32'sh3b7a9a07, 32'sh3b7847eb, 32'sh3b75f53c, 32'sh3b73a1fa, 32'sh3b714e25, 32'sh3b6ef9be, 
               32'sh3b6ca4c4, 32'sh3b6a4f38, 32'sh3b67f919, 32'sh3b65a268, 32'sh3b634b23, 32'sh3b60f34d, 32'sh3b5e9ae4, 32'sh3b5c41e8, 
               32'sh3b59e85a, 32'sh3b578e39, 32'sh3b553386, 32'sh3b52d841, 32'sh3b507c69, 32'sh3b4e1fff, 32'sh3b4bc303, 32'sh3b496574, 
               32'sh3b470753, 32'sh3b44a8a0, 32'sh3b42495a, 32'sh3b3fe982, 32'sh3b3d8918, 32'sh3b3b281c, 32'sh3b38c68e, 32'sh3b36646e, 
               32'sh3b3401bb, 32'sh3b319e77, 32'sh3b2f3aa0, 32'sh3b2cd637, 32'sh3b2a713d, 32'sh3b280bb0, 32'sh3b25a591, 32'sh3b233ee1, 
               32'sh3b20d79e, 32'sh3b1e6fca, 32'sh3b1c0764, 32'sh3b199e6c, 32'sh3b1734e2, 32'sh3b14cac6, 32'sh3b126019, 32'sh3b0ff4d9, 
               32'sh3b0d8909, 32'sh3b0b1ca6, 32'sh3b08afb2, 32'sh3b06422c, 32'sh3b03d414, 32'sh3b01656b, 32'sh3afef630, 32'sh3afc8663, 
               32'sh3afa1605, 32'sh3af7a516, 32'sh3af53395, 32'sh3af2c183, 32'sh3af04edf, 32'sh3aeddba9, 32'sh3aeb67e3, 32'sh3ae8f38b, 
               32'sh3ae67ea1, 32'sh3ae40926, 32'sh3ae1931a, 32'sh3adf1c7d, 32'sh3adca54e, 32'sh3ada2d8e, 32'sh3ad7b53d, 32'sh3ad53c5b, 
               32'sh3ad2c2e8, 32'sh3ad048e3, 32'sh3acdce4d, 32'sh3acb5327, 32'sh3ac8d76f, 32'sh3ac65b26, 32'sh3ac3de4c, 32'sh3ac160e1, 
               32'sh3abee2e5, 32'sh3abc6458, 32'sh3ab9e53a, 32'sh3ab7658c, 32'sh3ab4e54c, 32'sh3ab2647c, 32'sh3aafe31b, 32'sh3aad6129, 
               32'sh3aaadea6, 32'sh3aa85b92, 32'sh3aa5d7ee, 32'sh3aa353b9, 32'sh3aa0cef3, 32'sh3a9e499d, 32'sh3a9bc3b6, 32'sh3a993d3e, 
               32'sh3a96b636, 32'sh3a942e9d, 32'sh3a91a674, 32'sh3a8f1dba, 32'sh3a8c9470, 32'sh3a8a0a95, 32'sh3a87802a, 32'sh3a84f52f, 
               32'sh3a8269a3, 32'sh3a7fdd86, 32'sh3a7d50da, 32'sh3a7ac39d, 32'sh3a7835cf, 32'sh3a75a772, 32'sh3a731884, 32'sh3a708906, 
               32'sh3a6df8f8, 32'sh3a6b6859, 32'sh3a68d72b, 32'sh3a66456c, 32'sh3a63b31d, 32'sh3a61203e, 32'sh3a5e8cd0, 32'sh3a5bf8d1, 
               32'sh3a596442, 32'sh3a56cf23, 32'sh3a543974, 32'sh3a51a335, 32'sh3a4f0c67, 32'sh3a4c7508, 32'sh3a49dd1a, 32'sh3a47449c, 
               32'sh3a44ab8e, 32'sh3a4211f0, 32'sh3a3f77c3, 32'sh3a3cdd05, 32'sh3a3a41b9, 32'sh3a37a5dc, 32'sh3a350970, 32'sh3a326c74, 
               32'sh3a2fcee8, 32'sh3a2d30cd, 32'sh3a2a9223, 32'sh3a27f2e9, 32'sh3a25531f, 32'sh3a22b2c6, 32'sh3a2011de, 32'sh3a1d7066, 
               32'sh3a1ace5f, 32'sh3a182bc8, 32'sh3a1588a2, 32'sh3a12e4ed, 32'sh3a1040a8, 32'sh3a0d9bd4, 32'sh3a0af671, 32'sh3a08507f, 
               32'sh3a05a9fd, 32'sh3a0302ed, 32'sh3a005b4d, 32'sh39fdb31e, 32'sh39fb0a60, 32'sh39f86113, 32'sh39f5b737, 32'sh39f30ccc, 
               32'sh39f061d2, 32'sh39edb649, 32'sh39eb0a31, 32'sh39e85d8a, 32'sh39e5b054, 32'sh39e3028f, 32'sh39e0543c, 32'sh39dda55a, 
               32'sh39daf5e8, 32'sh39d845e9, 32'sh39d5955a, 32'sh39d2e43d, 32'sh39d03291, 32'sh39cd8056, 32'sh39cacd8d, 32'sh39c81a36, 
               32'sh39c5664f, 32'sh39c2b1da, 32'sh39bffcd7, 32'sh39bd4745, 32'sh39ba9125, 32'sh39b7da76, 32'sh39b52339, 32'sh39b26b6d, 
               32'sh39afb313, 32'sh39acfa2b, 32'sh39aa40b4, 32'sh39a786af, 32'sh39a4cc1c, 32'sh39a210fb, 32'sh399f554b, 32'sh399c990d, 
               32'sh3999dc42, 32'sh39971ee7, 32'sh399460ff, 32'sh3991a289, 32'sh398ee385, 32'sh398c23f3, 32'sh398963d2, 32'sh3986a324, 
               32'sh3983e1e8, 32'sh3981201e, 32'sh397e5dc6, 32'sh397b9ae0, 32'sh3978d76c, 32'sh3976136b, 32'sh39734edc, 32'sh397089bf, 
               32'sh396dc414, 32'sh396afddc, 32'sh39683715, 32'sh39656fc2, 32'sh3962a7e0, 32'sh395fdf71, 32'sh395d1675, 32'sh395a4ceb, 
               32'sh395782d3, 32'sh3954b82e, 32'sh3951ecfc, 32'sh394f213c, 32'sh394c54ee, 32'sh39498814, 32'sh3946baac, 32'sh3943ecb6, 
               32'sh39411e33, 32'sh393e4f23, 32'sh393b7f86, 32'sh3938af5c, 32'sh3935dea4, 32'sh39330d5f, 32'sh39303b8e, 32'sh392d692f, 
               32'sh392a9642, 32'sh3927c2c9, 32'sh3924eec3, 32'sh39221a30, 32'sh391f4510, 32'sh391c6f63, 32'sh39199929, 32'sh3916c262, 
               32'sh3913eb0e, 32'sh3911132d, 32'sh390e3ac0, 32'sh390b61c6, 32'sh3908883f, 32'sh3905ae2b, 32'sh3902d38b, 32'sh38fff85e, 
               32'sh38fd1ca4, 32'sh38fa405e, 32'sh38f7638b, 32'sh38f4862c, 32'sh38f1a840, 32'sh38eec9c7, 32'sh38ebeac2, 32'sh38e90b31, 
               32'sh38e62b13, 32'sh38e34a69, 32'sh38e06932, 32'sh38dd8770, 32'sh38daa520, 32'sh38d7c245, 32'sh38d4dedd, 32'sh38d1fae9, 
               32'sh38cf1669, 32'sh38cc315d, 32'sh38c94bc4, 32'sh38c665a0, 32'sh38c37eef, 32'sh38c097b2, 32'sh38bdafea, 32'sh38bac795, 
               32'sh38b7deb4, 32'sh38b4f547, 32'sh38b20b4f, 32'sh38af20ca, 32'sh38ac35ba, 32'sh38a94a1e, 32'sh38a65df6, 32'sh38a37142, 
               32'sh38a08402, 32'sh389d9637, 32'sh389aa7e0, 32'sh3897b8fe, 32'sh3894c98f, 32'sh3891d995, 32'sh388ee910, 32'sh388bf7ff, 
               32'sh38890663, 32'sh3886143b, 32'sh38832187, 32'sh38802e48, 32'sh387d3a7e, 32'sh387a4628, 32'sh38775147, 32'sh38745bdb, 
               32'sh387165e3, 32'sh386e6f60, 32'sh386b7852, 32'sh386880b8, 32'sh38658894, 32'sh38628fe4, 32'sh385f96a9, 32'sh385c9ce3, 
               32'sh3859a292, 32'sh3856a7b6, 32'sh3853ac4f, 32'sh3850b05d, 32'sh384db3e0, 32'sh384ab6d8, 32'sh3847b946, 32'sh3844bb28, 
               32'sh3841bc7f, 32'sh383ebd4c, 32'sh383bbd8e, 32'sh3838bd45, 32'sh3835bc71, 32'sh3832bb13, 32'sh382fb92a, 32'sh382cb6b7, 
               32'sh3829b3b9, 32'sh3826b030, 32'sh3823ac1d, 32'sh3820a77f, 32'sh381da256, 32'sh381a9ca4, 32'sh38179666, 32'sh38148f9f, 
               32'sh3811884d, 32'sh380e8071, 32'sh380b780a, 32'sh38086f19, 32'sh3805659e, 32'sh38025b98, 32'sh37ff5109, 32'sh37fc45ef, 
               32'sh37f93a4b, 32'sh37f62e1d, 32'sh37f32165, 32'sh37f01423, 32'sh37ed0657, 32'sh37e9f801, 32'sh37e6e921, 32'sh37e3d9b7, 
               32'sh37e0c9c3, 32'sh37ddb945, 32'sh37daa83d, 32'sh37d796ac, 32'sh37d48490, 32'sh37d171eb, 32'sh37ce5ebd, 32'sh37cb4b04, 
               32'sh37c836c2, 32'sh37c521f6, 32'sh37c20ca1, 32'sh37bef6c2, 32'sh37bbe05a, 32'sh37b8c968, 32'sh37b5b1ec, 32'sh37b299e7, 
               32'sh37af8159, 32'sh37ac6841, 32'sh37a94ea0, 32'sh37a63476, 32'sh37a319c2, 32'sh379ffe85, 32'sh379ce2be, 32'sh3799c66f, 
               32'sh3796a996, 32'sh37938c34, 32'sh37906e49, 32'sh378d4fd5, 32'sh378a30d8, 32'sh37871152, 32'sh3783f143, 32'sh3780d0aa, 
               32'sh377daf89, 32'sh377a8ddf, 32'sh37776bac, 32'sh377448f0, 32'sh377125ac, 32'sh376e01de, 32'sh376add88, 32'sh3767b8a9, 
               32'sh37649341, 32'sh37616d51, 32'sh375e46d8, 32'sh375b1fd7, 32'sh3757f84c, 32'sh3754d03a, 32'sh3751a79e, 32'sh374e7e7b, 
               32'sh374b54ce, 32'sh37482a9a, 32'sh3744ffdd, 32'sh3741d497, 32'sh373ea8ca, 32'sh373b7c73, 32'sh37384f95, 32'sh3735222f, 
               32'sh3731f440, 32'sh372ec5c9, 32'sh372b96ca, 32'sh37286742, 32'sh37253733, 32'sh3722069b, 32'sh371ed57c, 32'sh371ba3d4, 
               32'sh371871a5, 32'sh37153eee, 32'sh37120bae, 32'sh370ed7e7, 32'sh370ba398, 32'sh37086ec1, 32'sh37053962, 32'sh3702037c, 
               32'sh36fecd0e, 32'sh36fb9618, 32'sh36f85e9a, 32'sh36f52695, 32'sh36f1ee09, 32'sh36eeb4f4, 32'sh36eb7b58, 32'sh36e84135, 
               32'sh36e5068a, 32'sh36e1cb58, 32'sh36de8f9e, 32'sh36db535d, 32'sh36d81695, 32'sh36d4d945, 32'sh36d19b6e, 32'sh36ce5d10, 
               32'sh36cb1e2a, 32'sh36c7debd, 32'sh36c49ec9, 32'sh36c15e4e, 32'sh36be1d4c, 32'sh36badbc3, 32'sh36b799b3, 32'sh36b4571b, 
               32'sh36b113fd, 32'sh36add058, 32'sh36aa8c2c, 32'sh36a74779, 32'sh36a4023f, 32'sh36a0bc7e, 32'sh369d7637, 32'sh369a2f69, 
               32'sh3696e814, 32'sh3693a038, 32'sh369057d6, 32'sh368d0eed, 32'sh3689c57d, 32'sh36867b87, 32'sh3683310b, 32'sh367fe608, 
               32'sh367c9a7e, 32'sh36794e6e, 32'sh367601d7, 32'sh3672b4bb, 32'sh366f6717, 32'sh366c18ee, 32'sh3668ca3e, 32'sh36657b08, 
               32'sh36622b4c, 32'sh365edb09, 32'sh365b8a41, 32'sh365838f2, 32'sh3654e71d, 32'sh365194c3, 32'sh364e41e2, 32'sh364aee7b, 
               32'sh36479a8e, 32'sh3644461b, 32'sh3640f123, 32'sh363d9ba4, 32'sh363a45a0, 32'sh3636ef16, 32'sh36339806, 32'sh36304070, 
               32'sh362ce855, 32'sh36298fb4, 32'sh3626368d, 32'sh3622dce1, 32'sh361f82af, 32'sh361c27f7, 32'sh3618ccba, 32'sh361570f8, 
               32'sh361214b0, 32'sh360eb7e3, 32'sh360b5a90, 32'sh3607fcb8, 32'sh36049e5b, 32'sh36013f78, 32'sh35fde011, 32'sh35fa8023, 
               32'sh35f71fb1, 32'sh35f3beba, 32'sh35f05d3d, 32'sh35ecfb3c, 32'sh35e998b5, 32'sh35e635a9, 32'sh35e2d219, 32'sh35df6e03, 
               32'sh35dc0968, 32'sh35d8a449, 32'sh35d53ea5, 32'sh35d1d87c, 32'sh35ce71ce, 32'sh35cb0a9b, 32'sh35c7a2e3, 32'sh35c43aa7, 
               32'sh35c0d1e7, 32'sh35bd68a1, 32'sh35b9fed7, 32'sh35b69489, 32'sh35b329b5, 32'sh35afbe5e, 32'sh35ac5282, 32'sh35a8e621, 
               32'sh35a5793c, 32'sh35a20bd3, 32'sh359e9de5, 32'sh359b2f73, 32'sh3597c07d, 32'sh35945103, 32'sh3590e104, 32'sh358d7081, 
               32'sh3589ff7a, 32'sh35868def, 32'sh35831be0, 32'sh357fa94d, 32'sh357c3636, 32'sh3578c29b, 32'sh35754e7c, 32'sh3571d9d9, 
               32'sh356e64b2, 32'sh356aef08, 32'sh356778d9, 32'sh35640227, 32'sh35608af1, 32'sh355d1337, 32'sh35599afa, 32'sh35562239, 
               32'sh3552a8f4, 32'sh354f2f2c, 32'sh354bb4e1, 32'sh35483a11, 32'sh3544bebf, 32'sh354142e9, 32'sh353dc68f, 32'sh353a49b2, 
               32'sh3536cc52, 32'sh35334e6f, 32'sh352fd008, 32'sh352c511e, 32'sh3528d1b1, 32'sh352551c0, 32'sh3521d14d, 32'sh351e5056, 
               32'sh351acedd, 32'sh35174ce0, 32'sh3513ca60, 32'sh3510475e, 32'sh350cc3d8, 32'sh35093fd0, 32'sh3505bb44, 32'sh35023636, 
               32'sh34feb0a5, 32'sh34fb2a92, 32'sh34f7a3fb, 32'sh34f41ce2, 32'sh34f09546, 32'sh34ed0d28, 32'sh34e98487, 32'sh34e5fb63, 
               32'sh34e271bd, 32'sh34dee795, 32'sh34db5cea, 32'sh34d7d1bc, 32'sh34d4460c, 32'sh34d0b9da, 32'sh34cd2d26, 32'sh34c99fef, 
               32'sh34c61236, 32'sh34c283fb, 32'sh34bef53d, 32'sh34bb65fe, 32'sh34b7d63c, 32'sh34b445f8, 32'sh34b0b533, 32'sh34ad23eb, 
               32'sh34a99221, 32'sh34a5ffd5, 32'sh34a26d08, 32'sh349ed9b8, 32'sh349b45e7, 32'sh3497b194, 32'sh34941cbf, 32'sh34908768, 
               32'sh348cf190, 32'sh34895b36, 32'sh3485c45b, 32'sh34822cfd, 32'sh347e951f, 32'sh347afcbe, 32'sh347763dd, 32'sh3473ca79, 
               32'sh34703095, 32'sh346c962f, 32'sh3468fb47, 32'sh34655fdf, 32'sh3461c3f5, 32'sh345e2789, 32'sh345a8a9d, 32'sh3456ed2f, 
               32'sh34534f41, 32'sh344fb0d1, 32'sh344c11e0, 32'sh3448726e, 32'sh3444d27b, 32'sh34413207, 32'sh343d9112, 32'sh3439ef9c, 
               32'sh34364da6, 32'sh3432ab2e, 32'sh342f0836, 32'sh342b64bd, 32'sh3427c0c3, 32'sh34241c49, 32'sh3420774d, 32'sh341cd1d2, 
               32'sh34192bd5, 32'sh34158559, 32'sh3411de5b, 32'sh340e36dd, 32'sh340a8edf, 32'sh3406e660, 32'sh34033d61, 32'sh33ff93e2, 
               32'sh33fbe9e2, 32'sh33f83f62, 32'sh33f49462, 32'sh33f0e8e2, 32'sh33ed3ce1, 32'sh33e99061, 32'sh33e5e360, 32'sh33e235df, 
               32'sh33de87de, 32'sh33dad95e, 32'sh33d72a5d, 32'sh33d37adc, 32'sh33cfcadc, 32'sh33cc1a5b, 32'sh33c8695b, 32'sh33c4b7db, 
               32'sh33c105db, 32'sh33bd535c, 32'sh33b9a05d, 32'sh33b5ecde, 32'sh33b238e0, 32'sh33ae8462, 32'sh33aacf65, 32'sh33a719e8, 
               32'sh33a363ec, 32'sh339fad70, 32'sh339bf675, 32'sh33983efb, 32'sh33948701, 32'sh3390ce88, 32'sh338d1590, 32'sh33895c18, 
               32'sh3385a222, 32'sh3381e7ac, 32'sh337e2cb7, 32'sh337a7144, 32'sh3376b551, 32'sh3372f8df, 32'sh336f3bee, 32'sh336b7e7e, 
               32'sh3367c090, 32'sh33640223, 32'sh33604336, 32'sh335c83cb, 32'sh3358c3e2, 32'sh33550379, 32'sh33514292, 32'sh334d812d, 
               32'sh3349bf48, 32'sh3345fce6, 32'sh33423a04, 32'sh333e76a4, 32'sh333ab2c6, 32'sh3336ee6a, 32'sh3333298f, 32'sh332f6435, 
               32'sh332b9e5e, 32'sh3327d808, 32'sh33241134, 32'sh332049e1, 32'sh331c8211, 32'sh3318b9c2, 32'sh3314f0f6, 32'sh331127ab, 
               32'sh330d5de3, 32'sh3309939c, 32'sh3305c8d7, 32'sh3301fd95, 32'sh32fe31d5, 32'sh32fa6596, 32'sh32f698db, 32'sh32f2cba1, 
               32'sh32eefdea, 32'sh32eb2fb5, 32'sh32e76102, 32'sh32e391d2, 32'sh32dfc224, 32'sh32dbf1f8, 32'sh32d82150, 32'sh32d45029, 
               32'sh32d07e85, 32'sh32ccac64, 32'sh32c8d9c6, 32'sh32c506aa, 32'sh32c13311, 32'sh32bd5efb, 32'sh32b98a67, 32'sh32b5b557, 
               32'sh32b1dfc9, 32'sh32ae09be, 32'sh32aa3336, 32'sh32a65c32, 32'sh32a284b0, 32'sh329eacb1, 32'sh329ad435, 32'sh3296fb3d, 
               32'sh329321c7, 32'sh328f47d5, 32'sh328b6d66, 32'sh3287927b, 32'sh3283b712, 32'sh327fdb2d, 32'sh327bfecc, 32'sh327821ee, 
               32'sh32744493, 32'sh327066bc, 32'sh326c8868, 32'sh3268a998, 32'sh3264ca4c, 32'sh3260ea83, 32'sh325d0a3e, 32'sh3259297d, 
               32'sh32554840, 32'sh32516686, 32'sh324d8450, 32'sh3249a19e, 32'sh3245be70, 32'sh3241dac6, 32'sh323df6a0, 32'sh323a11fe, 
               32'sh32362ce0, 32'sh32324746, 32'sh322e6130, 32'sh322a7a9e, 32'sh32269391, 32'sh3222ac08, 32'sh321ec403, 32'sh321adb83, 
               32'sh3216f287, 32'sh3213090f, 32'sh320f1f1c, 32'sh320b34ad, 32'sh320749c3, 32'sh32035e5d, 32'sh31ff727c, 32'sh31fb8620, 
               32'sh31f79948, 32'sh31f3abf5, 32'sh31efbe27, 32'sh31ebcfdd, 32'sh31e7e118, 32'sh31e3f1d8, 32'sh31e0021e, 32'sh31dc11e8, 
               32'sh31d82137, 32'sh31d4300b, 32'sh31d03e64, 32'sh31cc4c42, 32'sh31c859a5, 32'sh31c4668d, 32'sh31c072fb, 32'sh31bc7eee, 
               32'sh31b88a66, 32'sh31b49564, 32'sh31b09fe7, 32'sh31aca9ef, 32'sh31a8b37c, 32'sh31a4bc90, 32'sh31a0c528, 32'sh319ccd46, 
               32'sh3198d4ea, 32'sh3194dc14, 32'sh3190e2c3, 32'sh318ce8f7, 32'sh3188eeb2, 32'sh3184f3f2, 32'sh3180f8b8, 32'sh317cfd04, 
               32'sh317900d6, 32'sh3175042e, 32'sh3171070c, 32'sh316d096f, 32'sh31690b59, 32'sh31650cc9, 32'sh31610dbf, 32'sh315d0e3b, 
               32'sh31590e3e, 32'sh31550dc6, 32'sh31510cd5, 32'sh314d0b6a, 32'sh31490986, 32'sh31450728, 32'sh31410450, 32'sh313d00ff, 
               32'sh3138fd35, 32'sh3134f8f1, 32'sh3130f433, 32'sh312ceefc, 32'sh3128e94c, 32'sh3124e322, 32'sh3120dc80, 32'sh311cd564, 
               32'sh3118cdcf, 32'sh3114c5c0, 32'sh3110bd39, 32'sh310cb438, 32'sh3108aabf, 32'sh3104a0cc, 32'sh31009661, 32'sh30fc8b7d, 
               32'sh30f8801f, 32'sh30f47449, 32'sh30f067fb, 32'sh30ec5b33, 32'sh30e84df3, 32'sh30e4403a, 32'sh30e03208, 32'sh30dc235e, 
               32'sh30d8143b, 32'sh30d404a0, 32'sh30cff48c, 32'sh30cbe400, 32'sh30c7d2fb, 32'sh30c3c17e, 32'sh30bfaf89, 32'sh30bb9d1c, 
               32'sh30b78a36, 32'sh30b376d8, 32'sh30af6302, 32'sh30ab4eb3, 32'sh30a739ed, 32'sh30a324af, 32'sh309f0ef8, 32'sh309af8ca, 
               32'sh3096e223, 32'sh3092cb05, 32'sh308eb36f, 32'sh308a9b61, 32'sh308682dc, 32'sh308269de, 32'sh307e5069, 32'sh307a367c, 
               32'sh30761c18, 32'sh3072013c, 32'sh306de5e9, 32'sh3069ca1e, 32'sh3065addb, 32'sh30619121, 32'sh305d73f0, 32'sh30595648, 
               32'sh30553828, 32'sh30511991, 32'sh304cfa83, 32'sh3048dafd, 32'sh3044bb00, 32'sh30409a8d, 32'sh303c79a2, 32'sh30385840, 
               32'sh30343667, 32'sh30301418, 32'sh302bf151, 32'sh3027ce14, 32'sh3023aa5f, 32'sh301f8634, 32'sh301b6193, 32'sh30173c7a, 
               32'sh301316eb, 32'sh300ef0e5, 32'sh300aca69, 32'sh3006a376, 32'sh30027c0c, 32'sh2ffe542d, 32'sh2ffa2bd6, 32'sh2ff6030a, 
               32'sh2ff1d9c7, 32'sh2fedb00d, 32'sh2fe985de, 32'sh2fe55b38, 32'sh2fe1301c, 32'sh2fdd048a, 32'sh2fd8d882, 32'sh2fd4ac04, 
               32'sh2fd07f0f, 32'sh2fcc51a5, 32'sh2fc823c5, 32'sh2fc3f56f, 32'sh2fbfc6a3, 32'sh2fbb9761, 32'sh2fb767aa, 32'sh2fb3377c, 
               32'sh2faf06da, 32'sh2faad5c1, 32'sh2fa6a433, 32'sh2fa2722f, 32'sh2f9e3fb6, 32'sh2f9a0cc7, 32'sh2f95d963, 32'sh2f91a589, 
               32'sh2f8d713a, 32'sh2f893c75, 32'sh2f85073c, 32'sh2f80d18d, 32'sh2f7c9b69, 32'sh2f7864cf, 32'sh2f742dc1, 32'sh2f6ff63d, 
               32'sh2f6bbe45, 32'sh2f6785d7, 32'sh2f634cf5, 32'sh2f5f139d, 32'sh2f5ad9d1, 32'sh2f569f90, 32'sh2f5264da, 32'sh2f4e29af, 
               32'sh2f49ee0f, 32'sh2f45b1fb, 32'sh2f417573, 32'sh2f3d3875, 32'sh2f38fb03, 32'sh2f34bd1d, 32'sh2f307ec2, 32'sh2f2c3ff2, 
               32'sh2f2800af, 32'sh2f23c0f6, 32'sh2f1f80ca, 32'sh2f1b4029, 32'sh2f16ff14, 32'sh2f12bd8b, 32'sh2f0e7b8e, 32'sh2f0a391d, 
               32'sh2f05f637, 32'sh2f01b2de, 32'sh2efd6f10, 32'sh2ef92acf, 32'sh2ef4e619, 32'sh2ef0a0f0, 32'sh2eec5b53, 32'sh2ee81543, 
               32'sh2ee3cebe, 32'sh2edf87c6, 32'sh2edb405a, 32'sh2ed6f87a, 32'sh2ed2b027, 32'sh2ece6761, 32'sh2eca1e27, 32'sh2ec5d479, 
               32'sh2ec18a58, 32'sh2ebd3fc4, 32'sh2eb8f4bc, 32'sh2eb4a942, 32'sh2eb05d53, 32'sh2eac10f2, 32'sh2ea7c41e, 32'sh2ea376d6, 
               32'sh2e9f291b, 32'sh2e9adaee, 32'sh2e968c4d, 32'sh2e923d39, 32'sh2e8dedb3, 32'sh2e899db9, 32'sh2e854d4d, 32'sh2e80fc6e, 
               32'sh2e7cab1c, 32'sh2e785958, 32'sh2e740720, 32'sh2e6fb477, 32'sh2e6b615a, 32'sh2e670dcb, 32'sh2e62b9ca, 32'sh2e5e6556, 
               32'sh2e5a1070, 32'sh2e55bb17, 32'sh2e51654c, 32'sh2e4d0f0f, 32'sh2e48b860, 32'sh2e44613e, 32'sh2e4009aa, 32'sh2e3bb1a4, 
               32'sh2e37592c, 32'sh2e330042, 32'sh2e2ea6e6, 32'sh2e2a4d18, 32'sh2e25f2d8, 32'sh2e219826, 32'sh2e1d3d03, 32'sh2e18e16d, 
               32'sh2e148566, 32'sh2e1028ed, 32'sh2e0bcc03, 32'sh2e076ea7, 32'sh2e0310d9, 32'sh2dfeb29a, 32'sh2dfa53e9, 32'sh2df5f4c7, 
               32'sh2df19534, 32'sh2ded352f, 32'sh2de8d4b8, 32'sh2de473d1, 32'sh2de01278, 32'sh2ddbb0ae, 32'sh2dd74e73, 32'sh2dd2ebc7, 
               32'sh2dce88aa, 32'sh2dca251c, 32'sh2dc5c11c, 32'sh2dc15cac, 32'sh2dbcf7cb, 32'sh2db89279, 32'sh2db42cb6, 32'sh2dafc683, 
               32'sh2dab5fdf, 32'sh2da6f8ca, 32'sh2da29144, 32'sh2d9e294e, 32'sh2d99c0e7, 32'sh2d955810, 32'sh2d90eec8, 32'sh2d8c8510, 
               32'sh2d881ae8, 32'sh2d83b04f, 32'sh2d7f4545, 32'sh2d7ad9cc, 32'sh2d766de2, 32'sh2d720189, 32'sh2d6d94bf, 32'sh2d692784, 
               32'sh2d64b9da, 32'sh2d604bc0, 32'sh2d5bdd36, 32'sh2d576e3c, 32'sh2d52fed2, 32'sh2d4e8ef9, 32'sh2d4a1eaf, 32'sh2d45adf6, 
               32'sh2d413ccd, 32'sh2d3ccb34, 32'sh2d38592c, 32'sh2d33e6b4, 32'sh2d2f73cd, 32'sh2d2b0076, 32'sh2d268cb0, 32'sh2d22187a, 
               32'sh2d1da3d5, 32'sh2d192ec1, 32'sh2d14b93d, 32'sh2d10434a, 32'sh2d0bcce8, 32'sh2d075617, 32'sh2d02ded7, 32'sh2cfe6728, 
               32'sh2cf9ef09, 32'sh2cf5767c, 32'sh2cf0fd80, 32'sh2cec8414, 32'sh2ce80a3a, 32'sh2ce38ff1, 32'sh2cdf153a, 32'sh2cda9a14, 
               32'sh2cd61e7f, 32'sh2cd1a27b, 32'sh2ccd2609, 32'sh2cc8a928, 32'sh2cc42bd9, 32'sh2cbfae1b, 32'sh2cbb2fef, 32'sh2cb6b155, 
               32'sh2cb2324c, 32'sh2cadb2d5, 32'sh2ca932ef, 32'sh2ca4b29c, 32'sh2ca031da, 32'sh2c9bb0ab, 32'sh2c972f0d, 32'sh2c92ad01, 
               32'sh2c8e2a87, 32'sh2c89a79f, 32'sh2c85244a, 32'sh2c80a086, 32'sh2c7c1c55, 32'sh2c7797b6, 32'sh2c7312a9, 32'sh2c6e8d2e, 
               32'sh2c6a0746, 32'sh2c6580f1, 32'sh2c60fa2d, 32'sh2c5c72fd, 32'sh2c57eb5e, 32'sh2c536353, 32'sh2c4edada, 32'sh2c4a51f3, 
               32'sh2c45c8a0, 32'sh2c413edf, 32'sh2c3cb4b1, 32'sh2c382a16, 32'sh2c339f0e, 32'sh2c2f1398, 32'sh2c2a87b6, 32'sh2c25fb66, 
               32'sh2c216eaa, 32'sh2c1ce181, 32'sh2c1853eb, 32'sh2c13c5e8, 32'sh2c0f3779, 32'sh2c0aa89c, 32'sh2c061953, 32'sh2c01899e, 
               32'sh2bfcf97c, 32'sh2bf868ed, 32'sh2bf3d7f2, 32'sh2bef468a, 32'sh2beab4b6, 32'sh2be62276, 32'sh2be18fc9, 32'sh2bdcfcb0, 
               32'sh2bd8692b, 32'sh2bd3d53a, 32'sh2bcf40dc, 32'sh2bcaac12, 32'sh2bc616dd, 32'sh2bc1813b, 32'sh2bbceb2d, 32'sh2bb854b4, 
               32'sh2bb3bdce, 32'sh2baf267d, 32'sh2baa8ec0, 32'sh2ba5f697, 32'sh2ba15e03, 32'sh2b9cc503, 32'sh2b982b97, 32'sh2b9391c0, 
               32'sh2b8ef77d, 32'sh2b8a5cce, 32'sh2b85c1b5, 32'sh2b812630, 32'sh2b7c8a3f, 32'sh2b77ede3, 32'sh2b73511c, 32'sh2b6eb3ea, 
               32'sh2b6a164d, 32'sh2b657844, 32'sh2b60d9d0, 32'sh2b5c3af2, 32'sh2b579ba8, 32'sh2b52fbf4, 32'sh2b4e5bd4, 32'sh2b49bb4a, 
               32'sh2b451a55, 32'sh2b4078f5, 32'sh2b3bd72a, 32'sh2b3734f5, 32'sh2b329255, 32'sh2b2def4b, 32'sh2b294bd5, 32'sh2b24a7f6, 
               32'sh2b2003ac, 32'sh2b1b5ef8, 32'sh2b16b9d9, 32'sh2b121450, 32'sh2b0d6e5c, 32'sh2b08c7ff, 32'sh2b042137, 32'sh2aff7a05, 
               32'sh2afad269, 32'sh2af62a63, 32'sh2af181f3, 32'sh2aecd919, 32'sh2ae82fd5, 32'sh2ae38627, 32'sh2adedc10, 32'sh2ada318e, 
               32'sh2ad586a3, 32'sh2ad0db4e, 32'sh2acc2f90, 32'sh2ac78368, 32'sh2ac2d6d6, 32'sh2abe29db, 32'sh2ab97c77, 32'sh2ab4cea9, 
               32'sh2ab02071, 32'sh2aab71d0, 32'sh2aa6c2c6, 32'sh2aa21353, 32'sh2a9d6377, 32'sh2a98b331, 32'sh2a940283, 32'sh2a8f516b, 
               32'sh2a8a9fea, 32'sh2a85ee00, 32'sh2a813bae, 32'sh2a7c88f2, 32'sh2a77d5ce, 32'sh2a732241, 32'sh2a6e6e4b, 32'sh2a69b9ec, 
               32'sh2a650525, 32'sh2a604ff5, 32'sh2a5b9a5d, 32'sh2a56e45c, 32'sh2a522df3, 32'sh2a4d7721, 32'sh2a48bfe7, 32'sh2a440844, 
               32'sh2a3f503a, 32'sh2a3a97c7, 32'sh2a35deeb, 32'sh2a3125a8, 32'sh2a2c6bfd, 32'sh2a27b1e9, 32'sh2a22f76e, 32'sh2a1e3c8a, 
               32'sh2a19813f, 32'sh2a14c58b, 32'sh2a100970, 32'sh2a0b4ced, 32'sh2a069003, 32'sh2a01d2b0, 32'sh29fd14f6, 32'sh29f856d5, 
               32'sh29f3984c, 32'sh29eed95b, 32'sh29ea1a03, 32'sh29e55a43, 32'sh29e09a1c, 32'sh29dbd98e, 32'sh29d71899, 32'sh29d2573c, 
               32'sh29cd9578, 32'sh29c8d34d, 32'sh29c410ba, 32'sh29bf4dc1, 32'sh29ba8a61, 32'sh29b5c69a, 32'sh29b1026c, 32'sh29ac3dd7, 
               32'sh29a778db, 32'sh29a2b378, 32'sh299dedaf, 32'sh2999277f, 32'sh299460e8, 32'sh298f99eb, 32'sh298ad287, 32'sh29860abd, 
               32'sh2981428c, 32'sh297c79f5, 32'sh2977b0f7, 32'sh2972e793, 32'sh296e1dc9, 32'sh29695399, 32'sh29648902, 32'sh295fbe06, 
               32'sh295af2a3, 32'sh295626da, 32'sh29515aab, 32'sh294c8e16, 32'sh2947c11c, 32'sh2942f3bb, 32'sh293e25f5, 32'sh293957c9, 
               32'sh29348937, 32'sh292fba40, 32'sh292aeae3, 32'sh29261b20, 32'sh29214af8, 32'sh291c7a6a, 32'sh2917a977, 32'sh2912d81f, 
               32'sh290e0661, 32'sh2909343e, 32'sh290461b5, 32'sh28ff8ec8, 32'sh28fabb75, 32'sh28f5e7bd, 32'sh28f113a0, 32'sh28ec3f1e, 
               32'sh28e76a37, 32'sh28e294eb, 32'sh28ddbf3b, 32'sh28d8e925, 32'sh28d412ab, 32'sh28cf3bcc, 32'sh28ca6488, 32'sh28c58cdf, 
               32'sh28c0b4d2, 32'sh28bbdc61, 32'sh28b7038b, 32'sh28b22a50, 32'sh28ad50b1, 32'sh28a876ae, 32'sh28a39c46, 32'sh289ec17a, 
               32'sh2899e64a, 32'sh28950ab6, 32'sh28902ebd, 32'sh288b5261, 32'sh288675a0, 32'sh2881987c, 32'sh287cbaf3, 32'sh2877dd07, 
               32'sh2872feb6, 32'sh286e2002, 32'sh286940ea, 32'sh2864616f, 32'sh285f8190, 32'sh285aa14d, 32'sh2855c0a6, 32'sh2850df9d, 
               32'sh284bfe2f, 32'sh28471c5e, 32'sh28423a2a, 32'sh283d5793, 32'sh28387498, 32'sh2833913a, 32'sh282ead78, 32'sh2829c954, 
               32'sh2824e4cc, 32'sh281fffe2, 32'sh281b1a94, 32'sh281634e4, 32'sh28114ed0, 32'sh280c685a, 32'sh28078181, 32'sh28029a45, 
               32'sh27fdb2a7, 32'sh27f8caa5, 32'sh27f3e241, 32'sh27eef97b, 32'sh27ea1052, 32'sh27e526c6, 32'sh27e03cd8, 32'sh27db5288, 
               32'sh27d667d5, 32'sh27d17cc1, 32'sh27cc9149, 32'sh27c7a570, 32'sh27c2b934, 32'sh27bdcc97, 32'sh27b8df97, 32'sh27b3f235, 
               32'sh27af0472, 32'sh27aa164c, 32'sh27a527c4, 32'sh27a038db, 32'sh279b4990, 32'sh279659e3, 32'sh279169d5, 32'sh278c7965, 
               32'sh27878893, 32'sh27829760, 32'sh277da5cb, 32'sh2778b3d5, 32'sh2773c17d, 32'sh276ecec5, 32'sh2769dbaa, 32'sh2764e82f, 
               32'sh275ff452, 32'sh275b0014, 32'sh27560b76, 32'sh27511676, 32'sh274c2115, 32'sh27472b53, 32'sh27423530, 32'sh273d3eac, 
               32'sh273847c8, 32'sh27335082, 32'sh272e58dc, 32'sh272960d6, 32'sh2724686e, 32'sh271f6fa6, 32'sh271a767e, 32'sh27157cf5, 
               32'sh2710830c, 32'sh270b88c2, 32'sh27068e18, 32'sh2701930e, 32'sh26fc97a3, 32'sh26f79bd8, 32'sh26f29fad, 32'sh26eda322, 
               32'sh26e8a637, 32'sh26e3a8ec, 32'sh26deab41, 32'sh26d9ad36, 32'sh26d4aecb, 32'sh26cfb000, 32'sh26cab0d6, 32'sh26c5b14c, 
               32'sh26c0b162, 32'sh26bbb119, 32'sh26b6b070, 32'sh26b1af67, 32'sh26acadff, 32'sh26a7ac38, 32'sh26a2aa11, 32'sh269da78b, 
               32'sh2698a4a6, 32'sh2693a161, 32'sh268e9dbd, 32'sh268999ba, 32'sh26849558, 32'sh267f9097, 32'sh267a8b77, 32'sh267585f8, 
               32'sh2670801a, 32'sh266b79dd, 32'sh26667342, 32'sh26616c48, 32'sh265c64ef, 32'sh26575d37, 32'sh26525521, 32'sh264d4cac, 
               32'sh264843d9, 32'sh26433aa7, 32'sh263e3117, 32'sh26392728, 32'sh26341cdb, 32'sh262f1230, 32'sh262a0727, 32'sh2624fbbf, 
               32'sh261feffa, 32'sh261ae3d6, 32'sh2615d754, 32'sh2610ca75, 32'sh260bbd37, 32'sh2606af9c, 32'sh2601a1a2, 32'sh25fc934b, 
               32'sh25f78497, 32'sh25f27584, 32'sh25ed6614, 32'sh25e85646, 32'sh25e3461b, 32'sh25de3592, 32'sh25d924ac, 32'sh25d41369, 
               32'sh25cf01c8, 32'sh25c9efca, 32'sh25c4dd6e, 32'sh25bfcab6, 32'sh25bab7a0, 32'sh25b5a42d, 32'sh25b0905d, 32'sh25ab7c30, 
               32'sh25a667a7, 32'sh25a152c0, 32'sh259c3d7c, 32'sh259727dc, 32'sh259211df, 32'sh258cfb85, 32'sh2587e4cf, 32'sh2582cdbc, 
               32'sh257db64c, 32'sh25789e80, 32'sh25738657, 32'sh256e6dd2, 32'sh256954f1, 32'sh25643bb3, 32'sh255f2219, 32'sh255a0823, 
               32'sh2554edd1, 32'sh254fd323, 32'sh254ab818, 32'sh25459cb2, 32'sh254080ef, 32'sh253b64d1, 32'sh25364857, 32'sh25312b81, 
               32'sh252c0e4f, 32'sh2526f0c1, 32'sh2521d2d8, 32'sh251cb493, 32'sh251795f3, 32'sh251276f7, 32'sh250d57a0, 32'sh250837ed, 
               32'sh250317df, 32'sh24fdf775, 32'sh24f8d6b0, 32'sh24f3b590, 32'sh24ee9415, 32'sh24e9723f, 32'sh24e4500e, 32'sh24df2d81, 
               32'sh24da0a9a, 32'sh24d4e757, 32'sh24cfc3ba, 32'sh24ca9fc2, 32'sh24c57b6f, 32'sh24c056c2, 32'sh24bb31ba, 32'sh24b60c57, 
               32'sh24b0e699, 32'sh24abc082, 32'sh24a69a0f, 32'sh24a17342, 32'sh249c4c1b, 32'sh24972499, 32'sh2491fcbe, 32'sh248cd487, 
               32'sh2487abf7, 32'sh2482830d, 32'sh247d59c8, 32'sh2478302a, 32'sh24730631, 32'sh246ddbdf, 32'sh2468b132, 32'sh2463862c, 
               32'sh245e5acc, 32'sh24592f13, 32'sh245402ff, 32'sh244ed692, 32'sh2449a9cc, 32'sh24447cac, 32'sh243f4f32, 32'sh243a215f, 
               32'sh2434f332, 32'sh242fc4ad, 32'sh242a95ce, 32'sh24256695, 32'sh24203704, 32'sh241b0719, 32'sh2415d6d5, 32'sh2410a639, 
               32'sh240b7543, 32'sh240643f4, 32'sh2401124d, 32'sh23fbe04c, 32'sh23f6adf3, 32'sh23f17b41, 32'sh23ec4837, 32'sh23e714d3, 
               32'sh23e1e117, 32'sh23dcad03, 32'sh23d77896, 32'sh23d243d1, 32'sh23cd0eb3, 32'sh23c7d93d, 32'sh23c2a36f, 32'sh23bd6d48, 
               32'sh23b836ca, 32'sh23b2fff3, 32'sh23adc8c4, 32'sh23a8913d, 32'sh23a3595e, 32'sh239e2127, 32'sh2398e898, 32'sh2393afb2, 
               32'sh238e7673, 32'sh23893cdd, 32'sh238402ef, 32'sh237ec8aa, 32'sh23798e0d, 32'sh23745318, 32'sh236f17cc, 32'sh2369dc29, 
               32'sh2364a02e, 32'sh235f63dc, 32'sh235a2733, 32'sh2354ea32, 32'sh234facda, 32'sh234a6f2b, 32'sh23453125, 32'sh233ff2c8, 
               32'sh233ab414, 32'sh23357509, 32'sh233035a7, 32'sh232af5ee, 32'sh2325b5df, 32'sh23207579, 32'sh231b34bc, 32'sh2315f3a8, 
               32'sh2310b23e, 32'sh230b707e, 32'sh23062e67, 32'sh2300ebf9, 32'sh22fba936, 32'sh22f6661c, 32'sh22f122ab, 32'sh22ebdee5, 
               32'sh22e69ac8, 32'sh22e15655, 32'sh22dc118c, 32'sh22d6cc6d, 32'sh22d186f8, 32'sh22cc412d, 32'sh22c6fb0c, 32'sh22c1b496, 
               32'sh22bc6dca, 32'sh22b726a8, 32'sh22b1df30, 32'sh22ac9763, 32'sh22a74f40, 32'sh22a206c8, 32'sh229cbdfa, 32'sh229774d7, 
               32'sh22922b5e, 32'sh228ce191, 32'sh2287976e, 32'sh22824cf5, 32'sh227d0228, 32'sh2277b705, 32'sh22726b8e, 32'sh226d1fc1, 
               32'sh2267d3a0, 32'sh22628729, 32'sh225d3a5e, 32'sh2257ed3e, 32'sh22529fca, 32'sh224d5200, 32'sh224803e2, 32'sh2242b56f, 
               32'sh223d66a8, 32'sh2238178d, 32'sh2232c81c, 32'sh222d7858, 32'sh2228283f, 32'sh2222d7d2, 32'sh221d8711, 32'sh221835fb, 
               32'sh2212e492, 32'sh220d92d4, 32'sh220840c2, 32'sh2202ee5d, 32'sh21fd9ba3, 32'sh21f84895, 32'sh21f2f534, 32'sh21eda17f, 
               32'sh21e84d76, 32'sh21e2f91a, 32'sh21dda46a, 32'sh21d84f66, 32'sh21d2fa0f, 32'sh21cda465, 32'sh21c84e67, 32'sh21c2f815, 
               32'sh21bda171, 32'sh21b84a79, 32'sh21b2f32e, 32'sh21ad9b8f, 32'sh21a8439e, 32'sh21a2eb5a, 32'sh219d92c2, 32'sh219839d8, 
               32'sh2192e09b, 32'sh218d870b, 32'sh21882d28, 32'sh2182d2f2, 32'sh217d786a, 32'sh21781d8f, 32'sh2172c262, 32'sh216d66e2, 
               32'sh21680b0f, 32'sh2162aeea, 32'sh215d5273, 32'sh2157f5a9, 32'sh2152988d, 32'sh214d3b1f, 32'sh2147dd5f, 32'sh21427f4d, 
               32'sh213d20e8, 32'sh2137c232, 32'sh21326329, 32'sh212d03cf, 32'sh2127a423, 32'sh21224425, 32'sh211ce3d5, 32'sh21178334, 
               32'sh21122240, 32'sh210cc0fc, 32'sh21075f65, 32'sh2101fd7e, 32'sh20fc9b44, 32'sh20f738ba, 32'sh20f1d5de, 32'sh20ec72b1, 
               32'sh20e70f32, 32'sh20e1ab63, 32'sh20dc4742, 32'sh20d6e2d0, 32'sh20d17e0d, 32'sh20cc18f9, 32'sh20c6b395, 32'sh20c14ddf, 
               32'sh20bbe7d8, 32'sh20b68181, 32'sh20b11ad9, 32'sh20abb3e1, 32'sh20a64c97, 32'sh20a0e4fe, 32'sh209b7d13, 32'sh209614d9, 
               32'sh2090ac4d, 32'sh208b4372, 32'sh2085da46, 32'sh208070ca, 32'sh207b06fe, 32'sh20759ce1, 32'sh20703275, 32'sh206ac7b8, 
               32'sh20655cac, 32'sh205ff14f, 32'sh205a85a3, 32'sh205519a7, 32'sh204fad5b, 32'sh204a40bf, 32'sh2044d3d4, 32'sh203f6699, 
               32'sh2039f90f, 32'sh20348b35, 32'sh202f1d0b, 32'sh2029ae92, 32'sh20243fca, 32'sh201ed0b2, 32'sh2019614c, 32'sh2013f196, 
               32'sh200e8190, 32'sh2009113c, 32'sh2003a099, 32'sh1ffe2fa6, 32'sh1ff8be65, 32'sh1ff34cd5, 32'sh1feddaf6, 32'sh1fe868c8, 
               32'sh1fe2f64c, 32'sh1fdd8381, 32'sh1fd81067, 32'sh1fd29cff, 32'sh1fcd2948, 32'sh1fc7b542, 32'sh1fc240ef, 32'sh1fbccc4d, 
               32'sh1fb7575c, 32'sh1fb1e21d, 32'sh1fac6c91, 32'sh1fa6f6b6, 32'sh1fa1808c, 32'sh1f9c0a15, 32'sh1f969350, 32'sh1f911c3d, 
               32'sh1f8ba4dc, 32'sh1f862d2d, 32'sh1f80b531, 32'sh1f7b3ce6, 32'sh1f75c44e, 32'sh1f704b69, 32'sh1f6ad235, 32'sh1f6558b5, 
               32'sh1f5fdee6, 32'sh1f5a64cb, 32'sh1f54ea62, 32'sh1f4f6fab, 32'sh1f49f4a8, 32'sh1f447957, 32'sh1f3efdb9, 32'sh1f3981ce, 
               32'sh1f340596, 32'sh1f2e8911, 32'sh1f290c3f, 32'sh1f238f20, 32'sh1f1e11b5, 32'sh1f1893fc, 32'sh1f1315f7, 32'sh1f0d97a5, 
               32'sh1f081907, 32'sh1f029a1c, 32'sh1efd1ae4, 32'sh1ef79b60, 32'sh1ef21b90, 32'sh1eec9b73, 32'sh1ee71b0a, 32'sh1ee19a54, 
               32'sh1edc1953, 32'sh1ed69805, 32'sh1ed1166b, 32'sh1ecb9486, 32'sh1ec61254, 32'sh1ec08fd6, 32'sh1ebb0d0d, 32'sh1eb589f7, 
               32'sh1eb00696, 32'sh1eaa82e9, 32'sh1ea4fef0, 32'sh1e9f7aac, 32'sh1e99f61d, 32'sh1e947141, 32'sh1e8eec1b, 32'sh1e8966a8, 
               32'sh1e83e0eb, 32'sh1e7e5ae2, 32'sh1e78d48e, 32'sh1e734def, 32'sh1e6dc705, 32'sh1e683fcf, 32'sh1e62b84f, 32'sh1e5d3084, 
               32'sh1e57a86d, 32'sh1e52200c, 32'sh1e4c9760, 32'sh1e470e69, 32'sh1e418528, 32'sh1e3bfb9c, 32'sh1e3671c5, 32'sh1e30e7a4, 
               32'sh1e2b5d38, 32'sh1e25d282, 32'sh1e204781, 32'sh1e1abc36, 32'sh1e1530a1, 32'sh1e0fa4c2, 32'sh1e0a1898, 32'sh1e048c24, 
               32'sh1dfeff67, 32'sh1df9725f, 32'sh1df3e50d, 32'sh1dee5771, 32'sh1de8c98c, 32'sh1de33b5d, 32'sh1dddace4, 32'sh1dd81e21, 
               32'sh1dd28f15, 32'sh1dccffbf, 32'sh1dc7701f, 32'sh1dc1e036, 32'sh1dbc5004, 32'sh1db6bf88, 32'sh1db12ec3, 32'sh1dab9db5, 
               32'sh1da60c5d, 32'sh1da07abc, 32'sh1d9ae8d2, 32'sh1d9556a0, 32'sh1d8fc424, 32'sh1d8a315f, 32'sh1d849e51, 32'sh1d7f0afb, 
               32'sh1d79775c, 32'sh1d73e374, 32'sh1d6e4f43, 32'sh1d68baca, 32'sh1d632608, 32'sh1d5d90fd, 32'sh1d57fbaa, 32'sh1d52660f, 
               32'sh1d4cd02c, 32'sh1d473a00, 32'sh1d41a38c, 32'sh1d3c0ccf, 32'sh1d3675cb, 32'sh1d30de7e, 32'sh1d2b46ea, 32'sh1d25af0d, 
               32'sh1d2016e9, 32'sh1d1a7e7d, 32'sh1d14e5c9, 32'sh1d0f4ccd, 32'sh1d09b389, 32'sh1d0419fe, 32'sh1cfe802b, 32'sh1cf8e611, 
               32'sh1cf34baf, 32'sh1cedb106, 32'sh1ce81615, 32'sh1ce27add, 32'sh1cdcdf5e, 32'sh1cd74397, 32'sh1cd1a78a, 32'sh1ccc0b35, 
               32'sh1cc66e99, 32'sh1cc0d1b6, 32'sh1cbb348d, 32'sh1cb5971c, 32'sh1caff965, 32'sh1caa5b66, 32'sh1ca4bd21, 32'sh1c9f1e96, 
               32'sh1c997fc4, 32'sh1c93e0ab, 32'sh1c8e414b, 32'sh1c88a1a6, 32'sh1c8301b9, 32'sh1c7d6187, 32'sh1c77c10e, 32'sh1c72204f, 
               32'sh1c6c7f4a, 32'sh1c66ddfe, 32'sh1c613c6d, 32'sh1c5b9a95, 32'sh1c55f878, 32'sh1c505614, 32'sh1c4ab36b, 32'sh1c45107c, 
               32'sh1c3f6d47, 32'sh1c39c9cd, 32'sh1c34260c, 32'sh1c2e8207, 32'sh1c28ddbb, 32'sh1c23392b, 32'sh1c1d9454, 32'sh1c17ef39, 
               32'sh1c1249d8, 32'sh1c0ca432, 32'sh1c06fe46, 32'sh1c015816, 32'sh1bfbb1a0, 32'sh1bf60ae6, 32'sh1bf063e6, 32'sh1beabca1, 
               32'sh1be51518, 32'sh1bdf6d4a, 32'sh1bd9c537, 32'sh1bd41cdf, 32'sh1bce7442, 32'sh1bc8cb61, 32'sh1bc3223c, 32'sh1bbd78d2, 
               32'sh1bb7cf23, 32'sh1bb22530, 32'sh1bac7af9, 32'sh1ba6d07d, 32'sh1ba125bd, 32'sh1b9b7ab9, 32'sh1b95cf71, 32'sh1b9023e5, 
               32'sh1b8a7815, 32'sh1b84cc01, 32'sh1b7f1fa9, 32'sh1b79730d, 32'sh1b73c62d, 32'sh1b6e190a, 32'sh1b686ba3, 32'sh1b62bdf8, 
               32'sh1b5d100a, 32'sh1b5761d8, 32'sh1b51b363, 32'sh1b4c04aa, 32'sh1b4655ae, 32'sh1b40a66f, 32'sh1b3af6ec, 32'sh1b354727, 
               32'sh1b2f971e, 32'sh1b29e6d2, 32'sh1b243643, 32'sh1b1e8571, 32'sh1b18d45c, 32'sh1b132304, 32'sh1b0d716a, 32'sh1b07bf8c, 
               32'sh1b020d6c, 32'sh1afc5b0a, 32'sh1af6a865, 32'sh1af0f57d, 32'sh1aeb4253, 32'sh1ae58ee6, 32'sh1adfdb37, 32'sh1ada2746, 
               32'sh1ad47312, 32'sh1acebe9d, 32'sh1ac909e5, 32'sh1ac354eb, 32'sh1abd9faf, 32'sh1ab7ea31, 32'sh1ab23471, 32'sh1aac7e6f, 
               32'sh1aa6c82b, 32'sh1aa111a6, 32'sh1a9b5adf, 32'sh1a95a3d6, 32'sh1a8fec8c, 32'sh1a8a3500, 32'sh1a847d33, 32'sh1a7ec524, 
               32'sh1a790cd4, 32'sh1a735442, 32'sh1a6d9b70, 32'sh1a67e25c, 32'sh1a622907, 32'sh1a5c6f70, 32'sh1a56b599, 32'sh1a50fb81, 
               32'sh1a4b4128, 32'sh1a45868e, 32'sh1a3fcbb3, 32'sh1a3a1097, 32'sh1a34553b, 32'sh1a2e999e, 32'sh1a28ddc0, 32'sh1a2321a2, 
               32'sh1a1d6544, 32'sh1a17a8a5, 32'sh1a11ebc5, 32'sh1a0c2ea5, 32'sh1a067145, 32'sh1a00b3a5, 32'sh19faf5c5, 32'sh19f537a4, 
               32'sh19ef7944, 32'sh19e9baa3, 32'sh19e3fbc3, 32'sh19de3ca2, 32'sh19d87d42, 32'sh19d2bda2, 32'sh19ccfdc2, 32'sh19c73da3, 
               32'sh19c17d44, 32'sh19bbbca6, 32'sh19b5fbc8, 32'sh19b03aaa, 32'sh19aa794d, 32'sh19a4b7b1, 32'sh199ef5d6, 32'sh199933bb, 
               32'sh19937161, 32'sh198daec8, 32'sh1987ebf0, 32'sh198228d9, 32'sh197c6584, 32'sh1976a1ef, 32'sh1970de1b, 32'sh196b1a09, 
               32'sh196555b8, 32'sh195f9128, 32'sh1959cc5a, 32'sh1954074d, 32'sh194e4201, 32'sh19487c77, 32'sh1942b6af, 32'sh193cf0a9, 
               32'sh19372a64, 32'sh193163e1, 32'sh192b9d1f, 32'sh1925d620, 32'sh19200ee3, 32'sh191a4767, 32'sh19147fae, 32'sh190eb7b7, 
               32'sh1908ef82, 32'sh1903270f, 32'sh18fd5e5f, 32'sh18f79571, 32'sh18f1cc45, 32'sh18ec02db, 32'sh18e63935, 32'sh18e06f50, 
               32'sh18daa52f, 32'sh18d4dad0, 32'sh18cf1034, 32'sh18c9455a, 32'sh18c37a44, 32'sh18bdaef0, 32'sh18b7e35f, 32'sh18b21791, 
               32'sh18ac4b87, 32'sh18a67f3f, 32'sh18a0b2bb, 32'sh189ae5fa, 32'sh189518fc, 32'sh188f4bc2, 32'sh18897e4a, 32'sh1883b097, 
               32'sh187de2a7, 32'sh1878147a, 32'sh18724611, 32'sh186c776c, 32'sh1866a88a, 32'sh1860d96d, 32'sh185b0a13, 32'sh18553a7d, 
               32'sh184f6aab, 32'sh18499a9d, 32'sh1843ca53, 32'sh183df9cd, 32'sh1838290c, 32'sh1832580e, 32'sh182c86d5, 32'sh1826b561, 
               32'sh1820e3b0, 32'sh181b11c4, 32'sh18153f9d, 32'sh180f6d3a, 32'sh18099a9c, 32'sh1803c7c3, 32'sh17fdf4ae, 32'sh17f8215e, 
               32'sh17f24dd3, 32'sh17ec7a0d, 32'sh17e6a60c, 32'sh17e0d1d0, 32'sh17dafd59, 32'sh17d528a7, 32'sh17cf53bb, 32'sh17c97e93, 
               32'sh17c3a931, 32'sh17bdd394, 32'sh17b7fdbd, 32'sh17b227ab, 32'sh17ac515f, 32'sh17a67ad8, 32'sh17a0a417, 32'sh179acd1c, 
               32'sh1794f5e6, 32'sh178f1e76, 32'sh178946cc, 32'sh17836ee8, 32'sh177d96ca, 32'sh1777be72, 32'sh1771e5e0, 32'sh176c0d15, 
               32'sh1766340f, 32'sh17605ad0, 32'sh175a8157, 32'sh1754a7a4, 32'sh174ecdb8, 32'sh1748f393, 32'sh17431933, 32'sh173d3e9b, 
               32'sh173763c9, 32'sh173188be, 32'sh172bad7a, 32'sh1725d1fc, 32'sh171ff646, 32'sh171a1a56, 32'sh17143e2d, 32'sh170e61cc, 
               32'sh17088531, 32'sh1702a85e, 32'sh16fccb51, 32'sh16f6ee0d, 32'sh16f1108f, 32'sh16eb32d9, 32'sh16e554ea, 32'sh16df76c3, 
               32'sh16d99864, 32'sh16d3b9cc, 32'sh16cddafb, 32'sh16c7fbf3, 32'sh16c21cb2, 32'sh16bc3d39, 32'sh16b65d88, 32'sh16b07d9f, 
               32'sh16aa9d7e, 32'sh16a4bd25, 32'sh169edc94, 32'sh1698fbcb, 32'sh16931acb, 32'sh168d3993, 32'sh16875823, 32'sh1681767c, 
               32'sh167b949d, 32'sh1675b286, 32'sh166fd039, 32'sh1669edb3, 32'sh16640af7, 32'sh165e2803, 32'sh165844d8, 32'sh16526176, 
               32'sh164c7ddd, 32'sh16469a0d, 32'sh1640b606, 32'sh163ad1c8, 32'sh1634ed53, 32'sh162f08a8, 32'sh162923c5, 32'sh16233eac, 
               32'sh161d595d, 32'sh161773d6, 32'sh16118e1a, 32'sh160ba826, 32'sh1605c1fd, 32'sh15ffdb9d, 32'sh15f9f507, 32'sh15f40e3a, 
               32'sh15ee2738, 32'sh15e83fff, 32'sh15e25890, 32'sh15dc70eb, 32'sh15d68911, 32'sh15d0a100, 32'sh15cab8ba, 32'sh15c4d03e, 
               32'sh15bee78c, 32'sh15b8fea4, 32'sh15b31587, 32'sh15ad2c34, 32'sh15a742ac, 32'sh15a158ee, 32'sh159b6efb, 32'sh159584d3, 
               32'sh158f9a76, 32'sh1589afe3, 32'sh1583c51b, 32'sh157dda1e, 32'sh1577eeec, 32'sh15720385, 32'sh156c17e9, 32'sh15662c18, 
               32'sh15604013, 32'sh155a53d9, 32'sh1554676a, 32'sh154e7ac6, 32'sh15488dee, 32'sh1542a0e1, 32'sh153cb3a0, 32'sh1536c62b, 
               32'sh1530d881, 32'sh152aeaa3, 32'sh1524fc90, 32'sh151f0e4a, 32'sh15191fcf, 32'sh15133120, 32'sh150d423d, 32'sh15075327, 
               32'sh150163dc, 32'sh14fb745e, 32'sh14f584ac, 32'sh14ef94c6, 32'sh14e9a4ac, 32'sh14e3b45f, 32'sh14ddc3de, 32'sh14d7d32a, 
               32'sh14d1e242, 32'sh14cbf127, 32'sh14c5ffd9, 32'sh14c00e58, 32'sh14ba1ca3, 32'sh14b42abb, 32'sh14ae38a0, 32'sh14a84652, 
               32'sh14a253d1, 32'sh149c611d, 32'sh14966e36, 32'sh14907b1d, 32'sh148a87d1, 32'sh14849452, 32'sh147ea0a0, 32'sh1478acbc, 
               32'sh1472b8a5, 32'sh146cc45c, 32'sh1466cfe1, 32'sh1460db33, 32'sh145ae653, 32'sh1454f140, 32'sh144efbfc, 32'sh14490685, 
               32'sh144310dd, 32'sh143d1b02, 32'sh143724f5, 32'sh14312eb7, 32'sh142b3846, 32'sh142541a4, 32'sh141f4ad1, 32'sh141953cb, 
               32'sh14135c94, 32'sh140d652c, 32'sh14076d91, 32'sh140175c6, 32'sh13fb7dc9, 32'sh13f5859b, 32'sh13ef8d3c, 32'sh13e994ab, 
               32'sh13e39be9, 32'sh13dda2f7, 32'sh13d7a9d3, 32'sh13d1b07e, 32'sh13cbb6f8, 32'sh13c5bd42, 32'sh13bfc35b, 32'sh13b9c943, 
               32'sh13b3cefa, 32'sh13add481, 32'sh13a7d9d7, 32'sh13a1defd, 32'sh139be3f2, 32'sh1395e8b7, 32'sh138fed4b, 32'sh1389f1af, 
               32'sh1383f5e3, 32'sh137df9e7, 32'sh1377fdbb, 32'sh1372015f, 32'sh136c04d2, 32'sh13660816, 32'sh13600b2a, 32'sh135a0e0e, 
               32'sh135410c3, 32'sh134e1348, 32'sh1348159d, 32'sh134217c2, 32'sh133c19b8, 32'sh13361b7f, 32'sh13301d16, 32'sh132a1e7e, 
               32'sh13241fb6, 32'sh131e20c0, 32'sh1318219a, 32'sh13122245, 32'sh130c22c1, 32'sh1306230d, 32'sh1300232c, 32'sh12fa231b, 
               32'sh12f422db, 32'sh12ee226c, 32'sh12e821cf, 32'sh12e22103, 32'sh12dc2009, 32'sh12d61ee0, 32'sh12d01d89, 32'sh12ca1c03, 
               32'sh12c41a4f, 32'sh12be186c, 32'sh12b8165b, 32'sh12b2141c, 32'sh12ac11af, 32'sh12a60f14, 32'sh12a00c4b, 32'sh129a0954, 
               32'sh1294062f, 32'sh128e02dc, 32'sh1287ff5b, 32'sh1281fbad, 32'sh127bf7d1, 32'sh1275f3c7, 32'sh126fef90, 32'sh1269eb2b, 
               32'sh1263e699, 32'sh125de1da, 32'sh1257dced, 32'sh1251d7d3, 32'sh124bd28c, 32'sh1245cd17, 32'sh123fc776, 32'sh1239c1a7, 
               32'sh1233bbac, 32'sh122db583, 32'sh1227af2e, 32'sh1221a8ac, 32'sh121ba1fd, 32'sh12159b22, 32'sh120f941a, 32'sh12098ce5, 
               32'sh12038584, 32'sh11fd7df6, 32'sh11f7763c, 32'sh11f16e56, 32'sh11eb6643, 32'sh11e55e04, 32'sh11df5599, 32'sh11d94d02, 
               32'sh11d3443f, 32'sh11cd3b50, 32'sh11c73235, 32'sh11c128ee, 32'sh11bb1f7c, 32'sh11b515dd, 32'sh11af0c13, 32'sh11a9021d, 
               32'sh11a2f7fc, 32'sh119cedaf, 32'sh1196e337, 32'sh1190d893, 32'sh118acdc4, 32'sh1184c2ca, 32'sh117eb7a4, 32'sh1178ac53, 
               32'sh1172a0d7, 32'sh116c9531, 32'sh1166895f, 32'sh11607d62, 32'sh115a713a, 32'sh115464e8, 32'sh114e586a, 32'sh11484bc2, 
               32'sh11423ef0, 32'sh113c31f3, 32'sh113624cb, 32'sh11301779, 32'sh112a09fc, 32'sh1123fc55, 32'sh111dee84, 32'sh1117e088, 
               32'sh1111d263, 32'sh110bc413, 32'sh1105b599, 32'sh10ffa6f5, 32'sh10f99827, 32'sh10f38930, 32'sh10ed7a0e, 32'sh10e76ac3, 
               32'sh10e15b4e, 32'sh10db4baf, 32'sh10d53be7, 32'sh10cf2bf6, 32'sh10c91bda, 32'sh10c30b96, 32'sh10bcfb28, 32'sh10b6ea90, 
               32'sh10b0d9d0, 32'sh10aac8e6, 32'sh10a4b7d3, 32'sh109ea697, 32'sh10989532, 32'sh109283a5, 32'sh108c71ee, 32'sh1086600e, 
               32'sh10804e06, 32'sh107a3bd5, 32'sh1074297b, 32'sh106e16f9, 32'sh1068044e, 32'sh1061f17b, 32'sh105bde7f, 32'sh1055cb5b, 
               32'sh104fb80e, 32'sh1049a49a, 32'sh104390fd, 32'sh103d7d38, 32'sh1037694b, 32'sh10315535, 32'sh102b40f8, 32'sh10252c94, 
               32'sh101f1807, 32'sh10190352, 32'sh1012ee76, 32'sh100cd972, 32'sh1006c446, 32'sh1000aef3, 32'sh0ffa9979, 32'sh0ff483d7, 
               32'sh0fee6e0d, 32'sh0fe8581d, 32'sh0fe24205, 32'sh0fdc2bc6, 32'sh0fd6155f, 32'sh0fcffed2, 32'sh0fc9e81e, 32'sh0fc3d143, 
               32'sh0fbdba40, 32'sh0fb7a317, 32'sh0fb18bc8, 32'sh0fab7451, 32'sh0fa55cb4, 32'sh0f9f44f0, 32'sh0f992d06, 32'sh0f9314f5, 
               32'sh0f8cfcbe, 32'sh0f86e460, 32'sh0f80cbdc, 32'sh0f7ab332, 32'sh0f749a61, 32'sh0f6e816b, 32'sh0f68684e, 32'sh0f624f0c, 
               32'sh0f5c35a3, 32'sh0f561c15, 32'sh0f500260, 32'sh0f49e886, 32'sh0f43ce86, 32'sh0f3db461, 32'sh0f379a16, 32'sh0f317fa5, 
               32'sh0f2b650f, 32'sh0f254a53, 32'sh0f1f2f73, 32'sh0f19146c, 32'sh0f12f941, 32'sh0f0cddf0, 32'sh0f06c27a, 32'sh0f00a6df, 
               32'sh0efa8b20, 32'sh0ef46f3b, 32'sh0eee5331, 32'sh0ee83702, 32'sh0ee21aaf, 32'sh0edbfe37, 32'sh0ed5e19a, 32'sh0ecfc4d9, 
               32'sh0ec9a7f3, 32'sh0ec38ae8, 32'sh0ebd6db9, 32'sh0eb75066, 32'sh0eb132ef, 32'sh0eab1553, 32'sh0ea4f793, 32'sh0e9ed9af, 
               32'sh0e98bba7, 32'sh0e929d7a, 32'sh0e8c7f2a, 32'sh0e8660b6, 32'sh0e80421e, 32'sh0e7a2363, 32'sh0e740483, 32'sh0e6de580, 
               32'sh0e67c65a, 32'sh0e61a70f, 32'sh0e5b87a2, 32'sh0e556811, 32'sh0e4f485c, 32'sh0e492884, 32'sh0e430889, 32'sh0e3ce86b, 
               32'sh0e36c82a, 32'sh0e30a7c5, 32'sh0e2a873e, 32'sh0e246693, 32'sh0e1e45c6, 32'sh0e1824d6, 32'sh0e1203c3, 32'sh0e0be28e, 
               32'sh0e05c135, 32'sh0dff9fba, 32'sh0df97e1d, 32'sh0df35c5d, 32'sh0ded3a7b, 32'sh0de71876, 32'sh0de0f64f, 32'sh0ddad406, 
               32'sh0dd4b19a, 32'sh0dce8f0d, 32'sh0dc86c5d, 32'sh0dc2498c, 32'sh0dbc2698, 32'sh0db60383, 32'sh0dafe04b, 32'sh0da9bcf2, 
               32'sh0da39978, 32'sh0d9d75db, 32'sh0d97521d, 32'sh0d912e3e, 32'sh0d8b0a3d, 32'sh0d84e61a, 32'sh0d7ec1d6, 32'sh0d789d71, 
               32'sh0d7278eb, 32'sh0d6c5443, 32'sh0d662f7b, 32'sh0d600a91, 32'sh0d59e586, 32'sh0d53c05b, 32'sh0d4d9b0e, 32'sh0d4775a1, 
               32'sh0d415013, 32'sh0d3b2a64, 32'sh0d350495, 32'sh0d2edea5, 32'sh0d28b894, 32'sh0d229263, 32'sh0d1c6c11, 32'sh0d1645a0, 
               32'sh0d101f0e, 32'sh0d09f85b, 32'sh0d03d189, 32'sh0cfdaa96, 32'sh0cf78383, 32'sh0cf15c51, 32'sh0ceb34fe, 32'sh0ce50d8c, 
               32'sh0cdee5f9, 32'sh0cd8be47, 32'sh0cd29676, 32'sh0ccc6e84, 32'sh0cc64673, 32'sh0cc01e43, 32'sh0cb9f5f3, 32'sh0cb3cd84, 
               32'sh0cada4f5, 32'sh0ca77c47, 32'sh0ca1537a, 32'sh0c9b2a8d, 32'sh0c950182, 32'sh0c8ed857, 32'sh0c88af0e, 32'sh0c8285a5, 
               32'sh0c7c5c1e, 32'sh0c763278, 32'sh0c7008b3, 32'sh0c69ded0, 32'sh0c63b4ce, 32'sh0c5d8aad, 32'sh0c57606e, 32'sh0c513610, 
               32'sh0c4b0b94, 32'sh0c44e0f9, 32'sh0c3eb641, 32'sh0c388b6a, 32'sh0c326075, 32'sh0c2c3562, 32'sh0c260a31, 32'sh0c1fdee1, 
               32'sh0c19b374, 32'sh0c1387e9, 32'sh0c0d5c41, 32'sh0c07307a, 32'sh0c010496, 32'sh0bfad894, 32'sh0bf4ac75, 32'sh0bee8038, 
               32'sh0be853de, 32'sh0be22766, 32'sh0bdbfad1, 32'sh0bd5ce1f, 32'sh0bcfa150, 32'sh0bc97463, 32'sh0bc34759, 32'sh0bbd1a33, 
               32'sh0bb6ecef, 32'sh0bb0bf8f, 32'sh0baa9211, 32'sh0ba46477, 32'sh0b9e36c0, 32'sh0b9808ed, 32'sh0b91dafc, 32'sh0b8bacf0, 
               32'sh0b857ec7, 32'sh0b7f5081, 32'sh0b79221f, 32'sh0b72f3a1, 32'sh0b6cc506, 32'sh0b66964f, 32'sh0b60677c, 32'sh0b5a388d, 
               32'sh0b540982, 32'sh0b4dda5c, 32'sh0b47ab19, 32'sh0b417bba, 32'sh0b3b4c40, 32'sh0b351caa, 32'sh0b2eecf8, 32'sh0b28bd2a, 
               32'sh0b228d42, 32'sh0b1c5d3d, 32'sh0b162d1d, 32'sh0b0ffce2, 32'sh0b09cc8c, 32'sh0b039c1a, 32'sh0afd6b8d, 32'sh0af73ae5, 
               32'sh0af10a22, 32'sh0aead944, 32'sh0ae4a84b, 32'sh0ade7737, 32'sh0ad84609, 32'sh0ad214bf, 32'sh0acbe35b, 32'sh0ac5b1dc, 
               32'sh0abf8043, 32'sh0ab94e8f, 32'sh0ab31cc1, 32'sh0aacead8, 32'sh0aa6b8d5, 32'sh0aa086b8, 32'sh0a9a5480, 32'sh0a94222f, 
               32'sh0a8defc3, 32'sh0a87bd3d, 32'sh0a818a9d, 32'sh0a7b57e3, 32'sh0a752510, 32'sh0a6ef222, 32'sh0a68bf1b, 32'sh0a628bfa, 
               32'sh0a5c58c0, 32'sh0a56256c, 32'sh0a4ff1fe, 32'sh0a49be77, 32'sh0a438ad7, 32'sh0a3d571d, 32'sh0a37234a, 32'sh0a30ef5e, 
               32'sh0a2abb59, 32'sh0a24873a, 32'sh0a1e5303, 32'sh0a181eb2, 32'sh0a11ea49, 32'sh0a0bb5c7, 32'sh0a05812c, 32'sh09ff4c78, 
               32'sh09f917ac, 32'sh09f2e2c7, 32'sh09ecadc9, 32'sh09e678b4, 32'sh09e04385, 32'sh09da0e3e, 32'sh09d3d8df, 32'sh09cda368, 
               32'sh09c76dd8, 32'sh09c13831, 32'sh09bb0271, 32'sh09b4cc99, 32'sh09ae96aa, 32'sh09a860a2, 32'sh09a22a83, 32'sh099bf44c, 
               32'sh0995bdfd, 32'sh098f8796, 32'sh09895118, 32'sh09831a82, 32'sh097ce3d5, 32'sh0976ad11, 32'sh09707635, 32'sh096a3f42, 
               32'sh09640837, 32'sh095dd116, 32'sh095799dd, 32'sh0951628d, 32'sh094b2b27, 32'sh0944f3a9, 32'sh093ebc14, 32'sh09388469, 
               32'sh09324ca7, 32'sh092c14ce, 32'sh0925dcdf, 32'sh091fa4d9, 32'sh09196cbc, 32'sh09133489, 32'sh090cfc40, 32'sh0906c3e0, 
               32'sh09008b6a, 32'sh08fa52de, 32'sh08f41a3c, 32'sh08ede184, 32'sh08e7a8b5, 32'sh08e16fd1, 32'sh08db36d6, 32'sh08d4fdc6, 
               32'sh08cec4a0, 32'sh08c88b65, 32'sh08c25213, 32'sh08bc18ac, 32'sh08b5df30, 32'sh08afa59e, 32'sh08a96bf6, 32'sh08a3323a, 
               32'sh089cf867, 32'sh0896be80, 32'sh08908483, 32'sh088a4a72, 32'sh0884104b, 32'sh087dd60f, 32'sh08779bbe, 32'sh08716159, 
               32'sh086b26de, 32'sh0864ec4f, 32'sh085eb1ab, 32'sh085876f3, 32'sh08523c25, 32'sh084c0144, 32'sh0845c64d, 32'sh083f8b43, 
               32'sh08395024, 32'sh083314f1, 32'sh082cd9a9, 32'sh08269e4d, 32'sh082062de, 32'sh081a275a, 32'sh0813ebc2, 32'sh080db016, 
               32'sh08077457, 32'sh08013883, 32'sh07fafc9c, 32'sh07f4c0a1, 32'sh07ee8493, 32'sh07e84871, 32'sh07e20c3b, 32'sh07dbcff2, 
               32'sh07d59396, 32'sh07cf5726, 32'sh07c91aa3, 32'sh07c2de0d, 32'sh07bca163, 32'sh07b664a7, 32'sh07b027d7, 32'sh07a9eaf5, 
               32'sh07a3adff, 32'sh079d70f7, 32'sh079733dc, 32'sh0790f6ae, 32'sh078ab96e, 32'sh07847c1b, 32'sh077e3eb5, 32'sh0778013d, 
               32'sh0771c3b3, 32'sh076b8616, 32'sh07654867, 32'sh075f0aa5, 32'sh0758ccd2, 32'sh07528eec, 32'sh074c50f4, 32'sh074612eb, 
               32'sh073fd4cf, 32'sh073996a1, 32'sh07335862, 32'sh072d1a10, 32'sh0726dbae, 32'sh07209d39, 32'sh071a5eb3, 32'sh0714201b, 
               32'sh070de172, 32'sh0707a2b7, 32'sh070163eb, 32'sh06fb250e, 32'sh06f4e620, 32'sh06eea720, 32'sh06e86810, 32'sh06e228ee, 
               32'sh06dbe9bb, 32'sh06d5aa77, 32'sh06cf6b23, 32'sh06c92bbe, 32'sh06c2ec48, 32'sh06bcacc1, 32'sh06b66d29, 32'sh06b02d81, 
               32'sh06a9edc9, 32'sh06a3ae00, 32'sh069d6e27, 32'sh06972e3d, 32'sh0690ee44, 32'sh068aae3a, 32'sh06846e1f, 32'sh067e2df5, 
               32'sh0677edbb, 32'sh0671ad71, 32'sh066b6d16, 32'sh06652cac, 32'sh065eec33, 32'sh0658aba9, 32'sh06526b10, 32'sh064c2a67, 
               32'sh0645e9af, 32'sh063fa8e7, 32'sh06396810, 32'sh0633272a, 32'sh062ce634, 32'sh0626a52f, 32'sh0620641a, 32'sh061a22f7, 
               32'sh0613e1c5, 32'sh060da083, 32'sh06075f33, 32'sh06011dd4, 32'sh05fadc66, 32'sh05f49ae9, 32'sh05ee595d, 32'sh05e817c3, 
               32'sh05e1d61b, 32'sh05db9463, 32'sh05d5529e, 32'sh05cf10ca, 32'sh05c8cee7, 32'sh05c28cf7, 32'sh05bc4af8, 32'sh05b608eb, 
               32'sh05afc6d0, 32'sh05a984a6, 32'sh05a3426f, 32'sh059d002a, 32'sh0596bdd7, 32'sh05907b77, 32'sh058a3908, 32'sh0583f68c, 
               32'sh057db403, 32'sh0577716b, 32'sh05712ec7, 32'sh056aec15, 32'sh0564a955, 32'sh055e6688, 32'sh055823ae, 32'sh0551e0c7, 
               32'sh054b9dd3, 32'sh05455ad1, 32'sh053f17c3, 32'sh0538d4a7, 32'sh0532917f, 32'sh052c4e4a, 32'sh05260b08, 32'sh051fc7b9, 
               32'sh0519845e, 32'sh051340f6, 32'sh050cfd82, 32'sh0506ba01, 32'sh05007674, 32'sh04fa32db, 32'sh04f3ef35, 32'sh04edab83, 
               32'sh04e767c5, 32'sh04e123fa, 32'sh04dae024, 32'sh04d49c42, 32'sh04ce5854, 32'sh04c81459, 32'sh04c1d054, 32'sh04bb8c42, 
               32'sh04b54825, 32'sh04af03fc, 32'sh04a8bfc7, 32'sh04a27b87, 32'sh049c373c, 32'sh0495f2e5, 32'sh048fae83, 32'sh04896a16, 
               32'sh0483259d, 32'sh047ce11a, 32'sh04769c8b, 32'sh047057f1, 32'sh046a134c, 32'sh0463ce9d, 32'sh045d89e2, 32'sh0457451d, 
               32'sh0451004d, 32'sh044abb73, 32'sh0444768d, 32'sh043e319e, 32'sh0437eca4, 32'sh0431a79f, 32'sh042b6290, 32'sh04251d77, 
               32'sh041ed854, 32'sh04189326, 32'sh04124dee, 32'sh040c08ad, 32'sh0405c361, 32'sh03ff7e0b, 32'sh03f938ac, 32'sh03f2f342, 
               32'sh03ecadcf, 32'sh03e66852, 32'sh03e022cc, 32'sh03d9dd3c, 32'sh03d397a3, 32'sh03cd5200, 32'sh03c70c54, 32'sh03c0c69e, 
               32'sh03ba80df, 32'sh03b43b17, 32'sh03adf546, 32'sh03a7af6c, 32'sh03a16988, 32'sh039b239c, 32'sh0394dda7, 32'sh038e97a9, 
               32'sh038851a2, 32'sh03820b93, 32'sh037bc57b, 32'sh03757f5a, 32'sh036f3931, 32'sh0368f2ff, 32'sh0362acc5, 32'sh035c6682, 
               32'sh03562038, 32'sh034fd9e5, 32'sh03499389, 32'sh03434d26, 32'sh033d06bb, 32'sh0336c047, 32'sh033079cc, 32'sh032a3349, 
               32'sh0323ecbe, 32'sh031da62b, 32'sh03175f91, 32'sh031118ef, 32'sh030ad245, 32'sh03048b94, 32'sh02fe44dc, 32'sh02f7fe1c, 
               32'sh02f1b755, 32'sh02eb7086, 32'sh02e529b0, 32'sh02dee2d4, 32'sh02d89bf0, 32'sh02d25505, 32'sh02cc0e13, 32'sh02c5c71a, 
               32'sh02bf801a, 32'sh02b93914, 32'sh02b2f207, 32'sh02acaaf3, 32'sh02a663d8, 32'sh02a01cb8, 32'sh0299d590, 32'sh02938e62, 
               32'sh028d472e, 32'sh0286fff3, 32'sh0280b8b3, 32'sh027a716c, 32'sh02742a1f, 32'sh026de2cc, 32'sh02679b73, 32'sh02615414, 
               32'sh025b0caf, 32'sh0254c544, 32'sh024e7dd4, 32'sh0248365d, 32'sh0241eee2, 32'sh023ba760, 32'sh02355fd9, 32'sh022f184d, 
               32'sh0228d0bb, 32'sh02228924, 32'sh021c4188, 32'sh0215f9e7, 32'sh020fb240, 32'sh02096a94, 32'sh020322e3, 32'sh01fcdb2e, 
               32'sh01f69373, 32'sh01f04bb4, 32'sh01ea03ef, 32'sh01e3bc26, 32'sh01dd7459, 32'sh01d72c87, 32'sh01d0e4b0, 32'sh01ca9cd4, 
               32'sh01c454f5, 32'sh01be0d11, 32'sh01b7c528, 32'sh01b17d3c, 32'sh01ab354b, 32'sh01a4ed56, 32'sh019ea55d, 32'sh01985d60, 
               32'sh0192155f, 32'sh018bcd5b, 32'sh01858552, 32'sh017f3d46, 32'sh0178f536, 32'sh0172ad22, 32'sh016c650b, 32'sh01661cf0, 
               32'sh015fd4d2, 32'sh01598cb1, 32'sh0153448c, 32'sh014cfc63, 32'sh0146b438, 32'sh01406c0a, 32'sh013a23d8, 32'sh0133dba3, 
               32'sh012d936c, 32'sh01274b31, 32'sh012102f4, 32'sh011abab4, 32'sh01147271, 32'sh010e2a2b, 32'sh0107e1e3, 32'sh01019998, 
               32'sh00fb514b, 32'sh00f508fc, 32'sh00eec0aa, 32'sh00e87856, 32'sh00e22fff, 32'sh00dbe7a6, 32'sh00d59f4c, 32'sh00cf56ef, 
               32'sh00c90e90, 32'sh00c2c62f, 32'sh00bc7dcc, 32'sh00b63568, 32'sh00afed02, 32'sh00a9a49a, 32'sh00a35c30, 32'sh009d13c5, 
               32'sh0096cb58, 32'sh009082ea, 32'sh008a3a7b, 32'sh0083f20a, 32'sh007da998, 32'sh00776125, 32'sh007118b0, 32'sh006ad03b, 
               32'sh006487c4, 32'sh005e3f4c, 32'sh0057f6d4, 32'sh0051ae5b, 32'sh004b65e1, 32'sh00451d66, 32'sh003ed4ea, 32'sh00388c6e, 
               32'sh003243f1, 32'sh002bfb74, 32'sh0025b2f7, 32'sh001f6a79, 32'sh001921fb, 32'sh0012d97c, 32'sh000c90fe, 32'sh0006487f, 
               32'sh00000000, 32'shfff9b781, 32'shfff36f02, 32'shffed2684, 32'shffe6de05, 32'shffe09587, 32'shffda4d09, 32'shffd4048c, 
               32'shffcdbc0f, 32'shffc77392, 32'shffc12b16, 32'shffbae29a, 32'shffb49a1f, 32'shffae51a5, 32'shffa8092c, 32'shffa1c0b4, 
               32'shff9b783c, 32'shff952fc5, 32'shff8ee750, 32'shff889edb, 32'shff825668, 32'shff7c0df6, 32'shff75c585, 32'shff6f7d16, 
               32'shff6934a8, 32'shff62ec3b, 32'shff5ca3d0, 32'shff565b66, 32'shff5012fe, 32'shff49ca98, 32'shff438234, 32'shff3d39d1, 
               32'shff36f170, 32'shff30a911, 32'shff2a60b4, 32'shff24185a, 32'shff1dd001, 32'shff1787aa, 32'shff113f56, 32'shff0af704, 
               32'shff04aeb5, 32'shfefe6668, 32'shfef81e1d, 32'shfef1d5d5, 32'shfeeb8d8f, 32'shfee5454c, 32'shfedefd0c, 32'shfed8b4cf, 
               32'shfed26c94, 32'shfecc245d, 32'shfec5dc28, 32'shfebf93f6, 32'shfeb94bc8, 32'shfeb3039d, 32'shfeacbb74, 32'shfea6734f, 
               32'shfea02b2e, 32'shfe99e310, 32'shfe939af5, 32'shfe8d52de, 32'shfe870aca, 32'shfe80c2ba, 32'shfe7a7aae, 32'shfe7432a5, 
               32'shfe6deaa1, 32'shfe67a2a0, 32'shfe615aa3, 32'shfe5b12aa, 32'shfe54cab5, 32'shfe4e82c4, 32'shfe483ad8, 32'shfe41f2ef, 
               32'shfe3bab0b, 32'shfe35632c, 32'shfe2f1b50, 32'shfe28d379, 32'shfe228ba7, 32'shfe1c43da, 32'shfe15fc11, 32'shfe0fb44c, 
               32'shfe096c8d, 32'shfe0324d2, 32'shfdfcdd1d, 32'shfdf6956c, 32'shfdf04dc0, 32'shfdea0619, 32'shfde3be78, 32'shfddd76dc, 
               32'shfdd72f45, 32'shfdd0e7b3, 32'shfdcaa027, 32'shfdc458a0, 32'shfdbe111e, 32'shfdb7c9a3, 32'shfdb1822c, 32'shfdab3abc, 
               32'shfda4f351, 32'shfd9eabec, 32'shfd98648d, 32'shfd921d34, 32'shfd8bd5e1, 32'shfd858e94, 32'shfd7f474d, 32'shfd79000d, 
               32'shfd72b8d2, 32'shfd6c719e, 32'shfd662a70, 32'shfd5fe348, 32'shfd599c28, 32'shfd53550d, 32'shfd4d0df9, 32'shfd46c6ec, 
               32'shfd407fe6, 32'shfd3a38e6, 32'shfd33f1ed, 32'shfd2daafb, 32'shfd276410, 32'shfd211d2c, 32'shfd1ad650, 32'shfd148f7a, 
               32'shfd0e48ab, 32'shfd0801e4, 32'shfd01bb24, 32'shfcfb746c, 32'shfcf52dbb, 32'shfceee711, 32'shfce8a06f, 32'shfce259d5, 
               32'shfcdc1342, 32'shfcd5ccb7, 32'shfccf8634, 32'shfcc93fb9, 32'shfcc2f945, 32'shfcbcb2da, 32'shfcb66c77, 32'shfcb0261b, 
               32'shfca9dfc8, 32'shfca3997e, 32'shfc9d533b, 32'shfc970d01, 32'shfc90c6cf, 32'shfc8a80a6, 32'shfc843a85, 32'shfc7df46d, 
               32'shfc77ae5e, 32'shfc716857, 32'shfc6b2259, 32'shfc64dc64, 32'shfc5e9678, 32'shfc585094, 32'shfc520aba, 32'shfc4bc4e9, 
               32'shfc457f21, 32'shfc3f3962, 32'shfc38f3ac, 32'shfc32ae00, 32'shfc2c685d, 32'shfc2622c4, 32'shfc1fdd34, 32'shfc1997ae, 
               32'shfc135231, 32'shfc0d0cbe, 32'shfc06c754, 32'shfc0081f5, 32'shfbfa3c9f, 32'shfbf3f753, 32'shfbedb212, 32'shfbe76cda, 
               32'shfbe127ac, 32'shfbdae289, 32'shfbd49d70, 32'shfbce5861, 32'shfbc8135c, 32'shfbc1ce62, 32'shfbbb8973, 32'shfbb5448d, 
               32'shfbaeffb3, 32'shfba8bae3, 32'shfba2761e, 32'shfb9c3163, 32'shfb95ecb4, 32'shfb8fa80f, 32'shfb896375, 32'shfb831ee6, 
               32'shfb7cda63, 32'shfb7695ea, 32'shfb70517d, 32'shfb6a0d1b, 32'shfb63c8c4, 32'shfb5d8479, 32'shfb574039, 32'shfb50fc04, 
               32'shfb4ab7db, 32'shfb4473be, 32'shfb3e2fac, 32'shfb37eba7, 32'shfb31a7ac, 32'shfb2b63be, 32'shfb251fdc, 32'shfb1edc06, 
               32'shfb18983b, 32'shfb12547d, 32'shfb0c10cb, 32'shfb05cd25, 32'shfaff898c, 32'shfaf945ff, 32'shfaf3027e, 32'shfaecbf0a, 
               32'shfae67ba2, 32'shfae03847, 32'shfad9f4f8, 32'shfad3b1b6, 32'shfacd6e81, 32'shfac72b59, 32'shfac0e83d, 32'shfabaa52f, 
               32'shfab4622d, 32'shfaae1f39, 32'shfaa7dc52, 32'shfaa19978, 32'shfa9b56ab, 32'shfa9513eb, 32'shfa8ed139, 32'shfa888e95, 
               32'shfa824bfd, 32'shfa7c0974, 32'shfa75c6f8, 32'shfa6f8489, 32'shfa694229, 32'shfa62ffd6, 32'shfa5cbd91, 32'shfa567b5a, 
               32'shfa503930, 32'shfa49f715, 32'shfa43b508, 32'shfa3d7309, 32'shfa373119, 32'shfa30ef36, 32'shfa2aad62, 32'shfa246b9d, 
               32'shfa1e29e5, 32'shfa17e83d, 32'shfa11a6a3, 32'shfa0b6517, 32'shfa05239a, 32'shf9fee22c, 32'shf9f8a0cd, 32'shf9f25f7d, 
               32'shf9ec1e3b, 32'shf9e5dd09, 32'shf9df9be6, 32'shf9d95ad1, 32'shf9d319cc, 32'shf9ccd8d6, 32'shf9c697f0, 32'shf9c05719, 
               32'shf9ba1651, 32'shf9b3d599, 32'shf9ad94f0, 32'shf9a75457, 32'shf9a113cd, 32'shf99ad354, 32'shf99492ea, 32'shf98e528f, 
               32'shf9881245, 32'shf981d20b, 32'shf97b91e1, 32'shf97551c6, 32'shf96f11bc, 32'shf968d1c3, 32'shf96291d9, 32'shf95c5200, 
               32'shf9561237, 32'shf94fd27f, 32'shf94992d7, 32'shf943533f, 32'shf93d13b8, 32'shf936d442, 32'shf93094dd, 32'shf92a5589, 
               32'shf9241645, 32'shf91dd712, 32'shf91797f0, 32'shf91158e0, 32'shf90b19e0, 32'shf904daf2, 32'shf8fe9c15, 32'shf8f85d49, 
               32'shf8f21e8e, 32'shf8ebdfe5, 32'shf8e5a14d, 32'shf8df62c7, 32'shf8d92452, 32'shf8d2e5f0, 32'shf8cca79e, 32'shf8c6695f, 
               32'shf8c02b31, 32'shf8b9ed15, 32'shf8b3af0c, 32'shf8ad7114, 32'shf8a7332e, 32'shf8a0f55b, 32'shf89ab799, 32'shf89479ea, 
               32'shf88e3c4d, 32'shf887fec3, 32'shf881c14b, 32'shf87b83e5, 32'shf8754692, 32'shf86f0952, 32'shf868cc24, 32'shf8628f09, 
               32'shf85c5201, 32'shf856150b, 32'shf84fd829, 32'shf8499b59, 32'shf8435e9d, 32'shf83d21f3, 32'shf836e55d, 32'shf830a8da, 
               32'shf82a6c6a, 32'shf824300e, 32'shf81df3c5, 32'shf817b78f, 32'shf8117b6d, 32'shf80b3f5f, 32'shf8050364, 32'shf7fec77d, 
               32'shf7f88ba9, 32'shf7f24fea, 32'shf7ec143e, 32'shf7e5d8a6, 32'shf7df9d22, 32'shf7d961b3, 32'shf7d32657, 32'shf7cceb0f, 
               32'shf7c6afdc, 32'shf7c074bd, 32'shf7ba39b3, 32'shf7b3febc, 32'shf7adc3db, 32'shf7a7890d, 32'shf7a14e55, 32'shf79b13b1, 
               32'shf794d922, 32'shf78e9ea7, 32'shf7886442, 32'shf78229f1, 32'shf77befb5, 32'shf775b58e, 32'shf76f7b7d, 32'shf7694180, 
               32'shf7630799, 32'shf75ccdc6, 32'shf756940a, 32'shf7505a62, 32'shf74a20d0, 32'shf743e754, 32'shf73daded, 32'shf737749b, 
               32'shf7313b60, 32'shf72b023a, 32'shf724c92a, 32'shf71e902f, 32'shf718574b, 32'shf7121e7c, 32'shf70be5c4, 32'shf705ad22, 
               32'shf6ff7496, 32'shf6f93c20, 32'shf6f303c0, 32'shf6eccb77, 32'shf6e69344, 32'shf6e05b27, 32'shf6da2321, 32'shf6d3eb32, 
               32'shf6cdb359, 32'shf6c77b97, 32'shf6c143ec, 32'shf6bb0c57, 32'shf6b4d4d9, 32'shf6ae9d73, 32'shf6a86623, 32'shf6a22eea, 
               32'shf69bf7c9, 32'shf695c0be, 32'shf68f89cb, 32'shf68952ef, 32'shf6831c2b, 32'shf67ce57e, 32'shf676aee8, 32'shf670786a, 
               32'shf66a4203, 32'shf6640bb4, 32'shf65dd57d, 32'shf6579f5e, 32'shf6516956, 32'shf64b3367, 32'shf644fd8f, 32'shf63ec7cf, 
               32'shf6389228, 32'shf6325c98, 32'shf62c2721, 32'shf625f1c2, 32'shf61fbc7b, 32'shf619874c, 32'shf6135237, 32'shf60d1d39, 
               32'shf606e854, 32'shf600b388, 32'shf5fa7ed4, 32'shf5f44a39, 32'shf5ee15b7, 32'shf5e7e14e, 32'shf5e1acfd, 32'shf5db78c6, 
               32'shf5d544a7, 32'shf5cf10a2, 32'shf5c8dcb6, 32'shf5c2a8e3, 32'shf5bc7529, 32'shf5b64189, 32'shf5b00e02, 32'shf5a9da94, 
               32'shf5a3a740, 32'shf59d7406, 32'shf59740e5, 32'shf5910dde, 32'shf58adaf0, 32'shf584a81d, 32'shf57e7563, 32'shf57842c3, 
               32'shf572103d, 32'shf56bddd1, 32'shf565ab80, 32'shf55f7948, 32'shf559472b, 32'shf5531528, 32'shf54ce33f, 32'shf546b171, 
               32'shf5407fbd, 32'shf53a4e24, 32'shf5341ca5, 32'shf52deb41, 32'shf527b9f7, 32'shf52188c9, 32'shf51b57b5, 32'shf51526bc, 
               32'shf50ef5de, 32'shf508c51b, 32'shf5029473, 32'shf4fc63e6, 32'shf4f63374, 32'shf4f0031e, 32'shf4e9d2e3, 32'shf4e3a2c3, 
               32'shf4dd72be, 32'shf4d742d6, 32'shf4d11308, 32'shf4cae356, 32'shf4c4b3c0, 32'shf4be8446, 32'shf4b854e7, 32'shf4b225a4, 
               32'shf4abf67e, 32'shf4a5c773, 32'shf49f9884, 32'shf49969b1, 32'shf4933afa, 32'shf48d0c5f, 32'shf486dde1, 32'shf480af7f, 
               32'shf47a8139, 32'shf4745310, 32'shf46e2504, 32'shf467f713, 32'shf461c940, 32'shf45b9b89, 32'shf4556def, 32'shf44f4071, 
               32'shf4491311, 32'shf442e5cd, 32'shf43cb8a7, 32'shf4368b9d, 32'shf4305eb0, 32'shf42a31e1, 32'shf424052f, 32'shf41dd89a, 
               32'shf417ac22, 32'shf4117fc8, 32'shf40b538b, 32'shf405276c, 32'shf3fefb6a, 32'shf3f8cf86, 32'shf3f2a3bf, 32'shf3ec7817, 
               32'shf3e64c8c, 32'shf3e0211f, 32'shf3d9f5cf, 32'shf3d3ca9e, 32'shf3cd9f8b, 32'shf3c77496, 32'shf3c149bf, 32'shf3bb1f07, 
               32'shf3b4f46c, 32'shf3aec9f0, 32'shf3a89f92, 32'shf3a27553, 32'shf39c4b32, 32'shf3962130, 32'shf38ff74d, 32'shf389cd88, 
               32'shf383a3e2, 32'shf37d7a5b, 32'shf37750f2, 32'shf37127a9, 32'shf36afe7e, 32'shf364d573, 32'shf35eac86, 32'shf35883b9, 
               32'shf3525b0b, 32'shf34c327c, 32'shf3460a0d, 32'shf33fe1bd, 32'shf339b98d, 32'shf333917c, 32'shf32d698a, 32'shf32741b9, 
               32'shf3211a07, 32'shf31af274, 32'shf314cb02, 32'shf30ea3af, 32'shf3087c7d, 32'shf302556a, 32'shf2fc2e77, 32'shf2f607a5, 
               32'shf2efe0f2, 32'shf2e9ba60, 32'shf2e393ef, 32'shf2dd6d9d, 32'shf2d7476c, 32'shf2d1215b, 32'shf2cafb6b, 32'shf2c4d59c, 
               32'shf2beafed, 32'shf2b88a5f, 32'shf2b264f2, 32'shf2ac3fa5, 32'shf2a61a7a, 32'shf29ff56f, 32'shf299d085, 32'shf293abbd, 
               32'shf28d8715, 32'shf287628f, 32'shf2813e2a, 32'shf27b19e6, 32'shf274f5c3, 32'shf26ed1c2, 32'shf268ade3, 32'shf2628a25, 
               32'shf25c6688, 32'shf256430e, 32'shf2501fb5, 32'shf249fc7d, 32'shf243d968, 32'shf23db674, 32'shf23793a3, 32'shf23170f3, 
               32'shf22b4e66, 32'shf2252bfa, 32'shf21f09b1, 32'shf218e78a, 32'shf212c585, 32'shf20ca3a3, 32'shf20681e3, 32'shf2006046, 
               32'shf1fa3ecb, 32'shf1f41d72, 32'shf1edfc3d, 32'shf1e7db2a, 32'shf1e1ba3a, 32'shf1db996d, 32'shf1d578c2, 32'shf1cf583b, 
               32'shf1c937d6, 32'shf1c31795, 32'shf1bcf777, 32'shf1b6d77c, 32'shf1b0b7a4, 32'shf1aa97ef, 32'shf1a4785e, 32'shf19e58f1, 
               32'shf19839a6, 32'shf1921a80, 32'shf18bfb7d, 32'shf185dc9d, 32'shf17fbde2, 32'shf1799f4a, 32'shf17380d6, 32'shf16d6286, 
               32'shf1674459, 32'shf1612651, 32'shf15b086d, 32'shf154eaad, 32'shf14ecd11, 32'shf148af9a, 32'shf1429247, 32'shf13c7518, 
               32'shf136580d, 32'shf1303b27, 32'shf12a1e66, 32'shf12401c9, 32'shf11de551, 32'shf117c8fe, 32'shf111accf, 32'shf10b90c5, 
               32'shf10574e0, 32'shf0ff5921, 32'shf0f93d86, 32'shf0f32210, 32'shf0ed06bf, 32'shf0e6eb94, 32'shf0e0d08d, 32'shf0dab5ad, 
               32'shf0d49af1, 32'shf0ce805b, 32'shf0c865ea, 32'shf0c24b9f, 32'shf0bc317a, 32'shf0b6177a, 32'shf0affda0, 32'shf0a9e3eb, 
               32'shf0a3ca5d, 32'shf09db0f4, 32'shf09797b2, 32'shf0917e95, 32'shf08b659f, 32'shf0854cce, 32'shf07f3424, 32'shf0791ba0, 
               32'shf0730342, 32'shf06ceb0b, 32'shf066d2fa, 32'shf060bb10, 32'shf05aa34c, 32'shf0548baf, 32'shf04e7438, 32'shf0485ce9, 
               32'shf04245c0, 32'shf03c2ebd, 32'shf03617e2, 32'shf030012e, 32'shf029eaa1, 32'shf023d43a, 32'shf01dbdfb, 32'shf017a7e3, 
               32'shf01191f3, 32'shf00b7c29, 32'shf0056687, 32'shefff510d, 32'sheff93bba, 32'sheff3268e, 32'shefed118a, 32'shefe6fcae, 
               32'shefe0e7f9, 32'shefdad36c, 32'shefd4bf08, 32'shefceaacb, 32'shefc896b5, 32'shefc282c8, 32'shefbc6f03, 32'shefb65b66, 
               32'shefb047f2, 32'shefaa34a5, 32'shefa42181, 32'shef9e0e85, 32'shef97fbb2, 32'shef91e907, 32'shef8bd685, 32'shef85c42b, 
               32'shef7fb1fa, 32'shef799ff2, 32'shef738e12, 32'shef6d7c5b, 32'shef676ace, 32'shef615969, 32'shef5b482d, 32'shef55371a, 
               32'shef4f2630, 32'shef491570, 32'shef4304d8, 32'shef3cf46a, 32'shef36e426, 32'shef30d40a, 32'shef2ac419, 32'shef24b451, 
               32'shef1ea4b2, 32'shef18953d, 32'shef1285f2, 32'shef0c76d0, 32'shef0667d9, 32'shef00590b, 32'sheefa4a67, 32'sheef43bed, 
               32'sheeee2d9d, 32'sheee81f78, 32'sheee2117c, 32'sheedc03ab, 32'sheed5f604, 32'sheecfe887, 32'sheec9db35, 32'sheec3ce0d, 
               32'sheebdc110, 32'sheeb7b43e, 32'sheeb1a796, 32'sheeab9b18, 32'sheea58ec6, 32'shee9f829e, 32'shee9976a1, 32'shee936acf, 
               32'shee8d5f29, 32'shee8753ad, 32'shee81485c, 32'shee7b3d36, 32'shee75323c, 32'shee6f276d, 32'shee691cc9, 32'shee631251, 
               32'shee5d0804, 32'shee56fde3, 32'shee50f3ed, 32'shee4aea23, 32'shee44e084, 32'shee3ed712, 32'shee38cdcb, 32'shee32c4b0, 
               32'shee2cbbc1, 32'shee26b2fe, 32'shee20aa67, 32'shee1aa1fc, 32'shee1499bd, 32'shee0e91aa, 32'shee0889c4, 32'shee02820a, 
               32'shedfc7a7c, 32'shedf6731b, 32'shedf06be6, 32'shedea64de, 32'shede45e03, 32'shedde5754, 32'shedd850d2, 32'shedd24a7d, 
               32'shedcc4454, 32'shedc63e59, 32'shedc0388a, 32'shedba32e9, 32'shedb42d74, 32'shedae282d, 32'sheda82313, 32'sheda21e26, 
               32'shed9c1967, 32'shed9614d5, 32'shed901070, 32'shed8a0c39, 32'shed84082f, 32'shed7e0453, 32'shed7800a5, 32'shed71fd24, 
               32'shed6bf9d1, 32'shed65f6ac, 32'shed5ff3b5, 32'shed59f0ec, 32'shed53ee51, 32'shed4debe4, 32'shed47e9a5, 32'shed41e794, 
               32'shed3be5b1, 32'shed35e3fd, 32'shed2fe277, 32'shed29e120, 32'shed23dff7, 32'shed1ddefd, 32'shed17de31, 32'shed11dd94, 
               32'shed0bdd25, 32'shed05dce5, 32'shecffdcd4, 32'shecf9dcf3, 32'shecf3dd3f, 32'shecedddbb, 32'shece7de66, 32'shece1df40, 
               32'shecdbe04a, 32'shecd5e182, 32'sheccfe2ea, 32'shecc9e481, 32'shecc3e648, 32'shecbde83e, 32'shecb7ea63, 32'shecb1ecb8, 
               32'shecabef3d, 32'sheca5f1f2, 32'shec9ff4d6, 32'shec99f7ea, 32'shec93fb2e, 32'shec8dfea1, 32'shec880245, 32'shec820619, 
               32'shec7c0a1d, 32'shec760e51, 32'shec7012b5, 32'shec6a1749, 32'shec641c0e, 32'shec5e2103, 32'shec582629, 32'shec522b7f, 
               32'shec4c3106, 32'shec4636bd, 32'shec403ca5, 32'shec3a42be, 32'shec344908, 32'shec2e4f82, 32'shec28562d, 32'shec225d09, 
               32'shec1c6417, 32'shec166b55, 32'shec1072c4, 32'shec0a7a65, 32'shec048237, 32'shebfe8a3a, 32'shebf8926f, 32'shebf29ad4, 
               32'shebeca36c, 32'shebe6ac35, 32'shebe0b52f, 32'shebdabe5c, 32'shebd4c7ba, 32'shebced149, 32'shebc8db0b, 32'shebc2e4fe, 
               32'shebbcef23, 32'shebb6f97b, 32'shebb10404, 32'shebab0ec0, 32'sheba519ad, 32'sheb9f24cd, 32'sheb99301f, 32'sheb933ba4, 
               32'sheb8d475b, 32'sheb875344, 32'sheb815f60, 32'sheb7b6bae, 32'sheb75782f, 32'sheb6f84e3, 32'sheb6991ca, 32'sheb639ee3, 
               32'sheb5dac2f, 32'sheb57b9ae, 32'sheb51c760, 32'sheb4bd545, 32'sheb45e35d, 32'sheb3ff1a8, 32'sheb3a0027, 32'sheb340ed9, 
               32'sheb2e1dbe, 32'sheb282cd6, 32'sheb223c22, 32'sheb1c4ba1, 32'sheb165b54, 32'sheb106b3a, 32'sheb0a7b54, 32'sheb048ba2, 
               32'sheafe9c24, 32'sheaf8acd9, 32'sheaf2bdc3, 32'sheaeccee0, 32'sheae6e031, 32'sheae0f1b6, 32'sheadb0370, 32'shead5155d, 
               32'sheacf277f, 32'sheac939d5, 32'sheac34c60, 32'sheabd5f1f, 32'sheab77212, 32'sheab1853a, 32'sheaab9896, 32'sheaa5ac27, 
               32'shea9fbfed, 32'shea99d3e8, 32'shea93e817, 32'shea8dfc7b, 32'shea881114, 32'shea8225e2, 32'shea7c3ae5, 32'shea76501d, 
               32'shea70658a, 32'shea6a7b2d, 32'shea649105, 32'shea5ea712, 32'shea58bd54, 32'shea52d3cc, 32'shea4cea79, 32'shea47015c, 
               32'shea411874, 32'shea3b2fc2, 32'shea354746, 32'shea2f5f00, 32'shea2976ef, 32'shea238f15, 32'shea1da770, 32'shea17c001, 
               32'shea11d8c8, 32'shea0bf1c6, 32'shea060af9, 32'shea002463, 32'she9fa3e03, 32'she9f457da, 32'she9ee71e6, 32'she9e88c2a, 
               32'she9e2a6a3, 32'she9dcc154, 32'she9d6dc3b, 32'she9d0f758, 32'she9cb12ad, 32'she9c52e38, 32'she9bf49fa, 32'she9b965f3, 
               32'she9b38223, 32'she9ad9e8a, 32'she9a7bb28, 32'she9a1d7fd, 32'she99bf509, 32'she996124d, 32'she9902fc7, 32'she98a4d7a, 
               32'she9846b63, 32'she97e8984, 32'she978a7dd, 32'she972c66d, 32'she96ce535, 32'she9670435, 32'she961236c, 32'she95b42db, 
               32'she9556282, 32'she94f8261, 32'she949a278, 32'she943c2c7, 32'she93de34e, 32'she938040d, 32'she9322505, 32'she92c4634, 
               32'she926679c, 32'she920893d, 32'she91aab16, 32'she914cd27, 32'she90eef71, 32'she90911f3, 32'she90334af, 32'she8fd57a2, 
               32'she8f77acf, 32'she8f19e34, 32'she8ebc1d3, 32'she8e5e5aa, 32'she8e009ba, 32'she8da2e04, 32'she8d45286, 32'she8ce7742, 
               32'she8c89c37, 32'she8c2c165, 32'she8bce6cd, 32'she8b70c6d, 32'she8b13248, 32'she8ab585c, 32'she8a57ea9, 32'she89fa530, 
               32'she899cbf1, 32'she893f2eb, 32'she88e1a20, 32'she888418e, 32'she8826936, 32'she87c9118, 32'she876b934, 32'she870e18a, 
               32'she86b0a1a, 32'she86532e4, 32'she85f5be9, 32'she8598528, 32'she853aea1, 32'she84dd855, 32'she8480243, 32'she8422c6c, 
               32'she83c56cf, 32'she836816d, 32'she830ac45, 32'she82ad759, 32'she82502a7, 32'she81f2e30, 32'she81959f4, 32'she81385f3, 
               32'she80db22d, 32'she807dea2, 32'she8020b52, 32'she7fc383d, 32'she7f66564, 32'she7f092c6, 32'she7eac063, 32'she7e4ee3c, 
               32'she7df1c50, 32'she7d94a9f, 32'she7d3792b, 32'she7cda7f2, 32'she7c7d6f4, 32'she7c20633, 32'she7bc35ad, 32'she7b66563, 
               32'she7b09555, 32'she7aac583, 32'she7a4f5ed, 32'she79f2693, 32'she7995776, 32'she7938894, 32'she78db9ef, 32'she787eb86, 
               32'she7821d59, 32'she77c4f69, 32'she77681b6, 32'she770b43e, 32'she76ae704, 32'she7651a06, 32'she75f4d45, 32'she75980c1, 
               32'she753b479, 32'she74de86f, 32'she7481ca1, 32'she7425110, 32'she73c85bc, 32'she736baa6, 32'she730efcc, 32'she72b2530, 
               32'she7255ad1, 32'she71f90b0, 32'she719c6cb, 32'she713fd25, 32'she70e33bb, 32'she7086a8f, 32'she702a1a1, 32'she6fcd8f1, 
               32'she6f7107e, 32'she6f14849, 32'she6eb8052, 32'she6e5b899, 32'she6dff11d, 32'she6da29e0, 32'she6d462e1, 32'she6ce9c1f, 
               32'she6c8d59c, 32'she6c30f57, 32'she6bd4951, 32'she6b78389, 32'she6b1bdff, 32'she6abf8b3, 32'she6a633a6, 32'she6a06ed8, 
               32'she69aaa48, 32'she694e5f7, 32'she68f21e5, 32'she6895e11, 32'she6839a7c, 32'she67dd727, 32'she6781410, 32'she6725138, 
               32'she66c8e9f, 32'she666cc45, 32'she6610a2a, 32'she65b484f, 32'she65586b3, 32'she64fc556, 32'she64a0438, 32'she644435a, 
               32'she63e82bc, 32'she638c25d, 32'she633023e, 32'she62d425e, 32'she62782be, 32'she621c35e, 32'she61c043d, 32'she616455d, 
               32'she61086bc, 32'she60ac85c, 32'she6050a3b, 32'she5ff4c5b, 32'she5f98ebb, 32'she5f3d15b, 32'she5ee143b, 32'she5e8575b, 
               32'she5e29abc, 32'she5dcde5e, 32'she5d72240, 32'she5d16662, 32'she5cbaac5, 32'she5c5ef69, 32'she5c0344d, 32'she5ba7972, 
               32'she5b4bed8, 32'she5af047f, 32'she5a94a67, 32'she5a39090, 32'she59dd6f9, 32'she5981da4, 32'she5926490, 32'she58cabbe, 
               32'she586f32c, 32'she5813adc, 32'she57b82cd, 32'she575cb00, 32'she5701374, 32'she56a5c2a, 32'she564a521, 32'she55eee5a, 
               32'she55937d5, 32'she5538191, 32'she54dcb8f, 32'she54815cf, 32'she5426051, 32'she53cab15, 32'she536f61b, 32'she5314163, 
               32'she52b8cee, 32'she525d8ba, 32'she52024c9, 32'she51a711a, 32'she514bdad, 32'she50f0a83, 32'she509579b, 32'she503a4f6, 
               32'she4fdf294, 32'she4f84074, 32'she4f28e96, 32'she4ecdcfc, 32'she4e72ba4, 32'she4e17a8f, 32'she4dbc9bd, 32'she4d6192e, 
               32'she4d068e2, 32'she4cab8d9, 32'she4c50914, 32'she4bf5991, 32'she4b9aa52, 32'she4b3fb56, 32'she4ae4c9d, 32'she4a89e28, 
               32'she4a2eff6, 32'she49d4208, 32'she497945d, 32'she491e6f6, 32'she48c39d3, 32'she4868cf3, 32'she480e057, 32'she47b33ff, 
               32'she47587eb, 32'she46fdc1b, 32'she46a308f, 32'she4648547, 32'she45eda43, 32'she4592f83, 32'she4538507, 32'she44ddad0, 
               32'she44830dd, 32'she442872e, 32'she43cddc4, 32'she437349f, 32'she4318bbe, 32'she42be321, 32'she4263ac9, 32'she42092b6, 
               32'she41aeae8, 32'she415435f, 32'she40f9c1a, 32'she409f51a, 32'she4044e60, 32'she3fea7ea, 32'she3f901ba, 32'she3f35bce, 
               32'she3edb628, 32'she3e810c7, 32'she3e26bac, 32'she3dcc6d5, 32'she3d72245, 32'she3d17df9, 32'she3cbd9f4, 32'she3c63633, 
               32'she3c092b9, 32'she3baef84, 32'she3b54c95, 32'she3afa9ec, 32'she3aa0788, 32'she3a4656b, 32'she39ec393, 32'she3992202, 
               32'she39380b6, 32'she38ddfb1, 32'she3883ef2, 32'she3829e79, 32'she37cfe47, 32'she3775e5a, 32'she371beb5, 32'she36c1f55, 
               32'she366803c, 32'she360e16a, 32'she35b42df, 32'she355a49a, 32'she350069b, 32'she34a68e4, 32'she344cb73, 32'she33f2e4a, 
               32'she3399167, 32'she333f4cb, 32'she32e5876, 32'she328bc69, 32'she32320a2, 32'she31d8523, 32'she317e9eb, 32'she3124efa, 
               32'she30cb451, 32'she30719ef, 32'she3017fd5, 32'she2fbe602, 32'she2f64c77, 32'she2f0b333, 32'she2eb1a37, 32'she2e58183, 
               32'she2dfe917, 32'she2da50f3, 32'she2d4b916, 32'she2cf2182, 32'she2c98a35, 32'she2c3f331, 32'she2be5c74, 32'she2b8c600, 
               32'she2b32fd4, 32'she2ad99f1, 32'she2a80456, 32'she2a26f03, 32'she29cd9f8, 32'she2974536, 32'she291b0bd, 32'she28c1c8c, 
               32'she28688a4, 32'she280f505, 32'she27b61af, 32'she275cea1, 32'she2703bdc, 32'she26aa960, 32'she265172e, 32'she25f8544, 
               32'she259f3a3, 32'she254624b, 32'she24ed13d, 32'she2494078, 32'she243affc, 32'she23e1fca, 32'she2388fe1, 32'she2330041, 
               32'she22d70eb, 32'she227e1df, 32'she222531c, 32'she21cc4a3, 32'she2173674, 32'she211a88f, 32'she20c1af3, 32'she2068da1, 
               32'she2010099, 32'she1fb73dc, 32'she1f5e768, 32'she1f05b3e, 32'she1eacf5f, 32'she1e543ca, 32'she1dfb87f, 32'she1da2d7e, 
               32'she1d4a2c8, 32'she1cf185c, 32'she1c98e3b, 32'she1c40464, 32'she1be7ad8, 32'she1b8f197, 32'she1b368a0, 32'she1addff4, 
               32'she1a85793, 32'she1a2cf7c, 32'she19d47b1, 32'she197c031, 32'she19238fb, 32'she18cb211, 32'she1872b72, 32'she181a51e, 
               32'she17c1f15, 32'she1769958, 32'she17113e5, 32'she16b8ebf, 32'she16609e3, 32'she1608554, 32'she15b0110, 32'she1557d17, 
               32'she14ff96a, 32'she14a7609, 32'she144f2f3, 32'she13f702a, 32'she139edac, 32'she1346b7a, 32'she12ee995, 32'she12967fb, 
               32'she123e6ad, 32'she11e65ac, 32'she118e4f6, 32'she113648d, 32'she10de470, 32'she10864a0, 32'she102e51c, 32'she0fd65e4, 
               32'she0f7e6f9, 32'she0f2685b, 32'she0ecea09, 32'she0e76c04, 32'she0e1ee4b, 32'she0dc70e0, 32'she0d6f3c1, 32'she0d176ef, 
               32'she0cbfa6a, 32'she0c67e32, 32'she0c10247, 32'she0bb86a9, 32'she0b60b58, 32'she0b09055, 32'she0ab159e, 32'she0a59b35, 
               32'she0a0211a, 32'she09aa74b, 32'she0952dcb, 32'she08fb497, 32'she08a3bb2, 32'she084c31a, 32'she07f4acf, 32'she079d2d3, 
               32'she0745b24, 32'she06ee3c3, 32'she0696cb0, 32'she063f5eb, 32'she05e7f74, 32'she059094a, 32'she053936f, 32'she04e1de3, 
               32'she048a8a4, 32'she04333b3, 32'she03dbf11, 32'she0384abe, 32'she032d6b8, 32'she02d6301, 32'she027ef99, 32'she0227c7f, 
               32'she01d09b4, 32'she0179738, 32'she012250a, 32'she00cb32b, 32'she007419b, 32'she001d05a, 32'shdffc5f67, 32'shdff6eec4, 
               32'shdff17e70, 32'shdfec0e6a, 32'shdfe69eb4, 32'shdfe12f4e, 32'shdfdbc036, 32'shdfd6516e, 32'shdfd0e2f5, 32'shdfcb74cb, 
               32'shdfc606f1, 32'shdfc09967, 32'shdfbb2c2c, 32'shdfb5bf41, 32'shdfb052a5, 32'shdfaae659, 32'shdfa57a5d, 32'shdfa00eb1, 
               32'shdf9aa354, 32'shdf953848, 32'shdf8fcd8b, 32'shdf8a631f, 32'shdf84f902, 32'shdf7f8f36, 32'shdf7a25ba, 32'shdf74bc8e, 
               32'shdf6f53b3, 32'shdf69eb27, 32'shdf6482ed, 32'shdf5f1b02, 32'shdf59b369, 32'shdf544c1f, 32'shdf4ee527, 32'shdf497e7f, 
               32'shdf441828, 32'shdf3eb221, 32'shdf394c6b, 32'shdf33e707, 32'shdf2e81f3, 32'shdf291d30, 32'shdf23b8be, 32'shdf1e549d, 
               32'shdf18f0ce, 32'shdf138d4f, 32'shdf0e2a22, 32'shdf08c746, 32'shdf0364bc, 32'shdefe0282, 32'shdef8a09b, 32'shdef33f04, 
               32'shdeedddc0, 32'shdee87ccc, 32'shdee31c2b, 32'shdeddbbdb, 32'shded85bdd, 32'shded2fc31, 32'shdecd9cd7, 32'shdec83dce, 
               32'shdec2df18, 32'shdebd80b3, 32'shdeb822a1, 32'shdeb2c4e1, 32'shdead6773, 32'shdea80a57, 32'shdea2ad8d, 32'shde9d5116, 
               32'shde97f4f1, 32'shde92991e, 32'shde8d3d9e, 32'shde87e271, 32'shde828796, 32'shde7d2d0e, 32'shde77d2d8, 32'shde7278f5, 
               32'shde6d1f65, 32'shde67c628, 32'shde626d3e, 32'shde5d14a6, 32'shde57bc62, 32'shde526471, 32'shde4d0cd2, 32'shde47b587, 
               32'shde425e8f, 32'shde3d07eb, 32'shde37b199, 32'shde325b9b, 32'shde2d05f1, 32'shde27b09a, 32'shde225b96, 32'shde1d06e6, 
               32'shde17b28a, 32'shde125e81, 32'shde0d0acc, 32'shde07b76b, 32'shde02645d, 32'shddfd11a3, 32'shddf7bf3e, 32'shddf26d2c, 
               32'shdded1b6e, 32'shdde7ca05, 32'shdde278ef, 32'shdddd282e, 32'shddd7d7c1, 32'shddd287a8, 32'shddcd37e4, 32'shddc7e873, 
               32'shddc29958, 32'shddbd4a91, 32'shddb7fc1e, 32'shddb2ae00, 32'shddad6036, 32'shdda812c2, 32'shdda2c5a2, 32'shdd9d78d7, 
               32'shdd982c60, 32'shdd92e03f, 32'shdd8d9472, 32'shdd8848fb, 32'shdd82fdd8, 32'shdd7db30b, 32'shdd786892, 32'shdd731e6f, 
               32'shdd6dd4a2, 32'shdd688b29, 32'shdd634206, 32'shdd5df938, 32'shdd58b0c0, 32'shdd53689d, 32'shdd4e20d0, 32'shdd48d958, 
               32'shdd439236, 32'shdd3e4b6a, 32'shdd3904f4, 32'shdd33bed3, 32'shdd2e7908, 32'shdd293393, 32'shdd23ee74, 32'shdd1ea9ab, 
               32'shdd196538, 32'shdd14211b, 32'shdd0edd55, 32'shdd0999e4, 32'shdd0456ca, 32'shdcff1407, 32'shdcf9d199, 32'shdcf48f82, 
               32'shdcef4dc2, 32'shdcea0c58, 32'shdce4cb44, 32'shdcdf8a87, 32'shdcda4a21, 32'shdcd50a12, 32'shdccfca59, 32'shdcca8af7, 
               32'shdcc54bec, 32'shdcc00d38, 32'shdcbacedb, 32'shdcb590d5, 32'shdcb05326, 32'shdcab15ce, 32'shdca5d8cd, 32'shdca09c24, 
               32'shdc9b5fd2, 32'shdc9623d7, 32'shdc90e834, 32'shdc8bace8, 32'shdc8671f3, 32'shdc813756, 32'shdc7bfd11, 32'shdc76c323, 
               32'shdc71898d, 32'shdc6c504e, 32'shdc671768, 32'shdc61ded9, 32'shdc5ca6a2, 32'shdc576ec3, 32'shdc52373c, 32'shdc4d000d, 
               32'shdc47c936, 32'shdc4292b8, 32'shdc3d5c91, 32'shdc3826c3, 32'shdc32f14d, 32'shdc2dbc2f, 32'shdc28876a, 32'shdc2352fd, 
               32'shdc1e1ee9, 32'shdc18eb2d, 32'shdc13b7c9, 32'shdc0e84bf, 32'shdc09520d, 32'shdc041fb4, 32'shdbfeedb3, 32'shdbf9bc0c, 
               32'shdbf48abd, 32'shdbef59c7, 32'shdbea292b, 32'shdbe4f8e7, 32'shdbdfc8fc, 32'shdbda996b, 32'shdbd56a32, 32'shdbd03b53, 
               32'shdbcb0cce, 32'shdbc5dea1, 32'shdbc0b0ce, 32'shdbbb8354, 32'shdbb65634, 32'shdbb1296e, 32'shdbabfd01, 32'shdba6d0ed, 
               32'shdba1a534, 32'shdb9c79d4, 32'shdb974ece, 32'shdb922421, 32'shdb8cf9cf, 32'shdb87cfd6, 32'shdb82a638, 32'shdb7d7cf3, 
               32'shdb785409, 32'shdb732b79, 32'shdb6e0342, 32'shdb68db67, 32'shdb63b3e5, 32'shdb5e8cbe, 32'shdb5965f1, 32'shdb543f7e, 
               32'shdb4f1967, 32'shdb49f3a9, 32'shdb44ce46, 32'shdb3fa93e, 32'shdb3a8491, 32'shdb35603e, 32'shdb303c46, 32'shdb2b18a9, 
               32'shdb25f566, 32'shdb20d27f, 32'shdb1baff2, 32'shdb168dc1, 32'shdb116beb, 32'shdb0c4a70, 32'shdb072950, 32'shdb02088b, 
               32'shdafce821, 32'shdaf7c813, 32'shdaf2a860, 32'shdaed8909, 32'shdae86a0d, 32'shdae34b6d, 32'shdade2d28, 32'shdad90f3f, 
               32'shdad3f1b1, 32'shdaced47f, 32'shdac9b7a9, 32'shdac49b2f, 32'shdabf7f11, 32'shdaba634e, 32'shdab547e8, 32'shdab02cdd, 
               32'shdaab122f, 32'shdaa5f7dd, 32'shdaa0dde7, 32'shda9bc44d, 32'shda96ab0f, 32'shda91922e, 32'shda8c79a9, 32'shda876180, 
               32'shda8249b4, 32'shda7d3244, 32'shda781b31, 32'shda73047b, 32'shda6dee21, 32'shda68d824, 32'shda63c284, 32'shda5ead40, 
               32'shda599859, 32'shda5483d0, 32'shda4f6fa3, 32'shda4a5bd3, 32'shda454860, 32'shda40354a, 32'shda3b2292, 32'shda361036, 
               32'shda30fe38, 32'shda2bec97, 32'shda26db54, 32'shda21ca6e, 32'shda1cb9e5, 32'shda17a9ba, 32'shda1299ec, 32'shda0d8a7c, 
               32'shda087b69, 32'shda036cb5, 32'shd9fe5e5e, 32'shd9f95064, 32'shd9f442c9, 32'shd9ef358b, 32'shd9ea28ac, 32'shd9e51c2a, 
               32'shd9e01006, 32'shd9db0441, 32'shd9d5f8d9, 32'shd9d0edd0, 32'shd9cbe325, 32'shd9c6d8d8, 32'shd9c1cee9, 32'shd9bcc559, 
               32'shd9b7bc27, 32'shd9b2b354, 32'shd9adaadf, 32'shd9a8a2c9, 32'shd9a39b11, 32'shd99e93b8, 32'shd9998cbe, 32'shd9948623, 
               32'shd98f7fe6, 32'shd98a7a08, 32'shd9857489, 32'shd9806f69, 32'shd97b6aa8, 32'shd9766646, 32'shd9716243, 32'shd96c5e9f, 
               32'shd9675b5a, 32'shd9625875, 32'shd95d55ef, 32'shd95853c8, 32'shd9535201, 32'shd94e5099, 32'shd9494f90, 32'shd9444ee7, 
               32'shd93f4e9e, 32'shd93a4eb4, 32'shd9354f2a, 32'shd9305000, 32'shd92b5135, 32'shd92652ca, 32'shd92154bf, 32'shd91c5714, 
               32'shd91759c9, 32'shd9125cde, 32'shd90d6053, 32'shd9086428, 32'shd903685d, 32'shd8fe6cf2, 32'shd8f971e8, 32'shd8f4773e, 
               32'shd8ef7cf4, 32'shd8ea830b, 32'shd8e58982, 32'shd8e0905a, 32'shd8db9792, 32'shd8d69f2a, 32'shd8d1a724, 32'shd8ccaf7e, 
               32'shd8c7b838, 32'shd8c2c154, 32'shd8bdcad0, 32'shd8b8d4ad, 32'shd8b3deeb, 32'shd8aee98a, 32'shd8a9f48a, 32'shd8a4ffec, 
               32'shd8a00bae, 32'shd89b17d1, 32'shd8962456, 32'shd891313b, 32'shd88c3e83, 32'shd8874c2b, 32'shd8825a35, 32'shd87d68a0, 
               32'shd878776d, 32'shd873869b, 32'shd86e962b, 32'shd869a61d, 32'shd864b670, 32'shd85fc725, 32'shd85ad83c, 32'shd855e9b4, 
               32'shd850fb8e, 32'shd84c0dcb, 32'shd8472069, 32'shd8423369, 32'shd83d46cc, 32'shd8385a90, 32'shd8336eb7, 32'shd82e833f, 
               32'shd829982b, 32'shd824ad78, 32'shd81fc328, 32'shd81ad93a, 32'shd815efae, 32'shd8110685, 32'shd80c1dbf, 32'shd807355b, 
               32'shd8024d59, 32'shd7fd65bb, 32'shd7f87e7f, 32'shd7f397a6, 32'shd7eeb130, 32'shd7e9cb1c, 32'shd7e4e56c, 32'shd7e0001e, 
               32'shd7db1b34, 32'shd7d636ac, 32'shd7d15288, 32'shd7cc6ec6, 32'shd7c78b68, 32'shd7c2a86d, 32'shd7bdc5d6, 32'shd7b8e3a2, 
               32'shd7b401d1, 32'shd7af2063, 32'shd7aa3f5a, 32'shd7a55eb3, 32'shd7a07e70, 32'shd79b9e91, 32'shd796bf16, 32'shd791dffe, 
               32'shd78d014a, 32'shd78822f9, 32'shd783450d, 32'shd77e6784, 32'shd7798a60, 32'shd774ad9f, 32'shd76fd143, 32'shd76af54a, 
               32'shd76619b6, 32'shd7613e86, 32'shd75c63ba, 32'shd7578952, 32'shd752af4f, 32'shd74dd5b0, 32'shd748fc75, 32'shd744239f, 
               32'shd73f4b2e, 32'shd73a7321, 32'shd7359b78, 32'shd730c434, 32'shd72bed55, 32'shd72716db, 32'shd72240c5, 32'shd71d6b15, 
               32'shd71895c9, 32'shd713c0e2, 32'shd70eec60, 32'shd70a1843, 32'shd705448b, 32'shd7007138, 32'shd6fb9e4b, 32'shd6f6cbc2, 
               32'shd6f1f99f, 32'shd6ed27e1, 32'shd6e85689, 32'shd6e38596, 32'shd6deb508, 32'shd6d9e4e0, 32'shd6d5151d, 32'shd6d045c0, 
               32'shd6cb76c9, 32'shd6c6a837, 32'shd6c1da0b, 32'shd6bd0c45, 32'shd6b83ee4, 32'shd6b371ea, 32'shd6aea555, 32'shd6a9d926, 
               32'shd6a50d5d, 32'shd6a041fa, 32'shd69b76fe, 32'shd696ac67, 32'shd691e237, 32'shd68d186d, 32'shd6884f09, 32'shd683860b, 
               32'shd67ebd74, 32'shd679f543, 32'shd6752d79, 32'shd6706615, 32'shd66b9f18, 32'shd666d881, 32'shd6621251, 32'shd65d4c88, 
               32'shd6588725, 32'shd653c229, 32'shd64efd94, 32'shd64a3966, 32'shd645759f, 32'shd640b23f, 32'shd63bef46, 32'shd6372cb3, 
               32'shd6326a88, 32'shd62da8c4, 32'shd628e767, 32'shd6242672, 32'shd61f65e4, 32'shd61aa5bd, 32'shd615e5fd, 32'shd61126a5, 
               32'shd60c67b4, 32'shd607a92b, 32'shd602eb0a, 32'shd5fe2d50, 32'shd5f96ffd, 32'shd5f4b313, 32'shd5eff690, 32'shd5eb3a75, 
               32'shd5e67ec1, 32'shd5e1c376, 32'shd5dd0892, 32'shd5d84e17, 32'shd5d39403, 32'shd5ceda58, 32'shd5ca2115, 32'shd5c56839, 
               32'shd5c0afc6, 32'shd5bbf7bc, 32'shd5b74019, 32'shd5b288df, 32'shd5add20d, 32'shd5a91ba4, 32'shd5a465a3, 32'shd59fb00b, 
               32'shd59afadb, 32'shd5964614, 32'shd59191b5, 32'shd58cddbf, 32'shd5882a32, 32'shd583770e, 32'shd57ec452, 32'shd57a1200, 
               32'shd5756016, 32'shd570ae95, 32'shd56bfd7d, 32'shd5674ccf, 32'shd5629c89, 32'shd55decad, 32'shd5593d3a, 32'shd5548e30, 
               32'shd54fdf8f, 32'shd54b3157, 32'shd5468389, 32'shd541d625, 32'shd53d292a, 32'shd5387c98, 32'shd533d070, 32'shd52f24b2, 
               32'shd52a795d, 32'shd525ce72, 32'shd52123f0, 32'shd51c79d9, 32'shd517d02b, 32'shd51326e7, 32'shd50e7e0d, 32'shd509d59d, 
               32'shd5052d97, 32'shd50085fb, 32'shd4fbdec9, 32'shd4f73801, 32'shd4f291a4, 32'shd4edebb0, 32'shd4e94627, 32'shd4e4a108, 
               32'shd4dffc54, 32'shd4db580a, 32'shd4d6b42b, 32'shd4d210b5, 32'shd4cd6dab, 32'shd4c8cb0b, 32'shd4c428d6, 32'shd4bf870b, 
               32'shd4bae5ab, 32'shd4b644b6, 32'shd4b1a42c, 32'shd4ad040c, 32'shd4a86458, 32'shd4a3c50e, 32'shd49f2630, 32'shd49a87bc, 
               32'shd495e9b3, 32'shd4914c16, 32'shd48caee4, 32'shd488121d, 32'shd48375c1, 32'shd47ed9d0, 32'shd47a3e4b, 32'shd475a332, 
               32'shd4710883, 32'shd46c6e40, 32'shd467d469, 32'shd4633afd, 32'shd45ea1fd, 32'shd45a0969, 32'shd4557140, 32'shd450d983, 
               32'shd44c4232, 32'shd447ab4c, 32'shd44314d3, 32'shd43e7ec5, 32'shd439e923, 32'shd43553ee, 32'shd430bf24, 32'shd42c2ac6, 
               32'shd42796d5, 32'shd4230350, 32'shd41e7037, 32'shd419dd8a, 32'shd4154b4a, 32'shd410b976, 32'shd40c280e, 32'shd4079713, 
               32'shd4030684, 32'shd3fe7662, 32'shd3f9e6ad, 32'shd3f55764, 32'shd3f0c887, 32'shd3ec3a18, 32'shd3e7ac15, 32'shd3e31e7f, 
               32'shd3de9156, 32'shd3da049a, 32'shd3d5784a, 32'shd3d0ec68, 32'shd3cc60f2, 32'shd3c7d5ea, 32'shd3c34b4f, 32'shd3bec121, 
               32'shd3ba3760, 32'shd3b5ae0d, 32'shd3b12526, 32'shd3ac9cad, 32'shd3a814a2, 32'shd3a38d03, 32'shd39f05d3, 32'shd39a7f0f, 
               32'shd395f8ba, 32'shd39172d2, 32'shd38ced57, 32'shd388684a, 32'shd383e3ab, 32'shd37f5f7a, 32'shd37adbb6, 32'shd3765861, 
               32'shd371d579, 32'shd36d52ff, 32'shd368d0f3, 32'shd3644f55, 32'shd35fce26, 32'shd35b4d64, 32'shd356cd11, 32'shd3524d2b, 
               32'shd34dcdb4, 32'shd3494eab, 32'shd344d011, 32'shd34051e5, 32'shd33bd427, 32'shd33756d8, 32'shd332d9f7, 32'shd32e5d85, 
               32'shd329e181, 32'shd32565ec, 32'shd320eac6, 32'shd31c700f, 32'shd317f5c6, 32'shd3137bec, 32'shd30f0280, 32'shd30a8984, 
               32'shd30610f7, 32'shd30198d8, 32'shd2fd2129, 32'shd2f8a9e9, 32'shd2f43318, 32'shd2efbcb6, 32'shd2eb46c3, 32'shd2e6d13f, 
               32'shd2e25c2b, 32'shd2dde786, 32'shd2d97350, 32'shd2d4ff8a, 32'shd2d08c33, 32'shd2cc194c, 32'shd2c7a6d4, 32'shd2c334cc, 
               32'shd2bec333, 32'shd2ba520a, 32'shd2b5e151, 32'shd2b17107, 32'shd2ad012e, 32'shd2a891c4, 32'shd2a422ca, 32'shd29fb440, 
               32'shd29b4626, 32'shd296d87c, 32'shd2926b41, 32'shd28dfe77, 32'shd289921e, 32'shd2852634, 32'shd280babb, 32'shd27c4fb1, 
               32'shd277e518, 32'shd2737af0, 32'shd26f1138, 32'shd26aa7f0, 32'shd2663f19, 32'shd261d6b2, 32'shd25d6ebc, 32'shd2590736, 
               32'shd254a021, 32'shd250397d, 32'shd24bd34a, 32'shd2476d87, 32'shd2430835, 32'shd23ea354, 32'shd23a3ee4, 32'shd235dae4, 
               32'shd2317756, 32'shd22d1439, 32'shd228b18d, 32'shd2244f52, 32'shd21fed88, 32'shd21b8c2f, 32'shd2172b48, 32'shd212cad1, 
               32'shd20e6acc, 32'shd20a0b39, 32'shd205ac17, 32'shd2014d66, 32'shd1fcef27, 32'shd1f89159, 32'shd1f433fd, 32'shd1efd713, 
               32'shd1eb7a9a, 32'shd1e71e93, 32'shd1e2c2fd, 32'shd1de67da, 32'shd1da0d28, 32'shd1d5b2e8, 32'shd1d1591a, 32'shd1ccffbe, 
               32'shd1c8a6d4, 32'shd1c44e5c, 32'shd1bff656, 32'shd1bb9ec2, 32'shd1b747a0, 32'shd1b2f0f1, 32'shd1ae9ab4, 32'shd1aa44e9, 
               32'shd1a5ef90, 32'shd1a19aaa, 32'shd19d4636, 32'shd198f235, 32'shd1949ea6, 32'shd1904b89, 32'shd18bf8e0, 32'shd187a6a8, 
               32'shd18354e4, 32'shd17f0392, 32'shd17ab2b3, 32'shd1766247, 32'shd172124d, 32'shd16dc2c7, 32'shd16973b3, 32'shd1652512, 
               32'shd160d6e5, 32'shd15c892a, 32'shd1583be2, 32'shd153ef0e, 32'shd14fa2ad, 32'shd14b56be, 32'shd1470b44, 32'shd142c03c, 
               32'shd13e75a8, 32'shd13a2b87, 32'shd135e1d9, 32'shd131989f, 32'shd12d4fd9, 32'shd1290786, 32'shd124bfa6, 32'shd120783a, 
               32'shd11c3142, 32'shd117eabd, 32'shd113a4ad, 32'shd10f5f10, 32'shd10b19e7, 32'shd106d531, 32'shd10290f0, 32'shd0fe4d22, 
               32'shd0fa09c9, 32'shd0f5c6e3, 32'shd0f18472, 32'shd0ed4275, 32'shd0e900ec, 32'shd0e4bfd7, 32'shd0e07f36, 32'shd0dc3f0a, 
               32'shd0d7ff51, 32'shd0d3c00e, 32'shd0cf813e, 32'shd0cb42e3, 32'shd0c704fd, 32'shd0c2c78b, 32'shd0be8a8d, 32'shd0ba4e05, 
               32'shd0b611f1, 32'shd0b1d651, 32'shd0ad9b26, 32'shd0a96070, 32'shd0a5262f, 32'shd0a0ec63, 32'shd09cb30b, 32'shd0987a29, 
               32'shd09441bb, 32'shd09009c3, 32'shd08bd23f, 32'shd0879b31, 32'shd0836497, 32'shd07f2e73, 32'shd07af8c4, 32'shd076c38b, 
               32'shd0728ec6, 32'shd06e5a77, 32'shd06a269d, 32'shd065f339, 32'shd061c04a, 32'shd05d8dd1, 32'shd0595bcd, 32'shd0552a3f, 
               32'shd050f926, 32'shd04cc884, 32'shd0489856, 32'shd044689f, 32'shd040395d, 32'shd03c0a91, 32'shd037dc3b, 32'shd033ae5b, 
               32'shd02f80f1, 32'shd02b53fc, 32'shd027277e, 32'shd022fb76, 32'shd01ecfe4, 32'shd01aa4c8, 32'shd0167a22, 32'shd0124ff3, 
               32'shd00e2639, 32'shd009fcf6, 32'shd005d42a, 32'shd001abd3, 32'shcffd83f4, 32'shcff95c8a, 32'shcff53597, 32'shcff10f1b, 
               32'shcfece915, 32'shcfe8c386, 32'shcfe49e6d, 32'shcfe079cc, 32'shcfdc55a1, 32'shcfd831ec, 32'shcfd40eaf, 32'shcfcfebe8, 
               32'shcfcbc999, 32'shcfc7a7c0, 32'shcfc3865e, 32'shcfbf6573, 32'shcfbb4500, 32'shcfb72503, 32'shcfb3057d, 32'shcfaee66f, 
               32'shcfaac7d8, 32'shcfa6a9b8, 32'shcfa28c10, 32'shcf9e6edf, 32'shcf9a5225, 32'shcf9635e2, 32'shcf921a17, 32'shcf8dfec4, 
               32'shcf89e3e8, 32'shcf85c984, 32'shcf81af97, 32'shcf7d9622, 32'shcf797d24, 32'shcf75649f, 32'shcf714c91, 32'shcf6d34fb, 
               32'shcf691ddd, 32'shcf650736, 32'shcf60f108, 32'shcf5cdb51, 32'shcf58c613, 32'shcf54b14d, 32'shcf509cfe, 32'shcf4c8928, 
               32'shcf4875ca, 32'shcf4462e4, 32'shcf405077, 32'shcf3c3e82, 32'shcf382d05, 32'shcf341c00, 32'shcf300b74, 32'shcf2bfb60, 
               32'shcf27ebc5, 32'shcf23dca2, 32'shcf1fcdf8, 32'shcf1bbfc6, 32'shcf17b20d, 32'shcf13a4cd, 32'shcf0f9805, 32'shcf0b8bb7, 
               32'shcf077fe1, 32'shcf037483, 32'shceff699f, 32'shcefb5f34, 32'shcef75541, 32'shcef34bc8, 32'shceef42c7, 32'shceeb3a40, 
               32'shcee73231, 32'shcee32a9c, 32'shcedf2380, 32'shcedb1cde, 32'shced716b4, 32'shced31104, 32'shcecf0bcd, 32'shcecb070f, 
               32'shcec702cb, 32'shcec2ff01, 32'shcebefbb0, 32'shcebaf8d8, 32'shceb6f67a, 32'shceb2f496, 32'shceaef32b, 32'shceaaf23a, 
               32'shcea6f1c2, 32'shcea2f1c5, 32'shce9ef241, 32'shce9af337, 32'shce96f4a7, 32'shce92f691, 32'shce8ef8f4, 32'shce8afbd2, 
               32'shce86ff2a, 32'shce8302fc, 32'shce7f0748, 32'shce7b0c0e, 32'shce77114e, 32'shce731709, 32'shce6f1d3d, 32'shce6b23ec, 
               32'shce672b16, 32'shce6332ba, 32'shce5f3ad8, 32'shce5b4370, 32'shce574c84, 32'shce535611, 32'shce4f6019, 32'shce4b6a9c, 
               32'shce47759a, 32'shce438112, 32'shce3f8d05, 32'shce3b9973, 32'shce37a65b, 32'shce33b3be, 32'shce2fc19c, 32'shce2bcff5, 
               32'shce27dec9, 32'shce23ee18, 32'shce1ffde2, 32'shce1c0e28, 32'shce181ee8, 32'shce143023, 32'shce1041d9, 32'shce0c540b, 
               32'shce0866b8, 32'shce0479e0, 32'shce008d84, 32'shcdfca1a3, 32'shcdf8b63d, 32'shcdf4cb53, 32'shcdf0e0e4, 32'shcdecf6f1, 
               32'shcde90d79, 32'shcde5247d, 32'shcde13bfd, 32'shcddd53f8, 32'shcdd96c6f, 32'shcdd58562, 32'shcdd19ed0, 32'shcdcdb8ba, 
               32'shcdc9d320, 32'shcdc5ee02, 32'shcdc20960, 32'shcdbe253a, 32'shcdba4190, 32'shcdb65e62, 32'shcdb27bb0, 32'shcdae997a, 
               32'shcdaab7c0, 32'shcda6d683, 32'shcda2f5c2, 32'shcd9f157d, 32'shcd9b35b4, 32'shcd975668, 32'shcd937798, 32'shcd8f9944, 
               32'shcd8bbb6d, 32'shcd87de12, 32'shcd840134, 32'shcd8024d3, 32'shcd7c48ee, 32'shcd786d85, 32'shcd74929a, 32'shcd70b82b, 
               32'shcd6cde39, 32'shcd6904c3, 32'shcd652bcb, 32'shcd61534f, 32'shcd5d7b50, 32'shcd59a3ce, 32'shcd55ccca, 32'shcd51f642, 
               32'shcd4e2037, 32'shcd4a4aa9, 32'shcd467599, 32'shcd42a105, 32'shcd3eccef, 32'shcd3af956, 32'shcd37263a, 32'shcd33539c, 
               32'shcd2f817b, 32'shcd2bafd7, 32'shcd27deb0, 32'shcd240e08, 32'shcd203ddc, 32'shcd1c6e2e, 32'shcd189efe, 32'shcd14d04b, 
               32'shcd110216, 32'shcd0d345f, 32'shcd096725, 32'shcd059a6a, 32'shcd01ce2b, 32'shccfe026b, 32'shccfa3729, 32'shccf66c64, 
               32'shccf2a21d, 32'shcceed855, 32'shcceb0f0a, 32'shcce7463e, 32'shcce37def, 32'shccdfb61f, 32'shccdbeecc, 32'shccd827f8, 
               32'shccd461a2, 32'shccd09bcb, 32'shccccd671, 32'shccc91196, 32'shccc54d3a, 32'shccc1895c, 32'shccbdc5fc, 32'shccba031a, 
               32'shccb640b8, 32'shccb27ed3, 32'shccaebd6e, 32'shccaafc87, 32'shcca73c1e, 32'shcca37c35, 32'shcc9fbcca, 32'shcc9bfddd, 
               32'shcc983f70, 32'shcc948182, 32'shcc90c412, 32'shcc8d0721, 32'shcc894aaf, 32'shcc858ebc, 32'shcc81d349, 32'shcc7e1854, 
               32'shcc7a5dde, 32'shcc76a3e8, 32'shcc72ea70, 32'shcc6f3178, 32'shcc6b78ff, 32'shcc67c105, 32'shcc64098b, 32'shcc605290, 
               32'shcc5c9c14, 32'shcc58e618, 32'shcc55309b, 32'shcc517b9e, 32'shcc4dc720, 32'shcc4a1322, 32'shcc465fa3, 32'shcc42aca4, 
               32'shcc3efa25, 32'shcc3b4825, 32'shcc3796a5, 32'shcc33e5a5, 32'shcc303524, 32'shcc2c8524, 32'shcc28d5a3, 32'shcc2526a2, 
               32'shcc217822, 32'shcc1dca21, 32'shcc1a1ca0, 32'shcc166f9f, 32'shcc12c31f, 32'shcc0f171e, 32'shcc0b6b9e, 32'shcc07c09e, 
               32'shcc04161e, 32'shcc006c1e, 32'shcbfcc29f, 32'shcbf919a0, 32'shcbf57121, 32'shcbf1c923, 32'shcbee21a5, 32'shcbea7aa7, 
               32'shcbe6d42b, 32'shcbe32e2e, 32'shcbdf88b3, 32'shcbdbe3b7, 32'shcbd83f3d, 32'shcbd49b43, 32'shcbd0f7ca, 32'shcbcd54d2, 
               32'shcbc9b25a, 32'shcbc61064, 32'shcbc26eee, 32'shcbbecdf9, 32'shcbbb2d85, 32'shcbb78d92, 32'shcbb3ee20, 32'shcbb04f2f, 
               32'shcbacb0bf, 32'shcba912d1, 32'shcba57563, 32'shcba1d877, 32'shcb9e3c0b, 32'shcb9aa021, 32'shcb9704b9, 32'shcb9369d1, 
               32'shcb8fcf6b, 32'shcb8c3587, 32'shcb889c23, 32'shcb850342, 32'shcb816ae1, 32'shcb7dd303, 32'shcb7a3ba5, 32'shcb76a4ca, 
               32'shcb730e70, 32'shcb6f7898, 32'shcb6be341, 32'shcb684e6c, 32'shcb64ba19, 32'shcb612648, 32'shcb5d92f8, 32'shcb5a002b, 
               32'shcb566ddf, 32'shcb52dc15, 32'shcb4f4acd, 32'shcb4bba08, 32'shcb4829c4, 32'shcb449a02, 32'shcb410ac3, 32'shcb3d7c05, 
               32'shcb39edca, 32'shcb366011, 32'shcb32d2da, 32'shcb2f4626, 32'shcb2bb9f4, 32'shcb282e44, 32'shcb24a316, 32'shcb21186b, 
               32'shcb1d8e43, 32'shcb1a049d, 32'shcb167b79, 32'shcb12f2d8, 32'shcb0f6aba, 32'shcb0be31e, 32'shcb085c05, 32'shcb04d56e, 
               32'shcb014f5b, 32'shcafdc9ca, 32'shcafa44bc, 32'shcaf6c030, 32'shcaf33c28, 32'shcaefb8a2, 32'shcaec35a0, 32'shcae8b320, 
               32'shcae53123, 32'shcae1afaa, 32'shcade2eb3, 32'shcadaae40, 32'shcad72e4f, 32'shcad3aee2, 32'shcad02ff8, 32'shcaccb191, 
               32'shcac933ae, 32'shcac5b64e, 32'shcac23971, 32'shcabebd17, 32'shcabb4141, 32'shcab7c5ef, 32'shcab44b1f, 32'shcab0d0d4, 
               32'shcaad570c, 32'shcaa9ddc7, 32'shcaa66506, 32'shcaa2ecc9, 32'shca9f750f, 32'shca9bfdd9, 32'shca988727, 32'shca9510f8, 
               32'shca919b4e, 32'shca8e2627, 32'shca8ab184, 32'shca873d65, 32'shca83c9ca, 32'shca8056b3, 32'shca7ce420, 32'shca797211, 
               32'shca760086, 32'shca728f7f, 32'shca6f1efc, 32'shca6baefd, 32'shca683f83, 32'shca64d08d, 32'shca61621b, 32'shca5df42d, 
               32'shca5a86c4, 32'shca5719df, 32'shca53ad7e, 32'shca5041a2, 32'shca4cd64b, 32'shca496b77, 32'shca460129, 32'shca42975f, 
               32'shca3f2e19, 32'shca3bc559, 32'shca385d1d, 32'shca34f565, 32'shca318e32, 32'shca2e2784, 32'shca2ac15b, 32'shca275bb7, 
               32'shca23f698, 32'shca2091fd, 32'shca1d2de7, 32'shca19ca57, 32'shca16674b, 32'shca1304c4, 32'shca0fa2c3, 32'shca0c4146, 
               32'shca08e04f, 32'shca057fdd, 32'shca021fef, 32'shc9fec088, 32'shc9fb61a5, 32'shc9f80348, 32'shc9f4a570, 32'shc9f1481d, 
               32'shc9edeb50, 32'shc9ea8f08, 32'shc9e73346, 32'shc9e3d809, 32'shc9e07d51, 32'shc9dd231f, 32'shc9d9c973, 32'shc9d6704c, 
               32'shc9d317ab, 32'shc9cfbf90, 32'shc9cc67fa, 32'shc9c910ea, 32'shc9c5ba60, 32'shc9c2645c, 32'shc9bf0edd, 32'shc9bbb9e5, 
               32'shc9b86572, 32'shc9b51185, 32'shc9b1be1e, 32'shc9ae6b3d, 32'shc9ab18e3, 32'shc9a7c70e, 32'shc9a475bf, 32'shc9a124f7, 
               32'shc99dd4b4, 32'shc99a84f8, 32'shc99735c2, 32'shc993e712, 32'shc99098e9, 32'shc98d4b45, 32'shc989fe29, 32'shc986b192, 
               32'shc9836582, 32'shc98019f8, 32'shc97ccef5, 32'shc9798479, 32'shc9763a83, 32'shc972f113, 32'shc96fa82a, 32'shc96c5fc8, 
               32'shc96917ec, 32'shc965d097, 32'shc96289c9, 32'shc95f4382, 32'shc95bfdc1, 32'shc958b887, 32'shc95573d4, 32'shc9522fa8, 
               32'shc94eec03, 32'shc94ba8e5, 32'shc948664d, 32'shc945243d, 32'shc941e2b4, 32'shc93ea1b2, 32'shc93b6137, 32'shc9382143, 
               32'shc934e1d6, 32'shc931a2f0, 32'shc92e6492, 32'shc92b26bb, 32'shc927e96b, 32'shc924aca3, 32'shc9217062, 32'shc91e34a8, 
               32'shc91af976, 32'shc917becb, 32'shc91484a8, 32'shc9114b0c, 32'shc90e11f7, 32'shc90ad96b, 32'shc907a166, 32'shc90469e8, 
               32'shc90132f2, 32'shc8fdfc84, 32'shc8fac69e, 32'shc8f7913f, 32'shc8f45c68, 32'shc8f12819, 32'shc8edf452, 32'shc8eac112, 
               32'shc8e78e5b, 32'shc8e45c2c, 32'shc8e12a84, 32'shc8ddf965, 32'shc8dac8cd, 32'shc8d798be, 32'shc8d46936, 32'shc8d13a37, 
               32'shc8ce0bc0, 32'shc8caddd1, 32'shc8c7b06b, 32'shc8c4838d, 32'shc8c15736, 32'shc8be2b69, 32'shc8bb0023, 32'shc8b7d566, 
               32'shc8b4ab32, 32'shc8b18185, 32'shc8ae5862, 32'shc8ab2fc6, 32'shc8a807b4, 32'shc8a4e029, 32'shc8a1b928, 32'shc89e92af, 
               32'shc89b6cbf, 32'shc8984757, 32'shc8952278, 32'shc891fe22, 32'shc88eda54, 32'shc88bb710, 32'shc8889454, 32'shc8857221, 
               32'shc8825077, 32'shc87f2f56, 32'shc87c0ebd, 32'shc878eeae, 32'shc875cf28, 32'shc872b02b, 32'shc86f91b7, 32'shc86c73cc, 
               32'shc869566a, 32'shc8663991, 32'shc8631d42, 32'shc860017b, 32'shc85ce63e, 32'shc859cb8a, 32'shc856b160, 32'shc85397bf, 
               32'shc8507ea7, 32'shc84d6619, 32'shc84a4e14, 32'shc8473698, 32'shc8441fa6, 32'shc841093e, 32'shc83df35f, 32'shc83ade0a, 
               32'shc837c93e, 32'shc834b4fc, 32'shc831a143, 32'shc82e8e15, 32'shc82b7b70, 32'shc8286954, 32'shc82557c3, 32'shc82246bb, 
               32'shc81f363d, 32'shc81c2649, 32'shc81916df, 32'shc81607ff, 32'shc812f9a9, 32'shc80febdd, 32'shc80cde9b, 32'shc809d1e3, 
               32'shc806c5b5, 32'shc803ba11, 32'shc800aef7, 32'shc7fda468, 32'shc7fa9a62, 32'shc7f790e7, 32'shc7f487f6, 32'shc7f17f8f, 
               32'shc7ee77b3, 32'shc7eb7061, 32'shc7e8699a, 32'shc7e5635c, 32'shc7e25daa, 32'shc7df5881, 32'shc7dc53e3, 32'shc7d94fd0, 
               32'shc7d64c47, 32'shc7d34949, 32'shc7d046d6, 32'shc7cd44ed, 32'shc7ca438f, 32'shc7c742bb, 32'shc7c44272, 32'shc7c142b4, 
               32'shc7be4381, 32'shc7bb44d8, 32'shc7b846ba, 32'shc7b54928, 32'shc7b24c20, 32'shc7af4fa3, 32'shc7ac53b1, 32'shc7a9584a, 
               32'shc7a65d6e, 32'shc7a3631d, 32'shc7a06957, 32'shc79d701c, 32'shc79a776c, 32'shc7977f48, 32'shc79487ae, 32'shc79190a0, 
               32'shc78e9a1d, 32'shc78ba425, 32'shc788aeb9, 32'shc785b9d8, 32'shc782c582, 32'shc77fd1b8, 32'shc77cde79, 32'shc779ebc5, 
               32'shc776f99d, 32'shc7740801, 32'shc77116f0, 32'shc76e266b, 32'shc76b3671, 32'shc7684702, 32'shc7655820, 32'shc76269c9, 
               32'shc75f7bfe, 32'shc75c8ebe, 32'shc759a20a, 32'shc756b5e2, 32'shc753ca46, 32'shc750df36, 32'shc74df4b1, 32'shc74b0ab9, 
               32'shc748214c, 32'shc745386b, 32'shc7425016, 32'shc73f684e, 32'shc73c8111, 32'shc7399a60, 32'shc736b43c, 32'shc733cea3, 
               32'shc730e997, 32'shc72e0517, 32'shc72b2123, 32'shc7283dbb, 32'shc7255ae0, 32'shc7227890, 32'shc71f96ce, 32'shc71cb597, 
               32'shc719d4ed, 32'shc716f4cf, 32'shc714153e, 32'shc7113639, 32'shc70e57c0, 32'shc70b79d4, 32'shc7089c75, 32'shc705bfa2, 
               32'shc702e35c, 32'shc70007a2, 32'shc6fd2c75, 32'shc6fa51d5, 32'shc6f777c1, 32'shc6f49e3a, 32'shc6f1c540, 32'shc6eeecd3, 
               32'shc6ec14f2, 32'shc6e93d9e, 32'shc6e666d7, 32'shc6e3909d, 32'shc6e0baf0, 32'shc6dde5d0, 32'shc6db113d, 32'shc6d83d37, 
               32'shc6d569be, 32'shc6d296d1, 32'shc6cfc472, 32'shc6ccf2a1, 32'shc6ca215c, 32'shc6c750a4, 32'shc6c4807a, 32'shc6c1b0dd, 
               32'shc6bee1cd, 32'shc6bc134a, 32'shc6b94554, 32'shc6b677ec, 32'shc6b3ab12, 32'shc6b0dec4, 32'shc6ae1304, 32'shc6ab47d2, 
               32'shc6a87d2d, 32'shc6a5b315, 32'shc6a2e98b, 32'shc6a0208f, 32'shc69d5820, 32'shc69a903e, 32'shc697c8eb, 32'shc6950224, 
               32'shc6923bec, 32'shc68f7641, 32'shc68cb124, 32'shc689ec95, 32'shc6872894, 32'shc6846520, 32'shc681a23a, 32'shc67edfe2, 
               32'shc67c1e18, 32'shc6795cdc, 32'shc6769c2e, 32'shc673dc0d, 32'shc6711c7b, 32'shc66e5d77, 32'shc66b9f01, 32'shc668e119, 
               32'shc66623be, 32'shc66366f3, 32'shc660aab5, 32'shc65def05, 32'shc65b33e4, 32'shc6587951, 32'shc655bf4c, 32'shc65305d5, 
               32'shc6504ced, 32'shc64d9493, 32'shc64adcc7, 32'shc648258a, 32'shc6456edb, 32'shc642b8bb, 32'shc6400329, 32'shc63d4e26, 
               32'shc63a99b1, 32'shc637e5ca, 32'shc6353273, 32'shc6327faa, 32'shc62fcd6f, 32'shc62d1bc3, 32'shc62a6aa6, 32'shc627ba17, 
               32'shc6250a18, 32'shc6225aa6, 32'shc61fabc4, 32'shc61cfd71, 32'shc61a4fac, 32'shc617a276, 32'shc614f5cf, 32'shc61249b7, 
               32'shc60f9e2e, 32'shc60cf334, 32'shc60a48c9, 32'shc6079eed, 32'shc604f5a0, 32'shc6024ce2, 32'shc5ffa4b3, 32'shc5fcfd13, 
               32'shc5fa5603, 32'shc5f7af81, 32'shc5f5098f, 32'shc5f2642c, 32'shc5efbf58, 32'shc5ed1b13, 32'shc5ea775e, 32'shc5e7d438, 
               32'shc5e531a1, 32'shc5e28f9a, 32'shc5dfee22, 32'shc5dd4d3a, 32'shc5daace1, 32'shc5d80d17, 32'shc5d56ddd, 32'shc5d2cf33, 
               32'shc5d03118, 32'shc5cd938c, 32'shc5caf690, 32'shc5c85a24, 32'shc5c5be47, 32'shc5c322fb, 32'shc5c0883d, 32'shc5bdee10, 
               32'shc5bb5472, 32'shc5b8bb64, 32'shc5b622e6, 32'shc5b38af8, 32'shc5b0f399, 32'shc5ae5ccb, 32'shc5abc68c, 32'shc5a930dd, 
               32'shc5a69bbe, 32'shc5a4072f, 32'shc5a17330, 32'shc59edfc2, 32'shc59c4ce3, 32'shc599ba94, 32'shc59728d5, 32'shc59497a7, 
               32'shc5920708, 32'shc58f76fa, 32'shc58ce77c, 32'shc58a588e, 32'shc587ca31, 32'shc5853c63, 32'shc582af26, 32'shc580227a, 
               32'shc57d965d, 32'shc57b0ad1, 32'shc5787fd6, 32'shc575f56b, 32'shc5736b90, 32'shc570e246, 32'shc56e598c, 32'shc56bd163, 
               32'shc56949ca, 32'shc566c2c2, 32'shc5643c4a, 32'shc561b663, 32'shc55f310d, 32'shc55cac47, 32'shc55a2812, 32'shc557a46e, 
               32'shc555215a, 32'shc5529ed7, 32'shc5501ce5, 32'shc54d9b84, 32'shc54b1ab4, 32'shc5489a74, 32'shc5461ac6, 32'shc5439ba8, 
               32'shc5411d1b, 32'shc53e9f1f, 32'shc53c21b4, 32'shc539a4da, 32'shc5372891, 32'shc534acd9, 32'shc53231b3, 32'shc52fb71d, 
               32'shc52d3d18, 32'shc52ac3a5, 32'shc5284ac3, 32'shc525d272, 32'shc5235ab2, 32'shc520e383, 32'shc51e6ce6, 32'shc51bf6da, 
               32'shc519815f, 32'shc5170c75, 32'shc514981d, 32'shc5122457, 32'shc50fb121, 32'shc50d3e7d, 32'shc50acc6b, 32'shc5085aea, 
               32'shc505e9fb, 32'shc503799d, 32'shc50109d0, 32'shc4fe9a95, 32'shc4fc2bec, 32'shc4f9bdd4, 32'shc4f7504e, 32'shc4f4e35a, 
               32'shc4f276f7, 32'shc4f00b27, 32'shc4ed9fe7, 32'shc4eb353a, 32'shc4e8cb1e, 32'shc4e66194, 32'shc4e3f89c, 32'shc4e19036, 
               32'shc4df2862, 32'shc4dcc11f, 32'shc4da5a6f, 32'shc4d7f450, 32'shc4d58ec3, 32'shc4d329c9, 32'shc4d0c560, 32'shc4ce6189, 
               32'shc4cbfe45, 32'shc4c99b92, 32'shc4c73972, 32'shc4c4d7e4, 32'shc4c276e8, 32'shc4c0167e, 32'shc4bdb6a6, 32'shc4bb5760, 
               32'shc4b8f8ad, 32'shc4b69a8c, 32'shc4b43cfd, 32'shc4b1e001, 32'shc4af8397, 32'shc4ad27bf, 32'shc4aacc7a, 32'shc4a871c7, 
               32'shc4a617a6, 32'shc4a3be18, 32'shc4a1651c, 32'shc49f0cb3, 32'shc49cb4dd, 32'shc49a5d98, 32'shc49806e7, 32'shc495b0c8, 
               32'shc4935b3c, 32'shc4910642, 32'shc48eb1db, 32'shc48c5e06, 32'shc48a0ac4, 32'shc487b815, 32'shc48565f9, 32'shc4831470, 
               32'shc480c379, 32'shc47e7315, 32'shc47c2344, 32'shc479d405, 32'shc477855a, 32'shc4753741, 32'shc472e9bc, 32'shc4709cc9, 
               32'shc46e5069, 32'shc46c049d, 32'shc469b963, 32'shc4676ebc, 32'shc46524a9, 32'shc462db28, 32'shc460923b, 32'shc45e49e0, 
               32'shc45c0219, 32'shc459bae5, 32'shc4577444, 32'shc4552e36, 32'shc452e8bc, 32'shc450a3d4, 32'shc44e5f80, 32'shc44c1bc0, 
               32'shc449d892, 32'shc44795f8, 32'shc44553f2, 32'shc443127e, 32'shc440d19e, 32'shc43e9152, 32'shc43c5199, 32'shc43a1273, 
               32'shc437d3e1, 32'shc43595e3, 32'shc4335877, 32'shc4311ba0, 32'shc42edf5c, 32'shc42ca3ac, 32'shc42a688f, 32'shc4282e06, 
               32'shc425f410, 32'shc423baae, 32'shc42181e0, 32'shc41f49a6, 32'shc41d11ff, 32'shc41adaed, 32'shc418a46d, 32'shc4166e82, 
               32'shc414392b, 32'shc4120467, 32'shc40fd037, 32'shc40d9c9c, 32'shc40b6994, 32'shc4093720, 32'shc4070540, 32'shc404d3f4, 
               32'shc402a33c, 32'shc4007318, 32'shc3fe4388, 32'shc3fc148c, 32'shc3f9e624, 32'shc3f7b850, 32'shc3f58b10, 32'shc3f35e65, 
               32'shc3f1324e, 32'shc3ef06cb, 32'shc3ecdbdc, 32'shc3eab181, 32'shc3e887bb, 32'shc3e65e88, 32'shc3e435ea, 32'shc3e20de1, 
               32'shc3dfe66c, 32'shc3ddbf8b, 32'shc3db993e, 32'shc3d97386, 32'shc3d74e62, 32'shc3d529d3, 32'shc3d305d8, 32'shc3d0e272, 
               32'shc3cebfa0, 32'shc3cc9d63, 32'shc3ca7bba, 32'shc3c85aa6, 32'shc3c63a26, 32'shc3c41a3b, 32'shc3c1fae5, 32'shc3bfdc23, 
               32'shc3bdbdf6, 32'shc3bba05e, 32'shc3b9835a, 32'shc3b766eb, 32'shc3b54b11, 32'shc3b32fcb, 32'shc3b1151b, 32'shc3aefaff, 
               32'shc3ace178, 32'shc3aac885, 32'shc3a8b028, 32'shc3a6985f, 32'shc3a4812c, 32'shc3a26a8d, 32'shc3a05484, 32'shc39e3f0f, 
               32'shc39c2a2f, 32'shc39a15e4, 32'shc398022f, 32'shc395ef0e, 32'shc393dc82, 32'shc391ca8c, 32'shc38fb92a, 32'shc38da85e, 
               32'shc38b9827, 32'shc3898885, 32'shc3877978, 32'shc3856b01, 32'shc3835d1e, 32'shc3814fd1, 32'shc37f4319, 32'shc37d36f7, 
               32'shc37b2b6a, 32'shc3792072, 32'shc377160f, 32'shc3750c42, 32'shc373030a, 32'shc370fa68, 32'shc36ef25b, 32'shc36ceae3, 
               32'shc36ae401, 32'shc368ddb4, 32'shc366d7fd, 32'shc364d2dc, 32'shc362ce50, 32'shc360ca59, 32'shc35ec6f8, 32'shc35cc42d, 
               32'shc35ac1f7, 32'shc358c057, 32'shc356bf4d, 32'shc354bed8, 32'shc352bef9, 32'shc350bfaf, 32'shc34ec0fc, 32'shc34cc2de, 
               32'shc34ac556, 32'shc348c864, 32'shc346cc07, 32'shc344d041, 32'shc342d510, 32'shc340da75, 32'shc33ee070, 32'shc33ce701, 
               32'shc33aee27, 32'shc338f5e4, 32'shc336fe37, 32'shc3350720, 32'shc333109e, 32'shc3311ab3, 32'shc32f255e, 32'shc32d309e, 
               32'shc32b3c75, 32'shc32948e2, 32'shc32755e5, 32'shc325637f, 32'shc32371ae, 32'shc3218073, 32'shc31f8fcf, 32'shc31d9fc1, 
               32'shc31bb049, 32'shc319c168, 32'shc317d31c, 32'shc315e567, 32'shc313f848, 32'shc3120bc0, 32'shc3101fce, 32'shc30e3472, 
               32'shc30c49ad, 32'shc30a5f7e, 32'shc30875e5, 32'shc3068ce3, 32'shc304a477, 32'shc302bca2, 32'shc300d563, 32'shc2feeebb, 
               32'shc2fd08a9, 32'shc2fb232e, 32'shc2f93e4a, 32'shc2f759fc, 32'shc2f57644, 32'shc2f39323, 32'shc2f1b099, 32'shc2efcea6, 
               32'shc2eded49, 32'shc2ec0c82, 32'shc2ea2c53, 32'shc2e84cba, 32'shc2e66db8, 32'shc2e48f4d, 32'shc2e2b178, 32'shc2e0d43b, 
               32'shc2def794, 32'shc2dd1b84, 32'shc2db400a, 32'shc2d96528, 32'shc2d78add, 32'shc2d5b128, 32'shc2d3d80a, 32'shc2d1ff84, 
               32'shc2d02794, 32'shc2ce503b, 32'shc2cc7979, 32'shc2caa34f, 32'shc2c8cdbb, 32'shc2c6f8be, 32'shc2c52459, 32'shc2c3508a, 
               32'shc2c17d52, 32'shc2bfaab2, 32'shc2bdd8a9, 32'shc2bc0737, 32'shc2ba365c, 32'shc2b86618, 32'shc2b6966c, 32'shc2b4c756, 
               32'shc2b2f8d8, 32'shc2b12af1, 32'shc2af5da2, 32'shc2ad90ea, 32'shc2abc4c9, 32'shc2a9f93f, 32'shc2a82e4d, 32'shc2a663f2, 
               32'shc2a49a2e, 32'shc2a2d102, 32'shc2a1086d, 32'shc29f4070, 32'shc29d790a, 32'shc29bb23c, 32'shc299ec05, 32'shc2982665, 
               32'shc296615d, 32'shc2949ced, 32'shc292d914, 32'shc29115d3, 32'shc28f5329, 32'shc28d9117, 32'shc28bcf9c, 32'shc28a0eb9, 
               32'shc2884e6e, 32'shc2868ebb, 32'shc284cf9f, 32'shc283111b, 32'shc281532e, 32'shc27f95d9, 32'shc27dd91c, 32'shc27c1cf7, 
               32'shc27a616a, 32'shc278a674, 32'shc276ec16, 32'shc2753250, 32'shc2737922, 32'shc271c08c, 32'shc270088e, 32'shc26e5127, 
               32'shc26c9a58, 32'shc26ae422, 32'shc2692e83, 32'shc267797c, 32'shc265c50e, 32'shc2641137, 32'shc2625df8, 32'shc260ab51, 
               32'shc25ef943, 32'shc25d47cc, 32'shc25b96ee, 32'shc259e6a7, 32'shc25836f9, 32'shc25687e3, 32'shc254d965, 32'shc2532b7f, 
               32'shc2517e31, 32'shc24fd17c, 32'shc24e255e, 32'shc24c79d9, 32'shc24aceed, 32'shc2492498, 32'shc2477adc, 32'shc245d1b8, 
               32'shc244292c, 32'shc2428139, 32'shc240d9de, 32'shc23f331b, 32'shc23d8cf1, 32'shc23be75f, 32'shc23a4265, 32'shc2389e04, 
               32'shc236fa3b, 32'shc235570b, 32'shc233b473, 32'shc2321274, 32'shc230710d, 32'shc22ed03f, 32'shc22d3009, 32'shc22b906c, 
               32'shc229f167, 32'shc22852fb, 32'shc226b528, 32'shc22517ed, 32'shc2237b4b, 32'shc221df41, 32'shc22043d0, 32'shc21ea8f8, 
               32'shc21d0eb8, 32'shc21b7511, 32'shc219dc03, 32'shc218438e, 32'shc216abb1, 32'shc215146d, 32'shc2137dc2, 32'shc211e7af, 
               32'shc2105236, 32'shc20ebd55, 32'shc20d290d, 32'shc20b955e, 32'shc20a0248, 32'shc2086fca, 32'shc206dde6, 32'shc2054c9b, 
               32'shc203bbe8, 32'shc2022bce, 32'shc2009c4e, 32'shc1ff0d66, 32'shc1fd7f17, 32'shc1fbf161, 32'shc1fa6445, 32'shc1f8d7c1, 
               32'shc1f74bd6, 32'shc1f5c085, 32'shc1f435cc, 32'shc1f2abad, 32'shc1f12227, 32'shc1ef9939, 32'shc1ee10e5, 32'shc1ec892b, 
               32'shc1eb0209, 32'shc1e97b80, 32'shc1e7f591, 32'shc1e6703b, 32'shc1e4eb7e, 32'shc1e3675a, 32'shc1e1e3d0, 32'shc1e060df, 
               32'shc1dede87, 32'shc1dd5cc8, 32'shc1dbdba3, 32'shc1da5b17, 32'shc1d8db25, 32'shc1d75bcb, 32'shc1d5dd0c, 32'shc1d45ee5, 
               32'shc1d2e158, 32'shc1d16464, 32'shc1cfe80a, 32'shc1ce6c49, 32'shc1ccf122, 32'shc1cb7694, 32'shc1c9fca0, 32'shc1c88345, 
               32'shc1c70a84, 32'shc1c5925c, 32'shc1c41ace, 32'shc1c2a3d9, 32'shc1c12d7e, 32'shc1bfb7bc, 32'shc1be4294, 32'shc1bcce06, 
               32'shc1bb5a11, 32'shc1b9e6b6, 32'shc1b873f5, 32'shc1b701cd, 32'shc1b5903f, 32'shc1b41f4a, 32'shc1b2aef0, 32'shc1b13f2f, 
               32'shc1afd007, 32'shc1ae617a, 32'shc1acf386, 32'shc1ab862c, 32'shc1aa196c, 32'shc1a8ad46, 32'shc1a741b9, 32'shc1a5d6c7, 
               32'shc1a46c6e, 32'shc1a302af, 32'shc1a1998a, 32'shc1a030ff, 32'shc19ec90d, 32'shc19d61b6, 32'shc19bfaf9, 32'shc19a94d5, 
               32'shc1992f4c, 32'shc197ca5c, 32'shc1966606, 32'shc195024b, 32'shc1939f29, 32'shc1923ca2, 32'shc190dab4, 32'shc18f7961, 
               32'shc18e18a7, 32'shc18cb888, 32'shc18b5903, 32'shc189fa17, 32'shc1889bc6, 32'shc1873e10, 32'shc185e0f3, 32'shc1848470, 
               32'shc1832888, 32'shc181cd3a, 32'shc1807285, 32'shc17f186c, 32'shc17dbeec, 32'shc17c6607, 32'shc17b0dbb, 32'shc179b60b, 
               32'shc1785ef4, 32'shc1770878, 32'shc175b296, 32'shc1745d4e, 32'shc17308a1, 32'shc171b48e, 32'shc1706115, 32'shc16f0e36, 
               32'shc16dbbf3, 32'shc16c6a49, 32'shc16b193a, 32'shc169c8c5, 32'shc16878eb, 32'shc16729ab, 32'shc165db05, 32'shc1648cfa, 
               32'shc1633f8a, 32'shc161f2b4, 32'shc160a678, 32'shc15f5ad7, 32'shc15e0fd1, 32'shc15cc565, 32'shc15b7b94, 32'shc15a325d, 
               32'shc158e9c1, 32'shc157a1bf, 32'shc1565a58, 32'shc155138c, 32'shc153cd5a, 32'shc15287c3, 32'shc15142c6, 32'shc14ffe64, 
               32'shc14eba9d, 32'shc14d7771, 32'shc14c34df, 32'shc14af2e8, 32'shc149b18b, 32'shc14870ca, 32'shc14730a3, 32'shc145f117, 
               32'shc144b225, 32'shc14373cf, 32'shc1423613, 32'shc140f8f2, 32'shc13fbc6c, 32'shc13e8081, 32'shc13d4530, 32'shc13c0a7b, 
               32'shc13ad060, 32'shc13996e0, 32'shc1385dfb, 32'shc13725b1, 32'shc135ee02, 32'shc134b6ee, 32'shc1338075, 32'shc1324a96, 
               32'shc1311553, 32'shc12fe0ab, 32'shc12eac9d, 32'shc12d792b, 32'shc12c4653, 32'shc12b1417, 32'shc129e276, 32'shc128b16f, 
               32'shc1278104, 32'shc1265134, 32'shc12521ff, 32'shc123f365, 32'shc122c566, 32'shc1219802, 32'shc1206b39, 32'shc11f3f0c, 
               32'shc11e1379, 32'shc11ce882, 32'shc11bbe26, 32'shc11a9465, 32'shc1196b3f, 32'shc11842b5, 32'shc1171ac6, 32'shc115f372, 
               32'shc114ccb9, 32'shc113a69b, 32'shc1128119, 32'shc1115c32, 32'shc11037e6, 32'shc10f1435, 32'shc10df120, 32'shc10ccea6, 
               32'shc10bacc8, 32'shc10a8b85, 32'shc1096add, 32'shc1084ad0, 32'shc1072b5f, 32'shc1060c89, 32'shc104ee4f, 32'shc103d0b0, 
               32'shc102b3ac, 32'shc1019744, 32'shc1007b77, 32'shc0ff6046, 32'shc0fe45b0, 32'shc0fd2bb6, 32'shc0fc1257, 32'shc0faf993, 
               32'shc0f9e16b, 32'shc0f8c9df, 32'shc0f7b2ee, 32'shc0f69c99, 32'shc0f586df, 32'shc0f471c1, 32'shc0f35d3e, 32'shc0f24957, 
               32'shc0f1360b, 32'shc0f0235b, 32'shc0ef1147, 32'shc0edffce, 32'shc0eceef1, 32'shc0ebdeaf, 32'shc0eacf09, 32'shc0e9bfff, 
               32'shc0e8b190, 32'shc0e7a3bd, 32'shc0e69686, 32'shc0e589eb, 32'shc0e47deb, 32'shc0e37287, 32'shc0e267be, 32'shc0e15d92, 
               32'shc0e05401, 32'shc0df4b0b, 32'shc0de42b2, 32'shc0dd3af4, 32'shc0dc33d2, 32'shc0db2d4c, 32'shc0da2762, 32'shc0d92214, 
               32'shc0d81d61, 32'shc0d7194a, 32'shc0d615cf, 32'shc0d512f0, 32'shc0d410ad, 32'shc0d30f05, 32'shc0d20dfa, 32'shc0d10d8a, 
               32'shc0d00db6, 32'shc0cf0e7f, 32'shc0ce0fe3, 32'shc0cd11e3, 32'shc0cc147f, 32'shc0cb17b7, 32'shc0ca1b8a, 32'shc0c91ffa, 
               32'shc0c82506, 32'shc0c72aae, 32'shc0c630f2, 32'shc0c537d1, 32'shc0c43f4d, 32'shc0c34765, 32'shc0c25019, 32'shc0c15969, 
               32'shc0c06355, 32'shc0bf6ddd, 32'shc0be7901, 32'shc0bd84c1, 32'shc0bc911d, 32'shc0bb9e15, 32'shc0baabaa, 32'shc0b9b9da, 
               32'shc0b8c8a7, 32'shc0b7d810, 32'shc0b6e815, 32'shc0b5f8b6, 32'shc0b509f3, 32'shc0b41bcd, 32'shc0b32e42, 32'shc0b24154, 
               32'shc0b15502, 32'shc0b0694c, 32'shc0af7e33, 32'shc0ae93b5, 32'shc0ada9d4, 32'shc0acc08f, 32'shc0abd7e6, 32'shc0aaefda, 
               32'shc0aa086a, 32'shc0a92196, 32'shc0a83b5e, 32'shc0a755c3, 32'shc0a670c4, 32'shc0a58c62, 32'shc0a4a89b, 32'shc0a3c571, 
               32'shc0a2e2e3, 32'shc0a200f2, 32'shc0a11f9d, 32'shc0a03ee4, 32'shc09f5ec8, 32'shc09e7f48, 32'shc09da065, 32'shc09cc21e, 
               32'shc09be473, 32'shc09b0765, 32'shc09a2af3, 32'shc0994f1d, 32'shc09873e4, 32'shc0979948, 32'shc096bf48, 32'shc095e5e4, 
               32'shc0950d1d, 32'shc09434f2, 32'shc0935d64, 32'shc0928672, 32'shc091b01d, 32'shc090da64, 32'shc0900548, 32'shc08f30c8, 
               32'shc08e5ce5, 32'shc08d899f, 32'shc08cb6f5, 32'shc08be4e7, 32'shc08b1376, 32'shc08a42a2, 32'shc089726a, 32'shc088a2cf, 
               32'shc087d3d0, 32'shc087056e, 32'shc08637a9, 32'shc0856a80, 32'shc0849df4, 32'shc083d204, 32'shc08306b2, 32'shc0823bfb, 
               32'shc08171e2, 32'shc080a865, 32'shc07fdf85, 32'shc07f1741, 32'shc07e4f9b, 32'shc07d8890, 32'shc07cc223, 32'shc07bfc52, 
               32'shc07b371e, 32'shc07a7287, 32'shc079ae8c, 32'shc078eb2f, 32'shc078286e, 32'shc0776649, 32'shc076a4c2, 32'shc075e3d7, 
               32'shc0752389, 32'shc07463d8, 32'shc073a4c3, 32'shc072e64c, 32'shc0722871, 32'shc0716b33, 32'shc070ae92, 32'shc06ff28e, 
               32'shc06f3726, 32'shc06e7c5b, 32'shc06dc22e, 32'shc06d089d, 32'shc06c4fa8, 32'shc06b9751, 32'shc06adf97, 32'shc06a2879, 
               32'shc06971f9, 32'shc068bc15, 32'shc06806ce, 32'shc0675225, 32'shc0669e18, 32'shc065eaa8, 32'shc06537d4, 32'shc064859e, 
               32'shc063d405, 32'shc0632309, 32'shc06272aa, 32'shc061c2e7, 32'shc06113c2, 32'shc060653a, 32'shc05fb74e, 32'shc05f0a00, 
               32'shc05e5d4e, 32'shc05db13a, 32'shc05d05c3, 32'shc05c5ae8, 32'shc05bb0ab, 32'shc05b070a, 32'shc05a5e07, 32'shc059b5a1, 
               32'shc0590dd8, 32'shc05866ac, 32'shc057c01d, 32'shc0571a2b, 32'shc05674d6, 32'shc055d01e, 32'shc0552c03, 32'shc0548885, 
               32'shc053e5a5, 32'shc0534361, 32'shc052a1bb, 32'shc05200b2, 32'shc0516045, 32'shc050c077, 32'shc0502145, 32'shc04f82b0, 
               32'shc04ee4b8, 32'shc04e475e, 32'shc04daaa1, 32'shc04d0e81, 32'shc04c72fe, 32'shc04bd818, 32'shc04b3dcf, 32'shc04aa424, 
               32'shc04a0b16, 32'shc04972a5, 32'shc048dad1, 32'shc048439b, 32'shc047ad01, 32'shc0471705, 32'shc04681a6, 32'shc045ece5, 
               32'shc04558c0, 32'shc044c539, 32'shc044324f, 32'shc043a002, 32'shc0430e53, 32'shc0427d41, 32'shc041eccc, 32'shc0415cf4, 
               32'shc040cdba, 32'shc0403f1d, 32'shc03fb11d, 32'shc03f23bb, 32'shc03e96f6, 32'shc03e0ace, 32'shc03d7f44, 32'shc03cf456, 
               32'shc03c6a07, 32'shc03be054, 32'shc03b573f, 32'shc03acec7, 32'shc03a46ed, 32'shc039bfaf, 32'shc0393910, 32'shc038b30d, 
               32'shc0382da8, 32'shc037a8e1, 32'shc03724b6, 32'shc036a129, 32'shc0361e3a, 32'shc0359be8, 32'shc0351a33, 32'shc034991c, 
               32'shc03418a2, 32'shc03398c5, 32'shc0331986, 32'shc0329ae4, 32'shc0321ce0, 32'shc0319f79, 32'shc03122b0, 32'shc030a684, 
               32'shc0302af5, 32'shc02fb004, 32'shc02f35b1, 32'shc02ebbfb, 32'shc02e42e2, 32'shc02dca67, 32'shc02d5289, 32'shc02cdb49, 
               32'shc02c64a6, 32'shc02beea1, 32'shc02b7939, 32'shc02b046f, 32'shc02a9042, 32'shc02a1cb2, 32'shc029a9c1, 32'shc029376c, 
               32'shc028c5b6, 32'shc028549c, 32'shc027e421, 32'shc0277442, 32'shc0270502, 32'shc026965f, 32'shc0262859, 32'shc025baf1, 
               32'shc0254e27, 32'shc024e1fa, 32'shc024766a, 32'shc0240b78, 32'shc023a124, 32'shc023376e, 32'shc022ce54, 32'shc02265d9, 
               32'shc021fdfb, 32'shc02196bb, 32'shc0213018, 32'shc020ca13, 32'shc02064ab, 32'shc01fffe1, 32'shc01f9bb5, 32'shc01f3826, 
               32'shc01ed535, 32'shc01e72e1, 32'shc01e112b, 32'shc01db013, 32'shc01d4f99, 32'shc01cefbb, 32'shc01c907c, 32'shc01c31da, 
               32'shc01bd3d6, 32'shc01b7670, 32'shc01b19a7, 32'shc01abd7c, 32'shc01a61ee, 32'shc01a06fe, 32'shc019acac, 32'shc01952f8, 
               32'shc018f9e1, 32'shc018a168, 32'shc018498c, 32'shc017f24e, 32'shc0179bae, 32'shc01745ac, 32'shc016f047, 32'shc0169b80, 
               32'shc0164757, 32'shc015f3cb, 32'shc015a0dd, 32'shc0154e8d, 32'shc014fcda, 32'shc014abc5, 32'shc0145b4e, 32'shc0140b75, 
               32'shc013bc39, 32'shc0136d9b, 32'shc0131f9b, 32'shc012d238, 32'shc0128574, 32'shc012394c, 32'shc011edc3, 32'shc011a2d8, 
               32'shc011588a, 32'shc0110eda, 32'shc010c5c7, 32'shc0107d53, 32'shc010357c, 32'shc00fee43, 32'shc00fa7a8, 32'shc00f61aa, 
               32'shc00f1c4a, 32'shc00ed788, 32'shc00e9364, 32'shc00e4fde, 32'shc00e0cf5, 32'shc00dcaaa, 32'shc00d88fd, 32'shc00d47ed, 
               32'shc00d077c, 32'shc00cc7a8, 32'shc00c8872, 32'shc00c49da, 32'shc00c0be0, 32'shc00bce83, 32'shc00b91c4, 32'shc00b55a3, 
               32'shc00b1a20, 32'shc00adf3b, 32'shc00aa4f3, 32'shc00a6b49, 32'shc00a323d, 32'shc009f9cf, 32'shc009c1ff, 32'shc0098acc, 
               32'shc0095438, 32'shc0091e41, 32'shc008e8e8, 32'shc008b42d, 32'shc008800f, 32'shc0084c90, 32'shc00819ae, 32'shc007e76a, 
               32'shc007b5c4, 32'shc00784bc, 32'shc0075452, 32'shc0072485, 32'shc006f556, 32'shc006c6c6, 32'shc00698d3, 32'shc0066b7d, 
               32'shc0063ec6, 32'shc00612ad, 32'shc005e731, 32'shc005bc54, 32'shc0059214, 32'shc0056872, 32'shc0053f6e, 32'shc0051707, 
               32'shc004ef3f, 32'shc004c814, 32'shc004a188, 32'shc0047b99, 32'shc0045648, 32'shc0043195, 32'shc0040d80, 32'shc003ea09, 
               32'shc003c72f, 32'shc003a4f4, 32'shc0038356, 32'shc0036256, 32'shc00341f4, 32'shc0032230, 32'shc003030a, 32'shc002e482, 
               32'shc002c697, 32'shc002a94b, 32'shc0028c9c, 32'shc002708c, 32'shc0025519, 32'shc0023a44, 32'shc002200d, 32'shc0020674, 
               32'shc001ed78, 32'shc001d51b, 32'shc001bd5c, 32'shc001a63a, 32'shc0018fb6, 32'shc00179d1, 32'shc0016489, 32'shc0014fdf, 
               32'shc0013bd3, 32'shc0012865, 32'shc0011594, 32'shc0010362, 32'shc000f1ce, 32'shc000e0d7, 32'shc000d07e, 32'shc000c0c4, 
               32'shc000b1a7, 32'shc000a328, 32'shc0009547, 32'shc0008804, 32'shc0007b5f, 32'shc0006f57, 32'shc00063ee, 32'shc0005922, 
               32'shc0004ef5, 32'shc0004565, 32'shc0003c74, 32'shc0003420, 32'shc0002c6a, 32'shc0002552, 32'shc0001ed8, 32'shc00018fb, 
               32'shc00013bd, 32'shc0000f1d, 32'shc0000b1a, 32'shc00007b6, 32'shc00004ef, 32'shc00002c7, 32'shc000013c, 32'shc000004f
            };

            reg signed [31:0] W_Im_table[8192] = '{
               32'sh00000000, 32'shfff9b781, 32'shfff36f02, 32'shffed2684, 32'shffe6de05, 32'shffe09587, 32'shffda4d09, 32'shffd4048c, 
               32'shffcdbc0f, 32'shffc77392, 32'shffc12b16, 32'shffbae29a, 32'shffb49a1f, 32'shffae51a5, 32'shffa8092c, 32'shffa1c0b4, 
               32'shff9b783c, 32'shff952fc5, 32'shff8ee750, 32'shff889edb, 32'shff825668, 32'shff7c0df6, 32'shff75c585, 32'shff6f7d16, 
               32'shff6934a8, 32'shff62ec3b, 32'shff5ca3d0, 32'shff565b66, 32'shff5012fe, 32'shff49ca98, 32'shff438234, 32'shff3d39d1, 
               32'shff36f170, 32'shff30a911, 32'shff2a60b4, 32'shff24185a, 32'shff1dd001, 32'shff1787aa, 32'shff113f56, 32'shff0af704, 
               32'shff04aeb5, 32'shfefe6668, 32'shfef81e1d, 32'shfef1d5d5, 32'shfeeb8d8f, 32'shfee5454c, 32'shfedefd0c, 32'shfed8b4cf, 
               32'shfed26c94, 32'shfecc245d, 32'shfec5dc28, 32'shfebf93f6, 32'shfeb94bc8, 32'shfeb3039d, 32'shfeacbb74, 32'shfea6734f, 
               32'shfea02b2e, 32'shfe99e310, 32'shfe939af5, 32'shfe8d52de, 32'shfe870aca, 32'shfe80c2ba, 32'shfe7a7aae, 32'shfe7432a5, 
               32'shfe6deaa1, 32'shfe67a2a0, 32'shfe615aa3, 32'shfe5b12aa, 32'shfe54cab5, 32'shfe4e82c4, 32'shfe483ad8, 32'shfe41f2ef, 
               32'shfe3bab0b, 32'shfe35632c, 32'shfe2f1b50, 32'shfe28d379, 32'shfe228ba7, 32'shfe1c43da, 32'shfe15fc11, 32'shfe0fb44c, 
               32'shfe096c8d, 32'shfe0324d2, 32'shfdfcdd1d, 32'shfdf6956c, 32'shfdf04dc0, 32'shfdea0619, 32'shfde3be78, 32'shfddd76dc, 
               32'shfdd72f45, 32'shfdd0e7b3, 32'shfdcaa027, 32'shfdc458a0, 32'shfdbe111e, 32'shfdb7c9a3, 32'shfdb1822c, 32'shfdab3abc, 
               32'shfda4f351, 32'shfd9eabec, 32'shfd98648d, 32'shfd921d34, 32'shfd8bd5e1, 32'shfd858e94, 32'shfd7f474d, 32'shfd79000d, 
               32'shfd72b8d2, 32'shfd6c719e, 32'shfd662a70, 32'shfd5fe348, 32'shfd599c28, 32'shfd53550d, 32'shfd4d0df9, 32'shfd46c6ec, 
               32'shfd407fe6, 32'shfd3a38e6, 32'shfd33f1ed, 32'shfd2daafb, 32'shfd276410, 32'shfd211d2c, 32'shfd1ad650, 32'shfd148f7a, 
               32'shfd0e48ab, 32'shfd0801e4, 32'shfd01bb24, 32'shfcfb746c, 32'shfcf52dbb, 32'shfceee711, 32'shfce8a06f, 32'shfce259d5, 
               32'shfcdc1342, 32'shfcd5ccb7, 32'shfccf8634, 32'shfcc93fb9, 32'shfcc2f945, 32'shfcbcb2da, 32'shfcb66c77, 32'shfcb0261b, 
               32'shfca9dfc8, 32'shfca3997e, 32'shfc9d533b, 32'shfc970d01, 32'shfc90c6cf, 32'shfc8a80a6, 32'shfc843a85, 32'shfc7df46d, 
               32'shfc77ae5e, 32'shfc716857, 32'shfc6b2259, 32'shfc64dc64, 32'shfc5e9678, 32'shfc585094, 32'shfc520aba, 32'shfc4bc4e9, 
               32'shfc457f21, 32'shfc3f3962, 32'shfc38f3ac, 32'shfc32ae00, 32'shfc2c685d, 32'shfc2622c4, 32'shfc1fdd34, 32'shfc1997ae, 
               32'shfc135231, 32'shfc0d0cbe, 32'shfc06c754, 32'shfc0081f5, 32'shfbfa3c9f, 32'shfbf3f753, 32'shfbedb212, 32'shfbe76cda, 
               32'shfbe127ac, 32'shfbdae289, 32'shfbd49d70, 32'shfbce5861, 32'shfbc8135c, 32'shfbc1ce62, 32'shfbbb8973, 32'shfbb5448d, 
               32'shfbaeffb3, 32'shfba8bae3, 32'shfba2761e, 32'shfb9c3163, 32'shfb95ecb4, 32'shfb8fa80f, 32'shfb896375, 32'shfb831ee6, 
               32'shfb7cda63, 32'shfb7695ea, 32'shfb70517d, 32'shfb6a0d1b, 32'shfb63c8c4, 32'shfb5d8479, 32'shfb574039, 32'shfb50fc04, 
               32'shfb4ab7db, 32'shfb4473be, 32'shfb3e2fac, 32'shfb37eba7, 32'shfb31a7ac, 32'shfb2b63be, 32'shfb251fdc, 32'shfb1edc06, 
               32'shfb18983b, 32'shfb12547d, 32'shfb0c10cb, 32'shfb05cd25, 32'shfaff898c, 32'shfaf945ff, 32'shfaf3027e, 32'shfaecbf0a, 
               32'shfae67ba2, 32'shfae03847, 32'shfad9f4f8, 32'shfad3b1b6, 32'shfacd6e81, 32'shfac72b59, 32'shfac0e83d, 32'shfabaa52f, 
               32'shfab4622d, 32'shfaae1f39, 32'shfaa7dc52, 32'shfaa19978, 32'shfa9b56ab, 32'shfa9513eb, 32'shfa8ed139, 32'shfa888e95, 
               32'shfa824bfd, 32'shfa7c0974, 32'shfa75c6f8, 32'shfa6f8489, 32'shfa694229, 32'shfa62ffd6, 32'shfa5cbd91, 32'shfa567b5a, 
               32'shfa503930, 32'shfa49f715, 32'shfa43b508, 32'shfa3d7309, 32'shfa373119, 32'shfa30ef36, 32'shfa2aad62, 32'shfa246b9d, 
               32'shfa1e29e5, 32'shfa17e83d, 32'shfa11a6a3, 32'shfa0b6517, 32'shfa05239a, 32'shf9fee22c, 32'shf9f8a0cd, 32'shf9f25f7d, 
               32'shf9ec1e3b, 32'shf9e5dd09, 32'shf9df9be6, 32'shf9d95ad1, 32'shf9d319cc, 32'shf9ccd8d6, 32'shf9c697f0, 32'shf9c05719, 
               32'shf9ba1651, 32'shf9b3d599, 32'shf9ad94f0, 32'shf9a75457, 32'shf9a113cd, 32'shf99ad354, 32'shf99492ea, 32'shf98e528f, 
               32'shf9881245, 32'shf981d20b, 32'shf97b91e1, 32'shf97551c6, 32'shf96f11bc, 32'shf968d1c3, 32'shf96291d9, 32'shf95c5200, 
               32'shf9561237, 32'shf94fd27f, 32'shf94992d7, 32'shf943533f, 32'shf93d13b8, 32'shf936d442, 32'shf93094dd, 32'shf92a5589, 
               32'shf9241645, 32'shf91dd712, 32'shf91797f0, 32'shf91158e0, 32'shf90b19e0, 32'shf904daf2, 32'shf8fe9c15, 32'shf8f85d49, 
               32'shf8f21e8e, 32'shf8ebdfe5, 32'shf8e5a14d, 32'shf8df62c7, 32'shf8d92452, 32'shf8d2e5f0, 32'shf8cca79e, 32'shf8c6695f, 
               32'shf8c02b31, 32'shf8b9ed15, 32'shf8b3af0c, 32'shf8ad7114, 32'shf8a7332e, 32'shf8a0f55b, 32'shf89ab799, 32'shf89479ea, 
               32'shf88e3c4d, 32'shf887fec3, 32'shf881c14b, 32'shf87b83e5, 32'shf8754692, 32'shf86f0952, 32'shf868cc24, 32'shf8628f09, 
               32'shf85c5201, 32'shf856150b, 32'shf84fd829, 32'shf8499b59, 32'shf8435e9d, 32'shf83d21f3, 32'shf836e55d, 32'shf830a8da, 
               32'shf82a6c6a, 32'shf824300e, 32'shf81df3c5, 32'shf817b78f, 32'shf8117b6d, 32'shf80b3f5f, 32'shf8050364, 32'shf7fec77d, 
               32'shf7f88ba9, 32'shf7f24fea, 32'shf7ec143e, 32'shf7e5d8a6, 32'shf7df9d22, 32'shf7d961b3, 32'shf7d32657, 32'shf7cceb0f, 
               32'shf7c6afdc, 32'shf7c074bd, 32'shf7ba39b3, 32'shf7b3febc, 32'shf7adc3db, 32'shf7a7890d, 32'shf7a14e55, 32'shf79b13b1, 
               32'shf794d922, 32'shf78e9ea7, 32'shf7886442, 32'shf78229f1, 32'shf77befb5, 32'shf775b58e, 32'shf76f7b7d, 32'shf7694180, 
               32'shf7630799, 32'shf75ccdc6, 32'shf756940a, 32'shf7505a62, 32'shf74a20d0, 32'shf743e754, 32'shf73daded, 32'shf737749b, 
               32'shf7313b60, 32'shf72b023a, 32'shf724c92a, 32'shf71e902f, 32'shf718574b, 32'shf7121e7c, 32'shf70be5c4, 32'shf705ad22, 
               32'shf6ff7496, 32'shf6f93c20, 32'shf6f303c0, 32'shf6eccb77, 32'shf6e69344, 32'shf6e05b27, 32'shf6da2321, 32'shf6d3eb32, 
               32'shf6cdb359, 32'shf6c77b97, 32'shf6c143ec, 32'shf6bb0c57, 32'shf6b4d4d9, 32'shf6ae9d73, 32'shf6a86623, 32'shf6a22eea, 
               32'shf69bf7c9, 32'shf695c0be, 32'shf68f89cb, 32'shf68952ef, 32'shf6831c2b, 32'shf67ce57e, 32'shf676aee8, 32'shf670786a, 
               32'shf66a4203, 32'shf6640bb4, 32'shf65dd57d, 32'shf6579f5e, 32'shf6516956, 32'shf64b3367, 32'shf644fd8f, 32'shf63ec7cf, 
               32'shf6389228, 32'shf6325c98, 32'shf62c2721, 32'shf625f1c2, 32'shf61fbc7b, 32'shf619874c, 32'shf6135237, 32'shf60d1d39, 
               32'shf606e854, 32'shf600b388, 32'shf5fa7ed4, 32'shf5f44a39, 32'shf5ee15b7, 32'shf5e7e14e, 32'shf5e1acfd, 32'shf5db78c6, 
               32'shf5d544a7, 32'shf5cf10a2, 32'shf5c8dcb6, 32'shf5c2a8e3, 32'shf5bc7529, 32'shf5b64189, 32'shf5b00e02, 32'shf5a9da94, 
               32'shf5a3a740, 32'shf59d7406, 32'shf59740e5, 32'shf5910dde, 32'shf58adaf0, 32'shf584a81d, 32'shf57e7563, 32'shf57842c3, 
               32'shf572103d, 32'shf56bddd1, 32'shf565ab80, 32'shf55f7948, 32'shf559472b, 32'shf5531528, 32'shf54ce33f, 32'shf546b171, 
               32'shf5407fbd, 32'shf53a4e24, 32'shf5341ca5, 32'shf52deb41, 32'shf527b9f7, 32'shf52188c9, 32'shf51b57b5, 32'shf51526bc, 
               32'shf50ef5de, 32'shf508c51b, 32'shf5029473, 32'shf4fc63e6, 32'shf4f63374, 32'shf4f0031e, 32'shf4e9d2e3, 32'shf4e3a2c3, 
               32'shf4dd72be, 32'shf4d742d6, 32'shf4d11308, 32'shf4cae356, 32'shf4c4b3c0, 32'shf4be8446, 32'shf4b854e7, 32'shf4b225a4, 
               32'shf4abf67e, 32'shf4a5c773, 32'shf49f9884, 32'shf49969b1, 32'shf4933afa, 32'shf48d0c5f, 32'shf486dde1, 32'shf480af7f, 
               32'shf47a8139, 32'shf4745310, 32'shf46e2504, 32'shf467f713, 32'shf461c940, 32'shf45b9b89, 32'shf4556def, 32'shf44f4071, 
               32'shf4491311, 32'shf442e5cd, 32'shf43cb8a7, 32'shf4368b9d, 32'shf4305eb0, 32'shf42a31e1, 32'shf424052f, 32'shf41dd89a, 
               32'shf417ac22, 32'shf4117fc8, 32'shf40b538b, 32'shf405276c, 32'shf3fefb6a, 32'shf3f8cf86, 32'shf3f2a3bf, 32'shf3ec7817, 
               32'shf3e64c8c, 32'shf3e0211f, 32'shf3d9f5cf, 32'shf3d3ca9e, 32'shf3cd9f8b, 32'shf3c77496, 32'shf3c149bf, 32'shf3bb1f07, 
               32'shf3b4f46c, 32'shf3aec9f0, 32'shf3a89f92, 32'shf3a27553, 32'shf39c4b32, 32'shf3962130, 32'shf38ff74d, 32'shf389cd88, 
               32'shf383a3e2, 32'shf37d7a5b, 32'shf37750f2, 32'shf37127a9, 32'shf36afe7e, 32'shf364d573, 32'shf35eac86, 32'shf35883b9, 
               32'shf3525b0b, 32'shf34c327c, 32'shf3460a0d, 32'shf33fe1bd, 32'shf339b98d, 32'shf333917c, 32'shf32d698a, 32'shf32741b9, 
               32'shf3211a07, 32'shf31af274, 32'shf314cb02, 32'shf30ea3af, 32'shf3087c7d, 32'shf302556a, 32'shf2fc2e77, 32'shf2f607a5, 
               32'shf2efe0f2, 32'shf2e9ba60, 32'shf2e393ef, 32'shf2dd6d9d, 32'shf2d7476c, 32'shf2d1215b, 32'shf2cafb6b, 32'shf2c4d59c, 
               32'shf2beafed, 32'shf2b88a5f, 32'shf2b264f2, 32'shf2ac3fa5, 32'shf2a61a7a, 32'shf29ff56f, 32'shf299d085, 32'shf293abbd, 
               32'shf28d8715, 32'shf287628f, 32'shf2813e2a, 32'shf27b19e6, 32'shf274f5c3, 32'shf26ed1c2, 32'shf268ade3, 32'shf2628a25, 
               32'shf25c6688, 32'shf256430e, 32'shf2501fb5, 32'shf249fc7d, 32'shf243d968, 32'shf23db674, 32'shf23793a3, 32'shf23170f3, 
               32'shf22b4e66, 32'shf2252bfa, 32'shf21f09b1, 32'shf218e78a, 32'shf212c585, 32'shf20ca3a3, 32'shf20681e3, 32'shf2006046, 
               32'shf1fa3ecb, 32'shf1f41d72, 32'shf1edfc3d, 32'shf1e7db2a, 32'shf1e1ba3a, 32'shf1db996d, 32'shf1d578c2, 32'shf1cf583b, 
               32'shf1c937d6, 32'shf1c31795, 32'shf1bcf777, 32'shf1b6d77c, 32'shf1b0b7a4, 32'shf1aa97ef, 32'shf1a4785e, 32'shf19e58f1, 
               32'shf19839a6, 32'shf1921a80, 32'shf18bfb7d, 32'shf185dc9d, 32'shf17fbde2, 32'shf1799f4a, 32'shf17380d6, 32'shf16d6286, 
               32'shf1674459, 32'shf1612651, 32'shf15b086d, 32'shf154eaad, 32'shf14ecd11, 32'shf148af9a, 32'shf1429247, 32'shf13c7518, 
               32'shf136580d, 32'shf1303b27, 32'shf12a1e66, 32'shf12401c9, 32'shf11de551, 32'shf117c8fe, 32'shf111accf, 32'shf10b90c5, 
               32'shf10574e0, 32'shf0ff5921, 32'shf0f93d86, 32'shf0f32210, 32'shf0ed06bf, 32'shf0e6eb94, 32'shf0e0d08d, 32'shf0dab5ad, 
               32'shf0d49af1, 32'shf0ce805b, 32'shf0c865ea, 32'shf0c24b9f, 32'shf0bc317a, 32'shf0b6177a, 32'shf0affda0, 32'shf0a9e3eb, 
               32'shf0a3ca5d, 32'shf09db0f4, 32'shf09797b2, 32'shf0917e95, 32'shf08b659f, 32'shf0854cce, 32'shf07f3424, 32'shf0791ba0, 
               32'shf0730342, 32'shf06ceb0b, 32'shf066d2fa, 32'shf060bb10, 32'shf05aa34c, 32'shf0548baf, 32'shf04e7438, 32'shf0485ce9, 
               32'shf04245c0, 32'shf03c2ebd, 32'shf03617e2, 32'shf030012e, 32'shf029eaa1, 32'shf023d43a, 32'shf01dbdfb, 32'shf017a7e3, 
               32'shf01191f3, 32'shf00b7c29, 32'shf0056687, 32'shefff510d, 32'sheff93bba, 32'sheff3268e, 32'shefed118a, 32'shefe6fcae, 
               32'shefe0e7f9, 32'shefdad36c, 32'shefd4bf08, 32'shefceaacb, 32'shefc896b5, 32'shefc282c8, 32'shefbc6f03, 32'shefb65b66, 
               32'shefb047f2, 32'shefaa34a5, 32'shefa42181, 32'shef9e0e85, 32'shef97fbb2, 32'shef91e907, 32'shef8bd685, 32'shef85c42b, 
               32'shef7fb1fa, 32'shef799ff2, 32'shef738e12, 32'shef6d7c5b, 32'shef676ace, 32'shef615969, 32'shef5b482d, 32'shef55371a, 
               32'shef4f2630, 32'shef491570, 32'shef4304d8, 32'shef3cf46a, 32'shef36e426, 32'shef30d40a, 32'shef2ac419, 32'shef24b451, 
               32'shef1ea4b2, 32'shef18953d, 32'shef1285f2, 32'shef0c76d0, 32'shef0667d9, 32'shef00590b, 32'sheefa4a67, 32'sheef43bed, 
               32'sheeee2d9d, 32'sheee81f78, 32'sheee2117c, 32'sheedc03ab, 32'sheed5f604, 32'sheecfe887, 32'sheec9db35, 32'sheec3ce0d, 
               32'sheebdc110, 32'sheeb7b43e, 32'sheeb1a796, 32'sheeab9b18, 32'sheea58ec6, 32'shee9f829e, 32'shee9976a1, 32'shee936acf, 
               32'shee8d5f29, 32'shee8753ad, 32'shee81485c, 32'shee7b3d36, 32'shee75323c, 32'shee6f276d, 32'shee691cc9, 32'shee631251, 
               32'shee5d0804, 32'shee56fde3, 32'shee50f3ed, 32'shee4aea23, 32'shee44e084, 32'shee3ed712, 32'shee38cdcb, 32'shee32c4b0, 
               32'shee2cbbc1, 32'shee26b2fe, 32'shee20aa67, 32'shee1aa1fc, 32'shee1499bd, 32'shee0e91aa, 32'shee0889c4, 32'shee02820a, 
               32'shedfc7a7c, 32'shedf6731b, 32'shedf06be6, 32'shedea64de, 32'shede45e03, 32'shedde5754, 32'shedd850d2, 32'shedd24a7d, 
               32'shedcc4454, 32'shedc63e59, 32'shedc0388a, 32'shedba32e9, 32'shedb42d74, 32'shedae282d, 32'sheda82313, 32'sheda21e26, 
               32'shed9c1967, 32'shed9614d5, 32'shed901070, 32'shed8a0c39, 32'shed84082f, 32'shed7e0453, 32'shed7800a5, 32'shed71fd24, 
               32'shed6bf9d1, 32'shed65f6ac, 32'shed5ff3b5, 32'shed59f0ec, 32'shed53ee51, 32'shed4debe4, 32'shed47e9a5, 32'shed41e794, 
               32'shed3be5b1, 32'shed35e3fd, 32'shed2fe277, 32'shed29e120, 32'shed23dff7, 32'shed1ddefd, 32'shed17de31, 32'shed11dd94, 
               32'shed0bdd25, 32'shed05dce5, 32'shecffdcd4, 32'shecf9dcf3, 32'shecf3dd3f, 32'shecedddbb, 32'shece7de66, 32'shece1df40, 
               32'shecdbe04a, 32'shecd5e182, 32'sheccfe2ea, 32'shecc9e481, 32'shecc3e648, 32'shecbde83e, 32'shecb7ea63, 32'shecb1ecb8, 
               32'shecabef3d, 32'sheca5f1f2, 32'shec9ff4d6, 32'shec99f7ea, 32'shec93fb2e, 32'shec8dfea1, 32'shec880245, 32'shec820619, 
               32'shec7c0a1d, 32'shec760e51, 32'shec7012b5, 32'shec6a1749, 32'shec641c0e, 32'shec5e2103, 32'shec582629, 32'shec522b7f, 
               32'shec4c3106, 32'shec4636bd, 32'shec403ca5, 32'shec3a42be, 32'shec344908, 32'shec2e4f82, 32'shec28562d, 32'shec225d09, 
               32'shec1c6417, 32'shec166b55, 32'shec1072c4, 32'shec0a7a65, 32'shec048237, 32'shebfe8a3a, 32'shebf8926f, 32'shebf29ad4, 
               32'shebeca36c, 32'shebe6ac35, 32'shebe0b52f, 32'shebdabe5c, 32'shebd4c7ba, 32'shebced149, 32'shebc8db0b, 32'shebc2e4fe, 
               32'shebbcef23, 32'shebb6f97b, 32'shebb10404, 32'shebab0ec0, 32'sheba519ad, 32'sheb9f24cd, 32'sheb99301f, 32'sheb933ba4, 
               32'sheb8d475b, 32'sheb875344, 32'sheb815f60, 32'sheb7b6bae, 32'sheb75782f, 32'sheb6f84e3, 32'sheb6991ca, 32'sheb639ee3, 
               32'sheb5dac2f, 32'sheb57b9ae, 32'sheb51c760, 32'sheb4bd545, 32'sheb45e35d, 32'sheb3ff1a8, 32'sheb3a0027, 32'sheb340ed9, 
               32'sheb2e1dbe, 32'sheb282cd6, 32'sheb223c22, 32'sheb1c4ba1, 32'sheb165b54, 32'sheb106b3a, 32'sheb0a7b54, 32'sheb048ba2, 
               32'sheafe9c24, 32'sheaf8acd9, 32'sheaf2bdc3, 32'sheaeccee0, 32'sheae6e031, 32'sheae0f1b6, 32'sheadb0370, 32'shead5155d, 
               32'sheacf277f, 32'sheac939d5, 32'sheac34c60, 32'sheabd5f1f, 32'sheab77212, 32'sheab1853a, 32'sheaab9896, 32'sheaa5ac27, 
               32'shea9fbfed, 32'shea99d3e8, 32'shea93e817, 32'shea8dfc7b, 32'shea881114, 32'shea8225e2, 32'shea7c3ae5, 32'shea76501d, 
               32'shea70658a, 32'shea6a7b2d, 32'shea649105, 32'shea5ea712, 32'shea58bd54, 32'shea52d3cc, 32'shea4cea79, 32'shea47015c, 
               32'shea411874, 32'shea3b2fc2, 32'shea354746, 32'shea2f5f00, 32'shea2976ef, 32'shea238f15, 32'shea1da770, 32'shea17c001, 
               32'shea11d8c8, 32'shea0bf1c6, 32'shea060af9, 32'shea002463, 32'she9fa3e03, 32'she9f457da, 32'she9ee71e6, 32'she9e88c2a, 
               32'she9e2a6a3, 32'she9dcc154, 32'she9d6dc3b, 32'she9d0f758, 32'she9cb12ad, 32'she9c52e38, 32'she9bf49fa, 32'she9b965f3, 
               32'she9b38223, 32'she9ad9e8a, 32'she9a7bb28, 32'she9a1d7fd, 32'she99bf509, 32'she996124d, 32'she9902fc7, 32'she98a4d7a, 
               32'she9846b63, 32'she97e8984, 32'she978a7dd, 32'she972c66d, 32'she96ce535, 32'she9670435, 32'she961236c, 32'she95b42db, 
               32'she9556282, 32'she94f8261, 32'she949a278, 32'she943c2c7, 32'she93de34e, 32'she938040d, 32'she9322505, 32'she92c4634, 
               32'she926679c, 32'she920893d, 32'she91aab16, 32'she914cd27, 32'she90eef71, 32'she90911f3, 32'she90334af, 32'she8fd57a2, 
               32'she8f77acf, 32'she8f19e34, 32'she8ebc1d3, 32'she8e5e5aa, 32'she8e009ba, 32'she8da2e04, 32'she8d45286, 32'she8ce7742, 
               32'she8c89c37, 32'she8c2c165, 32'she8bce6cd, 32'she8b70c6d, 32'she8b13248, 32'she8ab585c, 32'she8a57ea9, 32'she89fa530, 
               32'she899cbf1, 32'she893f2eb, 32'she88e1a20, 32'she888418e, 32'she8826936, 32'she87c9118, 32'she876b934, 32'she870e18a, 
               32'she86b0a1a, 32'she86532e4, 32'she85f5be9, 32'she8598528, 32'she853aea1, 32'she84dd855, 32'she8480243, 32'she8422c6c, 
               32'she83c56cf, 32'she836816d, 32'she830ac45, 32'she82ad759, 32'she82502a7, 32'she81f2e30, 32'she81959f4, 32'she81385f3, 
               32'she80db22d, 32'she807dea2, 32'she8020b52, 32'she7fc383d, 32'she7f66564, 32'she7f092c6, 32'she7eac063, 32'she7e4ee3c, 
               32'she7df1c50, 32'she7d94a9f, 32'she7d3792b, 32'she7cda7f2, 32'she7c7d6f4, 32'she7c20633, 32'she7bc35ad, 32'she7b66563, 
               32'she7b09555, 32'she7aac583, 32'she7a4f5ed, 32'she79f2693, 32'she7995776, 32'she7938894, 32'she78db9ef, 32'she787eb86, 
               32'she7821d59, 32'she77c4f69, 32'she77681b6, 32'she770b43e, 32'she76ae704, 32'she7651a06, 32'she75f4d45, 32'she75980c1, 
               32'she753b479, 32'she74de86f, 32'she7481ca1, 32'she7425110, 32'she73c85bc, 32'she736baa6, 32'she730efcc, 32'she72b2530, 
               32'she7255ad1, 32'she71f90b0, 32'she719c6cb, 32'she713fd25, 32'she70e33bb, 32'she7086a8f, 32'she702a1a1, 32'she6fcd8f1, 
               32'she6f7107e, 32'she6f14849, 32'she6eb8052, 32'she6e5b899, 32'she6dff11d, 32'she6da29e0, 32'she6d462e1, 32'she6ce9c1f, 
               32'she6c8d59c, 32'she6c30f57, 32'she6bd4951, 32'she6b78389, 32'she6b1bdff, 32'she6abf8b3, 32'she6a633a6, 32'she6a06ed8, 
               32'she69aaa48, 32'she694e5f7, 32'she68f21e5, 32'she6895e11, 32'she6839a7c, 32'she67dd727, 32'she6781410, 32'she6725138, 
               32'she66c8e9f, 32'she666cc45, 32'she6610a2a, 32'she65b484f, 32'she65586b3, 32'she64fc556, 32'she64a0438, 32'she644435a, 
               32'she63e82bc, 32'she638c25d, 32'she633023e, 32'she62d425e, 32'she62782be, 32'she621c35e, 32'she61c043d, 32'she616455d, 
               32'she61086bc, 32'she60ac85c, 32'she6050a3b, 32'she5ff4c5b, 32'she5f98ebb, 32'she5f3d15b, 32'she5ee143b, 32'she5e8575b, 
               32'she5e29abc, 32'she5dcde5e, 32'she5d72240, 32'she5d16662, 32'she5cbaac5, 32'she5c5ef69, 32'she5c0344d, 32'she5ba7972, 
               32'she5b4bed8, 32'she5af047f, 32'she5a94a67, 32'she5a39090, 32'she59dd6f9, 32'she5981da4, 32'she5926490, 32'she58cabbe, 
               32'she586f32c, 32'she5813adc, 32'she57b82cd, 32'she575cb00, 32'she5701374, 32'she56a5c2a, 32'she564a521, 32'she55eee5a, 
               32'she55937d5, 32'she5538191, 32'she54dcb8f, 32'she54815cf, 32'she5426051, 32'she53cab15, 32'she536f61b, 32'she5314163, 
               32'she52b8cee, 32'she525d8ba, 32'she52024c9, 32'she51a711a, 32'she514bdad, 32'she50f0a83, 32'she509579b, 32'she503a4f6, 
               32'she4fdf294, 32'she4f84074, 32'she4f28e96, 32'she4ecdcfc, 32'she4e72ba4, 32'she4e17a8f, 32'she4dbc9bd, 32'she4d6192e, 
               32'she4d068e2, 32'she4cab8d9, 32'she4c50914, 32'she4bf5991, 32'she4b9aa52, 32'she4b3fb56, 32'she4ae4c9d, 32'she4a89e28, 
               32'she4a2eff6, 32'she49d4208, 32'she497945d, 32'she491e6f6, 32'she48c39d3, 32'she4868cf3, 32'she480e057, 32'she47b33ff, 
               32'she47587eb, 32'she46fdc1b, 32'she46a308f, 32'she4648547, 32'she45eda43, 32'she4592f83, 32'she4538507, 32'she44ddad0, 
               32'she44830dd, 32'she442872e, 32'she43cddc4, 32'she437349f, 32'she4318bbe, 32'she42be321, 32'she4263ac9, 32'she42092b6, 
               32'she41aeae8, 32'she415435f, 32'she40f9c1a, 32'she409f51a, 32'she4044e60, 32'she3fea7ea, 32'she3f901ba, 32'she3f35bce, 
               32'she3edb628, 32'she3e810c7, 32'she3e26bac, 32'she3dcc6d5, 32'she3d72245, 32'she3d17df9, 32'she3cbd9f4, 32'she3c63633, 
               32'she3c092b9, 32'she3baef84, 32'she3b54c95, 32'she3afa9ec, 32'she3aa0788, 32'she3a4656b, 32'she39ec393, 32'she3992202, 
               32'she39380b6, 32'she38ddfb1, 32'she3883ef2, 32'she3829e79, 32'she37cfe47, 32'she3775e5a, 32'she371beb5, 32'she36c1f55, 
               32'she366803c, 32'she360e16a, 32'she35b42df, 32'she355a49a, 32'she350069b, 32'she34a68e4, 32'she344cb73, 32'she33f2e4a, 
               32'she3399167, 32'she333f4cb, 32'she32e5876, 32'she328bc69, 32'she32320a2, 32'she31d8523, 32'she317e9eb, 32'she3124efa, 
               32'she30cb451, 32'she30719ef, 32'she3017fd5, 32'she2fbe602, 32'she2f64c77, 32'she2f0b333, 32'she2eb1a37, 32'she2e58183, 
               32'she2dfe917, 32'she2da50f3, 32'she2d4b916, 32'she2cf2182, 32'she2c98a35, 32'she2c3f331, 32'she2be5c74, 32'she2b8c600, 
               32'she2b32fd4, 32'she2ad99f1, 32'she2a80456, 32'she2a26f03, 32'she29cd9f8, 32'she2974536, 32'she291b0bd, 32'she28c1c8c, 
               32'she28688a4, 32'she280f505, 32'she27b61af, 32'she275cea1, 32'she2703bdc, 32'she26aa960, 32'she265172e, 32'she25f8544, 
               32'she259f3a3, 32'she254624b, 32'she24ed13d, 32'she2494078, 32'she243affc, 32'she23e1fca, 32'she2388fe1, 32'she2330041, 
               32'she22d70eb, 32'she227e1df, 32'she222531c, 32'she21cc4a3, 32'she2173674, 32'she211a88f, 32'she20c1af3, 32'she2068da1, 
               32'she2010099, 32'she1fb73dc, 32'she1f5e768, 32'she1f05b3e, 32'she1eacf5f, 32'she1e543ca, 32'she1dfb87f, 32'she1da2d7e, 
               32'she1d4a2c8, 32'she1cf185c, 32'she1c98e3b, 32'she1c40464, 32'she1be7ad8, 32'she1b8f197, 32'she1b368a0, 32'she1addff4, 
               32'she1a85793, 32'she1a2cf7c, 32'she19d47b1, 32'she197c031, 32'she19238fb, 32'she18cb211, 32'she1872b72, 32'she181a51e, 
               32'she17c1f15, 32'she1769958, 32'she17113e5, 32'she16b8ebf, 32'she16609e3, 32'she1608554, 32'she15b0110, 32'she1557d17, 
               32'she14ff96a, 32'she14a7609, 32'she144f2f3, 32'she13f702a, 32'she139edac, 32'she1346b7a, 32'she12ee995, 32'she12967fb, 
               32'she123e6ad, 32'she11e65ac, 32'she118e4f6, 32'she113648d, 32'she10de470, 32'she10864a0, 32'she102e51c, 32'she0fd65e4, 
               32'she0f7e6f9, 32'she0f2685b, 32'she0ecea09, 32'she0e76c04, 32'she0e1ee4b, 32'she0dc70e0, 32'she0d6f3c1, 32'she0d176ef, 
               32'she0cbfa6a, 32'she0c67e32, 32'she0c10247, 32'she0bb86a9, 32'she0b60b58, 32'she0b09055, 32'she0ab159e, 32'she0a59b35, 
               32'she0a0211a, 32'she09aa74b, 32'she0952dcb, 32'she08fb497, 32'she08a3bb2, 32'she084c31a, 32'she07f4acf, 32'she079d2d3, 
               32'she0745b24, 32'she06ee3c3, 32'she0696cb0, 32'she063f5eb, 32'she05e7f74, 32'she059094a, 32'she053936f, 32'she04e1de3, 
               32'she048a8a4, 32'she04333b3, 32'she03dbf11, 32'she0384abe, 32'she032d6b8, 32'she02d6301, 32'she027ef99, 32'she0227c7f, 
               32'she01d09b4, 32'she0179738, 32'she012250a, 32'she00cb32b, 32'she007419b, 32'she001d05a, 32'shdffc5f67, 32'shdff6eec4, 
               32'shdff17e70, 32'shdfec0e6a, 32'shdfe69eb4, 32'shdfe12f4e, 32'shdfdbc036, 32'shdfd6516e, 32'shdfd0e2f5, 32'shdfcb74cb, 
               32'shdfc606f1, 32'shdfc09967, 32'shdfbb2c2c, 32'shdfb5bf41, 32'shdfb052a5, 32'shdfaae659, 32'shdfa57a5d, 32'shdfa00eb1, 
               32'shdf9aa354, 32'shdf953848, 32'shdf8fcd8b, 32'shdf8a631f, 32'shdf84f902, 32'shdf7f8f36, 32'shdf7a25ba, 32'shdf74bc8e, 
               32'shdf6f53b3, 32'shdf69eb27, 32'shdf6482ed, 32'shdf5f1b02, 32'shdf59b369, 32'shdf544c1f, 32'shdf4ee527, 32'shdf497e7f, 
               32'shdf441828, 32'shdf3eb221, 32'shdf394c6b, 32'shdf33e707, 32'shdf2e81f3, 32'shdf291d30, 32'shdf23b8be, 32'shdf1e549d, 
               32'shdf18f0ce, 32'shdf138d4f, 32'shdf0e2a22, 32'shdf08c746, 32'shdf0364bc, 32'shdefe0282, 32'shdef8a09b, 32'shdef33f04, 
               32'shdeedddc0, 32'shdee87ccc, 32'shdee31c2b, 32'shdeddbbdb, 32'shded85bdd, 32'shded2fc31, 32'shdecd9cd7, 32'shdec83dce, 
               32'shdec2df18, 32'shdebd80b3, 32'shdeb822a1, 32'shdeb2c4e1, 32'shdead6773, 32'shdea80a57, 32'shdea2ad8d, 32'shde9d5116, 
               32'shde97f4f1, 32'shde92991e, 32'shde8d3d9e, 32'shde87e271, 32'shde828796, 32'shde7d2d0e, 32'shde77d2d8, 32'shde7278f5, 
               32'shde6d1f65, 32'shde67c628, 32'shde626d3e, 32'shde5d14a6, 32'shde57bc62, 32'shde526471, 32'shde4d0cd2, 32'shde47b587, 
               32'shde425e8f, 32'shde3d07eb, 32'shde37b199, 32'shde325b9b, 32'shde2d05f1, 32'shde27b09a, 32'shde225b96, 32'shde1d06e6, 
               32'shde17b28a, 32'shde125e81, 32'shde0d0acc, 32'shde07b76b, 32'shde02645d, 32'shddfd11a3, 32'shddf7bf3e, 32'shddf26d2c, 
               32'shdded1b6e, 32'shdde7ca05, 32'shdde278ef, 32'shdddd282e, 32'shddd7d7c1, 32'shddd287a8, 32'shddcd37e4, 32'shddc7e873, 
               32'shddc29958, 32'shddbd4a91, 32'shddb7fc1e, 32'shddb2ae00, 32'shddad6036, 32'shdda812c2, 32'shdda2c5a2, 32'shdd9d78d7, 
               32'shdd982c60, 32'shdd92e03f, 32'shdd8d9472, 32'shdd8848fb, 32'shdd82fdd8, 32'shdd7db30b, 32'shdd786892, 32'shdd731e6f, 
               32'shdd6dd4a2, 32'shdd688b29, 32'shdd634206, 32'shdd5df938, 32'shdd58b0c0, 32'shdd53689d, 32'shdd4e20d0, 32'shdd48d958, 
               32'shdd439236, 32'shdd3e4b6a, 32'shdd3904f4, 32'shdd33bed3, 32'shdd2e7908, 32'shdd293393, 32'shdd23ee74, 32'shdd1ea9ab, 
               32'shdd196538, 32'shdd14211b, 32'shdd0edd55, 32'shdd0999e4, 32'shdd0456ca, 32'shdcff1407, 32'shdcf9d199, 32'shdcf48f82, 
               32'shdcef4dc2, 32'shdcea0c58, 32'shdce4cb44, 32'shdcdf8a87, 32'shdcda4a21, 32'shdcd50a12, 32'shdccfca59, 32'shdcca8af7, 
               32'shdcc54bec, 32'shdcc00d38, 32'shdcbacedb, 32'shdcb590d5, 32'shdcb05326, 32'shdcab15ce, 32'shdca5d8cd, 32'shdca09c24, 
               32'shdc9b5fd2, 32'shdc9623d7, 32'shdc90e834, 32'shdc8bace8, 32'shdc8671f3, 32'shdc813756, 32'shdc7bfd11, 32'shdc76c323, 
               32'shdc71898d, 32'shdc6c504e, 32'shdc671768, 32'shdc61ded9, 32'shdc5ca6a2, 32'shdc576ec3, 32'shdc52373c, 32'shdc4d000d, 
               32'shdc47c936, 32'shdc4292b8, 32'shdc3d5c91, 32'shdc3826c3, 32'shdc32f14d, 32'shdc2dbc2f, 32'shdc28876a, 32'shdc2352fd, 
               32'shdc1e1ee9, 32'shdc18eb2d, 32'shdc13b7c9, 32'shdc0e84bf, 32'shdc09520d, 32'shdc041fb4, 32'shdbfeedb3, 32'shdbf9bc0c, 
               32'shdbf48abd, 32'shdbef59c7, 32'shdbea292b, 32'shdbe4f8e7, 32'shdbdfc8fc, 32'shdbda996b, 32'shdbd56a32, 32'shdbd03b53, 
               32'shdbcb0cce, 32'shdbc5dea1, 32'shdbc0b0ce, 32'shdbbb8354, 32'shdbb65634, 32'shdbb1296e, 32'shdbabfd01, 32'shdba6d0ed, 
               32'shdba1a534, 32'shdb9c79d4, 32'shdb974ece, 32'shdb922421, 32'shdb8cf9cf, 32'shdb87cfd6, 32'shdb82a638, 32'shdb7d7cf3, 
               32'shdb785409, 32'shdb732b79, 32'shdb6e0342, 32'shdb68db67, 32'shdb63b3e5, 32'shdb5e8cbe, 32'shdb5965f1, 32'shdb543f7e, 
               32'shdb4f1967, 32'shdb49f3a9, 32'shdb44ce46, 32'shdb3fa93e, 32'shdb3a8491, 32'shdb35603e, 32'shdb303c46, 32'shdb2b18a9, 
               32'shdb25f566, 32'shdb20d27f, 32'shdb1baff2, 32'shdb168dc1, 32'shdb116beb, 32'shdb0c4a70, 32'shdb072950, 32'shdb02088b, 
               32'shdafce821, 32'shdaf7c813, 32'shdaf2a860, 32'shdaed8909, 32'shdae86a0d, 32'shdae34b6d, 32'shdade2d28, 32'shdad90f3f, 
               32'shdad3f1b1, 32'shdaced47f, 32'shdac9b7a9, 32'shdac49b2f, 32'shdabf7f11, 32'shdaba634e, 32'shdab547e8, 32'shdab02cdd, 
               32'shdaab122f, 32'shdaa5f7dd, 32'shdaa0dde7, 32'shda9bc44d, 32'shda96ab0f, 32'shda91922e, 32'shda8c79a9, 32'shda876180, 
               32'shda8249b4, 32'shda7d3244, 32'shda781b31, 32'shda73047b, 32'shda6dee21, 32'shda68d824, 32'shda63c284, 32'shda5ead40, 
               32'shda599859, 32'shda5483d0, 32'shda4f6fa3, 32'shda4a5bd3, 32'shda454860, 32'shda40354a, 32'shda3b2292, 32'shda361036, 
               32'shda30fe38, 32'shda2bec97, 32'shda26db54, 32'shda21ca6e, 32'shda1cb9e5, 32'shda17a9ba, 32'shda1299ec, 32'shda0d8a7c, 
               32'shda087b69, 32'shda036cb5, 32'shd9fe5e5e, 32'shd9f95064, 32'shd9f442c9, 32'shd9ef358b, 32'shd9ea28ac, 32'shd9e51c2a, 
               32'shd9e01006, 32'shd9db0441, 32'shd9d5f8d9, 32'shd9d0edd0, 32'shd9cbe325, 32'shd9c6d8d8, 32'shd9c1cee9, 32'shd9bcc559, 
               32'shd9b7bc27, 32'shd9b2b354, 32'shd9adaadf, 32'shd9a8a2c9, 32'shd9a39b11, 32'shd99e93b8, 32'shd9998cbe, 32'shd9948623, 
               32'shd98f7fe6, 32'shd98a7a08, 32'shd9857489, 32'shd9806f69, 32'shd97b6aa8, 32'shd9766646, 32'shd9716243, 32'shd96c5e9f, 
               32'shd9675b5a, 32'shd9625875, 32'shd95d55ef, 32'shd95853c8, 32'shd9535201, 32'shd94e5099, 32'shd9494f90, 32'shd9444ee7, 
               32'shd93f4e9e, 32'shd93a4eb4, 32'shd9354f2a, 32'shd9305000, 32'shd92b5135, 32'shd92652ca, 32'shd92154bf, 32'shd91c5714, 
               32'shd91759c9, 32'shd9125cde, 32'shd90d6053, 32'shd9086428, 32'shd903685d, 32'shd8fe6cf2, 32'shd8f971e8, 32'shd8f4773e, 
               32'shd8ef7cf4, 32'shd8ea830b, 32'shd8e58982, 32'shd8e0905a, 32'shd8db9792, 32'shd8d69f2a, 32'shd8d1a724, 32'shd8ccaf7e, 
               32'shd8c7b838, 32'shd8c2c154, 32'shd8bdcad0, 32'shd8b8d4ad, 32'shd8b3deeb, 32'shd8aee98a, 32'shd8a9f48a, 32'shd8a4ffec, 
               32'shd8a00bae, 32'shd89b17d1, 32'shd8962456, 32'shd891313b, 32'shd88c3e83, 32'shd8874c2b, 32'shd8825a35, 32'shd87d68a0, 
               32'shd878776d, 32'shd873869b, 32'shd86e962b, 32'shd869a61d, 32'shd864b670, 32'shd85fc725, 32'shd85ad83c, 32'shd855e9b4, 
               32'shd850fb8e, 32'shd84c0dcb, 32'shd8472069, 32'shd8423369, 32'shd83d46cc, 32'shd8385a90, 32'shd8336eb7, 32'shd82e833f, 
               32'shd829982b, 32'shd824ad78, 32'shd81fc328, 32'shd81ad93a, 32'shd815efae, 32'shd8110685, 32'shd80c1dbf, 32'shd807355b, 
               32'shd8024d59, 32'shd7fd65bb, 32'shd7f87e7f, 32'shd7f397a6, 32'shd7eeb130, 32'shd7e9cb1c, 32'shd7e4e56c, 32'shd7e0001e, 
               32'shd7db1b34, 32'shd7d636ac, 32'shd7d15288, 32'shd7cc6ec6, 32'shd7c78b68, 32'shd7c2a86d, 32'shd7bdc5d6, 32'shd7b8e3a2, 
               32'shd7b401d1, 32'shd7af2063, 32'shd7aa3f5a, 32'shd7a55eb3, 32'shd7a07e70, 32'shd79b9e91, 32'shd796bf16, 32'shd791dffe, 
               32'shd78d014a, 32'shd78822f9, 32'shd783450d, 32'shd77e6784, 32'shd7798a60, 32'shd774ad9f, 32'shd76fd143, 32'shd76af54a, 
               32'shd76619b6, 32'shd7613e86, 32'shd75c63ba, 32'shd7578952, 32'shd752af4f, 32'shd74dd5b0, 32'shd748fc75, 32'shd744239f, 
               32'shd73f4b2e, 32'shd73a7321, 32'shd7359b78, 32'shd730c434, 32'shd72bed55, 32'shd72716db, 32'shd72240c5, 32'shd71d6b15, 
               32'shd71895c9, 32'shd713c0e2, 32'shd70eec60, 32'shd70a1843, 32'shd705448b, 32'shd7007138, 32'shd6fb9e4b, 32'shd6f6cbc2, 
               32'shd6f1f99f, 32'shd6ed27e1, 32'shd6e85689, 32'shd6e38596, 32'shd6deb508, 32'shd6d9e4e0, 32'shd6d5151d, 32'shd6d045c0, 
               32'shd6cb76c9, 32'shd6c6a837, 32'shd6c1da0b, 32'shd6bd0c45, 32'shd6b83ee4, 32'shd6b371ea, 32'shd6aea555, 32'shd6a9d926, 
               32'shd6a50d5d, 32'shd6a041fa, 32'shd69b76fe, 32'shd696ac67, 32'shd691e237, 32'shd68d186d, 32'shd6884f09, 32'shd683860b, 
               32'shd67ebd74, 32'shd679f543, 32'shd6752d79, 32'shd6706615, 32'shd66b9f18, 32'shd666d881, 32'shd6621251, 32'shd65d4c88, 
               32'shd6588725, 32'shd653c229, 32'shd64efd94, 32'shd64a3966, 32'shd645759f, 32'shd640b23f, 32'shd63bef46, 32'shd6372cb3, 
               32'shd6326a88, 32'shd62da8c4, 32'shd628e767, 32'shd6242672, 32'shd61f65e4, 32'shd61aa5bd, 32'shd615e5fd, 32'shd61126a5, 
               32'shd60c67b4, 32'shd607a92b, 32'shd602eb0a, 32'shd5fe2d50, 32'shd5f96ffd, 32'shd5f4b313, 32'shd5eff690, 32'shd5eb3a75, 
               32'shd5e67ec1, 32'shd5e1c376, 32'shd5dd0892, 32'shd5d84e17, 32'shd5d39403, 32'shd5ceda58, 32'shd5ca2115, 32'shd5c56839, 
               32'shd5c0afc6, 32'shd5bbf7bc, 32'shd5b74019, 32'shd5b288df, 32'shd5add20d, 32'shd5a91ba4, 32'shd5a465a3, 32'shd59fb00b, 
               32'shd59afadb, 32'shd5964614, 32'shd59191b5, 32'shd58cddbf, 32'shd5882a32, 32'shd583770e, 32'shd57ec452, 32'shd57a1200, 
               32'shd5756016, 32'shd570ae95, 32'shd56bfd7d, 32'shd5674ccf, 32'shd5629c89, 32'shd55decad, 32'shd5593d3a, 32'shd5548e30, 
               32'shd54fdf8f, 32'shd54b3157, 32'shd5468389, 32'shd541d625, 32'shd53d292a, 32'shd5387c98, 32'shd533d070, 32'shd52f24b2, 
               32'shd52a795d, 32'shd525ce72, 32'shd52123f0, 32'shd51c79d9, 32'shd517d02b, 32'shd51326e7, 32'shd50e7e0d, 32'shd509d59d, 
               32'shd5052d97, 32'shd50085fb, 32'shd4fbdec9, 32'shd4f73801, 32'shd4f291a4, 32'shd4edebb0, 32'shd4e94627, 32'shd4e4a108, 
               32'shd4dffc54, 32'shd4db580a, 32'shd4d6b42b, 32'shd4d210b5, 32'shd4cd6dab, 32'shd4c8cb0b, 32'shd4c428d6, 32'shd4bf870b, 
               32'shd4bae5ab, 32'shd4b644b6, 32'shd4b1a42c, 32'shd4ad040c, 32'shd4a86458, 32'shd4a3c50e, 32'shd49f2630, 32'shd49a87bc, 
               32'shd495e9b3, 32'shd4914c16, 32'shd48caee4, 32'shd488121d, 32'shd48375c1, 32'shd47ed9d0, 32'shd47a3e4b, 32'shd475a332, 
               32'shd4710883, 32'shd46c6e40, 32'shd467d469, 32'shd4633afd, 32'shd45ea1fd, 32'shd45a0969, 32'shd4557140, 32'shd450d983, 
               32'shd44c4232, 32'shd447ab4c, 32'shd44314d3, 32'shd43e7ec5, 32'shd439e923, 32'shd43553ee, 32'shd430bf24, 32'shd42c2ac6, 
               32'shd42796d5, 32'shd4230350, 32'shd41e7037, 32'shd419dd8a, 32'shd4154b4a, 32'shd410b976, 32'shd40c280e, 32'shd4079713, 
               32'shd4030684, 32'shd3fe7662, 32'shd3f9e6ad, 32'shd3f55764, 32'shd3f0c887, 32'shd3ec3a18, 32'shd3e7ac15, 32'shd3e31e7f, 
               32'shd3de9156, 32'shd3da049a, 32'shd3d5784a, 32'shd3d0ec68, 32'shd3cc60f2, 32'shd3c7d5ea, 32'shd3c34b4f, 32'shd3bec121, 
               32'shd3ba3760, 32'shd3b5ae0d, 32'shd3b12526, 32'shd3ac9cad, 32'shd3a814a2, 32'shd3a38d03, 32'shd39f05d3, 32'shd39a7f0f, 
               32'shd395f8ba, 32'shd39172d2, 32'shd38ced57, 32'shd388684a, 32'shd383e3ab, 32'shd37f5f7a, 32'shd37adbb6, 32'shd3765861, 
               32'shd371d579, 32'shd36d52ff, 32'shd368d0f3, 32'shd3644f55, 32'shd35fce26, 32'shd35b4d64, 32'shd356cd11, 32'shd3524d2b, 
               32'shd34dcdb4, 32'shd3494eab, 32'shd344d011, 32'shd34051e5, 32'shd33bd427, 32'shd33756d8, 32'shd332d9f7, 32'shd32e5d85, 
               32'shd329e181, 32'shd32565ec, 32'shd320eac6, 32'shd31c700f, 32'shd317f5c6, 32'shd3137bec, 32'shd30f0280, 32'shd30a8984, 
               32'shd30610f7, 32'shd30198d8, 32'shd2fd2129, 32'shd2f8a9e9, 32'shd2f43318, 32'shd2efbcb6, 32'shd2eb46c3, 32'shd2e6d13f, 
               32'shd2e25c2b, 32'shd2dde786, 32'shd2d97350, 32'shd2d4ff8a, 32'shd2d08c33, 32'shd2cc194c, 32'shd2c7a6d4, 32'shd2c334cc, 
               32'shd2bec333, 32'shd2ba520a, 32'shd2b5e151, 32'shd2b17107, 32'shd2ad012e, 32'shd2a891c4, 32'shd2a422ca, 32'shd29fb440, 
               32'shd29b4626, 32'shd296d87c, 32'shd2926b41, 32'shd28dfe77, 32'shd289921e, 32'shd2852634, 32'shd280babb, 32'shd27c4fb1, 
               32'shd277e518, 32'shd2737af0, 32'shd26f1138, 32'shd26aa7f0, 32'shd2663f19, 32'shd261d6b2, 32'shd25d6ebc, 32'shd2590736, 
               32'shd254a021, 32'shd250397d, 32'shd24bd34a, 32'shd2476d87, 32'shd2430835, 32'shd23ea354, 32'shd23a3ee4, 32'shd235dae4, 
               32'shd2317756, 32'shd22d1439, 32'shd228b18d, 32'shd2244f52, 32'shd21fed88, 32'shd21b8c2f, 32'shd2172b48, 32'shd212cad1, 
               32'shd20e6acc, 32'shd20a0b39, 32'shd205ac17, 32'shd2014d66, 32'shd1fcef27, 32'shd1f89159, 32'shd1f433fd, 32'shd1efd713, 
               32'shd1eb7a9a, 32'shd1e71e93, 32'shd1e2c2fd, 32'shd1de67da, 32'shd1da0d28, 32'shd1d5b2e8, 32'shd1d1591a, 32'shd1ccffbe, 
               32'shd1c8a6d4, 32'shd1c44e5c, 32'shd1bff656, 32'shd1bb9ec2, 32'shd1b747a0, 32'shd1b2f0f1, 32'shd1ae9ab4, 32'shd1aa44e9, 
               32'shd1a5ef90, 32'shd1a19aaa, 32'shd19d4636, 32'shd198f235, 32'shd1949ea6, 32'shd1904b89, 32'shd18bf8e0, 32'shd187a6a8, 
               32'shd18354e4, 32'shd17f0392, 32'shd17ab2b3, 32'shd1766247, 32'shd172124d, 32'shd16dc2c7, 32'shd16973b3, 32'shd1652512, 
               32'shd160d6e5, 32'shd15c892a, 32'shd1583be2, 32'shd153ef0e, 32'shd14fa2ad, 32'shd14b56be, 32'shd1470b44, 32'shd142c03c, 
               32'shd13e75a8, 32'shd13a2b87, 32'shd135e1d9, 32'shd131989f, 32'shd12d4fd9, 32'shd1290786, 32'shd124bfa6, 32'shd120783a, 
               32'shd11c3142, 32'shd117eabd, 32'shd113a4ad, 32'shd10f5f10, 32'shd10b19e7, 32'shd106d531, 32'shd10290f0, 32'shd0fe4d22, 
               32'shd0fa09c9, 32'shd0f5c6e3, 32'shd0f18472, 32'shd0ed4275, 32'shd0e900ec, 32'shd0e4bfd7, 32'shd0e07f36, 32'shd0dc3f0a, 
               32'shd0d7ff51, 32'shd0d3c00e, 32'shd0cf813e, 32'shd0cb42e3, 32'shd0c704fd, 32'shd0c2c78b, 32'shd0be8a8d, 32'shd0ba4e05, 
               32'shd0b611f1, 32'shd0b1d651, 32'shd0ad9b26, 32'shd0a96070, 32'shd0a5262f, 32'shd0a0ec63, 32'shd09cb30b, 32'shd0987a29, 
               32'shd09441bb, 32'shd09009c3, 32'shd08bd23f, 32'shd0879b31, 32'shd0836497, 32'shd07f2e73, 32'shd07af8c4, 32'shd076c38b, 
               32'shd0728ec6, 32'shd06e5a77, 32'shd06a269d, 32'shd065f339, 32'shd061c04a, 32'shd05d8dd1, 32'shd0595bcd, 32'shd0552a3f, 
               32'shd050f926, 32'shd04cc884, 32'shd0489856, 32'shd044689f, 32'shd040395d, 32'shd03c0a91, 32'shd037dc3b, 32'shd033ae5b, 
               32'shd02f80f1, 32'shd02b53fc, 32'shd027277e, 32'shd022fb76, 32'shd01ecfe4, 32'shd01aa4c8, 32'shd0167a22, 32'shd0124ff3, 
               32'shd00e2639, 32'shd009fcf6, 32'shd005d42a, 32'shd001abd3, 32'shcffd83f4, 32'shcff95c8a, 32'shcff53597, 32'shcff10f1b, 
               32'shcfece915, 32'shcfe8c386, 32'shcfe49e6d, 32'shcfe079cc, 32'shcfdc55a1, 32'shcfd831ec, 32'shcfd40eaf, 32'shcfcfebe8, 
               32'shcfcbc999, 32'shcfc7a7c0, 32'shcfc3865e, 32'shcfbf6573, 32'shcfbb4500, 32'shcfb72503, 32'shcfb3057d, 32'shcfaee66f, 
               32'shcfaac7d8, 32'shcfa6a9b8, 32'shcfa28c10, 32'shcf9e6edf, 32'shcf9a5225, 32'shcf9635e2, 32'shcf921a17, 32'shcf8dfec4, 
               32'shcf89e3e8, 32'shcf85c984, 32'shcf81af97, 32'shcf7d9622, 32'shcf797d24, 32'shcf75649f, 32'shcf714c91, 32'shcf6d34fb, 
               32'shcf691ddd, 32'shcf650736, 32'shcf60f108, 32'shcf5cdb51, 32'shcf58c613, 32'shcf54b14d, 32'shcf509cfe, 32'shcf4c8928, 
               32'shcf4875ca, 32'shcf4462e4, 32'shcf405077, 32'shcf3c3e82, 32'shcf382d05, 32'shcf341c00, 32'shcf300b74, 32'shcf2bfb60, 
               32'shcf27ebc5, 32'shcf23dca2, 32'shcf1fcdf8, 32'shcf1bbfc6, 32'shcf17b20d, 32'shcf13a4cd, 32'shcf0f9805, 32'shcf0b8bb7, 
               32'shcf077fe1, 32'shcf037483, 32'shceff699f, 32'shcefb5f34, 32'shcef75541, 32'shcef34bc8, 32'shceef42c7, 32'shceeb3a40, 
               32'shcee73231, 32'shcee32a9c, 32'shcedf2380, 32'shcedb1cde, 32'shced716b4, 32'shced31104, 32'shcecf0bcd, 32'shcecb070f, 
               32'shcec702cb, 32'shcec2ff01, 32'shcebefbb0, 32'shcebaf8d8, 32'shceb6f67a, 32'shceb2f496, 32'shceaef32b, 32'shceaaf23a, 
               32'shcea6f1c2, 32'shcea2f1c5, 32'shce9ef241, 32'shce9af337, 32'shce96f4a7, 32'shce92f691, 32'shce8ef8f4, 32'shce8afbd2, 
               32'shce86ff2a, 32'shce8302fc, 32'shce7f0748, 32'shce7b0c0e, 32'shce77114e, 32'shce731709, 32'shce6f1d3d, 32'shce6b23ec, 
               32'shce672b16, 32'shce6332ba, 32'shce5f3ad8, 32'shce5b4370, 32'shce574c84, 32'shce535611, 32'shce4f6019, 32'shce4b6a9c, 
               32'shce47759a, 32'shce438112, 32'shce3f8d05, 32'shce3b9973, 32'shce37a65b, 32'shce33b3be, 32'shce2fc19c, 32'shce2bcff5, 
               32'shce27dec9, 32'shce23ee18, 32'shce1ffde2, 32'shce1c0e28, 32'shce181ee8, 32'shce143023, 32'shce1041d9, 32'shce0c540b, 
               32'shce0866b8, 32'shce0479e0, 32'shce008d84, 32'shcdfca1a3, 32'shcdf8b63d, 32'shcdf4cb53, 32'shcdf0e0e4, 32'shcdecf6f1, 
               32'shcde90d79, 32'shcde5247d, 32'shcde13bfd, 32'shcddd53f8, 32'shcdd96c6f, 32'shcdd58562, 32'shcdd19ed0, 32'shcdcdb8ba, 
               32'shcdc9d320, 32'shcdc5ee02, 32'shcdc20960, 32'shcdbe253a, 32'shcdba4190, 32'shcdb65e62, 32'shcdb27bb0, 32'shcdae997a, 
               32'shcdaab7c0, 32'shcda6d683, 32'shcda2f5c2, 32'shcd9f157d, 32'shcd9b35b4, 32'shcd975668, 32'shcd937798, 32'shcd8f9944, 
               32'shcd8bbb6d, 32'shcd87de12, 32'shcd840134, 32'shcd8024d3, 32'shcd7c48ee, 32'shcd786d85, 32'shcd74929a, 32'shcd70b82b, 
               32'shcd6cde39, 32'shcd6904c3, 32'shcd652bcb, 32'shcd61534f, 32'shcd5d7b50, 32'shcd59a3ce, 32'shcd55ccca, 32'shcd51f642, 
               32'shcd4e2037, 32'shcd4a4aa9, 32'shcd467599, 32'shcd42a105, 32'shcd3eccef, 32'shcd3af956, 32'shcd37263a, 32'shcd33539c, 
               32'shcd2f817b, 32'shcd2bafd7, 32'shcd27deb0, 32'shcd240e08, 32'shcd203ddc, 32'shcd1c6e2e, 32'shcd189efe, 32'shcd14d04b, 
               32'shcd110216, 32'shcd0d345f, 32'shcd096725, 32'shcd059a6a, 32'shcd01ce2b, 32'shccfe026b, 32'shccfa3729, 32'shccf66c64, 
               32'shccf2a21d, 32'shcceed855, 32'shcceb0f0a, 32'shcce7463e, 32'shcce37def, 32'shccdfb61f, 32'shccdbeecc, 32'shccd827f8, 
               32'shccd461a2, 32'shccd09bcb, 32'shccccd671, 32'shccc91196, 32'shccc54d3a, 32'shccc1895c, 32'shccbdc5fc, 32'shccba031a, 
               32'shccb640b8, 32'shccb27ed3, 32'shccaebd6e, 32'shccaafc87, 32'shcca73c1e, 32'shcca37c35, 32'shcc9fbcca, 32'shcc9bfddd, 
               32'shcc983f70, 32'shcc948182, 32'shcc90c412, 32'shcc8d0721, 32'shcc894aaf, 32'shcc858ebc, 32'shcc81d349, 32'shcc7e1854, 
               32'shcc7a5dde, 32'shcc76a3e8, 32'shcc72ea70, 32'shcc6f3178, 32'shcc6b78ff, 32'shcc67c105, 32'shcc64098b, 32'shcc605290, 
               32'shcc5c9c14, 32'shcc58e618, 32'shcc55309b, 32'shcc517b9e, 32'shcc4dc720, 32'shcc4a1322, 32'shcc465fa3, 32'shcc42aca4, 
               32'shcc3efa25, 32'shcc3b4825, 32'shcc3796a5, 32'shcc33e5a5, 32'shcc303524, 32'shcc2c8524, 32'shcc28d5a3, 32'shcc2526a2, 
               32'shcc217822, 32'shcc1dca21, 32'shcc1a1ca0, 32'shcc166f9f, 32'shcc12c31f, 32'shcc0f171e, 32'shcc0b6b9e, 32'shcc07c09e, 
               32'shcc04161e, 32'shcc006c1e, 32'shcbfcc29f, 32'shcbf919a0, 32'shcbf57121, 32'shcbf1c923, 32'shcbee21a5, 32'shcbea7aa7, 
               32'shcbe6d42b, 32'shcbe32e2e, 32'shcbdf88b3, 32'shcbdbe3b7, 32'shcbd83f3d, 32'shcbd49b43, 32'shcbd0f7ca, 32'shcbcd54d2, 
               32'shcbc9b25a, 32'shcbc61064, 32'shcbc26eee, 32'shcbbecdf9, 32'shcbbb2d85, 32'shcbb78d92, 32'shcbb3ee20, 32'shcbb04f2f, 
               32'shcbacb0bf, 32'shcba912d1, 32'shcba57563, 32'shcba1d877, 32'shcb9e3c0b, 32'shcb9aa021, 32'shcb9704b9, 32'shcb9369d1, 
               32'shcb8fcf6b, 32'shcb8c3587, 32'shcb889c23, 32'shcb850342, 32'shcb816ae1, 32'shcb7dd303, 32'shcb7a3ba5, 32'shcb76a4ca, 
               32'shcb730e70, 32'shcb6f7898, 32'shcb6be341, 32'shcb684e6c, 32'shcb64ba19, 32'shcb612648, 32'shcb5d92f8, 32'shcb5a002b, 
               32'shcb566ddf, 32'shcb52dc15, 32'shcb4f4acd, 32'shcb4bba08, 32'shcb4829c4, 32'shcb449a02, 32'shcb410ac3, 32'shcb3d7c05, 
               32'shcb39edca, 32'shcb366011, 32'shcb32d2da, 32'shcb2f4626, 32'shcb2bb9f4, 32'shcb282e44, 32'shcb24a316, 32'shcb21186b, 
               32'shcb1d8e43, 32'shcb1a049d, 32'shcb167b79, 32'shcb12f2d8, 32'shcb0f6aba, 32'shcb0be31e, 32'shcb085c05, 32'shcb04d56e, 
               32'shcb014f5b, 32'shcafdc9ca, 32'shcafa44bc, 32'shcaf6c030, 32'shcaf33c28, 32'shcaefb8a2, 32'shcaec35a0, 32'shcae8b320, 
               32'shcae53123, 32'shcae1afaa, 32'shcade2eb3, 32'shcadaae40, 32'shcad72e4f, 32'shcad3aee2, 32'shcad02ff8, 32'shcaccb191, 
               32'shcac933ae, 32'shcac5b64e, 32'shcac23971, 32'shcabebd17, 32'shcabb4141, 32'shcab7c5ef, 32'shcab44b1f, 32'shcab0d0d4, 
               32'shcaad570c, 32'shcaa9ddc7, 32'shcaa66506, 32'shcaa2ecc9, 32'shca9f750f, 32'shca9bfdd9, 32'shca988727, 32'shca9510f8, 
               32'shca919b4e, 32'shca8e2627, 32'shca8ab184, 32'shca873d65, 32'shca83c9ca, 32'shca8056b3, 32'shca7ce420, 32'shca797211, 
               32'shca760086, 32'shca728f7f, 32'shca6f1efc, 32'shca6baefd, 32'shca683f83, 32'shca64d08d, 32'shca61621b, 32'shca5df42d, 
               32'shca5a86c4, 32'shca5719df, 32'shca53ad7e, 32'shca5041a2, 32'shca4cd64b, 32'shca496b77, 32'shca460129, 32'shca42975f, 
               32'shca3f2e19, 32'shca3bc559, 32'shca385d1d, 32'shca34f565, 32'shca318e32, 32'shca2e2784, 32'shca2ac15b, 32'shca275bb7, 
               32'shca23f698, 32'shca2091fd, 32'shca1d2de7, 32'shca19ca57, 32'shca16674b, 32'shca1304c4, 32'shca0fa2c3, 32'shca0c4146, 
               32'shca08e04f, 32'shca057fdd, 32'shca021fef, 32'shc9fec088, 32'shc9fb61a5, 32'shc9f80348, 32'shc9f4a570, 32'shc9f1481d, 
               32'shc9edeb50, 32'shc9ea8f08, 32'shc9e73346, 32'shc9e3d809, 32'shc9e07d51, 32'shc9dd231f, 32'shc9d9c973, 32'shc9d6704c, 
               32'shc9d317ab, 32'shc9cfbf90, 32'shc9cc67fa, 32'shc9c910ea, 32'shc9c5ba60, 32'shc9c2645c, 32'shc9bf0edd, 32'shc9bbb9e5, 
               32'shc9b86572, 32'shc9b51185, 32'shc9b1be1e, 32'shc9ae6b3d, 32'shc9ab18e3, 32'shc9a7c70e, 32'shc9a475bf, 32'shc9a124f7, 
               32'shc99dd4b4, 32'shc99a84f8, 32'shc99735c2, 32'shc993e712, 32'shc99098e9, 32'shc98d4b45, 32'shc989fe29, 32'shc986b192, 
               32'shc9836582, 32'shc98019f8, 32'shc97ccef5, 32'shc9798479, 32'shc9763a83, 32'shc972f113, 32'shc96fa82a, 32'shc96c5fc8, 
               32'shc96917ec, 32'shc965d097, 32'shc96289c9, 32'shc95f4382, 32'shc95bfdc1, 32'shc958b887, 32'shc95573d4, 32'shc9522fa8, 
               32'shc94eec03, 32'shc94ba8e5, 32'shc948664d, 32'shc945243d, 32'shc941e2b4, 32'shc93ea1b2, 32'shc93b6137, 32'shc9382143, 
               32'shc934e1d6, 32'shc931a2f0, 32'shc92e6492, 32'shc92b26bb, 32'shc927e96b, 32'shc924aca3, 32'shc9217062, 32'shc91e34a8, 
               32'shc91af976, 32'shc917becb, 32'shc91484a8, 32'shc9114b0c, 32'shc90e11f7, 32'shc90ad96b, 32'shc907a166, 32'shc90469e8, 
               32'shc90132f2, 32'shc8fdfc84, 32'shc8fac69e, 32'shc8f7913f, 32'shc8f45c68, 32'shc8f12819, 32'shc8edf452, 32'shc8eac112, 
               32'shc8e78e5b, 32'shc8e45c2c, 32'shc8e12a84, 32'shc8ddf965, 32'shc8dac8cd, 32'shc8d798be, 32'shc8d46936, 32'shc8d13a37, 
               32'shc8ce0bc0, 32'shc8caddd1, 32'shc8c7b06b, 32'shc8c4838d, 32'shc8c15736, 32'shc8be2b69, 32'shc8bb0023, 32'shc8b7d566, 
               32'shc8b4ab32, 32'shc8b18185, 32'shc8ae5862, 32'shc8ab2fc6, 32'shc8a807b4, 32'shc8a4e029, 32'shc8a1b928, 32'shc89e92af, 
               32'shc89b6cbf, 32'shc8984757, 32'shc8952278, 32'shc891fe22, 32'shc88eda54, 32'shc88bb710, 32'shc8889454, 32'shc8857221, 
               32'shc8825077, 32'shc87f2f56, 32'shc87c0ebd, 32'shc878eeae, 32'shc875cf28, 32'shc872b02b, 32'shc86f91b7, 32'shc86c73cc, 
               32'shc869566a, 32'shc8663991, 32'shc8631d42, 32'shc860017b, 32'shc85ce63e, 32'shc859cb8a, 32'shc856b160, 32'shc85397bf, 
               32'shc8507ea7, 32'shc84d6619, 32'shc84a4e14, 32'shc8473698, 32'shc8441fa6, 32'shc841093e, 32'shc83df35f, 32'shc83ade0a, 
               32'shc837c93e, 32'shc834b4fc, 32'shc831a143, 32'shc82e8e15, 32'shc82b7b70, 32'shc8286954, 32'shc82557c3, 32'shc82246bb, 
               32'shc81f363d, 32'shc81c2649, 32'shc81916df, 32'shc81607ff, 32'shc812f9a9, 32'shc80febdd, 32'shc80cde9b, 32'shc809d1e3, 
               32'shc806c5b5, 32'shc803ba11, 32'shc800aef7, 32'shc7fda468, 32'shc7fa9a62, 32'shc7f790e7, 32'shc7f487f6, 32'shc7f17f8f, 
               32'shc7ee77b3, 32'shc7eb7061, 32'shc7e8699a, 32'shc7e5635c, 32'shc7e25daa, 32'shc7df5881, 32'shc7dc53e3, 32'shc7d94fd0, 
               32'shc7d64c47, 32'shc7d34949, 32'shc7d046d6, 32'shc7cd44ed, 32'shc7ca438f, 32'shc7c742bb, 32'shc7c44272, 32'shc7c142b4, 
               32'shc7be4381, 32'shc7bb44d8, 32'shc7b846ba, 32'shc7b54928, 32'shc7b24c20, 32'shc7af4fa3, 32'shc7ac53b1, 32'shc7a9584a, 
               32'shc7a65d6e, 32'shc7a3631d, 32'shc7a06957, 32'shc79d701c, 32'shc79a776c, 32'shc7977f48, 32'shc79487ae, 32'shc79190a0, 
               32'shc78e9a1d, 32'shc78ba425, 32'shc788aeb9, 32'shc785b9d8, 32'shc782c582, 32'shc77fd1b8, 32'shc77cde79, 32'shc779ebc5, 
               32'shc776f99d, 32'shc7740801, 32'shc77116f0, 32'shc76e266b, 32'shc76b3671, 32'shc7684702, 32'shc7655820, 32'shc76269c9, 
               32'shc75f7bfe, 32'shc75c8ebe, 32'shc759a20a, 32'shc756b5e2, 32'shc753ca46, 32'shc750df36, 32'shc74df4b1, 32'shc74b0ab9, 
               32'shc748214c, 32'shc745386b, 32'shc7425016, 32'shc73f684e, 32'shc73c8111, 32'shc7399a60, 32'shc736b43c, 32'shc733cea3, 
               32'shc730e997, 32'shc72e0517, 32'shc72b2123, 32'shc7283dbb, 32'shc7255ae0, 32'shc7227890, 32'shc71f96ce, 32'shc71cb597, 
               32'shc719d4ed, 32'shc716f4cf, 32'shc714153e, 32'shc7113639, 32'shc70e57c0, 32'shc70b79d4, 32'shc7089c75, 32'shc705bfa2, 
               32'shc702e35c, 32'shc70007a2, 32'shc6fd2c75, 32'shc6fa51d5, 32'shc6f777c1, 32'shc6f49e3a, 32'shc6f1c540, 32'shc6eeecd3, 
               32'shc6ec14f2, 32'shc6e93d9e, 32'shc6e666d7, 32'shc6e3909d, 32'shc6e0baf0, 32'shc6dde5d0, 32'shc6db113d, 32'shc6d83d37, 
               32'shc6d569be, 32'shc6d296d1, 32'shc6cfc472, 32'shc6ccf2a1, 32'shc6ca215c, 32'shc6c750a4, 32'shc6c4807a, 32'shc6c1b0dd, 
               32'shc6bee1cd, 32'shc6bc134a, 32'shc6b94554, 32'shc6b677ec, 32'shc6b3ab12, 32'shc6b0dec4, 32'shc6ae1304, 32'shc6ab47d2, 
               32'shc6a87d2d, 32'shc6a5b315, 32'shc6a2e98b, 32'shc6a0208f, 32'shc69d5820, 32'shc69a903e, 32'shc697c8eb, 32'shc6950224, 
               32'shc6923bec, 32'shc68f7641, 32'shc68cb124, 32'shc689ec95, 32'shc6872894, 32'shc6846520, 32'shc681a23a, 32'shc67edfe2, 
               32'shc67c1e18, 32'shc6795cdc, 32'shc6769c2e, 32'shc673dc0d, 32'shc6711c7b, 32'shc66e5d77, 32'shc66b9f01, 32'shc668e119, 
               32'shc66623be, 32'shc66366f3, 32'shc660aab5, 32'shc65def05, 32'shc65b33e4, 32'shc6587951, 32'shc655bf4c, 32'shc65305d5, 
               32'shc6504ced, 32'shc64d9493, 32'shc64adcc7, 32'shc648258a, 32'shc6456edb, 32'shc642b8bb, 32'shc6400329, 32'shc63d4e26, 
               32'shc63a99b1, 32'shc637e5ca, 32'shc6353273, 32'shc6327faa, 32'shc62fcd6f, 32'shc62d1bc3, 32'shc62a6aa6, 32'shc627ba17, 
               32'shc6250a18, 32'shc6225aa6, 32'shc61fabc4, 32'shc61cfd71, 32'shc61a4fac, 32'shc617a276, 32'shc614f5cf, 32'shc61249b7, 
               32'shc60f9e2e, 32'shc60cf334, 32'shc60a48c9, 32'shc6079eed, 32'shc604f5a0, 32'shc6024ce2, 32'shc5ffa4b3, 32'shc5fcfd13, 
               32'shc5fa5603, 32'shc5f7af81, 32'shc5f5098f, 32'shc5f2642c, 32'shc5efbf58, 32'shc5ed1b13, 32'shc5ea775e, 32'shc5e7d438, 
               32'shc5e531a1, 32'shc5e28f9a, 32'shc5dfee22, 32'shc5dd4d3a, 32'shc5daace1, 32'shc5d80d17, 32'shc5d56ddd, 32'shc5d2cf33, 
               32'shc5d03118, 32'shc5cd938c, 32'shc5caf690, 32'shc5c85a24, 32'shc5c5be47, 32'shc5c322fb, 32'shc5c0883d, 32'shc5bdee10, 
               32'shc5bb5472, 32'shc5b8bb64, 32'shc5b622e6, 32'shc5b38af8, 32'shc5b0f399, 32'shc5ae5ccb, 32'shc5abc68c, 32'shc5a930dd, 
               32'shc5a69bbe, 32'shc5a4072f, 32'shc5a17330, 32'shc59edfc2, 32'shc59c4ce3, 32'shc599ba94, 32'shc59728d5, 32'shc59497a7, 
               32'shc5920708, 32'shc58f76fa, 32'shc58ce77c, 32'shc58a588e, 32'shc587ca31, 32'shc5853c63, 32'shc582af26, 32'shc580227a, 
               32'shc57d965d, 32'shc57b0ad1, 32'shc5787fd6, 32'shc575f56b, 32'shc5736b90, 32'shc570e246, 32'shc56e598c, 32'shc56bd163, 
               32'shc56949ca, 32'shc566c2c2, 32'shc5643c4a, 32'shc561b663, 32'shc55f310d, 32'shc55cac47, 32'shc55a2812, 32'shc557a46e, 
               32'shc555215a, 32'shc5529ed7, 32'shc5501ce5, 32'shc54d9b84, 32'shc54b1ab4, 32'shc5489a74, 32'shc5461ac6, 32'shc5439ba8, 
               32'shc5411d1b, 32'shc53e9f1f, 32'shc53c21b4, 32'shc539a4da, 32'shc5372891, 32'shc534acd9, 32'shc53231b3, 32'shc52fb71d, 
               32'shc52d3d18, 32'shc52ac3a5, 32'shc5284ac3, 32'shc525d272, 32'shc5235ab2, 32'shc520e383, 32'shc51e6ce6, 32'shc51bf6da, 
               32'shc519815f, 32'shc5170c75, 32'shc514981d, 32'shc5122457, 32'shc50fb121, 32'shc50d3e7d, 32'shc50acc6b, 32'shc5085aea, 
               32'shc505e9fb, 32'shc503799d, 32'shc50109d0, 32'shc4fe9a95, 32'shc4fc2bec, 32'shc4f9bdd4, 32'shc4f7504e, 32'shc4f4e35a, 
               32'shc4f276f7, 32'shc4f00b27, 32'shc4ed9fe7, 32'shc4eb353a, 32'shc4e8cb1e, 32'shc4e66194, 32'shc4e3f89c, 32'shc4e19036, 
               32'shc4df2862, 32'shc4dcc11f, 32'shc4da5a6f, 32'shc4d7f450, 32'shc4d58ec3, 32'shc4d329c9, 32'shc4d0c560, 32'shc4ce6189, 
               32'shc4cbfe45, 32'shc4c99b92, 32'shc4c73972, 32'shc4c4d7e4, 32'shc4c276e8, 32'shc4c0167e, 32'shc4bdb6a6, 32'shc4bb5760, 
               32'shc4b8f8ad, 32'shc4b69a8c, 32'shc4b43cfd, 32'shc4b1e001, 32'shc4af8397, 32'shc4ad27bf, 32'shc4aacc7a, 32'shc4a871c7, 
               32'shc4a617a6, 32'shc4a3be18, 32'shc4a1651c, 32'shc49f0cb3, 32'shc49cb4dd, 32'shc49a5d98, 32'shc49806e7, 32'shc495b0c8, 
               32'shc4935b3c, 32'shc4910642, 32'shc48eb1db, 32'shc48c5e06, 32'shc48a0ac4, 32'shc487b815, 32'shc48565f9, 32'shc4831470, 
               32'shc480c379, 32'shc47e7315, 32'shc47c2344, 32'shc479d405, 32'shc477855a, 32'shc4753741, 32'shc472e9bc, 32'shc4709cc9, 
               32'shc46e5069, 32'shc46c049d, 32'shc469b963, 32'shc4676ebc, 32'shc46524a9, 32'shc462db28, 32'shc460923b, 32'shc45e49e0, 
               32'shc45c0219, 32'shc459bae5, 32'shc4577444, 32'shc4552e36, 32'shc452e8bc, 32'shc450a3d4, 32'shc44e5f80, 32'shc44c1bc0, 
               32'shc449d892, 32'shc44795f8, 32'shc44553f2, 32'shc443127e, 32'shc440d19e, 32'shc43e9152, 32'shc43c5199, 32'shc43a1273, 
               32'shc437d3e1, 32'shc43595e3, 32'shc4335877, 32'shc4311ba0, 32'shc42edf5c, 32'shc42ca3ac, 32'shc42a688f, 32'shc4282e06, 
               32'shc425f410, 32'shc423baae, 32'shc42181e0, 32'shc41f49a6, 32'shc41d11ff, 32'shc41adaed, 32'shc418a46d, 32'shc4166e82, 
               32'shc414392b, 32'shc4120467, 32'shc40fd037, 32'shc40d9c9c, 32'shc40b6994, 32'shc4093720, 32'shc4070540, 32'shc404d3f4, 
               32'shc402a33c, 32'shc4007318, 32'shc3fe4388, 32'shc3fc148c, 32'shc3f9e624, 32'shc3f7b850, 32'shc3f58b10, 32'shc3f35e65, 
               32'shc3f1324e, 32'shc3ef06cb, 32'shc3ecdbdc, 32'shc3eab181, 32'shc3e887bb, 32'shc3e65e88, 32'shc3e435ea, 32'shc3e20de1, 
               32'shc3dfe66c, 32'shc3ddbf8b, 32'shc3db993e, 32'shc3d97386, 32'shc3d74e62, 32'shc3d529d3, 32'shc3d305d8, 32'shc3d0e272, 
               32'shc3cebfa0, 32'shc3cc9d63, 32'shc3ca7bba, 32'shc3c85aa6, 32'shc3c63a26, 32'shc3c41a3b, 32'shc3c1fae5, 32'shc3bfdc23, 
               32'shc3bdbdf6, 32'shc3bba05e, 32'shc3b9835a, 32'shc3b766eb, 32'shc3b54b11, 32'shc3b32fcb, 32'shc3b1151b, 32'shc3aefaff, 
               32'shc3ace178, 32'shc3aac885, 32'shc3a8b028, 32'shc3a6985f, 32'shc3a4812c, 32'shc3a26a8d, 32'shc3a05484, 32'shc39e3f0f, 
               32'shc39c2a2f, 32'shc39a15e4, 32'shc398022f, 32'shc395ef0e, 32'shc393dc82, 32'shc391ca8c, 32'shc38fb92a, 32'shc38da85e, 
               32'shc38b9827, 32'shc3898885, 32'shc3877978, 32'shc3856b01, 32'shc3835d1e, 32'shc3814fd1, 32'shc37f4319, 32'shc37d36f7, 
               32'shc37b2b6a, 32'shc3792072, 32'shc377160f, 32'shc3750c42, 32'shc373030a, 32'shc370fa68, 32'shc36ef25b, 32'shc36ceae3, 
               32'shc36ae401, 32'shc368ddb4, 32'shc366d7fd, 32'shc364d2dc, 32'shc362ce50, 32'shc360ca59, 32'shc35ec6f8, 32'shc35cc42d, 
               32'shc35ac1f7, 32'shc358c057, 32'shc356bf4d, 32'shc354bed8, 32'shc352bef9, 32'shc350bfaf, 32'shc34ec0fc, 32'shc34cc2de, 
               32'shc34ac556, 32'shc348c864, 32'shc346cc07, 32'shc344d041, 32'shc342d510, 32'shc340da75, 32'shc33ee070, 32'shc33ce701, 
               32'shc33aee27, 32'shc338f5e4, 32'shc336fe37, 32'shc3350720, 32'shc333109e, 32'shc3311ab3, 32'shc32f255e, 32'shc32d309e, 
               32'shc32b3c75, 32'shc32948e2, 32'shc32755e5, 32'shc325637f, 32'shc32371ae, 32'shc3218073, 32'shc31f8fcf, 32'shc31d9fc1, 
               32'shc31bb049, 32'shc319c168, 32'shc317d31c, 32'shc315e567, 32'shc313f848, 32'shc3120bc0, 32'shc3101fce, 32'shc30e3472, 
               32'shc30c49ad, 32'shc30a5f7e, 32'shc30875e5, 32'shc3068ce3, 32'shc304a477, 32'shc302bca2, 32'shc300d563, 32'shc2feeebb, 
               32'shc2fd08a9, 32'shc2fb232e, 32'shc2f93e4a, 32'shc2f759fc, 32'shc2f57644, 32'shc2f39323, 32'shc2f1b099, 32'shc2efcea6, 
               32'shc2eded49, 32'shc2ec0c82, 32'shc2ea2c53, 32'shc2e84cba, 32'shc2e66db8, 32'shc2e48f4d, 32'shc2e2b178, 32'shc2e0d43b, 
               32'shc2def794, 32'shc2dd1b84, 32'shc2db400a, 32'shc2d96528, 32'shc2d78add, 32'shc2d5b128, 32'shc2d3d80a, 32'shc2d1ff84, 
               32'shc2d02794, 32'shc2ce503b, 32'shc2cc7979, 32'shc2caa34f, 32'shc2c8cdbb, 32'shc2c6f8be, 32'shc2c52459, 32'shc2c3508a, 
               32'shc2c17d52, 32'shc2bfaab2, 32'shc2bdd8a9, 32'shc2bc0737, 32'shc2ba365c, 32'shc2b86618, 32'shc2b6966c, 32'shc2b4c756, 
               32'shc2b2f8d8, 32'shc2b12af1, 32'shc2af5da2, 32'shc2ad90ea, 32'shc2abc4c9, 32'shc2a9f93f, 32'shc2a82e4d, 32'shc2a663f2, 
               32'shc2a49a2e, 32'shc2a2d102, 32'shc2a1086d, 32'shc29f4070, 32'shc29d790a, 32'shc29bb23c, 32'shc299ec05, 32'shc2982665, 
               32'shc296615d, 32'shc2949ced, 32'shc292d914, 32'shc29115d3, 32'shc28f5329, 32'shc28d9117, 32'shc28bcf9c, 32'shc28a0eb9, 
               32'shc2884e6e, 32'shc2868ebb, 32'shc284cf9f, 32'shc283111b, 32'shc281532e, 32'shc27f95d9, 32'shc27dd91c, 32'shc27c1cf7, 
               32'shc27a616a, 32'shc278a674, 32'shc276ec16, 32'shc2753250, 32'shc2737922, 32'shc271c08c, 32'shc270088e, 32'shc26e5127, 
               32'shc26c9a58, 32'shc26ae422, 32'shc2692e83, 32'shc267797c, 32'shc265c50e, 32'shc2641137, 32'shc2625df8, 32'shc260ab51, 
               32'shc25ef943, 32'shc25d47cc, 32'shc25b96ee, 32'shc259e6a7, 32'shc25836f9, 32'shc25687e3, 32'shc254d965, 32'shc2532b7f, 
               32'shc2517e31, 32'shc24fd17c, 32'shc24e255e, 32'shc24c79d9, 32'shc24aceed, 32'shc2492498, 32'shc2477adc, 32'shc245d1b8, 
               32'shc244292c, 32'shc2428139, 32'shc240d9de, 32'shc23f331b, 32'shc23d8cf1, 32'shc23be75f, 32'shc23a4265, 32'shc2389e04, 
               32'shc236fa3b, 32'shc235570b, 32'shc233b473, 32'shc2321274, 32'shc230710d, 32'shc22ed03f, 32'shc22d3009, 32'shc22b906c, 
               32'shc229f167, 32'shc22852fb, 32'shc226b528, 32'shc22517ed, 32'shc2237b4b, 32'shc221df41, 32'shc22043d0, 32'shc21ea8f8, 
               32'shc21d0eb8, 32'shc21b7511, 32'shc219dc03, 32'shc218438e, 32'shc216abb1, 32'shc215146d, 32'shc2137dc2, 32'shc211e7af, 
               32'shc2105236, 32'shc20ebd55, 32'shc20d290d, 32'shc20b955e, 32'shc20a0248, 32'shc2086fca, 32'shc206dde6, 32'shc2054c9b, 
               32'shc203bbe8, 32'shc2022bce, 32'shc2009c4e, 32'shc1ff0d66, 32'shc1fd7f17, 32'shc1fbf161, 32'shc1fa6445, 32'shc1f8d7c1, 
               32'shc1f74bd6, 32'shc1f5c085, 32'shc1f435cc, 32'shc1f2abad, 32'shc1f12227, 32'shc1ef9939, 32'shc1ee10e5, 32'shc1ec892b, 
               32'shc1eb0209, 32'shc1e97b80, 32'shc1e7f591, 32'shc1e6703b, 32'shc1e4eb7e, 32'shc1e3675a, 32'shc1e1e3d0, 32'shc1e060df, 
               32'shc1dede87, 32'shc1dd5cc8, 32'shc1dbdba3, 32'shc1da5b17, 32'shc1d8db25, 32'shc1d75bcb, 32'shc1d5dd0c, 32'shc1d45ee5, 
               32'shc1d2e158, 32'shc1d16464, 32'shc1cfe80a, 32'shc1ce6c49, 32'shc1ccf122, 32'shc1cb7694, 32'shc1c9fca0, 32'shc1c88345, 
               32'shc1c70a84, 32'shc1c5925c, 32'shc1c41ace, 32'shc1c2a3d9, 32'shc1c12d7e, 32'shc1bfb7bc, 32'shc1be4294, 32'shc1bcce06, 
               32'shc1bb5a11, 32'shc1b9e6b6, 32'shc1b873f5, 32'shc1b701cd, 32'shc1b5903f, 32'shc1b41f4a, 32'shc1b2aef0, 32'shc1b13f2f, 
               32'shc1afd007, 32'shc1ae617a, 32'shc1acf386, 32'shc1ab862c, 32'shc1aa196c, 32'shc1a8ad46, 32'shc1a741b9, 32'shc1a5d6c7, 
               32'shc1a46c6e, 32'shc1a302af, 32'shc1a1998a, 32'shc1a030ff, 32'shc19ec90d, 32'shc19d61b6, 32'shc19bfaf9, 32'shc19a94d5, 
               32'shc1992f4c, 32'shc197ca5c, 32'shc1966606, 32'shc195024b, 32'shc1939f29, 32'shc1923ca2, 32'shc190dab4, 32'shc18f7961, 
               32'shc18e18a7, 32'shc18cb888, 32'shc18b5903, 32'shc189fa17, 32'shc1889bc6, 32'shc1873e10, 32'shc185e0f3, 32'shc1848470, 
               32'shc1832888, 32'shc181cd3a, 32'shc1807285, 32'shc17f186c, 32'shc17dbeec, 32'shc17c6607, 32'shc17b0dbb, 32'shc179b60b, 
               32'shc1785ef4, 32'shc1770878, 32'shc175b296, 32'shc1745d4e, 32'shc17308a1, 32'shc171b48e, 32'shc1706115, 32'shc16f0e36, 
               32'shc16dbbf3, 32'shc16c6a49, 32'shc16b193a, 32'shc169c8c5, 32'shc16878eb, 32'shc16729ab, 32'shc165db05, 32'shc1648cfa, 
               32'shc1633f8a, 32'shc161f2b4, 32'shc160a678, 32'shc15f5ad7, 32'shc15e0fd1, 32'shc15cc565, 32'shc15b7b94, 32'shc15a325d, 
               32'shc158e9c1, 32'shc157a1bf, 32'shc1565a58, 32'shc155138c, 32'shc153cd5a, 32'shc15287c3, 32'shc15142c6, 32'shc14ffe64, 
               32'shc14eba9d, 32'shc14d7771, 32'shc14c34df, 32'shc14af2e8, 32'shc149b18b, 32'shc14870ca, 32'shc14730a3, 32'shc145f117, 
               32'shc144b225, 32'shc14373cf, 32'shc1423613, 32'shc140f8f2, 32'shc13fbc6c, 32'shc13e8081, 32'shc13d4530, 32'shc13c0a7b, 
               32'shc13ad060, 32'shc13996e0, 32'shc1385dfb, 32'shc13725b1, 32'shc135ee02, 32'shc134b6ee, 32'shc1338075, 32'shc1324a96, 
               32'shc1311553, 32'shc12fe0ab, 32'shc12eac9d, 32'shc12d792b, 32'shc12c4653, 32'shc12b1417, 32'shc129e276, 32'shc128b16f, 
               32'shc1278104, 32'shc1265134, 32'shc12521ff, 32'shc123f365, 32'shc122c566, 32'shc1219802, 32'shc1206b39, 32'shc11f3f0c, 
               32'shc11e1379, 32'shc11ce882, 32'shc11bbe26, 32'shc11a9465, 32'shc1196b3f, 32'shc11842b5, 32'shc1171ac6, 32'shc115f372, 
               32'shc114ccb9, 32'shc113a69b, 32'shc1128119, 32'shc1115c32, 32'shc11037e6, 32'shc10f1435, 32'shc10df120, 32'shc10ccea6, 
               32'shc10bacc8, 32'shc10a8b85, 32'shc1096add, 32'shc1084ad0, 32'shc1072b5f, 32'shc1060c89, 32'shc104ee4f, 32'shc103d0b0, 
               32'shc102b3ac, 32'shc1019744, 32'shc1007b77, 32'shc0ff6046, 32'shc0fe45b0, 32'shc0fd2bb6, 32'shc0fc1257, 32'shc0faf993, 
               32'shc0f9e16b, 32'shc0f8c9df, 32'shc0f7b2ee, 32'shc0f69c99, 32'shc0f586df, 32'shc0f471c1, 32'shc0f35d3e, 32'shc0f24957, 
               32'shc0f1360b, 32'shc0f0235b, 32'shc0ef1147, 32'shc0edffce, 32'shc0eceef1, 32'shc0ebdeaf, 32'shc0eacf09, 32'shc0e9bfff, 
               32'shc0e8b190, 32'shc0e7a3bd, 32'shc0e69686, 32'shc0e589eb, 32'shc0e47deb, 32'shc0e37287, 32'shc0e267be, 32'shc0e15d92, 
               32'shc0e05401, 32'shc0df4b0b, 32'shc0de42b2, 32'shc0dd3af4, 32'shc0dc33d2, 32'shc0db2d4c, 32'shc0da2762, 32'shc0d92214, 
               32'shc0d81d61, 32'shc0d7194a, 32'shc0d615cf, 32'shc0d512f0, 32'shc0d410ad, 32'shc0d30f05, 32'shc0d20dfa, 32'shc0d10d8a, 
               32'shc0d00db6, 32'shc0cf0e7f, 32'shc0ce0fe3, 32'shc0cd11e3, 32'shc0cc147f, 32'shc0cb17b7, 32'shc0ca1b8a, 32'shc0c91ffa, 
               32'shc0c82506, 32'shc0c72aae, 32'shc0c630f2, 32'shc0c537d1, 32'shc0c43f4d, 32'shc0c34765, 32'shc0c25019, 32'shc0c15969, 
               32'shc0c06355, 32'shc0bf6ddd, 32'shc0be7901, 32'shc0bd84c1, 32'shc0bc911d, 32'shc0bb9e15, 32'shc0baabaa, 32'shc0b9b9da, 
               32'shc0b8c8a7, 32'shc0b7d810, 32'shc0b6e815, 32'shc0b5f8b6, 32'shc0b509f3, 32'shc0b41bcd, 32'shc0b32e42, 32'shc0b24154, 
               32'shc0b15502, 32'shc0b0694c, 32'shc0af7e33, 32'shc0ae93b5, 32'shc0ada9d4, 32'shc0acc08f, 32'shc0abd7e6, 32'shc0aaefda, 
               32'shc0aa086a, 32'shc0a92196, 32'shc0a83b5e, 32'shc0a755c3, 32'shc0a670c4, 32'shc0a58c62, 32'shc0a4a89b, 32'shc0a3c571, 
               32'shc0a2e2e3, 32'shc0a200f2, 32'shc0a11f9d, 32'shc0a03ee4, 32'shc09f5ec8, 32'shc09e7f48, 32'shc09da065, 32'shc09cc21e, 
               32'shc09be473, 32'shc09b0765, 32'shc09a2af3, 32'shc0994f1d, 32'shc09873e4, 32'shc0979948, 32'shc096bf48, 32'shc095e5e4, 
               32'shc0950d1d, 32'shc09434f2, 32'shc0935d64, 32'shc0928672, 32'shc091b01d, 32'shc090da64, 32'shc0900548, 32'shc08f30c8, 
               32'shc08e5ce5, 32'shc08d899f, 32'shc08cb6f5, 32'shc08be4e7, 32'shc08b1376, 32'shc08a42a2, 32'shc089726a, 32'shc088a2cf, 
               32'shc087d3d0, 32'shc087056e, 32'shc08637a9, 32'shc0856a80, 32'shc0849df4, 32'shc083d204, 32'shc08306b2, 32'shc0823bfb, 
               32'shc08171e2, 32'shc080a865, 32'shc07fdf85, 32'shc07f1741, 32'shc07e4f9b, 32'shc07d8890, 32'shc07cc223, 32'shc07bfc52, 
               32'shc07b371e, 32'shc07a7287, 32'shc079ae8c, 32'shc078eb2f, 32'shc078286e, 32'shc0776649, 32'shc076a4c2, 32'shc075e3d7, 
               32'shc0752389, 32'shc07463d8, 32'shc073a4c3, 32'shc072e64c, 32'shc0722871, 32'shc0716b33, 32'shc070ae92, 32'shc06ff28e, 
               32'shc06f3726, 32'shc06e7c5b, 32'shc06dc22e, 32'shc06d089d, 32'shc06c4fa8, 32'shc06b9751, 32'shc06adf97, 32'shc06a2879, 
               32'shc06971f9, 32'shc068bc15, 32'shc06806ce, 32'shc0675225, 32'shc0669e18, 32'shc065eaa8, 32'shc06537d4, 32'shc064859e, 
               32'shc063d405, 32'shc0632309, 32'shc06272aa, 32'shc061c2e7, 32'shc06113c2, 32'shc060653a, 32'shc05fb74e, 32'shc05f0a00, 
               32'shc05e5d4e, 32'shc05db13a, 32'shc05d05c3, 32'shc05c5ae8, 32'shc05bb0ab, 32'shc05b070a, 32'shc05a5e07, 32'shc059b5a1, 
               32'shc0590dd8, 32'shc05866ac, 32'shc057c01d, 32'shc0571a2b, 32'shc05674d6, 32'shc055d01e, 32'shc0552c03, 32'shc0548885, 
               32'shc053e5a5, 32'shc0534361, 32'shc052a1bb, 32'shc05200b2, 32'shc0516045, 32'shc050c077, 32'shc0502145, 32'shc04f82b0, 
               32'shc04ee4b8, 32'shc04e475e, 32'shc04daaa1, 32'shc04d0e81, 32'shc04c72fe, 32'shc04bd818, 32'shc04b3dcf, 32'shc04aa424, 
               32'shc04a0b16, 32'shc04972a5, 32'shc048dad1, 32'shc048439b, 32'shc047ad01, 32'shc0471705, 32'shc04681a6, 32'shc045ece5, 
               32'shc04558c0, 32'shc044c539, 32'shc044324f, 32'shc043a002, 32'shc0430e53, 32'shc0427d41, 32'shc041eccc, 32'shc0415cf4, 
               32'shc040cdba, 32'shc0403f1d, 32'shc03fb11d, 32'shc03f23bb, 32'shc03e96f6, 32'shc03e0ace, 32'shc03d7f44, 32'shc03cf456, 
               32'shc03c6a07, 32'shc03be054, 32'shc03b573f, 32'shc03acec7, 32'shc03a46ed, 32'shc039bfaf, 32'shc0393910, 32'shc038b30d, 
               32'shc0382da8, 32'shc037a8e1, 32'shc03724b6, 32'shc036a129, 32'shc0361e3a, 32'shc0359be8, 32'shc0351a33, 32'shc034991c, 
               32'shc03418a2, 32'shc03398c5, 32'shc0331986, 32'shc0329ae4, 32'shc0321ce0, 32'shc0319f79, 32'shc03122b0, 32'shc030a684, 
               32'shc0302af5, 32'shc02fb004, 32'shc02f35b1, 32'shc02ebbfb, 32'shc02e42e2, 32'shc02dca67, 32'shc02d5289, 32'shc02cdb49, 
               32'shc02c64a6, 32'shc02beea1, 32'shc02b7939, 32'shc02b046f, 32'shc02a9042, 32'shc02a1cb2, 32'shc029a9c1, 32'shc029376c, 
               32'shc028c5b6, 32'shc028549c, 32'shc027e421, 32'shc0277442, 32'shc0270502, 32'shc026965f, 32'shc0262859, 32'shc025baf1, 
               32'shc0254e27, 32'shc024e1fa, 32'shc024766a, 32'shc0240b78, 32'shc023a124, 32'shc023376e, 32'shc022ce54, 32'shc02265d9, 
               32'shc021fdfb, 32'shc02196bb, 32'shc0213018, 32'shc020ca13, 32'shc02064ab, 32'shc01fffe1, 32'shc01f9bb5, 32'shc01f3826, 
               32'shc01ed535, 32'shc01e72e1, 32'shc01e112b, 32'shc01db013, 32'shc01d4f99, 32'shc01cefbb, 32'shc01c907c, 32'shc01c31da, 
               32'shc01bd3d6, 32'shc01b7670, 32'shc01b19a7, 32'shc01abd7c, 32'shc01a61ee, 32'shc01a06fe, 32'shc019acac, 32'shc01952f8, 
               32'shc018f9e1, 32'shc018a168, 32'shc018498c, 32'shc017f24e, 32'shc0179bae, 32'shc01745ac, 32'shc016f047, 32'shc0169b80, 
               32'shc0164757, 32'shc015f3cb, 32'shc015a0dd, 32'shc0154e8d, 32'shc014fcda, 32'shc014abc5, 32'shc0145b4e, 32'shc0140b75, 
               32'shc013bc39, 32'shc0136d9b, 32'shc0131f9b, 32'shc012d238, 32'shc0128574, 32'shc012394c, 32'shc011edc3, 32'shc011a2d8, 
               32'shc011588a, 32'shc0110eda, 32'shc010c5c7, 32'shc0107d53, 32'shc010357c, 32'shc00fee43, 32'shc00fa7a8, 32'shc00f61aa, 
               32'shc00f1c4a, 32'shc00ed788, 32'shc00e9364, 32'shc00e4fde, 32'shc00e0cf5, 32'shc00dcaaa, 32'shc00d88fd, 32'shc00d47ed, 
               32'shc00d077c, 32'shc00cc7a8, 32'shc00c8872, 32'shc00c49da, 32'shc00c0be0, 32'shc00bce83, 32'shc00b91c4, 32'shc00b55a3, 
               32'shc00b1a20, 32'shc00adf3b, 32'shc00aa4f3, 32'shc00a6b49, 32'shc00a323d, 32'shc009f9cf, 32'shc009c1ff, 32'shc0098acc, 
               32'shc0095438, 32'shc0091e41, 32'shc008e8e8, 32'shc008b42d, 32'shc008800f, 32'shc0084c90, 32'shc00819ae, 32'shc007e76a, 
               32'shc007b5c4, 32'shc00784bc, 32'shc0075452, 32'shc0072485, 32'shc006f556, 32'shc006c6c6, 32'shc00698d3, 32'shc0066b7d, 
               32'shc0063ec6, 32'shc00612ad, 32'shc005e731, 32'shc005bc54, 32'shc0059214, 32'shc0056872, 32'shc0053f6e, 32'shc0051707, 
               32'shc004ef3f, 32'shc004c814, 32'shc004a188, 32'shc0047b99, 32'shc0045648, 32'shc0043195, 32'shc0040d80, 32'shc003ea09, 
               32'shc003c72f, 32'shc003a4f4, 32'shc0038356, 32'shc0036256, 32'shc00341f4, 32'shc0032230, 32'shc003030a, 32'shc002e482, 
               32'shc002c697, 32'shc002a94b, 32'shc0028c9c, 32'shc002708c, 32'shc0025519, 32'shc0023a44, 32'shc002200d, 32'shc0020674, 
               32'shc001ed78, 32'shc001d51b, 32'shc001bd5c, 32'shc001a63a, 32'shc0018fb6, 32'shc00179d1, 32'shc0016489, 32'shc0014fdf, 
               32'shc0013bd3, 32'shc0012865, 32'shc0011594, 32'shc0010362, 32'shc000f1ce, 32'shc000e0d7, 32'shc000d07e, 32'shc000c0c4, 
               32'shc000b1a7, 32'shc000a328, 32'shc0009547, 32'shc0008804, 32'shc0007b5f, 32'shc0006f57, 32'shc00063ee, 32'shc0005922, 
               32'shc0004ef5, 32'shc0004565, 32'shc0003c74, 32'shc0003420, 32'shc0002c6a, 32'shc0002552, 32'shc0001ed8, 32'shc00018fb, 
               32'shc00013bd, 32'shc0000f1d, 32'shc0000b1a, 32'shc00007b6, 32'shc00004ef, 32'shc00002c7, 32'shc000013c, 32'shc000004f, 
               32'shc0000000, 32'shc000004f, 32'shc000013c, 32'shc00002c7, 32'shc00004ef, 32'shc00007b6, 32'shc0000b1a, 32'shc0000f1d, 
               32'shc00013bd, 32'shc00018fb, 32'shc0001ed8, 32'shc0002552, 32'shc0002c6a, 32'shc0003420, 32'shc0003c74, 32'shc0004565, 
               32'shc0004ef5, 32'shc0005922, 32'shc00063ee, 32'shc0006f57, 32'shc0007b5f, 32'shc0008804, 32'shc0009547, 32'shc000a328, 
               32'shc000b1a7, 32'shc000c0c4, 32'shc000d07e, 32'shc000e0d7, 32'shc000f1ce, 32'shc0010362, 32'shc0011594, 32'shc0012865, 
               32'shc0013bd3, 32'shc0014fdf, 32'shc0016489, 32'shc00179d1, 32'shc0018fb6, 32'shc001a63a, 32'shc001bd5c, 32'shc001d51b, 
               32'shc001ed78, 32'shc0020674, 32'shc002200d, 32'shc0023a44, 32'shc0025519, 32'shc002708c, 32'shc0028c9c, 32'shc002a94b, 
               32'shc002c697, 32'shc002e482, 32'shc003030a, 32'shc0032230, 32'shc00341f4, 32'shc0036256, 32'shc0038356, 32'shc003a4f4, 
               32'shc003c72f, 32'shc003ea09, 32'shc0040d80, 32'shc0043195, 32'shc0045648, 32'shc0047b99, 32'shc004a188, 32'shc004c814, 
               32'shc004ef3f, 32'shc0051707, 32'shc0053f6e, 32'shc0056872, 32'shc0059214, 32'shc005bc54, 32'shc005e731, 32'shc00612ad, 
               32'shc0063ec6, 32'shc0066b7d, 32'shc00698d3, 32'shc006c6c6, 32'shc006f556, 32'shc0072485, 32'shc0075452, 32'shc00784bc, 
               32'shc007b5c4, 32'shc007e76a, 32'shc00819ae, 32'shc0084c90, 32'shc008800f, 32'shc008b42d, 32'shc008e8e8, 32'shc0091e41, 
               32'shc0095438, 32'shc0098acc, 32'shc009c1ff, 32'shc009f9cf, 32'shc00a323d, 32'shc00a6b49, 32'shc00aa4f3, 32'shc00adf3b, 
               32'shc00b1a20, 32'shc00b55a3, 32'shc00b91c4, 32'shc00bce83, 32'shc00c0be0, 32'shc00c49da, 32'shc00c8872, 32'shc00cc7a8, 
               32'shc00d077c, 32'shc00d47ed, 32'shc00d88fd, 32'shc00dcaaa, 32'shc00e0cf5, 32'shc00e4fde, 32'shc00e9364, 32'shc00ed788, 
               32'shc00f1c4a, 32'shc00f61aa, 32'shc00fa7a8, 32'shc00fee43, 32'shc010357c, 32'shc0107d53, 32'shc010c5c7, 32'shc0110eda, 
               32'shc011588a, 32'shc011a2d8, 32'shc011edc3, 32'shc012394c, 32'shc0128574, 32'shc012d238, 32'shc0131f9b, 32'shc0136d9b, 
               32'shc013bc39, 32'shc0140b75, 32'shc0145b4e, 32'shc014abc5, 32'shc014fcda, 32'shc0154e8d, 32'shc015a0dd, 32'shc015f3cb, 
               32'shc0164757, 32'shc0169b80, 32'shc016f047, 32'shc01745ac, 32'shc0179bae, 32'shc017f24e, 32'shc018498c, 32'shc018a168, 
               32'shc018f9e1, 32'shc01952f8, 32'shc019acac, 32'shc01a06fe, 32'shc01a61ee, 32'shc01abd7c, 32'shc01b19a7, 32'shc01b7670, 
               32'shc01bd3d6, 32'shc01c31da, 32'shc01c907c, 32'shc01cefbb, 32'shc01d4f99, 32'shc01db013, 32'shc01e112b, 32'shc01e72e1, 
               32'shc01ed535, 32'shc01f3826, 32'shc01f9bb5, 32'shc01fffe1, 32'shc02064ab, 32'shc020ca13, 32'shc0213018, 32'shc02196bb, 
               32'shc021fdfb, 32'shc02265d9, 32'shc022ce54, 32'shc023376e, 32'shc023a124, 32'shc0240b78, 32'shc024766a, 32'shc024e1fa, 
               32'shc0254e27, 32'shc025baf1, 32'shc0262859, 32'shc026965f, 32'shc0270502, 32'shc0277442, 32'shc027e421, 32'shc028549c, 
               32'shc028c5b6, 32'shc029376c, 32'shc029a9c1, 32'shc02a1cb2, 32'shc02a9042, 32'shc02b046f, 32'shc02b7939, 32'shc02beea1, 
               32'shc02c64a6, 32'shc02cdb49, 32'shc02d5289, 32'shc02dca67, 32'shc02e42e2, 32'shc02ebbfb, 32'shc02f35b1, 32'shc02fb004, 
               32'shc0302af5, 32'shc030a684, 32'shc03122b0, 32'shc0319f79, 32'shc0321ce0, 32'shc0329ae4, 32'shc0331986, 32'shc03398c5, 
               32'shc03418a2, 32'shc034991c, 32'shc0351a33, 32'shc0359be8, 32'shc0361e3a, 32'shc036a129, 32'shc03724b6, 32'shc037a8e1, 
               32'shc0382da8, 32'shc038b30d, 32'shc0393910, 32'shc039bfaf, 32'shc03a46ed, 32'shc03acec7, 32'shc03b573f, 32'shc03be054, 
               32'shc03c6a07, 32'shc03cf456, 32'shc03d7f44, 32'shc03e0ace, 32'shc03e96f6, 32'shc03f23bb, 32'shc03fb11d, 32'shc0403f1d, 
               32'shc040cdba, 32'shc0415cf4, 32'shc041eccc, 32'shc0427d41, 32'shc0430e53, 32'shc043a002, 32'shc044324f, 32'shc044c539, 
               32'shc04558c0, 32'shc045ece5, 32'shc04681a6, 32'shc0471705, 32'shc047ad01, 32'shc048439b, 32'shc048dad1, 32'shc04972a5, 
               32'shc04a0b16, 32'shc04aa424, 32'shc04b3dcf, 32'shc04bd818, 32'shc04c72fe, 32'shc04d0e81, 32'shc04daaa1, 32'shc04e475e, 
               32'shc04ee4b8, 32'shc04f82b0, 32'shc0502145, 32'shc050c077, 32'shc0516045, 32'shc05200b2, 32'shc052a1bb, 32'shc0534361, 
               32'shc053e5a5, 32'shc0548885, 32'shc0552c03, 32'shc055d01e, 32'shc05674d6, 32'shc0571a2b, 32'shc057c01d, 32'shc05866ac, 
               32'shc0590dd8, 32'shc059b5a1, 32'shc05a5e07, 32'shc05b070a, 32'shc05bb0ab, 32'shc05c5ae8, 32'shc05d05c3, 32'shc05db13a, 
               32'shc05e5d4e, 32'shc05f0a00, 32'shc05fb74e, 32'shc060653a, 32'shc06113c2, 32'shc061c2e7, 32'shc06272aa, 32'shc0632309, 
               32'shc063d405, 32'shc064859e, 32'shc06537d4, 32'shc065eaa8, 32'shc0669e18, 32'shc0675225, 32'shc06806ce, 32'shc068bc15, 
               32'shc06971f9, 32'shc06a2879, 32'shc06adf97, 32'shc06b9751, 32'shc06c4fa8, 32'shc06d089d, 32'shc06dc22e, 32'shc06e7c5b, 
               32'shc06f3726, 32'shc06ff28e, 32'shc070ae92, 32'shc0716b33, 32'shc0722871, 32'shc072e64c, 32'shc073a4c3, 32'shc07463d8, 
               32'shc0752389, 32'shc075e3d7, 32'shc076a4c2, 32'shc0776649, 32'shc078286e, 32'shc078eb2f, 32'shc079ae8c, 32'shc07a7287, 
               32'shc07b371e, 32'shc07bfc52, 32'shc07cc223, 32'shc07d8890, 32'shc07e4f9b, 32'shc07f1741, 32'shc07fdf85, 32'shc080a865, 
               32'shc08171e2, 32'shc0823bfb, 32'shc08306b2, 32'shc083d204, 32'shc0849df4, 32'shc0856a80, 32'shc08637a9, 32'shc087056e, 
               32'shc087d3d0, 32'shc088a2cf, 32'shc089726a, 32'shc08a42a2, 32'shc08b1376, 32'shc08be4e7, 32'shc08cb6f5, 32'shc08d899f, 
               32'shc08e5ce5, 32'shc08f30c8, 32'shc0900548, 32'shc090da64, 32'shc091b01d, 32'shc0928672, 32'shc0935d64, 32'shc09434f2, 
               32'shc0950d1d, 32'shc095e5e4, 32'shc096bf48, 32'shc0979948, 32'shc09873e4, 32'shc0994f1d, 32'shc09a2af3, 32'shc09b0765, 
               32'shc09be473, 32'shc09cc21e, 32'shc09da065, 32'shc09e7f48, 32'shc09f5ec8, 32'shc0a03ee4, 32'shc0a11f9d, 32'shc0a200f2, 
               32'shc0a2e2e3, 32'shc0a3c571, 32'shc0a4a89b, 32'shc0a58c62, 32'shc0a670c4, 32'shc0a755c3, 32'shc0a83b5e, 32'shc0a92196, 
               32'shc0aa086a, 32'shc0aaefda, 32'shc0abd7e6, 32'shc0acc08f, 32'shc0ada9d4, 32'shc0ae93b5, 32'shc0af7e33, 32'shc0b0694c, 
               32'shc0b15502, 32'shc0b24154, 32'shc0b32e42, 32'shc0b41bcd, 32'shc0b509f3, 32'shc0b5f8b6, 32'shc0b6e815, 32'shc0b7d810, 
               32'shc0b8c8a7, 32'shc0b9b9da, 32'shc0baabaa, 32'shc0bb9e15, 32'shc0bc911d, 32'shc0bd84c1, 32'shc0be7901, 32'shc0bf6ddd, 
               32'shc0c06355, 32'shc0c15969, 32'shc0c25019, 32'shc0c34765, 32'shc0c43f4d, 32'shc0c537d1, 32'shc0c630f2, 32'shc0c72aae, 
               32'shc0c82506, 32'shc0c91ffa, 32'shc0ca1b8a, 32'shc0cb17b7, 32'shc0cc147f, 32'shc0cd11e3, 32'shc0ce0fe3, 32'shc0cf0e7f, 
               32'shc0d00db6, 32'shc0d10d8a, 32'shc0d20dfa, 32'shc0d30f05, 32'shc0d410ad, 32'shc0d512f0, 32'shc0d615cf, 32'shc0d7194a, 
               32'shc0d81d61, 32'shc0d92214, 32'shc0da2762, 32'shc0db2d4c, 32'shc0dc33d2, 32'shc0dd3af4, 32'shc0de42b2, 32'shc0df4b0b, 
               32'shc0e05401, 32'shc0e15d92, 32'shc0e267be, 32'shc0e37287, 32'shc0e47deb, 32'shc0e589eb, 32'shc0e69686, 32'shc0e7a3bd, 
               32'shc0e8b190, 32'shc0e9bfff, 32'shc0eacf09, 32'shc0ebdeaf, 32'shc0eceef1, 32'shc0edffce, 32'shc0ef1147, 32'shc0f0235b, 
               32'shc0f1360b, 32'shc0f24957, 32'shc0f35d3e, 32'shc0f471c1, 32'shc0f586df, 32'shc0f69c99, 32'shc0f7b2ee, 32'shc0f8c9df, 
               32'shc0f9e16b, 32'shc0faf993, 32'shc0fc1257, 32'shc0fd2bb6, 32'shc0fe45b0, 32'shc0ff6046, 32'shc1007b77, 32'shc1019744, 
               32'shc102b3ac, 32'shc103d0b0, 32'shc104ee4f, 32'shc1060c89, 32'shc1072b5f, 32'shc1084ad0, 32'shc1096add, 32'shc10a8b85, 
               32'shc10bacc8, 32'shc10ccea6, 32'shc10df120, 32'shc10f1435, 32'shc11037e6, 32'shc1115c32, 32'shc1128119, 32'shc113a69b, 
               32'shc114ccb9, 32'shc115f372, 32'shc1171ac6, 32'shc11842b5, 32'shc1196b3f, 32'shc11a9465, 32'shc11bbe26, 32'shc11ce882, 
               32'shc11e1379, 32'shc11f3f0c, 32'shc1206b39, 32'shc1219802, 32'shc122c566, 32'shc123f365, 32'shc12521ff, 32'shc1265134, 
               32'shc1278104, 32'shc128b16f, 32'shc129e276, 32'shc12b1417, 32'shc12c4653, 32'shc12d792b, 32'shc12eac9d, 32'shc12fe0ab, 
               32'shc1311553, 32'shc1324a96, 32'shc1338075, 32'shc134b6ee, 32'shc135ee02, 32'shc13725b1, 32'shc1385dfb, 32'shc13996e0, 
               32'shc13ad060, 32'shc13c0a7b, 32'shc13d4530, 32'shc13e8081, 32'shc13fbc6c, 32'shc140f8f2, 32'shc1423613, 32'shc14373cf, 
               32'shc144b225, 32'shc145f117, 32'shc14730a3, 32'shc14870ca, 32'shc149b18b, 32'shc14af2e8, 32'shc14c34df, 32'shc14d7771, 
               32'shc14eba9d, 32'shc14ffe64, 32'shc15142c6, 32'shc15287c3, 32'shc153cd5a, 32'shc155138c, 32'shc1565a58, 32'shc157a1bf, 
               32'shc158e9c1, 32'shc15a325d, 32'shc15b7b94, 32'shc15cc565, 32'shc15e0fd1, 32'shc15f5ad7, 32'shc160a678, 32'shc161f2b4, 
               32'shc1633f8a, 32'shc1648cfa, 32'shc165db05, 32'shc16729ab, 32'shc16878eb, 32'shc169c8c5, 32'shc16b193a, 32'shc16c6a49, 
               32'shc16dbbf3, 32'shc16f0e36, 32'shc1706115, 32'shc171b48e, 32'shc17308a1, 32'shc1745d4e, 32'shc175b296, 32'shc1770878, 
               32'shc1785ef4, 32'shc179b60b, 32'shc17b0dbb, 32'shc17c6607, 32'shc17dbeec, 32'shc17f186c, 32'shc1807285, 32'shc181cd3a, 
               32'shc1832888, 32'shc1848470, 32'shc185e0f3, 32'shc1873e10, 32'shc1889bc6, 32'shc189fa17, 32'shc18b5903, 32'shc18cb888, 
               32'shc18e18a7, 32'shc18f7961, 32'shc190dab4, 32'shc1923ca2, 32'shc1939f29, 32'shc195024b, 32'shc1966606, 32'shc197ca5c, 
               32'shc1992f4c, 32'shc19a94d5, 32'shc19bfaf9, 32'shc19d61b6, 32'shc19ec90d, 32'shc1a030ff, 32'shc1a1998a, 32'shc1a302af, 
               32'shc1a46c6e, 32'shc1a5d6c7, 32'shc1a741b9, 32'shc1a8ad46, 32'shc1aa196c, 32'shc1ab862c, 32'shc1acf386, 32'shc1ae617a, 
               32'shc1afd007, 32'shc1b13f2f, 32'shc1b2aef0, 32'shc1b41f4a, 32'shc1b5903f, 32'shc1b701cd, 32'shc1b873f5, 32'shc1b9e6b6, 
               32'shc1bb5a11, 32'shc1bcce06, 32'shc1be4294, 32'shc1bfb7bc, 32'shc1c12d7e, 32'shc1c2a3d9, 32'shc1c41ace, 32'shc1c5925c, 
               32'shc1c70a84, 32'shc1c88345, 32'shc1c9fca0, 32'shc1cb7694, 32'shc1ccf122, 32'shc1ce6c49, 32'shc1cfe80a, 32'shc1d16464, 
               32'shc1d2e158, 32'shc1d45ee5, 32'shc1d5dd0c, 32'shc1d75bcb, 32'shc1d8db25, 32'shc1da5b17, 32'shc1dbdba3, 32'shc1dd5cc8, 
               32'shc1dede87, 32'shc1e060df, 32'shc1e1e3d0, 32'shc1e3675a, 32'shc1e4eb7e, 32'shc1e6703b, 32'shc1e7f591, 32'shc1e97b80, 
               32'shc1eb0209, 32'shc1ec892b, 32'shc1ee10e5, 32'shc1ef9939, 32'shc1f12227, 32'shc1f2abad, 32'shc1f435cc, 32'shc1f5c085, 
               32'shc1f74bd6, 32'shc1f8d7c1, 32'shc1fa6445, 32'shc1fbf161, 32'shc1fd7f17, 32'shc1ff0d66, 32'shc2009c4e, 32'shc2022bce, 
               32'shc203bbe8, 32'shc2054c9b, 32'shc206dde6, 32'shc2086fca, 32'shc20a0248, 32'shc20b955e, 32'shc20d290d, 32'shc20ebd55, 
               32'shc2105236, 32'shc211e7af, 32'shc2137dc2, 32'shc215146d, 32'shc216abb1, 32'shc218438e, 32'shc219dc03, 32'shc21b7511, 
               32'shc21d0eb8, 32'shc21ea8f8, 32'shc22043d0, 32'shc221df41, 32'shc2237b4b, 32'shc22517ed, 32'shc226b528, 32'shc22852fb, 
               32'shc229f167, 32'shc22b906c, 32'shc22d3009, 32'shc22ed03f, 32'shc230710d, 32'shc2321274, 32'shc233b473, 32'shc235570b, 
               32'shc236fa3b, 32'shc2389e04, 32'shc23a4265, 32'shc23be75f, 32'shc23d8cf1, 32'shc23f331b, 32'shc240d9de, 32'shc2428139, 
               32'shc244292c, 32'shc245d1b8, 32'shc2477adc, 32'shc2492498, 32'shc24aceed, 32'shc24c79d9, 32'shc24e255e, 32'shc24fd17c, 
               32'shc2517e31, 32'shc2532b7f, 32'shc254d965, 32'shc25687e3, 32'shc25836f9, 32'shc259e6a7, 32'shc25b96ee, 32'shc25d47cc, 
               32'shc25ef943, 32'shc260ab51, 32'shc2625df8, 32'shc2641137, 32'shc265c50e, 32'shc267797c, 32'shc2692e83, 32'shc26ae422, 
               32'shc26c9a58, 32'shc26e5127, 32'shc270088e, 32'shc271c08c, 32'shc2737922, 32'shc2753250, 32'shc276ec16, 32'shc278a674, 
               32'shc27a616a, 32'shc27c1cf7, 32'shc27dd91c, 32'shc27f95d9, 32'shc281532e, 32'shc283111b, 32'shc284cf9f, 32'shc2868ebb, 
               32'shc2884e6e, 32'shc28a0eb9, 32'shc28bcf9c, 32'shc28d9117, 32'shc28f5329, 32'shc29115d3, 32'shc292d914, 32'shc2949ced, 
               32'shc296615d, 32'shc2982665, 32'shc299ec05, 32'shc29bb23c, 32'shc29d790a, 32'shc29f4070, 32'shc2a1086d, 32'shc2a2d102, 
               32'shc2a49a2e, 32'shc2a663f2, 32'shc2a82e4d, 32'shc2a9f93f, 32'shc2abc4c9, 32'shc2ad90ea, 32'shc2af5da2, 32'shc2b12af1, 
               32'shc2b2f8d8, 32'shc2b4c756, 32'shc2b6966c, 32'shc2b86618, 32'shc2ba365c, 32'shc2bc0737, 32'shc2bdd8a9, 32'shc2bfaab2, 
               32'shc2c17d52, 32'shc2c3508a, 32'shc2c52459, 32'shc2c6f8be, 32'shc2c8cdbb, 32'shc2caa34f, 32'shc2cc7979, 32'shc2ce503b, 
               32'shc2d02794, 32'shc2d1ff84, 32'shc2d3d80a, 32'shc2d5b128, 32'shc2d78add, 32'shc2d96528, 32'shc2db400a, 32'shc2dd1b84, 
               32'shc2def794, 32'shc2e0d43b, 32'shc2e2b178, 32'shc2e48f4d, 32'shc2e66db8, 32'shc2e84cba, 32'shc2ea2c53, 32'shc2ec0c82, 
               32'shc2eded49, 32'shc2efcea6, 32'shc2f1b099, 32'shc2f39323, 32'shc2f57644, 32'shc2f759fc, 32'shc2f93e4a, 32'shc2fb232e, 
               32'shc2fd08a9, 32'shc2feeebb, 32'shc300d563, 32'shc302bca2, 32'shc304a477, 32'shc3068ce3, 32'shc30875e5, 32'shc30a5f7e, 
               32'shc30c49ad, 32'shc30e3472, 32'shc3101fce, 32'shc3120bc0, 32'shc313f848, 32'shc315e567, 32'shc317d31c, 32'shc319c168, 
               32'shc31bb049, 32'shc31d9fc1, 32'shc31f8fcf, 32'shc3218073, 32'shc32371ae, 32'shc325637f, 32'shc32755e5, 32'shc32948e2, 
               32'shc32b3c75, 32'shc32d309e, 32'shc32f255e, 32'shc3311ab3, 32'shc333109e, 32'shc3350720, 32'shc336fe37, 32'shc338f5e4, 
               32'shc33aee27, 32'shc33ce701, 32'shc33ee070, 32'shc340da75, 32'shc342d510, 32'shc344d041, 32'shc346cc07, 32'shc348c864, 
               32'shc34ac556, 32'shc34cc2de, 32'shc34ec0fc, 32'shc350bfaf, 32'shc352bef9, 32'shc354bed8, 32'shc356bf4d, 32'shc358c057, 
               32'shc35ac1f7, 32'shc35cc42d, 32'shc35ec6f8, 32'shc360ca59, 32'shc362ce50, 32'shc364d2dc, 32'shc366d7fd, 32'shc368ddb4, 
               32'shc36ae401, 32'shc36ceae3, 32'shc36ef25b, 32'shc370fa68, 32'shc373030a, 32'shc3750c42, 32'shc377160f, 32'shc3792072, 
               32'shc37b2b6a, 32'shc37d36f7, 32'shc37f4319, 32'shc3814fd1, 32'shc3835d1e, 32'shc3856b01, 32'shc3877978, 32'shc3898885, 
               32'shc38b9827, 32'shc38da85e, 32'shc38fb92a, 32'shc391ca8c, 32'shc393dc82, 32'shc395ef0e, 32'shc398022f, 32'shc39a15e4, 
               32'shc39c2a2f, 32'shc39e3f0f, 32'shc3a05484, 32'shc3a26a8d, 32'shc3a4812c, 32'shc3a6985f, 32'shc3a8b028, 32'shc3aac885, 
               32'shc3ace178, 32'shc3aefaff, 32'shc3b1151b, 32'shc3b32fcb, 32'shc3b54b11, 32'shc3b766eb, 32'shc3b9835a, 32'shc3bba05e, 
               32'shc3bdbdf6, 32'shc3bfdc23, 32'shc3c1fae5, 32'shc3c41a3b, 32'shc3c63a26, 32'shc3c85aa6, 32'shc3ca7bba, 32'shc3cc9d63, 
               32'shc3cebfa0, 32'shc3d0e272, 32'shc3d305d8, 32'shc3d529d3, 32'shc3d74e62, 32'shc3d97386, 32'shc3db993e, 32'shc3ddbf8b, 
               32'shc3dfe66c, 32'shc3e20de1, 32'shc3e435ea, 32'shc3e65e88, 32'shc3e887bb, 32'shc3eab181, 32'shc3ecdbdc, 32'shc3ef06cb, 
               32'shc3f1324e, 32'shc3f35e65, 32'shc3f58b10, 32'shc3f7b850, 32'shc3f9e624, 32'shc3fc148c, 32'shc3fe4388, 32'shc4007318, 
               32'shc402a33c, 32'shc404d3f4, 32'shc4070540, 32'shc4093720, 32'shc40b6994, 32'shc40d9c9c, 32'shc40fd037, 32'shc4120467, 
               32'shc414392b, 32'shc4166e82, 32'shc418a46d, 32'shc41adaed, 32'shc41d11ff, 32'shc41f49a6, 32'shc42181e0, 32'shc423baae, 
               32'shc425f410, 32'shc4282e06, 32'shc42a688f, 32'shc42ca3ac, 32'shc42edf5c, 32'shc4311ba0, 32'shc4335877, 32'shc43595e3, 
               32'shc437d3e1, 32'shc43a1273, 32'shc43c5199, 32'shc43e9152, 32'shc440d19e, 32'shc443127e, 32'shc44553f2, 32'shc44795f8, 
               32'shc449d892, 32'shc44c1bc0, 32'shc44e5f80, 32'shc450a3d4, 32'shc452e8bc, 32'shc4552e36, 32'shc4577444, 32'shc459bae5, 
               32'shc45c0219, 32'shc45e49e0, 32'shc460923b, 32'shc462db28, 32'shc46524a9, 32'shc4676ebc, 32'shc469b963, 32'shc46c049d, 
               32'shc46e5069, 32'shc4709cc9, 32'shc472e9bc, 32'shc4753741, 32'shc477855a, 32'shc479d405, 32'shc47c2344, 32'shc47e7315, 
               32'shc480c379, 32'shc4831470, 32'shc48565f9, 32'shc487b815, 32'shc48a0ac4, 32'shc48c5e06, 32'shc48eb1db, 32'shc4910642, 
               32'shc4935b3c, 32'shc495b0c8, 32'shc49806e7, 32'shc49a5d98, 32'shc49cb4dd, 32'shc49f0cb3, 32'shc4a1651c, 32'shc4a3be18, 
               32'shc4a617a6, 32'shc4a871c7, 32'shc4aacc7a, 32'shc4ad27bf, 32'shc4af8397, 32'shc4b1e001, 32'shc4b43cfd, 32'shc4b69a8c, 
               32'shc4b8f8ad, 32'shc4bb5760, 32'shc4bdb6a6, 32'shc4c0167e, 32'shc4c276e8, 32'shc4c4d7e4, 32'shc4c73972, 32'shc4c99b92, 
               32'shc4cbfe45, 32'shc4ce6189, 32'shc4d0c560, 32'shc4d329c9, 32'shc4d58ec3, 32'shc4d7f450, 32'shc4da5a6f, 32'shc4dcc11f, 
               32'shc4df2862, 32'shc4e19036, 32'shc4e3f89c, 32'shc4e66194, 32'shc4e8cb1e, 32'shc4eb353a, 32'shc4ed9fe7, 32'shc4f00b27, 
               32'shc4f276f7, 32'shc4f4e35a, 32'shc4f7504e, 32'shc4f9bdd4, 32'shc4fc2bec, 32'shc4fe9a95, 32'shc50109d0, 32'shc503799d, 
               32'shc505e9fb, 32'shc5085aea, 32'shc50acc6b, 32'shc50d3e7d, 32'shc50fb121, 32'shc5122457, 32'shc514981d, 32'shc5170c75, 
               32'shc519815f, 32'shc51bf6da, 32'shc51e6ce6, 32'shc520e383, 32'shc5235ab2, 32'shc525d272, 32'shc5284ac3, 32'shc52ac3a5, 
               32'shc52d3d18, 32'shc52fb71d, 32'shc53231b3, 32'shc534acd9, 32'shc5372891, 32'shc539a4da, 32'shc53c21b4, 32'shc53e9f1f, 
               32'shc5411d1b, 32'shc5439ba8, 32'shc5461ac6, 32'shc5489a74, 32'shc54b1ab4, 32'shc54d9b84, 32'shc5501ce5, 32'shc5529ed7, 
               32'shc555215a, 32'shc557a46e, 32'shc55a2812, 32'shc55cac47, 32'shc55f310d, 32'shc561b663, 32'shc5643c4a, 32'shc566c2c2, 
               32'shc56949ca, 32'shc56bd163, 32'shc56e598c, 32'shc570e246, 32'shc5736b90, 32'shc575f56b, 32'shc5787fd6, 32'shc57b0ad1, 
               32'shc57d965d, 32'shc580227a, 32'shc582af26, 32'shc5853c63, 32'shc587ca31, 32'shc58a588e, 32'shc58ce77c, 32'shc58f76fa, 
               32'shc5920708, 32'shc59497a7, 32'shc59728d5, 32'shc599ba94, 32'shc59c4ce3, 32'shc59edfc2, 32'shc5a17330, 32'shc5a4072f, 
               32'shc5a69bbe, 32'shc5a930dd, 32'shc5abc68c, 32'shc5ae5ccb, 32'shc5b0f399, 32'shc5b38af8, 32'shc5b622e6, 32'shc5b8bb64, 
               32'shc5bb5472, 32'shc5bdee10, 32'shc5c0883d, 32'shc5c322fb, 32'shc5c5be47, 32'shc5c85a24, 32'shc5caf690, 32'shc5cd938c, 
               32'shc5d03118, 32'shc5d2cf33, 32'shc5d56ddd, 32'shc5d80d17, 32'shc5daace1, 32'shc5dd4d3a, 32'shc5dfee22, 32'shc5e28f9a, 
               32'shc5e531a1, 32'shc5e7d438, 32'shc5ea775e, 32'shc5ed1b13, 32'shc5efbf58, 32'shc5f2642c, 32'shc5f5098f, 32'shc5f7af81, 
               32'shc5fa5603, 32'shc5fcfd13, 32'shc5ffa4b3, 32'shc6024ce2, 32'shc604f5a0, 32'shc6079eed, 32'shc60a48c9, 32'shc60cf334, 
               32'shc60f9e2e, 32'shc61249b7, 32'shc614f5cf, 32'shc617a276, 32'shc61a4fac, 32'shc61cfd71, 32'shc61fabc4, 32'shc6225aa6, 
               32'shc6250a18, 32'shc627ba17, 32'shc62a6aa6, 32'shc62d1bc3, 32'shc62fcd6f, 32'shc6327faa, 32'shc6353273, 32'shc637e5ca, 
               32'shc63a99b1, 32'shc63d4e26, 32'shc6400329, 32'shc642b8bb, 32'shc6456edb, 32'shc648258a, 32'shc64adcc7, 32'shc64d9493, 
               32'shc6504ced, 32'shc65305d5, 32'shc655bf4c, 32'shc6587951, 32'shc65b33e4, 32'shc65def05, 32'shc660aab5, 32'shc66366f3, 
               32'shc66623be, 32'shc668e119, 32'shc66b9f01, 32'shc66e5d77, 32'shc6711c7b, 32'shc673dc0d, 32'shc6769c2e, 32'shc6795cdc, 
               32'shc67c1e18, 32'shc67edfe2, 32'shc681a23a, 32'shc6846520, 32'shc6872894, 32'shc689ec95, 32'shc68cb124, 32'shc68f7641, 
               32'shc6923bec, 32'shc6950224, 32'shc697c8eb, 32'shc69a903e, 32'shc69d5820, 32'shc6a0208f, 32'shc6a2e98b, 32'shc6a5b315, 
               32'shc6a87d2d, 32'shc6ab47d2, 32'shc6ae1304, 32'shc6b0dec4, 32'shc6b3ab12, 32'shc6b677ec, 32'shc6b94554, 32'shc6bc134a, 
               32'shc6bee1cd, 32'shc6c1b0dd, 32'shc6c4807a, 32'shc6c750a4, 32'shc6ca215c, 32'shc6ccf2a1, 32'shc6cfc472, 32'shc6d296d1, 
               32'shc6d569be, 32'shc6d83d37, 32'shc6db113d, 32'shc6dde5d0, 32'shc6e0baf0, 32'shc6e3909d, 32'shc6e666d7, 32'shc6e93d9e, 
               32'shc6ec14f2, 32'shc6eeecd3, 32'shc6f1c540, 32'shc6f49e3a, 32'shc6f777c1, 32'shc6fa51d5, 32'shc6fd2c75, 32'shc70007a2, 
               32'shc702e35c, 32'shc705bfa2, 32'shc7089c75, 32'shc70b79d4, 32'shc70e57c0, 32'shc7113639, 32'shc714153e, 32'shc716f4cf, 
               32'shc719d4ed, 32'shc71cb597, 32'shc71f96ce, 32'shc7227890, 32'shc7255ae0, 32'shc7283dbb, 32'shc72b2123, 32'shc72e0517, 
               32'shc730e997, 32'shc733cea3, 32'shc736b43c, 32'shc7399a60, 32'shc73c8111, 32'shc73f684e, 32'shc7425016, 32'shc745386b, 
               32'shc748214c, 32'shc74b0ab9, 32'shc74df4b1, 32'shc750df36, 32'shc753ca46, 32'shc756b5e2, 32'shc759a20a, 32'shc75c8ebe, 
               32'shc75f7bfe, 32'shc76269c9, 32'shc7655820, 32'shc7684702, 32'shc76b3671, 32'shc76e266b, 32'shc77116f0, 32'shc7740801, 
               32'shc776f99d, 32'shc779ebc5, 32'shc77cde79, 32'shc77fd1b8, 32'shc782c582, 32'shc785b9d8, 32'shc788aeb9, 32'shc78ba425, 
               32'shc78e9a1d, 32'shc79190a0, 32'shc79487ae, 32'shc7977f48, 32'shc79a776c, 32'shc79d701c, 32'shc7a06957, 32'shc7a3631d, 
               32'shc7a65d6e, 32'shc7a9584a, 32'shc7ac53b1, 32'shc7af4fa3, 32'shc7b24c20, 32'shc7b54928, 32'shc7b846ba, 32'shc7bb44d8, 
               32'shc7be4381, 32'shc7c142b4, 32'shc7c44272, 32'shc7c742bb, 32'shc7ca438f, 32'shc7cd44ed, 32'shc7d046d6, 32'shc7d34949, 
               32'shc7d64c47, 32'shc7d94fd0, 32'shc7dc53e3, 32'shc7df5881, 32'shc7e25daa, 32'shc7e5635c, 32'shc7e8699a, 32'shc7eb7061, 
               32'shc7ee77b3, 32'shc7f17f8f, 32'shc7f487f6, 32'shc7f790e7, 32'shc7fa9a62, 32'shc7fda468, 32'shc800aef7, 32'shc803ba11, 
               32'shc806c5b5, 32'shc809d1e3, 32'shc80cde9b, 32'shc80febdd, 32'shc812f9a9, 32'shc81607ff, 32'shc81916df, 32'shc81c2649, 
               32'shc81f363d, 32'shc82246bb, 32'shc82557c3, 32'shc8286954, 32'shc82b7b70, 32'shc82e8e15, 32'shc831a143, 32'shc834b4fc, 
               32'shc837c93e, 32'shc83ade0a, 32'shc83df35f, 32'shc841093e, 32'shc8441fa6, 32'shc8473698, 32'shc84a4e14, 32'shc84d6619, 
               32'shc8507ea7, 32'shc85397bf, 32'shc856b160, 32'shc859cb8a, 32'shc85ce63e, 32'shc860017b, 32'shc8631d42, 32'shc8663991, 
               32'shc869566a, 32'shc86c73cc, 32'shc86f91b7, 32'shc872b02b, 32'shc875cf28, 32'shc878eeae, 32'shc87c0ebd, 32'shc87f2f56, 
               32'shc8825077, 32'shc8857221, 32'shc8889454, 32'shc88bb710, 32'shc88eda54, 32'shc891fe22, 32'shc8952278, 32'shc8984757, 
               32'shc89b6cbf, 32'shc89e92af, 32'shc8a1b928, 32'shc8a4e029, 32'shc8a807b4, 32'shc8ab2fc6, 32'shc8ae5862, 32'shc8b18185, 
               32'shc8b4ab32, 32'shc8b7d566, 32'shc8bb0023, 32'shc8be2b69, 32'shc8c15736, 32'shc8c4838d, 32'shc8c7b06b, 32'shc8caddd1, 
               32'shc8ce0bc0, 32'shc8d13a37, 32'shc8d46936, 32'shc8d798be, 32'shc8dac8cd, 32'shc8ddf965, 32'shc8e12a84, 32'shc8e45c2c, 
               32'shc8e78e5b, 32'shc8eac112, 32'shc8edf452, 32'shc8f12819, 32'shc8f45c68, 32'shc8f7913f, 32'shc8fac69e, 32'shc8fdfc84, 
               32'shc90132f2, 32'shc90469e8, 32'shc907a166, 32'shc90ad96b, 32'shc90e11f7, 32'shc9114b0c, 32'shc91484a8, 32'shc917becb, 
               32'shc91af976, 32'shc91e34a8, 32'shc9217062, 32'shc924aca3, 32'shc927e96b, 32'shc92b26bb, 32'shc92e6492, 32'shc931a2f0, 
               32'shc934e1d6, 32'shc9382143, 32'shc93b6137, 32'shc93ea1b2, 32'shc941e2b4, 32'shc945243d, 32'shc948664d, 32'shc94ba8e5, 
               32'shc94eec03, 32'shc9522fa8, 32'shc95573d4, 32'shc958b887, 32'shc95bfdc1, 32'shc95f4382, 32'shc96289c9, 32'shc965d097, 
               32'shc96917ec, 32'shc96c5fc8, 32'shc96fa82a, 32'shc972f113, 32'shc9763a83, 32'shc9798479, 32'shc97ccef5, 32'shc98019f8, 
               32'shc9836582, 32'shc986b192, 32'shc989fe29, 32'shc98d4b45, 32'shc99098e9, 32'shc993e712, 32'shc99735c2, 32'shc99a84f8, 
               32'shc99dd4b4, 32'shc9a124f7, 32'shc9a475bf, 32'shc9a7c70e, 32'shc9ab18e3, 32'shc9ae6b3d, 32'shc9b1be1e, 32'shc9b51185, 
               32'shc9b86572, 32'shc9bbb9e5, 32'shc9bf0edd, 32'shc9c2645c, 32'shc9c5ba60, 32'shc9c910ea, 32'shc9cc67fa, 32'shc9cfbf90, 
               32'shc9d317ab, 32'shc9d6704c, 32'shc9d9c973, 32'shc9dd231f, 32'shc9e07d51, 32'shc9e3d809, 32'shc9e73346, 32'shc9ea8f08, 
               32'shc9edeb50, 32'shc9f1481d, 32'shc9f4a570, 32'shc9f80348, 32'shc9fb61a5, 32'shc9fec088, 32'shca021fef, 32'shca057fdd, 
               32'shca08e04f, 32'shca0c4146, 32'shca0fa2c3, 32'shca1304c4, 32'shca16674b, 32'shca19ca57, 32'shca1d2de7, 32'shca2091fd, 
               32'shca23f698, 32'shca275bb7, 32'shca2ac15b, 32'shca2e2784, 32'shca318e32, 32'shca34f565, 32'shca385d1d, 32'shca3bc559, 
               32'shca3f2e19, 32'shca42975f, 32'shca460129, 32'shca496b77, 32'shca4cd64b, 32'shca5041a2, 32'shca53ad7e, 32'shca5719df, 
               32'shca5a86c4, 32'shca5df42d, 32'shca61621b, 32'shca64d08d, 32'shca683f83, 32'shca6baefd, 32'shca6f1efc, 32'shca728f7f, 
               32'shca760086, 32'shca797211, 32'shca7ce420, 32'shca8056b3, 32'shca83c9ca, 32'shca873d65, 32'shca8ab184, 32'shca8e2627, 
               32'shca919b4e, 32'shca9510f8, 32'shca988727, 32'shca9bfdd9, 32'shca9f750f, 32'shcaa2ecc9, 32'shcaa66506, 32'shcaa9ddc7, 
               32'shcaad570c, 32'shcab0d0d4, 32'shcab44b1f, 32'shcab7c5ef, 32'shcabb4141, 32'shcabebd17, 32'shcac23971, 32'shcac5b64e, 
               32'shcac933ae, 32'shcaccb191, 32'shcad02ff8, 32'shcad3aee2, 32'shcad72e4f, 32'shcadaae40, 32'shcade2eb3, 32'shcae1afaa, 
               32'shcae53123, 32'shcae8b320, 32'shcaec35a0, 32'shcaefb8a2, 32'shcaf33c28, 32'shcaf6c030, 32'shcafa44bc, 32'shcafdc9ca, 
               32'shcb014f5b, 32'shcb04d56e, 32'shcb085c05, 32'shcb0be31e, 32'shcb0f6aba, 32'shcb12f2d8, 32'shcb167b79, 32'shcb1a049d, 
               32'shcb1d8e43, 32'shcb21186b, 32'shcb24a316, 32'shcb282e44, 32'shcb2bb9f4, 32'shcb2f4626, 32'shcb32d2da, 32'shcb366011, 
               32'shcb39edca, 32'shcb3d7c05, 32'shcb410ac3, 32'shcb449a02, 32'shcb4829c4, 32'shcb4bba08, 32'shcb4f4acd, 32'shcb52dc15, 
               32'shcb566ddf, 32'shcb5a002b, 32'shcb5d92f8, 32'shcb612648, 32'shcb64ba19, 32'shcb684e6c, 32'shcb6be341, 32'shcb6f7898, 
               32'shcb730e70, 32'shcb76a4ca, 32'shcb7a3ba5, 32'shcb7dd303, 32'shcb816ae1, 32'shcb850342, 32'shcb889c23, 32'shcb8c3587, 
               32'shcb8fcf6b, 32'shcb9369d1, 32'shcb9704b9, 32'shcb9aa021, 32'shcb9e3c0b, 32'shcba1d877, 32'shcba57563, 32'shcba912d1, 
               32'shcbacb0bf, 32'shcbb04f2f, 32'shcbb3ee20, 32'shcbb78d92, 32'shcbbb2d85, 32'shcbbecdf9, 32'shcbc26eee, 32'shcbc61064, 
               32'shcbc9b25a, 32'shcbcd54d2, 32'shcbd0f7ca, 32'shcbd49b43, 32'shcbd83f3d, 32'shcbdbe3b7, 32'shcbdf88b3, 32'shcbe32e2e, 
               32'shcbe6d42b, 32'shcbea7aa7, 32'shcbee21a5, 32'shcbf1c923, 32'shcbf57121, 32'shcbf919a0, 32'shcbfcc29f, 32'shcc006c1e, 
               32'shcc04161e, 32'shcc07c09e, 32'shcc0b6b9e, 32'shcc0f171e, 32'shcc12c31f, 32'shcc166f9f, 32'shcc1a1ca0, 32'shcc1dca21, 
               32'shcc217822, 32'shcc2526a2, 32'shcc28d5a3, 32'shcc2c8524, 32'shcc303524, 32'shcc33e5a5, 32'shcc3796a5, 32'shcc3b4825, 
               32'shcc3efa25, 32'shcc42aca4, 32'shcc465fa3, 32'shcc4a1322, 32'shcc4dc720, 32'shcc517b9e, 32'shcc55309b, 32'shcc58e618, 
               32'shcc5c9c14, 32'shcc605290, 32'shcc64098b, 32'shcc67c105, 32'shcc6b78ff, 32'shcc6f3178, 32'shcc72ea70, 32'shcc76a3e8, 
               32'shcc7a5dde, 32'shcc7e1854, 32'shcc81d349, 32'shcc858ebc, 32'shcc894aaf, 32'shcc8d0721, 32'shcc90c412, 32'shcc948182, 
               32'shcc983f70, 32'shcc9bfddd, 32'shcc9fbcca, 32'shcca37c35, 32'shcca73c1e, 32'shccaafc87, 32'shccaebd6e, 32'shccb27ed3, 
               32'shccb640b8, 32'shccba031a, 32'shccbdc5fc, 32'shccc1895c, 32'shccc54d3a, 32'shccc91196, 32'shccccd671, 32'shccd09bcb, 
               32'shccd461a2, 32'shccd827f8, 32'shccdbeecc, 32'shccdfb61f, 32'shcce37def, 32'shcce7463e, 32'shcceb0f0a, 32'shcceed855, 
               32'shccf2a21d, 32'shccf66c64, 32'shccfa3729, 32'shccfe026b, 32'shcd01ce2b, 32'shcd059a6a, 32'shcd096725, 32'shcd0d345f, 
               32'shcd110216, 32'shcd14d04b, 32'shcd189efe, 32'shcd1c6e2e, 32'shcd203ddc, 32'shcd240e08, 32'shcd27deb0, 32'shcd2bafd7, 
               32'shcd2f817b, 32'shcd33539c, 32'shcd37263a, 32'shcd3af956, 32'shcd3eccef, 32'shcd42a105, 32'shcd467599, 32'shcd4a4aa9, 
               32'shcd4e2037, 32'shcd51f642, 32'shcd55ccca, 32'shcd59a3ce, 32'shcd5d7b50, 32'shcd61534f, 32'shcd652bcb, 32'shcd6904c3, 
               32'shcd6cde39, 32'shcd70b82b, 32'shcd74929a, 32'shcd786d85, 32'shcd7c48ee, 32'shcd8024d3, 32'shcd840134, 32'shcd87de12, 
               32'shcd8bbb6d, 32'shcd8f9944, 32'shcd937798, 32'shcd975668, 32'shcd9b35b4, 32'shcd9f157d, 32'shcda2f5c2, 32'shcda6d683, 
               32'shcdaab7c0, 32'shcdae997a, 32'shcdb27bb0, 32'shcdb65e62, 32'shcdba4190, 32'shcdbe253a, 32'shcdc20960, 32'shcdc5ee02, 
               32'shcdc9d320, 32'shcdcdb8ba, 32'shcdd19ed0, 32'shcdd58562, 32'shcdd96c6f, 32'shcddd53f8, 32'shcde13bfd, 32'shcde5247d, 
               32'shcde90d79, 32'shcdecf6f1, 32'shcdf0e0e4, 32'shcdf4cb53, 32'shcdf8b63d, 32'shcdfca1a3, 32'shce008d84, 32'shce0479e0, 
               32'shce0866b8, 32'shce0c540b, 32'shce1041d9, 32'shce143023, 32'shce181ee8, 32'shce1c0e28, 32'shce1ffde2, 32'shce23ee18, 
               32'shce27dec9, 32'shce2bcff5, 32'shce2fc19c, 32'shce33b3be, 32'shce37a65b, 32'shce3b9973, 32'shce3f8d05, 32'shce438112, 
               32'shce47759a, 32'shce4b6a9c, 32'shce4f6019, 32'shce535611, 32'shce574c84, 32'shce5b4370, 32'shce5f3ad8, 32'shce6332ba, 
               32'shce672b16, 32'shce6b23ec, 32'shce6f1d3d, 32'shce731709, 32'shce77114e, 32'shce7b0c0e, 32'shce7f0748, 32'shce8302fc, 
               32'shce86ff2a, 32'shce8afbd2, 32'shce8ef8f4, 32'shce92f691, 32'shce96f4a7, 32'shce9af337, 32'shce9ef241, 32'shcea2f1c5, 
               32'shcea6f1c2, 32'shceaaf23a, 32'shceaef32b, 32'shceb2f496, 32'shceb6f67a, 32'shcebaf8d8, 32'shcebefbb0, 32'shcec2ff01, 
               32'shcec702cb, 32'shcecb070f, 32'shcecf0bcd, 32'shced31104, 32'shced716b4, 32'shcedb1cde, 32'shcedf2380, 32'shcee32a9c, 
               32'shcee73231, 32'shceeb3a40, 32'shceef42c7, 32'shcef34bc8, 32'shcef75541, 32'shcefb5f34, 32'shceff699f, 32'shcf037483, 
               32'shcf077fe1, 32'shcf0b8bb7, 32'shcf0f9805, 32'shcf13a4cd, 32'shcf17b20d, 32'shcf1bbfc6, 32'shcf1fcdf8, 32'shcf23dca2, 
               32'shcf27ebc5, 32'shcf2bfb60, 32'shcf300b74, 32'shcf341c00, 32'shcf382d05, 32'shcf3c3e82, 32'shcf405077, 32'shcf4462e4, 
               32'shcf4875ca, 32'shcf4c8928, 32'shcf509cfe, 32'shcf54b14d, 32'shcf58c613, 32'shcf5cdb51, 32'shcf60f108, 32'shcf650736, 
               32'shcf691ddd, 32'shcf6d34fb, 32'shcf714c91, 32'shcf75649f, 32'shcf797d24, 32'shcf7d9622, 32'shcf81af97, 32'shcf85c984, 
               32'shcf89e3e8, 32'shcf8dfec4, 32'shcf921a17, 32'shcf9635e2, 32'shcf9a5225, 32'shcf9e6edf, 32'shcfa28c10, 32'shcfa6a9b8, 
               32'shcfaac7d8, 32'shcfaee66f, 32'shcfb3057d, 32'shcfb72503, 32'shcfbb4500, 32'shcfbf6573, 32'shcfc3865e, 32'shcfc7a7c0, 
               32'shcfcbc999, 32'shcfcfebe8, 32'shcfd40eaf, 32'shcfd831ec, 32'shcfdc55a1, 32'shcfe079cc, 32'shcfe49e6d, 32'shcfe8c386, 
               32'shcfece915, 32'shcff10f1b, 32'shcff53597, 32'shcff95c8a, 32'shcffd83f4, 32'shd001abd3, 32'shd005d42a, 32'shd009fcf6, 
               32'shd00e2639, 32'shd0124ff3, 32'shd0167a22, 32'shd01aa4c8, 32'shd01ecfe4, 32'shd022fb76, 32'shd027277e, 32'shd02b53fc, 
               32'shd02f80f1, 32'shd033ae5b, 32'shd037dc3b, 32'shd03c0a91, 32'shd040395d, 32'shd044689f, 32'shd0489856, 32'shd04cc884, 
               32'shd050f926, 32'shd0552a3f, 32'shd0595bcd, 32'shd05d8dd1, 32'shd061c04a, 32'shd065f339, 32'shd06a269d, 32'shd06e5a77, 
               32'shd0728ec6, 32'shd076c38b, 32'shd07af8c4, 32'shd07f2e73, 32'shd0836497, 32'shd0879b31, 32'shd08bd23f, 32'shd09009c3, 
               32'shd09441bb, 32'shd0987a29, 32'shd09cb30b, 32'shd0a0ec63, 32'shd0a5262f, 32'shd0a96070, 32'shd0ad9b26, 32'shd0b1d651, 
               32'shd0b611f1, 32'shd0ba4e05, 32'shd0be8a8d, 32'shd0c2c78b, 32'shd0c704fd, 32'shd0cb42e3, 32'shd0cf813e, 32'shd0d3c00e, 
               32'shd0d7ff51, 32'shd0dc3f0a, 32'shd0e07f36, 32'shd0e4bfd7, 32'shd0e900ec, 32'shd0ed4275, 32'shd0f18472, 32'shd0f5c6e3, 
               32'shd0fa09c9, 32'shd0fe4d22, 32'shd10290f0, 32'shd106d531, 32'shd10b19e7, 32'shd10f5f10, 32'shd113a4ad, 32'shd117eabd, 
               32'shd11c3142, 32'shd120783a, 32'shd124bfa6, 32'shd1290786, 32'shd12d4fd9, 32'shd131989f, 32'shd135e1d9, 32'shd13a2b87, 
               32'shd13e75a8, 32'shd142c03c, 32'shd1470b44, 32'shd14b56be, 32'shd14fa2ad, 32'shd153ef0e, 32'shd1583be2, 32'shd15c892a, 
               32'shd160d6e5, 32'shd1652512, 32'shd16973b3, 32'shd16dc2c7, 32'shd172124d, 32'shd1766247, 32'shd17ab2b3, 32'shd17f0392, 
               32'shd18354e4, 32'shd187a6a8, 32'shd18bf8e0, 32'shd1904b89, 32'shd1949ea6, 32'shd198f235, 32'shd19d4636, 32'shd1a19aaa, 
               32'shd1a5ef90, 32'shd1aa44e9, 32'shd1ae9ab4, 32'shd1b2f0f1, 32'shd1b747a0, 32'shd1bb9ec2, 32'shd1bff656, 32'shd1c44e5c, 
               32'shd1c8a6d4, 32'shd1ccffbe, 32'shd1d1591a, 32'shd1d5b2e8, 32'shd1da0d28, 32'shd1de67da, 32'shd1e2c2fd, 32'shd1e71e93, 
               32'shd1eb7a9a, 32'shd1efd713, 32'shd1f433fd, 32'shd1f89159, 32'shd1fcef27, 32'shd2014d66, 32'shd205ac17, 32'shd20a0b39, 
               32'shd20e6acc, 32'shd212cad1, 32'shd2172b48, 32'shd21b8c2f, 32'shd21fed88, 32'shd2244f52, 32'shd228b18d, 32'shd22d1439, 
               32'shd2317756, 32'shd235dae4, 32'shd23a3ee4, 32'shd23ea354, 32'shd2430835, 32'shd2476d87, 32'shd24bd34a, 32'shd250397d, 
               32'shd254a021, 32'shd2590736, 32'shd25d6ebc, 32'shd261d6b2, 32'shd2663f19, 32'shd26aa7f0, 32'shd26f1138, 32'shd2737af0, 
               32'shd277e518, 32'shd27c4fb1, 32'shd280babb, 32'shd2852634, 32'shd289921e, 32'shd28dfe77, 32'shd2926b41, 32'shd296d87c, 
               32'shd29b4626, 32'shd29fb440, 32'shd2a422ca, 32'shd2a891c4, 32'shd2ad012e, 32'shd2b17107, 32'shd2b5e151, 32'shd2ba520a, 
               32'shd2bec333, 32'shd2c334cc, 32'shd2c7a6d4, 32'shd2cc194c, 32'shd2d08c33, 32'shd2d4ff8a, 32'shd2d97350, 32'shd2dde786, 
               32'shd2e25c2b, 32'shd2e6d13f, 32'shd2eb46c3, 32'shd2efbcb6, 32'shd2f43318, 32'shd2f8a9e9, 32'shd2fd2129, 32'shd30198d8, 
               32'shd30610f7, 32'shd30a8984, 32'shd30f0280, 32'shd3137bec, 32'shd317f5c6, 32'shd31c700f, 32'shd320eac6, 32'shd32565ec, 
               32'shd329e181, 32'shd32e5d85, 32'shd332d9f7, 32'shd33756d8, 32'shd33bd427, 32'shd34051e5, 32'shd344d011, 32'shd3494eab, 
               32'shd34dcdb4, 32'shd3524d2b, 32'shd356cd11, 32'shd35b4d64, 32'shd35fce26, 32'shd3644f55, 32'shd368d0f3, 32'shd36d52ff, 
               32'shd371d579, 32'shd3765861, 32'shd37adbb6, 32'shd37f5f7a, 32'shd383e3ab, 32'shd388684a, 32'shd38ced57, 32'shd39172d2, 
               32'shd395f8ba, 32'shd39a7f0f, 32'shd39f05d3, 32'shd3a38d03, 32'shd3a814a2, 32'shd3ac9cad, 32'shd3b12526, 32'shd3b5ae0d, 
               32'shd3ba3760, 32'shd3bec121, 32'shd3c34b4f, 32'shd3c7d5ea, 32'shd3cc60f2, 32'shd3d0ec68, 32'shd3d5784a, 32'shd3da049a, 
               32'shd3de9156, 32'shd3e31e7f, 32'shd3e7ac15, 32'shd3ec3a18, 32'shd3f0c887, 32'shd3f55764, 32'shd3f9e6ad, 32'shd3fe7662, 
               32'shd4030684, 32'shd4079713, 32'shd40c280e, 32'shd410b976, 32'shd4154b4a, 32'shd419dd8a, 32'shd41e7037, 32'shd4230350, 
               32'shd42796d5, 32'shd42c2ac6, 32'shd430bf24, 32'shd43553ee, 32'shd439e923, 32'shd43e7ec5, 32'shd44314d3, 32'shd447ab4c, 
               32'shd44c4232, 32'shd450d983, 32'shd4557140, 32'shd45a0969, 32'shd45ea1fd, 32'shd4633afd, 32'shd467d469, 32'shd46c6e40, 
               32'shd4710883, 32'shd475a332, 32'shd47a3e4b, 32'shd47ed9d0, 32'shd48375c1, 32'shd488121d, 32'shd48caee4, 32'shd4914c16, 
               32'shd495e9b3, 32'shd49a87bc, 32'shd49f2630, 32'shd4a3c50e, 32'shd4a86458, 32'shd4ad040c, 32'shd4b1a42c, 32'shd4b644b6, 
               32'shd4bae5ab, 32'shd4bf870b, 32'shd4c428d6, 32'shd4c8cb0b, 32'shd4cd6dab, 32'shd4d210b5, 32'shd4d6b42b, 32'shd4db580a, 
               32'shd4dffc54, 32'shd4e4a108, 32'shd4e94627, 32'shd4edebb0, 32'shd4f291a4, 32'shd4f73801, 32'shd4fbdec9, 32'shd50085fb, 
               32'shd5052d97, 32'shd509d59d, 32'shd50e7e0d, 32'shd51326e7, 32'shd517d02b, 32'shd51c79d9, 32'shd52123f0, 32'shd525ce72, 
               32'shd52a795d, 32'shd52f24b2, 32'shd533d070, 32'shd5387c98, 32'shd53d292a, 32'shd541d625, 32'shd5468389, 32'shd54b3157, 
               32'shd54fdf8f, 32'shd5548e30, 32'shd5593d3a, 32'shd55decad, 32'shd5629c89, 32'shd5674ccf, 32'shd56bfd7d, 32'shd570ae95, 
               32'shd5756016, 32'shd57a1200, 32'shd57ec452, 32'shd583770e, 32'shd5882a32, 32'shd58cddbf, 32'shd59191b5, 32'shd5964614, 
               32'shd59afadb, 32'shd59fb00b, 32'shd5a465a3, 32'shd5a91ba4, 32'shd5add20d, 32'shd5b288df, 32'shd5b74019, 32'shd5bbf7bc, 
               32'shd5c0afc6, 32'shd5c56839, 32'shd5ca2115, 32'shd5ceda58, 32'shd5d39403, 32'shd5d84e17, 32'shd5dd0892, 32'shd5e1c376, 
               32'shd5e67ec1, 32'shd5eb3a75, 32'shd5eff690, 32'shd5f4b313, 32'shd5f96ffd, 32'shd5fe2d50, 32'shd602eb0a, 32'shd607a92b, 
               32'shd60c67b4, 32'shd61126a5, 32'shd615e5fd, 32'shd61aa5bd, 32'shd61f65e4, 32'shd6242672, 32'shd628e767, 32'shd62da8c4, 
               32'shd6326a88, 32'shd6372cb3, 32'shd63bef46, 32'shd640b23f, 32'shd645759f, 32'shd64a3966, 32'shd64efd94, 32'shd653c229, 
               32'shd6588725, 32'shd65d4c88, 32'shd6621251, 32'shd666d881, 32'shd66b9f18, 32'shd6706615, 32'shd6752d79, 32'shd679f543, 
               32'shd67ebd74, 32'shd683860b, 32'shd6884f09, 32'shd68d186d, 32'shd691e237, 32'shd696ac67, 32'shd69b76fe, 32'shd6a041fa, 
               32'shd6a50d5d, 32'shd6a9d926, 32'shd6aea555, 32'shd6b371ea, 32'shd6b83ee4, 32'shd6bd0c45, 32'shd6c1da0b, 32'shd6c6a837, 
               32'shd6cb76c9, 32'shd6d045c0, 32'shd6d5151d, 32'shd6d9e4e0, 32'shd6deb508, 32'shd6e38596, 32'shd6e85689, 32'shd6ed27e1, 
               32'shd6f1f99f, 32'shd6f6cbc2, 32'shd6fb9e4b, 32'shd7007138, 32'shd705448b, 32'shd70a1843, 32'shd70eec60, 32'shd713c0e2, 
               32'shd71895c9, 32'shd71d6b15, 32'shd72240c5, 32'shd72716db, 32'shd72bed55, 32'shd730c434, 32'shd7359b78, 32'shd73a7321, 
               32'shd73f4b2e, 32'shd744239f, 32'shd748fc75, 32'shd74dd5b0, 32'shd752af4f, 32'shd7578952, 32'shd75c63ba, 32'shd7613e86, 
               32'shd76619b6, 32'shd76af54a, 32'shd76fd143, 32'shd774ad9f, 32'shd7798a60, 32'shd77e6784, 32'shd783450d, 32'shd78822f9, 
               32'shd78d014a, 32'shd791dffe, 32'shd796bf16, 32'shd79b9e91, 32'shd7a07e70, 32'shd7a55eb3, 32'shd7aa3f5a, 32'shd7af2063, 
               32'shd7b401d1, 32'shd7b8e3a2, 32'shd7bdc5d6, 32'shd7c2a86d, 32'shd7c78b68, 32'shd7cc6ec6, 32'shd7d15288, 32'shd7d636ac, 
               32'shd7db1b34, 32'shd7e0001e, 32'shd7e4e56c, 32'shd7e9cb1c, 32'shd7eeb130, 32'shd7f397a6, 32'shd7f87e7f, 32'shd7fd65bb, 
               32'shd8024d59, 32'shd807355b, 32'shd80c1dbf, 32'shd8110685, 32'shd815efae, 32'shd81ad93a, 32'shd81fc328, 32'shd824ad78, 
               32'shd829982b, 32'shd82e833f, 32'shd8336eb7, 32'shd8385a90, 32'shd83d46cc, 32'shd8423369, 32'shd8472069, 32'shd84c0dcb, 
               32'shd850fb8e, 32'shd855e9b4, 32'shd85ad83c, 32'shd85fc725, 32'shd864b670, 32'shd869a61d, 32'shd86e962b, 32'shd873869b, 
               32'shd878776d, 32'shd87d68a0, 32'shd8825a35, 32'shd8874c2b, 32'shd88c3e83, 32'shd891313b, 32'shd8962456, 32'shd89b17d1, 
               32'shd8a00bae, 32'shd8a4ffec, 32'shd8a9f48a, 32'shd8aee98a, 32'shd8b3deeb, 32'shd8b8d4ad, 32'shd8bdcad0, 32'shd8c2c154, 
               32'shd8c7b838, 32'shd8ccaf7e, 32'shd8d1a724, 32'shd8d69f2a, 32'shd8db9792, 32'shd8e0905a, 32'shd8e58982, 32'shd8ea830b, 
               32'shd8ef7cf4, 32'shd8f4773e, 32'shd8f971e8, 32'shd8fe6cf2, 32'shd903685d, 32'shd9086428, 32'shd90d6053, 32'shd9125cde, 
               32'shd91759c9, 32'shd91c5714, 32'shd92154bf, 32'shd92652ca, 32'shd92b5135, 32'shd9305000, 32'shd9354f2a, 32'shd93a4eb4, 
               32'shd93f4e9e, 32'shd9444ee7, 32'shd9494f90, 32'shd94e5099, 32'shd9535201, 32'shd95853c8, 32'shd95d55ef, 32'shd9625875, 
               32'shd9675b5a, 32'shd96c5e9f, 32'shd9716243, 32'shd9766646, 32'shd97b6aa8, 32'shd9806f69, 32'shd9857489, 32'shd98a7a08, 
               32'shd98f7fe6, 32'shd9948623, 32'shd9998cbe, 32'shd99e93b8, 32'shd9a39b11, 32'shd9a8a2c9, 32'shd9adaadf, 32'shd9b2b354, 
               32'shd9b7bc27, 32'shd9bcc559, 32'shd9c1cee9, 32'shd9c6d8d8, 32'shd9cbe325, 32'shd9d0edd0, 32'shd9d5f8d9, 32'shd9db0441, 
               32'shd9e01006, 32'shd9e51c2a, 32'shd9ea28ac, 32'shd9ef358b, 32'shd9f442c9, 32'shd9f95064, 32'shd9fe5e5e, 32'shda036cb5, 
               32'shda087b69, 32'shda0d8a7c, 32'shda1299ec, 32'shda17a9ba, 32'shda1cb9e5, 32'shda21ca6e, 32'shda26db54, 32'shda2bec97, 
               32'shda30fe38, 32'shda361036, 32'shda3b2292, 32'shda40354a, 32'shda454860, 32'shda4a5bd3, 32'shda4f6fa3, 32'shda5483d0, 
               32'shda599859, 32'shda5ead40, 32'shda63c284, 32'shda68d824, 32'shda6dee21, 32'shda73047b, 32'shda781b31, 32'shda7d3244, 
               32'shda8249b4, 32'shda876180, 32'shda8c79a9, 32'shda91922e, 32'shda96ab0f, 32'shda9bc44d, 32'shdaa0dde7, 32'shdaa5f7dd, 
               32'shdaab122f, 32'shdab02cdd, 32'shdab547e8, 32'shdaba634e, 32'shdabf7f11, 32'shdac49b2f, 32'shdac9b7a9, 32'shdaced47f, 
               32'shdad3f1b1, 32'shdad90f3f, 32'shdade2d28, 32'shdae34b6d, 32'shdae86a0d, 32'shdaed8909, 32'shdaf2a860, 32'shdaf7c813, 
               32'shdafce821, 32'shdb02088b, 32'shdb072950, 32'shdb0c4a70, 32'shdb116beb, 32'shdb168dc1, 32'shdb1baff2, 32'shdb20d27f, 
               32'shdb25f566, 32'shdb2b18a9, 32'shdb303c46, 32'shdb35603e, 32'shdb3a8491, 32'shdb3fa93e, 32'shdb44ce46, 32'shdb49f3a9, 
               32'shdb4f1967, 32'shdb543f7e, 32'shdb5965f1, 32'shdb5e8cbe, 32'shdb63b3e5, 32'shdb68db67, 32'shdb6e0342, 32'shdb732b79, 
               32'shdb785409, 32'shdb7d7cf3, 32'shdb82a638, 32'shdb87cfd6, 32'shdb8cf9cf, 32'shdb922421, 32'shdb974ece, 32'shdb9c79d4, 
               32'shdba1a534, 32'shdba6d0ed, 32'shdbabfd01, 32'shdbb1296e, 32'shdbb65634, 32'shdbbb8354, 32'shdbc0b0ce, 32'shdbc5dea1, 
               32'shdbcb0cce, 32'shdbd03b53, 32'shdbd56a32, 32'shdbda996b, 32'shdbdfc8fc, 32'shdbe4f8e7, 32'shdbea292b, 32'shdbef59c7, 
               32'shdbf48abd, 32'shdbf9bc0c, 32'shdbfeedb3, 32'shdc041fb4, 32'shdc09520d, 32'shdc0e84bf, 32'shdc13b7c9, 32'shdc18eb2d, 
               32'shdc1e1ee9, 32'shdc2352fd, 32'shdc28876a, 32'shdc2dbc2f, 32'shdc32f14d, 32'shdc3826c3, 32'shdc3d5c91, 32'shdc4292b8, 
               32'shdc47c936, 32'shdc4d000d, 32'shdc52373c, 32'shdc576ec3, 32'shdc5ca6a2, 32'shdc61ded9, 32'shdc671768, 32'shdc6c504e, 
               32'shdc71898d, 32'shdc76c323, 32'shdc7bfd11, 32'shdc813756, 32'shdc8671f3, 32'shdc8bace8, 32'shdc90e834, 32'shdc9623d7, 
               32'shdc9b5fd2, 32'shdca09c24, 32'shdca5d8cd, 32'shdcab15ce, 32'shdcb05326, 32'shdcb590d5, 32'shdcbacedb, 32'shdcc00d38, 
               32'shdcc54bec, 32'shdcca8af7, 32'shdccfca59, 32'shdcd50a12, 32'shdcda4a21, 32'shdcdf8a87, 32'shdce4cb44, 32'shdcea0c58, 
               32'shdcef4dc2, 32'shdcf48f82, 32'shdcf9d199, 32'shdcff1407, 32'shdd0456ca, 32'shdd0999e4, 32'shdd0edd55, 32'shdd14211b, 
               32'shdd196538, 32'shdd1ea9ab, 32'shdd23ee74, 32'shdd293393, 32'shdd2e7908, 32'shdd33bed3, 32'shdd3904f4, 32'shdd3e4b6a, 
               32'shdd439236, 32'shdd48d958, 32'shdd4e20d0, 32'shdd53689d, 32'shdd58b0c0, 32'shdd5df938, 32'shdd634206, 32'shdd688b29, 
               32'shdd6dd4a2, 32'shdd731e6f, 32'shdd786892, 32'shdd7db30b, 32'shdd82fdd8, 32'shdd8848fb, 32'shdd8d9472, 32'shdd92e03f, 
               32'shdd982c60, 32'shdd9d78d7, 32'shdda2c5a2, 32'shdda812c2, 32'shddad6036, 32'shddb2ae00, 32'shddb7fc1e, 32'shddbd4a91, 
               32'shddc29958, 32'shddc7e873, 32'shddcd37e4, 32'shddd287a8, 32'shddd7d7c1, 32'shdddd282e, 32'shdde278ef, 32'shdde7ca05, 
               32'shdded1b6e, 32'shddf26d2c, 32'shddf7bf3e, 32'shddfd11a3, 32'shde02645d, 32'shde07b76b, 32'shde0d0acc, 32'shde125e81, 
               32'shde17b28a, 32'shde1d06e6, 32'shde225b96, 32'shde27b09a, 32'shde2d05f1, 32'shde325b9b, 32'shde37b199, 32'shde3d07eb, 
               32'shde425e8f, 32'shde47b587, 32'shde4d0cd2, 32'shde526471, 32'shde57bc62, 32'shde5d14a6, 32'shde626d3e, 32'shde67c628, 
               32'shde6d1f65, 32'shde7278f5, 32'shde77d2d8, 32'shde7d2d0e, 32'shde828796, 32'shde87e271, 32'shde8d3d9e, 32'shde92991e, 
               32'shde97f4f1, 32'shde9d5116, 32'shdea2ad8d, 32'shdea80a57, 32'shdead6773, 32'shdeb2c4e1, 32'shdeb822a1, 32'shdebd80b3, 
               32'shdec2df18, 32'shdec83dce, 32'shdecd9cd7, 32'shded2fc31, 32'shded85bdd, 32'shdeddbbdb, 32'shdee31c2b, 32'shdee87ccc, 
               32'shdeedddc0, 32'shdef33f04, 32'shdef8a09b, 32'shdefe0282, 32'shdf0364bc, 32'shdf08c746, 32'shdf0e2a22, 32'shdf138d4f, 
               32'shdf18f0ce, 32'shdf1e549d, 32'shdf23b8be, 32'shdf291d30, 32'shdf2e81f3, 32'shdf33e707, 32'shdf394c6b, 32'shdf3eb221, 
               32'shdf441828, 32'shdf497e7f, 32'shdf4ee527, 32'shdf544c1f, 32'shdf59b369, 32'shdf5f1b02, 32'shdf6482ed, 32'shdf69eb27, 
               32'shdf6f53b3, 32'shdf74bc8e, 32'shdf7a25ba, 32'shdf7f8f36, 32'shdf84f902, 32'shdf8a631f, 32'shdf8fcd8b, 32'shdf953848, 
               32'shdf9aa354, 32'shdfa00eb1, 32'shdfa57a5d, 32'shdfaae659, 32'shdfb052a5, 32'shdfb5bf41, 32'shdfbb2c2c, 32'shdfc09967, 
               32'shdfc606f1, 32'shdfcb74cb, 32'shdfd0e2f5, 32'shdfd6516e, 32'shdfdbc036, 32'shdfe12f4e, 32'shdfe69eb4, 32'shdfec0e6a, 
               32'shdff17e70, 32'shdff6eec4, 32'shdffc5f67, 32'she001d05a, 32'she007419b, 32'she00cb32b, 32'she012250a, 32'she0179738, 
               32'she01d09b4, 32'she0227c7f, 32'she027ef99, 32'she02d6301, 32'she032d6b8, 32'she0384abe, 32'she03dbf11, 32'she04333b3, 
               32'she048a8a4, 32'she04e1de3, 32'she053936f, 32'she059094a, 32'she05e7f74, 32'she063f5eb, 32'she0696cb0, 32'she06ee3c3, 
               32'she0745b24, 32'she079d2d3, 32'she07f4acf, 32'she084c31a, 32'she08a3bb2, 32'she08fb497, 32'she0952dcb, 32'she09aa74b, 
               32'she0a0211a, 32'she0a59b35, 32'she0ab159e, 32'she0b09055, 32'she0b60b58, 32'she0bb86a9, 32'she0c10247, 32'she0c67e32, 
               32'she0cbfa6a, 32'she0d176ef, 32'she0d6f3c1, 32'she0dc70e0, 32'she0e1ee4b, 32'she0e76c04, 32'she0ecea09, 32'she0f2685b, 
               32'she0f7e6f9, 32'she0fd65e4, 32'she102e51c, 32'she10864a0, 32'she10de470, 32'she113648d, 32'she118e4f6, 32'she11e65ac, 
               32'she123e6ad, 32'she12967fb, 32'she12ee995, 32'she1346b7a, 32'she139edac, 32'she13f702a, 32'she144f2f3, 32'she14a7609, 
               32'she14ff96a, 32'she1557d17, 32'she15b0110, 32'she1608554, 32'she16609e3, 32'she16b8ebf, 32'she17113e5, 32'she1769958, 
               32'she17c1f15, 32'she181a51e, 32'she1872b72, 32'she18cb211, 32'she19238fb, 32'she197c031, 32'she19d47b1, 32'she1a2cf7c, 
               32'she1a85793, 32'she1addff4, 32'she1b368a0, 32'she1b8f197, 32'she1be7ad8, 32'she1c40464, 32'she1c98e3b, 32'she1cf185c, 
               32'she1d4a2c8, 32'she1da2d7e, 32'she1dfb87f, 32'she1e543ca, 32'she1eacf5f, 32'she1f05b3e, 32'she1f5e768, 32'she1fb73dc, 
               32'she2010099, 32'she2068da1, 32'she20c1af3, 32'she211a88f, 32'she2173674, 32'she21cc4a3, 32'she222531c, 32'she227e1df, 
               32'she22d70eb, 32'she2330041, 32'she2388fe1, 32'she23e1fca, 32'she243affc, 32'she2494078, 32'she24ed13d, 32'she254624b, 
               32'she259f3a3, 32'she25f8544, 32'she265172e, 32'she26aa960, 32'she2703bdc, 32'she275cea1, 32'she27b61af, 32'she280f505, 
               32'she28688a4, 32'she28c1c8c, 32'she291b0bd, 32'she2974536, 32'she29cd9f8, 32'she2a26f03, 32'she2a80456, 32'she2ad99f1, 
               32'she2b32fd4, 32'she2b8c600, 32'she2be5c74, 32'she2c3f331, 32'she2c98a35, 32'she2cf2182, 32'she2d4b916, 32'she2da50f3, 
               32'she2dfe917, 32'she2e58183, 32'she2eb1a37, 32'she2f0b333, 32'she2f64c77, 32'she2fbe602, 32'she3017fd5, 32'she30719ef, 
               32'she30cb451, 32'she3124efa, 32'she317e9eb, 32'she31d8523, 32'she32320a2, 32'she328bc69, 32'she32e5876, 32'she333f4cb, 
               32'she3399167, 32'she33f2e4a, 32'she344cb73, 32'she34a68e4, 32'she350069b, 32'she355a49a, 32'she35b42df, 32'she360e16a, 
               32'she366803c, 32'she36c1f55, 32'she371beb5, 32'she3775e5a, 32'she37cfe47, 32'she3829e79, 32'she3883ef2, 32'she38ddfb1, 
               32'she39380b6, 32'she3992202, 32'she39ec393, 32'she3a4656b, 32'she3aa0788, 32'she3afa9ec, 32'she3b54c95, 32'she3baef84, 
               32'she3c092b9, 32'she3c63633, 32'she3cbd9f4, 32'she3d17df9, 32'she3d72245, 32'she3dcc6d5, 32'she3e26bac, 32'she3e810c7, 
               32'she3edb628, 32'she3f35bce, 32'she3f901ba, 32'she3fea7ea, 32'she4044e60, 32'she409f51a, 32'she40f9c1a, 32'she415435f, 
               32'she41aeae8, 32'she42092b6, 32'she4263ac9, 32'she42be321, 32'she4318bbe, 32'she437349f, 32'she43cddc4, 32'she442872e, 
               32'she44830dd, 32'she44ddad0, 32'she4538507, 32'she4592f83, 32'she45eda43, 32'she4648547, 32'she46a308f, 32'she46fdc1b, 
               32'she47587eb, 32'she47b33ff, 32'she480e057, 32'she4868cf3, 32'she48c39d3, 32'she491e6f6, 32'she497945d, 32'she49d4208, 
               32'she4a2eff6, 32'she4a89e28, 32'she4ae4c9d, 32'she4b3fb56, 32'she4b9aa52, 32'she4bf5991, 32'she4c50914, 32'she4cab8d9, 
               32'she4d068e2, 32'she4d6192e, 32'she4dbc9bd, 32'she4e17a8f, 32'she4e72ba4, 32'she4ecdcfc, 32'she4f28e96, 32'she4f84074, 
               32'she4fdf294, 32'she503a4f6, 32'she509579b, 32'she50f0a83, 32'she514bdad, 32'she51a711a, 32'she52024c9, 32'she525d8ba, 
               32'she52b8cee, 32'she5314163, 32'she536f61b, 32'she53cab15, 32'she5426051, 32'she54815cf, 32'she54dcb8f, 32'she5538191, 
               32'she55937d5, 32'she55eee5a, 32'she564a521, 32'she56a5c2a, 32'she5701374, 32'she575cb00, 32'she57b82cd, 32'she5813adc, 
               32'she586f32c, 32'she58cabbe, 32'she5926490, 32'she5981da4, 32'she59dd6f9, 32'she5a39090, 32'she5a94a67, 32'she5af047f, 
               32'she5b4bed8, 32'she5ba7972, 32'she5c0344d, 32'she5c5ef69, 32'she5cbaac5, 32'she5d16662, 32'she5d72240, 32'she5dcde5e, 
               32'she5e29abc, 32'she5e8575b, 32'she5ee143b, 32'she5f3d15b, 32'she5f98ebb, 32'she5ff4c5b, 32'she6050a3b, 32'she60ac85c, 
               32'she61086bc, 32'she616455d, 32'she61c043d, 32'she621c35e, 32'she62782be, 32'she62d425e, 32'she633023e, 32'she638c25d, 
               32'she63e82bc, 32'she644435a, 32'she64a0438, 32'she64fc556, 32'she65586b3, 32'she65b484f, 32'she6610a2a, 32'she666cc45, 
               32'she66c8e9f, 32'she6725138, 32'she6781410, 32'she67dd727, 32'she6839a7c, 32'she6895e11, 32'she68f21e5, 32'she694e5f7, 
               32'she69aaa48, 32'she6a06ed8, 32'she6a633a6, 32'she6abf8b3, 32'she6b1bdff, 32'she6b78389, 32'she6bd4951, 32'she6c30f57, 
               32'she6c8d59c, 32'she6ce9c1f, 32'she6d462e1, 32'she6da29e0, 32'she6dff11d, 32'she6e5b899, 32'she6eb8052, 32'she6f14849, 
               32'she6f7107e, 32'she6fcd8f1, 32'she702a1a1, 32'she7086a8f, 32'she70e33bb, 32'she713fd25, 32'she719c6cb, 32'she71f90b0, 
               32'she7255ad1, 32'she72b2530, 32'she730efcc, 32'she736baa6, 32'she73c85bc, 32'she7425110, 32'she7481ca1, 32'she74de86f, 
               32'she753b479, 32'she75980c1, 32'she75f4d45, 32'she7651a06, 32'she76ae704, 32'she770b43e, 32'she77681b6, 32'she77c4f69, 
               32'she7821d59, 32'she787eb86, 32'she78db9ef, 32'she7938894, 32'she7995776, 32'she79f2693, 32'she7a4f5ed, 32'she7aac583, 
               32'she7b09555, 32'she7b66563, 32'she7bc35ad, 32'she7c20633, 32'she7c7d6f4, 32'she7cda7f2, 32'she7d3792b, 32'she7d94a9f, 
               32'she7df1c50, 32'she7e4ee3c, 32'she7eac063, 32'she7f092c6, 32'she7f66564, 32'she7fc383d, 32'she8020b52, 32'she807dea2, 
               32'she80db22d, 32'she81385f3, 32'she81959f4, 32'she81f2e30, 32'she82502a7, 32'she82ad759, 32'she830ac45, 32'she836816d, 
               32'she83c56cf, 32'she8422c6c, 32'she8480243, 32'she84dd855, 32'she853aea1, 32'she8598528, 32'she85f5be9, 32'she86532e4, 
               32'she86b0a1a, 32'she870e18a, 32'she876b934, 32'she87c9118, 32'she8826936, 32'she888418e, 32'she88e1a20, 32'she893f2eb, 
               32'she899cbf1, 32'she89fa530, 32'she8a57ea9, 32'she8ab585c, 32'she8b13248, 32'she8b70c6d, 32'she8bce6cd, 32'she8c2c165, 
               32'she8c89c37, 32'she8ce7742, 32'she8d45286, 32'she8da2e04, 32'she8e009ba, 32'she8e5e5aa, 32'she8ebc1d3, 32'she8f19e34, 
               32'she8f77acf, 32'she8fd57a2, 32'she90334af, 32'she90911f3, 32'she90eef71, 32'she914cd27, 32'she91aab16, 32'she920893d, 
               32'she926679c, 32'she92c4634, 32'she9322505, 32'she938040d, 32'she93de34e, 32'she943c2c7, 32'she949a278, 32'she94f8261, 
               32'she9556282, 32'she95b42db, 32'she961236c, 32'she9670435, 32'she96ce535, 32'she972c66d, 32'she978a7dd, 32'she97e8984, 
               32'she9846b63, 32'she98a4d7a, 32'she9902fc7, 32'she996124d, 32'she99bf509, 32'she9a1d7fd, 32'she9a7bb28, 32'she9ad9e8a, 
               32'she9b38223, 32'she9b965f3, 32'she9bf49fa, 32'she9c52e38, 32'she9cb12ad, 32'she9d0f758, 32'she9d6dc3b, 32'she9dcc154, 
               32'she9e2a6a3, 32'she9e88c2a, 32'she9ee71e6, 32'she9f457da, 32'she9fa3e03, 32'shea002463, 32'shea060af9, 32'shea0bf1c6, 
               32'shea11d8c8, 32'shea17c001, 32'shea1da770, 32'shea238f15, 32'shea2976ef, 32'shea2f5f00, 32'shea354746, 32'shea3b2fc2, 
               32'shea411874, 32'shea47015c, 32'shea4cea79, 32'shea52d3cc, 32'shea58bd54, 32'shea5ea712, 32'shea649105, 32'shea6a7b2d, 
               32'shea70658a, 32'shea76501d, 32'shea7c3ae5, 32'shea8225e2, 32'shea881114, 32'shea8dfc7b, 32'shea93e817, 32'shea99d3e8, 
               32'shea9fbfed, 32'sheaa5ac27, 32'sheaab9896, 32'sheab1853a, 32'sheab77212, 32'sheabd5f1f, 32'sheac34c60, 32'sheac939d5, 
               32'sheacf277f, 32'shead5155d, 32'sheadb0370, 32'sheae0f1b6, 32'sheae6e031, 32'sheaeccee0, 32'sheaf2bdc3, 32'sheaf8acd9, 
               32'sheafe9c24, 32'sheb048ba2, 32'sheb0a7b54, 32'sheb106b3a, 32'sheb165b54, 32'sheb1c4ba1, 32'sheb223c22, 32'sheb282cd6, 
               32'sheb2e1dbe, 32'sheb340ed9, 32'sheb3a0027, 32'sheb3ff1a8, 32'sheb45e35d, 32'sheb4bd545, 32'sheb51c760, 32'sheb57b9ae, 
               32'sheb5dac2f, 32'sheb639ee3, 32'sheb6991ca, 32'sheb6f84e3, 32'sheb75782f, 32'sheb7b6bae, 32'sheb815f60, 32'sheb875344, 
               32'sheb8d475b, 32'sheb933ba4, 32'sheb99301f, 32'sheb9f24cd, 32'sheba519ad, 32'shebab0ec0, 32'shebb10404, 32'shebb6f97b, 
               32'shebbcef23, 32'shebc2e4fe, 32'shebc8db0b, 32'shebced149, 32'shebd4c7ba, 32'shebdabe5c, 32'shebe0b52f, 32'shebe6ac35, 
               32'shebeca36c, 32'shebf29ad4, 32'shebf8926f, 32'shebfe8a3a, 32'shec048237, 32'shec0a7a65, 32'shec1072c4, 32'shec166b55, 
               32'shec1c6417, 32'shec225d09, 32'shec28562d, 32'shec2e4f82, 32'shec344908, 32'shec3a42be, 32'shec403ca5, 32'shec4636bd, 
               32'shec4c3106, 32'shec522b7f, 32'shec582629, 32'shec5e2103, 32'shec641c0e, 32'shec6a1749, 32'shec7012b5, 32'shec760e51, 
               32'shec7c0a1d, 32'shec820619, 32'shec880245, 32'shec8dfea1, 32'shec93fb2e, 32'shec99f7ea, 32'shec9ff4d6, 32'sheca5f1f2, 
               32'shecabef3d, 32'shecb1ecb8, 32'shecb7ea63, 32'shecbde83e, 32'shecc3e648, 32'shecc9e481, 32'sheccfe2ea, 32'shecd5e182, 
               32'shecdbe04a, 32'shece1df40, 32'shece7de66, 32'shecedddbb, 32'shecf3dd3f, 32'shecf9dcf3, 32'shecffdcd4, 32'shed05dce5, 
               32'shed0bdd25, 32'shed11dd94, 32'shed17de31, 32'shed1ddefd, 32'shed23dff7, 32'shed29e120, 32'shed2fe277, 32'shed35e3fd, 
               32'shed3be5b1, 32'shed41e794, 32'shed47e9a5, 32'shed4debe4, 32'shed53ee51, 32'shed59f0ec, 32'shed5ff3b5, 32'shed65f6ac, 
               32'shed6bf9d1, 32'shed71fd24, 32'shed7800a5, 32'shed7e0453, 32'shed84082f, 32'shed8a0c39, 32'shed901070, 32'shed9614d5, 
               32'shed9c1967, 32'sheda21e26, 32'sheda82313, 32'shedae282d, 32'shedb42d74, 32'shedba32e9, 32'shedc0388a, 32'shedc63e59, 
               32'shedcc4454, 32'shedd24a7d, 32'shedd850d2, 32'shedde5754, 32'shede45e03, 32'shedea64de, 32'shedf06be6, 32'shedf6731b, 
               32'shedfc7a7c, 32'shee02820a, 32'shee0889c4, 32'shee0e91aa, 32'shee1499bd, 32'shee1aa1fc, 32'shee20aa67, 32'shee26b2fe, 
               32'shee2cbbc1, 32'shee32c4b0, 32'shee38cdcb, 32'shee3ed712, 32'shee44e084, 32'shee4aea23, 32'shee50f3ed, 32'shee56fde3, 
               32'shee5d0804, 32'shee631251, 32'shee691cc9, 32'shee6f276d, 32'shee75323c, 32'shee7b3d36, 32'shee81485c, 32'shee8753ad, 
               32'shee8d5f29, 32'shee936acf, 32'shee9976a1, 32'shee9f829e, 32'sheea58ec6, 32'sheeab9b18, 32'sheeb1a796, 32'sheeb7b43e, 
               32'sheebdc110, 32'sheec3ce0d, 32'sheec9db35, 32'sheecfe887, 32'sheed5f604, 32'sheedc03ab, 32'sheee2117c, 32'sheee81f78, 
               32'sheeee2d9d, 32'sheef43bed, 32'sheefa4a67, 32'shef00590b, 32'shef0667d9, 32'shef0c76d0, 32'shef1285f2, 32'shef18953d, 
               32'shef1ea4b2, 32'shef24b451, 32'shef2ac419, 32'shef30d40a, 32'shef36e426, 32'shef3cf46a, 32'shef4304d8, 32'shef491570, 
               32'shef4f2630, 32'shef55371a, 32'shef5b482d, 32'shef615969, 32'shef676ace, 32'shef6d7c5b, 32'shef738e12, 32'shef799ff2, 
               32'shef7fb1fa, 32'shef85c42b, 32'shef8bd685, 32'shef91e907, 32'shef97fbb2, 32'shef9e0e85, 32'shefa42181, 32'shefaa34a5, 
               32'shefb047f2, 32'shefb65b66, 32'shefbc6f03, 32'shefc282c8, 32'shefc896b5, 32'shefceaacb, 32'shefd4bf08, 32'shefdad36c, 
               32'shefe0e7f9, 32'shefe6fcae, 32'shefed118a, 32'sheff3268e, 32'sheff93bba, 32'shefff510d, 32'shf0056687, 32'shf00b7c29, 
               32'shf01191f3, 32'shf017a7e3, 32'shf01dbdfb, 32'shf023d43a, 32'shf029eaa1, 32'shf030012e, 32'shf03617e2, 32'shf03c2ebd, 
               32'shf04245c0, 32'shf0485ce9, 32'shf04e7438, 32'shf0548baf, 32'shf05aa34c, 32'shf060bb10, 32'shf066d2fa, 32'shf06ceb0b, 
               32'shf0730342, 32'shf0791ba0, 32'shf07f3424, 32'shf0854cce, 32'shf08b659f, 32'shf0917e95, 32'shf09797b2, 32'shf09db0f4, 
               32'shf0a3ca5d, 32'shf0a9e3eb, 32'shf0affda0, 32'shf0b6177a, 32'shf0bc317a, 32'shf0c24b9f, 32'shf0c865ea, 32'shf0ce805b, 
               32'shf0d49af1, 32'shf0dab5ad, 32'shf0e0d08d, 32'shf0e6eb94, 32'shf0ed06bf, 32'shf0f32210, 32'shf0f93d86, 32'shf0ff5921, 
               32'shf10574e0, 32'shf10b90c5, 32'shf111accf, 32'shf117c8fe, 32'shf11de551, 32'shf12401c9, 32'shf12a1e66, 32'shf1303b27, 
               32'shf136580d, 32'shf13c7518, 32'shf1429247, 32'shf148af9a, 32'shf14ecd11, 32'shf154eaad, 32'shf15b086d, 32'shf1612651, 
               32'shf1674459, 32'shf16d6286, 32'shf17380d6, 32'shf1799f4a, 32'shf17fbde2, 32'shf185dc9d, 32'shf18bfb7d, 32'shf1921a80, 
               32'shf19839a6, 32'shf19e58f1, 32'shf1a4785e, 32'shf1aa97ef, 32'shf1b0b7a4, 32'shf1b6d77c, 32'shf1bcf777, 32'shf1c31795, 
               32'shf1c937d6, 32'shf1cf583b, 32'shf1d578c2, 32'shf1db996d, 32'shf1e1ba3a, 32'shf1e7db2a, 32'shf1edfc3d, 32'shf1f41d72, 
               32'shf1fa3ecb, 32'shf2006046, 32'shf20681e3, 32'shf20ca3a3, 32'shf212c585, 32'shf218e78a, 32'shf21f09b1, 32'shf2252bfa, 
               32'shf22b4e66, 32'shf23170f3, 32'shf23793a3, 32'shf23db674, 32'shf243d968, 32'shf249fc7d, 32'shf2501fb5, 32'shf256430e, 
               32'shf25c6688, 32'shf2628a25, 32'shf268ade3, 32'shf26ed1c2, 32'shf274f5c3, 32'shf27b19e6, 32'shf2813e2a, 32'shf287628f, 
               32'shf28d8715, 32'shf293abbd, 32'shf299d085, 32'shf29ff56f, 32'shf2a61a7a, 32'shf2ac3fa5, 32'shf2b264f2, 32'shf2b88a5f, 
               32'shf2beafed, 32'shf2c4d59c, 32'shf2cafb6b, 32'shf2d1215b, 32'shf2d7476c, 32'shf2dd6d9d, 32'shf2e393ef, 32'shf2e9ba60, 
               32'shf2efe0f2, 32'shf2f607a5, 32'shf2fc2e77, 32'shf302556a, 32'shf3087c7d, 32'shf30ea3af, 32'shf314cb02, 32'shf31af274, 
               32'shf3211a07, 32'shf32741b9, 32'shf32d698a, 32'shf333917c, 32'shf339b98d, 32'shf33fe1bd, 32'shf3460a0d, 32'shf34c327c, 
               32'shf3525b0b, 32'shf35883b9, 32'shf35eac86, 32'shf364d573, 32'shf36afe7e, 32'shf37127a9, 32'shf37750f2, 32'shf37d7a5b, 
               32'shf383a3e2, 32'shf389cd88, 32'shf38ff74d, 32'shf3962130, 32'shf39c4b32, 32'shf3a27553, 32'shf3a89f92, 32'shf3aec9f0, 
               32'shf3b4f46c, 32'shf3bb1f07, 32'shf3c149bf, 32'shf3c77496, 32'shf3cd9f8b, 32'shf3d3ca9e, 32'shf3d9f5cf, 32'shf3e0211f, 
               32'shf3e64c8c, 32'shf3ec7817, 32'shf3f2a3bf, 32'shf3f8cf86, 32'shf3fefb6a, 32'shf405276c, 32'shf40b538b, 32'shf4117fc8, 
               32'shf417ac22, 32'shf41dd89a, 32'shf424052f, 32'shf42a31e1, 32'shf4305eb0, 32'shf4368b9d, 32'shf43cb8a7, 32'shf442e5cd, 
               32'shf4491311, 32'shf44f4071, 32'shf4556def, 32'shf45b9b89, 32'shf461c940, 32'shf467f713, 32'shf46e2504, 32'shf4745310, 
               32'shf47a8139, 32'shf480af7f, 32'shf486dde1, 32'shf48d0c5f, 32'shf4933afa, 32'shf49969b1, 32'shf49f9884, 32'shf4a5c773, 
               32'shf4abf67e, 32'shf4b225a4, 32'shf4b854e7, 32'shf4be8446, 32'shf4c4b3c0, 32'shf4cae356, 32'shf4d11308, 32'shf4d742d6, 
               32'shf4dd72be, 32'shf4e3a2c3, 32'shf4e9d2e3, 32'shf4f0031e, 32'shf4f63374, 32'shf4fc63e6, 32'shf5029473, 32'shf508c51b, 
               32'shf50ef5de, 32'shf51526bc, 32'shf51b57b5, 32'shf52188c9, 32'shf527b9f7, 32'shf52deb41, 32'shf5341ca5, 32'shf53a4e24, 
               32'shf5407fbd, 32'shf546b171, 32'shf54ce33f, 32'shf5531528, 32'shf559472b, 32'shf55f7948, 32'shf565ab80, 32'shf56bddd1, 
               32'shf572103d, 32'shf57842c3, 32'shf57e7563, 32'shf584a81d, 32'shf58adaf0, 32'shf5910dde, 32'shf59740e5, 32'shf59d7406, 
               32'shf5a3a740, 32'shf5a9da94, 32'shf5b00e02, 32'shf5b64189, 32'shf5bc7529, 32'shf5c2a8e3, 32'shf5c8dcb6, 32'shf5cf10a2, 
               32'shf5d544a7, 32'shf5db78c6, 32'shf5e1acfd, 32'shf5e7e14e, 32'shf5ee15b7, 32'shf5f44a39, 32'shf5fa7ed4, 32'shf600b388, 
               32'shf606e854, 32'shf60d1d39, 32'shf6135237, 32'shf619874c, 32'shf61fbc7b, 32'shf625f1c2, 32'shf62c2721, 32'shf6325c98, 
               32'shf6389228, 32'shf63ec7cf, 32'shf644fd8f, 32'shf64b3367, 32'shf6516956, 32'shf6579f5e, 32'shf65dd57d, 32'shf6640bb4, 
               32'shf66a4203, 32'shf670786a, 32'shf676aee8, 32'shf67ce57e, 32'shf6831c2b, 32'shf68952ef, 32'shf68f89cb, 32'shf695c0be, 
               32'shf69bf7c9, 32'shf6a22eea, 32'shf6a86623, 32'shf6ae9d73, 32'shf6b4d4d9, 32'shf6bb0c57, 32'shf6c143ec, 32'shf6c77b97, 
               32'shf6cdb359, 32'shf6d3eb32, 32'shf6da2321, 32'shf6e05b27, 32'shf6e69344, 32'shf6eccb77, 32'shf6f303c0, 32'shf6f93c20, 
               32'shf6ff7496, 32'shf705ad22, 32'shf70be5c4, 32'shf7121e7c, 32'shf718574b, 32'shf71e902f, 32'shf724c92a, 32'shf72b023a, 
               32'shf7313b60, 32'shf737749b, 32'shf73daded, 32'shf743e754, 32'shf74a20d0, 32'shf7505a62, 32'shf756940a, 32'shf75ccdc6, 
               32'shf7630799, 32'shf7694180, 32'shf76f7b7d, 32'shf775b58e, 32'shf77befb5, 32'shf78229f1, 32'shf7886442, 32'shf78e9ea7, 
               32'shf794d922, 32'shf79b13b1, 32'shf7a14e55, 32'shf7a7890d, 32'shf7adc3db, 32'shf7b3febc, 32'shf7ba39b3, 32'shf7c074bd, 
               32'shf7c6afdc, 32'shf7cceb0f, 32'shf7d32657, 32'shf7d961b3, 32'shf7df9d22, 32'shf7e5d8a6, 32'shf7ec143e, 32'shf7f24fea, 
               32'shf7f88ba9, 32'shf7fec77d, 32'shf8050364, 32'shf80b3f5f, 32'shf8117b6d, 32'shf817b78f, 32'shf81df3c5, 32'shf824300e, 
               32'shf82a6c6a, 32'shf830a8da, 32'shf836e55d, 32'shf83d21f3, 32'shf8435e9d, 32'shf8499b59, 32'shf84fd829, 32'shf856150b, 
               32'shf85c5201, 32'shf8628f09, 32'shf868cc24, 32'shf86f0952, 32'shf8754692, 32'shf87b83e5, 32'shf881c14b, 32'shf887fec3, 
               32'shf88e3c4d, 32'shf89479ea, 32'shf89ab799, 32'shf8a0f55b, 32'shf8a7332e, 32'shf8ad7114, 32'shf8b3af0c, 32'shf8b9ed15, 
               32'shf8c02b31, 32'shf8c6695f, 32'shf8cca79e, 32'shf8d2e5f0, 32'shf8d92452, 32'shf8df62c7, 32'shf8e5a14d, 32'shf8ebdfe5, 
               32'shf8f21e8e, 32'shf8f85d49, 32'shf8fe9c15, 32'shf904daf2, 32'shf90b19e0, 32'shf91158e0, 32'shf91797f0, 32'shf91dd712, 
               32'shf9241645, 32'shf92a5589, 32'shf93094dd, 32'shf936d442, 32'shf93d13b8, 32'shf943533f, 32'shf94992d7, 32'shf94fd27f, 
               32'shf9561237, 32'shf95c5200, 32'shf96291d9, 32'shf968d1c3, 32'shf96f11bc, 32'shf97551c6, 32'shf97b91e1, 32'shf981d20b, 
               32'shf9881245, 32'shf98e528f, 32'shf99492ea, 32'shf99ad354, 32'shf9a113cd, 32'shf9a75457, 32'shf9ad94f0, 32'shf9b3d599, 
               32'shf9ba1651, 32'shf9c05719, 32'shf9c697f0, 32'shf9ccd8d6, 32'shf9d319cc, 32'shf9d95ad1, 32'shf9df9be6, 32'shf9e5dd09, 
               32'shf9ec1e3b, 32'shf9f25f7d, 32'shf9f8a0cd, 32'shf9fee22c, 32'shfa05239a, 32'shfa0b6517, 32'shfa11a6a3, 32'shfa17e83d, 
               32'shfa1e29e5, 32'shfa246b9d, 32'shfa2aad62, 32'shfa30ef36, 32'shfa373119, 32'shfa3d7309, 32'shfa43b508, 32'shfa49f715, 
               32'shfa503930, 32'shfa567b5a, 32'shfa5cbd91, 32'shfa62ffd6, 32'shfa694229, 32'shfa6f8489, 32'shfa75c6f8, 32'shfa7c0974, 
               32'shfa824bfd, 32'shfa888e95, 32'shfa8ed139, 32'shfa9513eb, 32'shfa9b56ab, 32'shfaa19978, 32'shfaa7dc52, 32'shfaae1f39, 
               32'shfab4622d, 32'shfabaa52f, 32'shfac0e83d, 32'shfac72b59, 32'shfacd6e81, 32'shfad3b1b6, 32'shfad9f4f8, 32'shfae03847, 
               32'shfae67ba2, 32'shfaecbf0a, 32'shfaf3027e, 32'shfaf945ff, 32'shfaff898c, 32'shfb05cd25, 32'shfb0c10cb, 32'shfb12547d, 
               32'shfb18983b, 32'shfb1edc06, 32'shfb251fdc, 32'shfb2b63be, 32'shfb31a7ac, 32'shfb37eba7, 32'shfb3e2fac, 32'shfb4473be, 
               32'shfb4ab7db, 32'shfb50fc04, 32'shfb574039, 32'shfb5d8479, 32'shfb63c8c4, 32'shfb6a0d1b, 32'shfb70517d, 32'shfb7695ea, 
               32'shfb7cda63, 32'shfb831ee6, 32'shfb896375, 32'shfb8fa80f, 32'shfb95ecb4, 32'shfb9c3163, 32'shfba2761e, 32'shfba8bae3, 
               32'shfbaeffb3, 32'shfbb5448d, 32'shfbbb8973, 32'shfbc1ce62, 32'shfbc8135c, 32'shfbce5861, 32'shfbd49d70, 32'shfbdae289, 
               32'shfbe127ac, 32'shfbe76cda, 32'shfbedb212, 32'shfbf3f753, 32'shfbfa3c9f, 32'shfc0081f5, 32'shfc06c754, 32'shfc0d0cbe, 
               32'shfc135231, 32'shfc1997ae, 32'shfc1fdd34, 32'shfc2622c4, 32'shfc2c685d, 32'shfc32ae00, 32'shfc38f3ac, 32'shfc3f3962, 
               32'shfc457f21, 32'shfc4bc4e9, 32'shfc520aba, 32'shfc585094, 32'shfc5e9678, 32'shfc64dc64, 32'shfc6b2259, 32'shfc716857, 
               32'shfc77ae5e, 32'shfc7df46d, 32'shfc843a85, 32'shfc8a80a6, 32'shfc90c6cf, 32'shfc970d01, 32'shfc9d533b, 32'shfca3997e, 
               32'shfca9dfc8, 32'shfcb0261b, 32'shfcb66c77, 32'shfcbcb2da, 32'shfcc2f945, 32'shfcc93fb9, 32'shfccf8634, 32'shfcd5ccb7, 
               32'shfcdc1342, 32'shfce259d5, 32'shfce8a06f, 32'shfceee711, 32'shfcf52dbb, 32'shfcfb746c, 32'shfd01bb24, 32'shfd0801e4, 
               32'shfd0e48ab, 32'shfd148f7a, 32'shfd1ad650, 32'shfd211d2c, 32'shfd276410, 32'shfd2daafb, 32'shfd33f1ed, 32'shfd3a38e6, 
               32'shfd407fe6, 32'shfd46c6ec, 32'shfd4d0df9, 32'shfd53550d, 32'shfd599c28, 32'shfd5fe348, 32'shfd662a70, 32'shfd6c719e, 
               32'shfd72b8d2, 32'shfd79000d, 32'shfd7f474d, 32'shfd858e94, 32'shfd8bd5e1, 32'shfd921d34, 32'shfd98648d, 32'shfd9eabec, 
               32'shfda4f351, 32'shfdab3abc, 32'shfdb1822c, 32'shfdb7c9a3, 32'shfdbe111e, 32'shfdc458a0, 32'shfdcaa027, 32'shfdd0e7b3, 
               32'shfdd72f45, 32'shfddd76dc, 32'shfde3be78, 32'shfdea0619, 32'shfdf04dc0, 32'shfdf6956c, 32'shfdfcdd1d, 32'shfe0324d2, 
               32'shfe096c8d, 32'shfe0fb44c, 32'shfe15fc11, 32'shfe1c43da, 32'shfe228ba7, 32'shfe28d379, 32'shfe2f1b50, 32'shfe35632c, 
               32'shfe3bab0b, 32'shfe41f2ef, 32'shfe483ad8, 32'shfe4e82c4, 32'shfe54cab5, 32'shfe5b12aa, 32'shfe615aa3, 32'shfe67a2a0, 
               32'shfe6deaa1, 32'shfe7432a5, 32'shfe7a7aae, 32'shfe80c2ba, 32'shfe870aca, 32'shfe8d52de, 32'shfe939af5, 32'shfe99e310, 
               32'shfea02b2e, 32'shfea6734f, 32'shfeacbb74, 32'shfeb3039d, 32'shfeb94bc8, 32'shfebf93f6, 32'shfec5dc28, 32'shfecc245d, 
               32'shfed26c94, 32'shfed8b4cf, 32'shfedefd0c, 32'shfee5454c, 32'shfeeb8d8f, 32'shfef1d5d5, 32'shfef81e1d, 32'shfefe6668, 
               32'shff04aeb5, 32'shff0af704, 32'shff113f56, 32'shff1787aa, 32'shff1dd001, 32'shff24185a, 32'shff2a60b4, 32'shff30a911, 
               32'shff36f170, 32'shff3d39d1, 32'shff438234, 32'shff49ca98, 32'shff5012fe, 32'shff565b66, 32'shff5ca3d0, 32'shff62ec3b, 
               32'shff6934a8, 32'shff6f7d16, 32'shff75c585, 32'shff7c0df6, 32'shff825668, 32'shff889edb, 32'shff8ee750, 32'shff952fc5, 
               32'shff9b783c, 32'shffa1c0b4, 32'shffa8092c, 32'shffae51a5, 32'shffb49a1f, 32'shffbae29a, 32'shffc12b16, 32'shffc77392, 
               32'shffcdbc0f, 32'shffd4048c, 32'shffda4d09, 32'shffe09587, 32'shffe6de05, 32'shffed2684, 32'shfff36f02, 32'shfff9b781
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 15)
         begin
            reg signed [31:0] W_Re_table[16384] = '{
               32'sh40000000, 32'sh3fffffec, 32'sh3fffffb1, 32'sh3fffff4e, 32'sh3ffffec4, 32'sh3ffffe13, 32'sh3ffffd39, 32'sh3ffffc39, 
               32'sh3ffffb11, 32'sh3ffff9c1, 32'sh3ffff84a, 32'sh3ffff6ac, 32'sh3ffff4e6, 32'sh3ffff2f8, 32'sh3ffff0e3, 32'sh3fffeea7, 
               32'sh3fffec43, 32'sh3fffe9b7, 32'sh3fffe705, 32'sh3fffe42a, 32'sh3fffe128, 32'sh3fffddff, 32'sh3fffdaae, 32'sh3fffd736, 
               32'sh3fffd396, 32'sh3fffcfcf, 32'sh3fffcbe0, 32'sh3fffc7ca, 32'sh3fffc38c, 32'sh3fffbf27, 32'sh3fffba9b, 32'sh3fffb5e7, 
               32'sh3fffb10b, 32'sh3fffac08, 32'sh3fffa6de, 32'sh3fffa18c, 32'sh3fff9c12, 32'sh3fff9671, 32'sh3fff90a9, 32'sh3fff8ab9, 
               32'sh3fff84a1, 32'sh3fff7e63, 32'sh3fff77fc, 32'sh3fff716e, 32'sh3fff6ab9, 32'sh3fff63dc, 32'sh3fff5cd8, 32'sh3fff55ac, 
               32'sh3fff4e59, 32'sh3fff46df, 32'sh3fff3f3c, 32'sh3fff3773, 32'sh3fff2f82, 32'sh3fff2769, 32'sh3fff1f29, 32'sh3fff16c1, 
               32'sh3fff0e32, 32'sh3fff057c, 32'sh3ffefc9e, 32'sh3ffef399, 32'sh3ffeea6c, 32'sh3ffee117, 32'sh3ffed79b, 32'sh3ffecdf8, 
               32'sh3ffec42d, 32'sh3ffeba3b, 32'sh3ffeb021, 32'sh3ffea5e0, 32'sh3ffe9b77, 32'sh3ffe90e7, 32'sh3ffe862f, 32'sh3ffe7b50, 
               32'sh3ffe704a, 32'sh3ffe651b, 32'sh3ffe59c6, 32'sh3ffe4e49, 32'sh3ffe42a4, 32'sh3ffe36d8, 32'sh3ffe2ae5, 32'sh3ffe1eca, 
               32'sh3ffe1288, 32'sh3ffe061e, 32'sh3ffdf98c, 32'sh3ffdecd3, 32'sh3ffddff3, 32'sh3ffdd2eb, 32'sh3ffdc5bc, 32'sh3ffdb865, 
               32'sh3ffdaae7, 32'sh3ffd9d42, 32'sh3ffd8f74, 32'sh3ffd8180, 32'sh3ffd7364, 32'sh3ffd6520, 32'sh3ffd56b5, 32'sh3ffd4823, 
               32'sh3ffd3969, 32'sh3ffd2a87, 32'sh3ffd1b7e, 32'sh3ffd0c4e, 32'sh3ffcfcf6, 32'sh3ffced77, 32'sh3ffcddd0, 32'sh3ffcce02, 
               32'sh3ffcbe0c, 32'sh3ffcadef, 32'sh3ffc9daa, 32'sh3ffc8d3e, 32'sh3ffc7caa, 32'sh3ffc6bef, 32'sh3ffc5b0c, 32'sh3ffc4a02, 
               32'sh3ffc38d1, 32'sh3ffc2778, 32'sh3ffc15f7, 32'sh3ffc0450, 32'sh3ffbf280, 32'sh3ffbe089, 32'sh3ffbce6b, 32'sh3ffbbc25, 
               32'sh3ffba9b8, 32'sh3ffb9723, 32'sh3ffb8467, 32'sh3ffb7183, 32'sh3ffb5e78, 32'sh3ffb4b46, 32'sh3ffb37ec, 32'sh3ffb246a, 
               32'sh3ffb10c1, 32'sh3ffafcf1, 32'sh3ffae8f9, 32'sh3ffad4d9, 32'sh3ffac092, 32'sh3ffaac24, 32'sh3ffa978e, 32'sh3ffa82d1, 
               32'sh3ffa6dec, 32'sh3ffa58e0, 32'sh3ffa43ac, 32'sh3ffa2e51, 32'sh3ffa18cf, 32'sh3ffa0325, 32'sh3ff9ed53, 32'sh3ff9d75a, 
               32'sh3ff9c13a, 32'sh3ff9aaf2, 32'sh3ff99483, 32'sh3ff97dec, 32'sh3ff9672d, 32'sh3ff95048, 32'sh3ff9393a, 32'sh3ff92206, 
               32'sh3ff90aaa, 32'sh3ff8f326, 32'sh3ff8db7b, 32'sh3ff8c3a8, 32'sh3ff8abae, 32'sh3ff8938d, 32'sh3ff87b44, 32'sh3ff862d4, 
               32'sh3ff84a3c, 32'sh3ff8317d, 32'sh3ff81896, 32'sh3ff7ff88, 32'sh3ff7e652, 32'sh3ff7ccf5, 32'sh3ff7b370, 32'sh3ff799c4, 
               32'sh3ff77ff1, 32'sh3ff765f6, 32'sh3ff74bd3, 32'sh3ff7318a, 32'sh3ff71718, 32'sh3ff6fc7f, 32'sh3ff6e1bf, 32'sh3ff6c6d7, 
               32'sh3ff6abc8, 32'sh3ff69092, 32'sh3ff67534, 32'sh3ff659ae, 32'sh3ff63e01, 32'sh3ff6222d, 32'sh3ff60631, 32'sh3ff5ea0d, 
               32'sh3ff5cdc3, 32'sh3ff5b150, 32'sh3ff594b7, 32'sh3ff577f6, 32'sh3ff55b0d, 32'sh3ff53dfd, 32'sh3ff520c5, 32'sh3ff50366, 
               32'sh3ff4e5e0, 32'sh3ff4c832, 32'sh3ff4aa5d, 32'sh3ff48c60, 32'sh3ff46e3c, 32'sh3ff44ff0, 32'sh3ff4317d, 32'sh3ff412e2, 
               32'sh3ff3f420, 32'sh3ff3d537, 32'sh3ff3b626, 32'sh3ff396ee, 32'sh3ff3778e, 32'sh3ff35807, 32'sh3ff33858, 32'sh3ff31882, 
               32'sh3ff2f884, 32'sh3ff2d85f, 32'sh3ff2b813, 32'sh3ff2979f, 32'sh3ff27703, 32'sh3ff25640, 32'sh3ff23556, 32'sh3ff21444, 
               32'sh3ff1f30b, 32'sh3ff1d1aa, 32'sh3ff1b022, 32'sh3ff18e73, 32'sh3ff16c9c, 32'sh3ff14a9e, 32'sh3ff12878, 32'sh3ff1062a, 
               32'sh3ff0e3b6, 32'sh3ff0c11a, 32'sh3ff09e56, 32'sh3ff07b6b, 32'sh3ff05858, 32'sh3ff0351e, 32'sh3ff011bd, 32'sh3fefee34, 
               32'sh3fefca84, 32'sh3fefa6ac, 32'sh3fef82ad, 32'sh3fef5e87, 32'sh3fef3a39, 32'sh3fef15c3, 32'sh3feef126, 32'sh3feecc62, 
               32'sh3feea776, 32'sh3fee8263, 32'sh3fee5d28, 32'sh3fee37c6, 32'sh3fee123d, 32'sh3fedec8c, 32'sh3fedc6b4, 32'sh3feda0b4, 
               32'sh3fed7a8c, 32'sh3fed543e, 32'sh3fed2dc8, 32'sh3fed072a, 32'sh3fece065, 32'sh3fecb979, 32'sh3fec9265, 32'sh3fec6b2a, 
               32'sh3fec43c7, 32'sh3fec1c3d, 32'sh3febf48b, 32'sh3febccb2, 32'sh3feba4b2, 32'sh3feb7c8a, 32'sh3feb543b, 32'sh3feb2bc4, 
               32'sh3feb0326, 32'sh3feada60, 32'sh3feab173, 32'sh3fea885f, 32'sh3fea5f23, 32'sh3fea35c0, 32'sh3fea0c35, 32'sh3fe9e283, 
               32'sh3fe9b8a9, 32'sh3fe98ea8, 32'sh3fe96480, 32'sh3fe93a30, 32'sh3fe90fb9, 32'sh3fe8e51a, 32'sh3fe8ba54, 32'sh3fe88f67, 
               32'sh3fe86452, 32'sh3fe83915, 32'sh3fe80db2, 32'sh3fe7e226, 32'sh3fe7b674, 32'sh3fe78a9a, 32'sh3fe75e98, 32'sh3fe7326f, 
               32'sh3fe7061f, 32'sh3fe6d9a7, 32'sh3fe6ad08, 32'sh3fe68042, 32'sh3fe65354, 32'sh3fe6263e, 32'sh3fe5f902, 32'sh3fe5cb9d, 
               32'sh3fe59e12, 32'sh3fe5705f, 32'sh3fe54284, 32'sh3fe51482, 32'sh3fe4e659, 32'sh3fe4b808, 32'sh3fe48990, 32'sh3fe45af1, 
               32'sh3fe42c2a, 32'sh3fe3fd3b, 32'sh3fe3ce26, 32'sh3fe39ee8, 32'sh3fe36f84, 32'sh3fe33ff8, 32'sh3fe31045, 32'sh3fe2e06a, 
               32'sh3fe2b067, 32'sh3fe2803e, 32'sh3fe24fed, 32'sh3fe21f74, 32'sh3fe1eed5, 32'sh3fe1be0d, 32'sh3fe18d1f, 32'sh3fe15c09, 
               32'sh3fe12acb, 32'sh3fe0f966, 32'sh3fe0c7da, 32'sh3fe09626, 32'sh3fe0644b, 32'sh3fe03249, 32'sh3fe0001f, 32'sh3fdfcdce, 
               32'sh3fdf9b55, 32'sh3fdf68b5, 32'sh3fdf35ed, 32'sh3fdf02fe, 32'sh3fdecfe8, 32'sh3fde9caa, 32'sh3fde6945, 32'sh3fde35b9, 
               32'sh3fde0205, 32'sh3fddce2a, 32'sh3fdd9a27, 32'sh3fdd65fd, 32'sh3fdd31ac, 32'sh3fdcfd33, 32'sh3fdcc892, 32'sh3fdc93cb, 
               32'sh3fdc5edc, 32'sh3fdc29c5, 32'sh3fdbf488, 32'sh3fdbbf22, 32'sh3fdb8996, 32'sh3fdb53e2, 32'sh3fdb1e06, 32'sh3fdae804, 
               32'sh3fdab1d9, 32'sh3fda7b88, 32'sh3fda450f, 32'sh3fda0e6f, 32'sh3fd9d7a7, 32'sh3fd9a0b8, 32'sh3fd969a1, 32'sh3fd93263, 
               32'sh3fd8fafe, 32'sh3fd8c372, 32'sh3fd88bbe, 32'sh3fd853e2, 32'sh3fd81bdf, 32'sh3fd7e3b5, 32'sh3fd7ab64, 32'sh3fd772eb, 
               32'sh3fd73a4a, 32'sh3fd70183, 32'sh3fd6c894, 32'sh3fd68f7d, 32'sh3fd6563f, 32'sh3fd61cda, 32'sh3fd5e34e, 32'sh3fd5a99a, 
               32'sh3fd56fbe, 32'sh3fd535bc, 32'sh3fd4fb91, 32'sh3fd4c140, 32'sh3fd486c7, 32'sh3fd44c27, 32'sh3fd4115f, 32'sh3fd3d670, 
               32'sh3fd39b5a, 32'sh3fd3601c, 32'sh3fd324b7, 32'sh3fd2e92b, 32'sh3fd2ad77, 32'sh3fd2719c, 32'sh3fd23599, 32'sh3fd1f96f, 
               32'sh3fd1bd1e, 32'sh3fd180a5, 32'sh3fd14405, 32'sh3fd1073e, 32'sh3fd0ca4f, 32'sh3fd08d39, 32'sh3fd04ffc, 32'sh3fd01297, 
               32'sh3fcfd50b, 32'sh3fcf9757, 32'sh3fcf597c, 32'sh3fcf1b7a, 32'sh3fcedd50, 32'sh3fce9eff, 32'sh3fce6087, 32'sh3fce21e7, 
               32'sh3fcde320, 32'sh3fcda431, 32'sh3fcd651c, 32'sh3fcd25de, 32'sh3fcce67a, 32'sh3fcca6ee, 32'sh3fcc673b, 32'sh3fcc2760, 
               32'sh3fcbe75e, 32'sh3fcba735, 32'sh3fcb66e4, 32'sh3fcb266c, 32'sh3fcae5cd, 32'sh3fcaa506, 32'sh3fca6418, 32'sh3fca2303, 
               32'sh3fc9e1c6, 32'sh3fc9a062, 32'sh3fc95ed7, 32'sh3fc91d24, 32'sh3fc8db4a, 32'sh3fc89948, 32'sh3fc8571f, 32'sh3fc814cf, 
               32'sh3fc7d258, 32'sh3fc78fb9, 32'sh3fc74cf3, 32'sh3fc70a05, 32'sh3fc6c6f0, 32'sh3fc683b4, 32'sh3fc64051, 32'sh3fc5fcc6, 
               32'sh3fc5b913, 32'sh3fc5753a, 32'sh3fc53139, 32'sh3fc4ed11, 32'sh3fc4a8c1, 32'sh3fc4644a, 32'sh3fc41fac, 32'sh3fc3dae6, 
               32'sh3fc395f9, 32'sh3fc350e5, 32'sh3fc30baa, 32'sh3fc2c647, 32'sh3fc280bc, 32'sh3fc23b0b, 32'sh3fc1f532, 32'sh3fc1af32, 
               32'sh3fc1690a, 32'sh3fc122bb, 32'sh3fc0dc45, 32'sh3fc095a8, 32'sh3fc04ee3, 32'sh3fc007f6, 32'sh3fbfc0e3, 32'sh3fbf79a8, 
               32'sh3fbf3246, 32'sh3fbeeabc, 32'sh3fbea30c, 32'sh3fbe5b33, 32'sh3fbe1334, 32'sh3fbdcb0d, 32'sh3fbd82bf, 32'sh3fbd3a4a, 
               32'sh3fbcf1ad, 32'sh3fbca8e9, 32'sh3fbc5ffe, 32'sh3fbc16eb, 32'sh3fbbcdb1, 32'sh3fbb8450, 32'sh3fbb3ac7, 32'sh3fbaf117, 
               32'sh3fbaa740, 32'sh3fba5d41, 32'sh3fba131b, 32'sh3fb9c8ce, 32'sh3fb97e5a, 32'sh3fb933be, 32'sh3fb8e8fb, 32'sh3fb89e11, 
               32'sh3fb852ff, 32'sh3fb807c6, 32'sh3fb7bc65, 32'sh3fb770de, 32'sh3fb7252f, 32'sh3fb6d959, 32'sh3fb68d5b, 32'sh3fb64136, 
               32'sh3fb5f4ea, 32'sh3fb5a877, 32'sh3fb55bdc, 32'sh3fb50f1a, 32'sh3fb4c231, 32'sh3fb47520, 32'sh3fb427e8, 32'sh3fb3da89, 
               32'sh3fb38d02, 32'sh3fb33f54, 32'sh3fb2f17f, 32'sh3fb2a383, 32'sh3fb2555f, 32'sh3fb20714, 32'sh3fb1b8a2, 32'sh3fb16a08, 
               32'sh3fb11b48, 32'sh3fb0cc5f, 32'sh3fb07d50, 32'sh3fb02e19, 32'sh3fafdebb, 32'sh3faf8f36, 32'sh3faf3f89, 32'sh3faeefb6, 
               32'sh3fae9fbb, 32'sh3fae4f98, 32'sh3fadff4e, 32'sh3fadaedd, 32'sh3fad5e45, 32'sh3fad0d86, 32'sh3facbc9f, 32'sh3fac6b91, 
               32'sh3fac1a5b, 32'sh3fabc8ff, 32'sh3fab777b, 32'sh3fab25d0, 32'sh3faad3fd, 32'sh3faa8203, 32'sh3faa2fe2, 32'sh3fa9dd9a, 
               32'sh3fa98b2a, 32'sh3fa93894, 32'sh3fa8e5d5, 32'sh3fa892f0, 32'sh3fa83fe3, 32'sh3fa7ecb0, 32'sh3fa79954, 32'sh3fa745d2, 
               32'sh3fa6f228, 32'sh3fa69e57, 32'sh3fa64a5f, 32'sh3fa5f640, 32'sh3fa5a1f9, 32'sh3fa54d8b, 32'sh3fa4f8f6, 32'sh3fa4a439, 
               32'sh3fa44f55, 32'sh3fa3fa4a, 32'sh3fa3a518, 32'sh3fa34fbe, 32'sh3fa2fa3d, 32'sh3fa2a495, 32'sh3fa24ec6, 32'sh3fa1f8d0, 
               32'sh3fa1a2b2, 32'sh3fa14c6d, 32'sh3fa0f600, 32'sh3fa09f6d, 32'sh3fa048b2, 32'sh3f9ff1d0, 32'sh3f9f9ac6, 32'sh3f9f4396, 
               32'sh3f9eec3e, 32'sh3f9e94bf, 32'sh3f9e3d19, 32'sh3f9de54b, 32'sh3f9d8d56, 32'sh3f9d353a, 32'sh3f9cdcf7, 32'sh3f9c848d, 
               32'sh3f9c2bfb, 32'sh3f9bd342, 32'sh3f9b7a62, 32'sh3f9b215a, 32'sh3f9ac82c, 32'sh3f9a6ed6, 32'sh3f9a1558, 32'sh3f99bbb4, 
               32'sh3f9961e8, 32'sh3f9907f6, 32'sh3f98addb, 32'sh3f98539a, 32'sh3f97f932, 32'sh3f979ea2, 32'sh3f9743eb, 32'sh3f96e90d, 
               32'sh3f968e07, 32'sh3f9632da, 32'sh3f95d787, 32'sh3f957c0b, 32'sh3f952069, 32'sh3f94c4a0, 32'sh3f9468af, 32'sh3f940c97, 
               32'sh3f93b058, 32'sh3f9353f1, 32'sh3f92f763, 32'sh3f929aaf, 32'sh3f923dd2, 32'sh3f91e0cf, 32'sh3f9183a5, 32'sh3f912653, 
               32'sh3f90c8da, 32'sh3f906b3a, 32'sh3f900d72, 32'sh3f8faf84, 32'sh3f8f516e, 32'sh3f8ef331, 32'sh3f8e94cd, 32'sh3f8e3642, 
               32'sh3f8dd78f, 32'sh3f8d78b5, 32'sh3f8d19b4, 32'sh3f8cba8c, 32'sh3f8c5b3d, 32'sh3f8bfbc6, 32'sh3f8b9c28, 32'sh3f8b3c63, 
               32'sh3f8adc77, 32'sh3f8a7c64, 32'sh3f8a1c29, 32'sh3f89bbc7, 32'sh3f895b3e, 32'sh3f88fa8e, 32'sh3f8899b7, 32'sh3f8838b8, 
               32'sh3f87d792, 32'sh3f877645, 32'sh3f8714d1, 32'sh3f86b336, 32'sh3f865174, 32'sh3f85ef8a, 32'sh3f858d79, 32'sh3f852b41, 
               32'sh3f84c8e2, 32'sh3f84665b, 32'sh3f8403ae, 32'sh3f83a0d9, 32'sh3f833ddd, 32'sh3f82daba, 32'sh3f827770, 32'sh3f8213fe, 
               32'sh3f81b065, 32'sh3f814ca6, 32'sh3f80e8bf, 32'sh3f8084b0, 32'sh3f80207b, 32'sh3f7fbc1f, 32'sh3f7f579b, 32'sh3f7ef2f0, 
               32'sh3f7e8e1e, 32'sh3f7e2925, 32'sh3f7dc405, 32'sh3f7d5ebd, 32'sh3f7cf94e, 32'sh3f7c93b9, 32'sh3f7c2dfc, 32'sh3f7bc817, 
               32'sh3f7b620c, 32'sh3f7afbda, 32'sh3f7a9580, 32'sh3f7a2eff, 32'sh3f79c857, 32'sh3f796188, 32'sh3f78fa92, 32'sh3f789374, 
               32'sh3f782c30, 32'sh3f77c4c4, 32'sh3f775d31, 32'sh3f76f577, 32'sh3f768d96, 32'sh3f76258e, 32'sh3f75bd5e, 32'sh3f755508, 
               32'sh3f74ec8a, 32'sh3f7483e5, 32'sh3f741b19, 32'sh3f73b226, 32'sh3f73490b, 32'sh3f72dfca, 32'sh3f727661, 32'sh3f720cd2, 
               32'sh3f71a31b, 32'sh3f71393d, 32'sh3f70cf38, 32'sh3f70650b, 32'sh3f6ffab8, 32'sh3f6f903d, 32'sh3f6f259c, 32'sh3f6ebad3, 
               32'sh3f6e4fe3, 32'sh3f6de4cc, 32'sh3f6d798e, 32'sh3f6d0e29, 32'sh3f6ca29c, 32'sh3f6c36e9, 32'sh3f6bcb0e, 32'sh3f6b5f0c, 
               32'sh3f6af2e3, 32'sh3f6a8693, 32'sh3f6a1a1c, 32'sh3f69ad7e, 32'sh3f6940b8, 32'sh3f68d3cc, 32'sh3f6866b8, 32'sh3f67f97d, 
               32'sh3f678c1c, 32'sh3f671e93, 32'sh3f66b0e3, 32'sh3f66430b, 32'sh3f65d50d, 32'sh3f6566e8, 32'sh3f64f89b, 32'sh3f648a28, 
               32'sh3f641b8d, 32'sh3f63accb, 32'sh3f633de2, 32'sh3f62ced2, 32'sh3f625f9b, 32'sh3f61f03d, 32'sh3f6180b8, 32'sh3f61110b, 
               32'sh3f60a138, 32'sh3f60313d, 32'sh3f5fc11c, 32'sh3f5f50d3, 32'sh3f5ee063, 32'sh3f5e6fcc, 32'sh3f5dff0e, 32'sh3f5d8e29, 
               32'sh3f5d1d1d, 32'sh3f5cabe9, 32'sh3f5c3a8f, 32'sh3f5bc90d, 32'sh3f5b5765, 32'sh3f5ae595, 32'sh3f5a739e, 32'sh3f5a0181, 
               32'sh3f598f3c, 32'sh3f591cd0, 32'sh3f58aa3d, 32'sh3f583783, 32'sh3f57c4a2, 32'sh3f575199, 32'sh3f56de6a, 32'sh3f566b14, 
               32'sh3f55f796, 32'sh3f5583f2, 32'sh3f551026, 32'sh3f549c33, 32'sh3f54281a, 32'sh3f53b3d9, 32'sh3f533f71, 32'sh3f52cae2, 
               32'sh3f52562c, 32'sh3f51e14f, 32'sh3f516c4b, 32'sh3f50f720, 32'sh3f5081cd, 32'sh3f500c54, 32'sh3f4f96b4, 32'sh3f4f20ed, 
               32'sh3f4eaafe, 32'sh3f4e34e9, 32'sh3f4dbeac, 32'sh3f4d4848, 32'sh3f4cd1be, 32'sh3f4c5b0c, 32'sh3f4be433, 32'sh3f4b6d34, 
               32'sh3f4af60d, 32'sh3f4a7ebf, 32'sh3f4a074a, 32'sh3f498fae, 32'sh3f4917eb, 32'sh3f48a001, 32'sh3f4827f0, 32'sh3f47afb8, 
               32'sh3f473759, 32'sh3f46bed3, 32'sh3f464626, 32'sh3f45cd51, 32'sh3f455456, 32'sh3f44db34, 32'sh3f4461eb, 32'sh3f43e87a, 
               32'sh3f436ee3, 32'sh3f42f525, 32'sh3f427b3f, 32'sh3f420133, 32'sh3f4186ff, 32'sh3f410ca5, 32'sh3f409223, 32'sh3f40177b, 
               32'sh3f3f9cab, 32'sh3f3f21b5, 32'sh3f3ea697, 32'sh3f3e2b53, 32'sh3f3dafe7, 32'sh3f3d3455, 32'sh3f3cb89b, 32'sh3f3c3cba, 
               32'sh3f3bc0b3, 32'sh3f3b4484, 32'sh3f3ac82f, 32'sh3f3a4bb2, 32'sh3f39cf0e, 32'sh3f395244, 32'sh3f38d552, 32'sh3f38583a, 
               32'sh3f37dafa, 32'sh3f375d93, 32'sh3f36e006, 32'sh3f366251, 32'sh3f35e476, 32'sh3f356673, 32'sh3f34e849, 32'sh3f3469f9, 
               32'sh3f33eb81, 32'sh3f336ce3, 32'sh3f32ee1d, 32'sh3f326f31, 32'sh3f31f01d, 32'sh3f3170e3, 32'sh3f30f181, 32'sh3f3071f9, 
               32'sh3f2ff24a, 32'sh3f2f7273, 32'sh3f2ef276, 32'sh3f2e7252, 32'sh3f2df206, 32'sh3f2d7194, 32'sh3f2cf0fb, 32'sh3f2c703a, 
               32'sh3f2bef53, 32'sh3f2b6e45, 32'sh3f2aed10, 32'sh3f2a6bb4, 32'sh3f29ea31, 32'sh3f296887, 32'sh3f28e6b6, 32'sh3f2864be, 
               32'sh3f27e29f, 32'sh3f276059, 32'sh3f26ddec, 32'sh3f265b59, 32'sh3f25d89e, 32'sh3f2555bc, 32'sh3f24d2b4, 32'sh3f244f84, 
               32'sh3f23cc2e, 32'sh3f2348b0, 32'sh3f22c50c, 32'sh3f224140, 32'sh3f21bd4e, 32'sh3f213935, 32'sh3f20b4f5, 32'sh3f20308d, 
               32'sh3f1fabff, 32'sh3f1f274a, 32'sh3f1ea26e, 32'sh3f1e1d6c, 32'sh3f1d9842, 32'sh3f1d12f1, 32'sh3f1c8d79, 32'sh3f1c07db, 
               32'sh3f1b8215, 32'sh3f1afc29, 32'sh3f1a7615, 32'sh3f19efdb, 32'sh3f19697a, 32'sh3f18e2f2, 32'sh3f185c43, 32'sh3f17d56d, 
               32'sh3f174e70, 32'sh3f16c74c, 32'sh3f164001, 32'sh3f15b88f, 32'sh3f1530f7, 32'sh3f14a937, 32'sh3f142151, 32'sh3f139944, 
               32'sh3f13110f, 32'sh3f1288b4, 32'sh3f120032, 32'sh3f117789, 32'sh3f10eeb9, 32'sh3f1065c3, 32'sh3f0fdca5, 32'sh3f0f5360, 
               32'sh3f0ec9f5, 32'sh3f0e4063, 32'sh3f0db6a9, 32'sh3f0d2cc9, 32'sh3f0ca2c2, 32'sh3f0c1894, 32'sh3f0b8e3f, 32'sh3f0b03c4, 
               32'sh3f0a7921, 32'sh3f09ee58, 32'sh3f096367, 32'sh3f08d850, 32'sh3f084d12, 32'sh3f07c1ad, 32'sh3f073621, 32'sh3f06aa6e, 
               32'sh3f061e95, 32'sh3f059294, 32'sh3f05066d, 32'sh3f047a1e, 32'sh3f03eda9, 32'sh3f03610d, 32'sh3f02d44a, 32'sh3f024760, 
               32'sh3f01ba50, 32'sh3f012d18, 32'sh3f009fba, 32'sh3f001235, 32'sh3eff8489, 32'sh3efef6b6, 32'sh3efe68bc, 32'sh3efdda9b, 
               32'sh3efd4c54, 32'sh3efcbde5, 32'sh3efc2f50, 32'sh3efba094, 32'sh3efb11b1, 32'sh3efa82a7, 32'sh3ef9f377, 32'sh3ef9641f, 
               32'sh3ef8d4a1, 32'sh3ef844fc, 32'sh3ef7b530, 32'sh3ef7253d, 32'sh3ef69523, 32'sh3ef604e3, 32'sh3ef5747b, 32'sh3ef4e3ed, 
               32'sh3ef45338, 32'sh3ef3c25c, 32'sh3ef3315a, 32'sh3ef2a030, 32'sh3ef20ee0, 32'sh3ef17d69, 32'sh3ef0ebcb, 32'sh3ef05a06, 
               32'sh3eefc81a, 32'sh3eef3608, 32'sh3eeea3ce, 32'sh3eee116e, 32'sh3eed7ee7, 32'sh3eecec39, 32'sh3eec5965, 32'sh3eebc669, 
               32'sh3eeb3347, 32'sh3eea9ffe, 32'sh3eea0c8e, 32'sh3ee978f8, 32'sh3ee8e53a, 32'sh3ee85156, 32'sh3ee7bd4b, 32'sh3ee72919, 
               32'sh3ee694c1, 32'sh3ee60041, 32'sh3ee56b9b, 32'sh3ee4d6ce, 32'sh3ee441da, 32'sh3ee3acbf, 32'sh3ee3177e, 32'sh3ee28216, 
               32'sh3ee1ec87, 32'sh3ee156d1, 32'sh3ee0c0f4, 32'sh3ee02af1, 32'sh3edf94c7, 32'sh3edefe76, 32'sh3ede67fe, 32'sh3eddd15f, 
               32'sh3edd3a9a, 32'sh3edca3ae, 32'sh3edc0c9b, 32'sh3edb7562, 32'sh3edade01, 32'sh3eda467a, 32'sh3ed9aecc, 32'sh3ed916f7, 
               32'sh3ed87efc, 32'sh3ed7e6da, 32'sh3ed74e91, 32'sh3ed6b621, 32'sh3ed61d8a, 32'sh3ed584cd, 32'sh3ed4ebe9, 32'sh3ed452de, 
               32'sh3ed3b9ad, 32'sh3ed32054, 32'sh3ed286d5, 32'sh3ed1ed2f, 32'sh3ed15363, 32'sh3ed0b970, 32'sh3ed01f55, 32'sh3ecf8515, 
               32'sh3eceeaad, 32'sh3ece501f, 32'sh3ecdb56a, 32'sh3ecd1a8e, 32'sh3ecc7f8b, 32'sh3ecbe462, 32'sh3ecb4912, 32'sh3ecaad9b, 
               32'sh3eca11fe, 32'sh3ec9763a, 32'sh3ec8da4f, 32'sh3ec83e3d, 32'sh3ec7a205, 32'sh3ec705a6, 32'sh3ec66920, 32'sh3ec5cc73, 
               32'sh3ec52fa0, 32'sh3ec492a6, 32'sh3ec3f585, 32'sh3ec3583e, 32'sh3ec2bad0, 32'sh3ec21d3b, 32'sh3ec17f7f, 32'sh3ec0e19d, 
               32'sh3ec04394, 32'sh3ebfa564, 32'sh3ebf070e, 32'sh3ebe6891, 32'sh3ebdc9ed, 32'sh3ebd2b22, 32'sh3ebc8c31, 32'sh3ebbed19, 
               32'sh3ebb4ddb, 32'sh3ebaae75, 32'sh3eba0ee9, 32'sh3eb96f36, 32'sh3eb8cf5d, 32'sh3eb82f5d, 32'sh3eb78f36, 32'sh3eb6eee9, 
               32'sh3eb64e75, 32'sh3eb5adda, 32'sh3eb50d18, 32'sh3eb46c30, 32'sh3eb3cb21, 32'sh3eb329ec, 32'sh3eb2888f, 32'sh3eb1e70d, 
               32'sh3eb14563, 32'sh3eb0a393, 32'sh3eb0019c, 32'sh3eaf5f7e, 32'sh3eaebd3a, 32'sh3eae1acf, 32'sh3ead783d, 32'sh3eacd585, 
               32'sh3eac32a6, 32'sh3eab8fa1, 32'sh3eaaec74, 32'sh3eaa4922, 32'sh3ea9a5a8, 32'sh3ea90208, 32'sh3ea85e41, 32'sh3ea7ba54, 
               32'sh3ea7163f, 32'sh3ea67205, 32'sh3ea5cda3, 32'sh3ea5291b, 32'sh3ea4846c, 32'sh3ea3df97, 32'sh3ea33a9b, 32'sh3ea29578, 
               32'sh3ea1f02f, 32'sh3ea14abf, 32'sh3ea0a529, 32'sh3e9fff6b, 32'sh3e9f5988, 32'sh3e9eb37d, 32'sh3e9e0d4c, 32'sh3e9d66f4, 
               32'sh3e9cc076, 32'sh3e9c19d1, 32'sh3e9b7306, 32'sh3e9acc13, 32'sh3e9a24fb, 32'sh3e997dbb, 32'sh3e98d655, 32'sh3e982ec9, 
               32'sh3e978715, 32'sh3e96df3b, 32'sh3e96373b, 32'sh3e958f14, 32'sh3e94e6c6, 32'sh3e943e52, 32'sh3e9395b7, 32'sh3e92ecf6, 
               32'sh3e92440d, 32'sh3e919aff, 32'sh3e90f1ca, 32'sh3e90486e, 32'sh3e8f9eeb, 32'sh3e8ef542, 32'sh3e8e4b72, 32'sh3e8da17c, 
               32'sh3e8cf75f, 32'sh3e8c4d1c, 32'sh3e8ba2b2, 32'sh3e8af821, 32'sh3e8a4d6a, 32'sh3e89a28d, 32'sh3e88f788, 32'sh3e884c5d, 
               32'sh3e87a10c, 32'sh3e86f594, 32'sh3e8649f5, 32'sh3e859e30, 32'sh3e84f245, 32'sh3e844632, 32'sh3e8399f9, 32'sh3e82ed9a, 
               32'sh3e824114, 32'sh3e819467, 32'sh3e80e794, 32'sh3e803a9b, 32'sh3e7f8d7b, 32'sh3e7ee034, 32'sh3e7e32c6, 32'sh3e7d8533, 
               32'sh3e7cd778, 32'sh3e7c2997, 32'sh3e7b7b90, 32'sh3e7acd62, 32'sh3e7a1f0d, 32'sh3e797092, 32'sh3e78c1f0, 32'sh3e781328, 
               32'sh3e77643a, 32'sh3e76b524, 32'sh3e7605e9, 32'sh3e755686, 32'sh3e74a6fd, 32'sh3e73f74e, 32'sh3e734778, 32'sh3e72977c, 
               32'sh3e71e759, 32'sh3e71370f, 32'sh3e70869f, 32'sh3e6fd609, 32'sh3e6f254c, 32'sh3e6e7468, 32'sh3e6dc35e, 32'sh3e6d122e, 
               32'sh3e6c60d7, 32'sh3e6baf59, 32'sh3e6afdb5, 32'sh3e6a4beb, 32'sh3e6999fa, 32'sh3e68e7e2, 32'sh3e6835a4, 32'sh3e67833f, 
               32'sh3e66d0b4, 32'sh3e661e03, 32'sh3e656b2b, 32'sh3e64b82c, 32'sh3e640507, 32'sh3e6351bc, 32'sh3e629e4a, 32'sh3e61eab2, 
               32'sh3e6136f3, 32'sh3e60830d, 32'sh3e5fcf01, 32'sh3e5f1acf, 32'sh3e5e6676, 32'sh3e5db1f7, 32'sh3e5cfd51, 32'sh3e5c4885, 
               32'sh3e5b9392, 32'sh3e5ade79, 32'sh3e5a2939, 32'sh3e5973d3, 32'sh3e58be47, 32'sh3e580894, 32'sh3e5752ba, 32'sh3e569cba, 
               32'sh3e55e694, 32'sh3e553047, 32'sh3e5479d4, 32'sh3e53c33a, 32'sh3e530c7a, 32'sh3e525593, 32'sh3e519e86, 32'sh3e50e752, 
               32'sh3e502ff9, 32'sh3e4f7878, 32'sh3e4ec0d1, 32'sh3e4e0904, 32'sh3e4d5110, 32'sh3e4c98f6, 32'sh3e4be0b6, 32'sh3e4b284f, 
               32'sh3e4a6fc1, 32'sh3e49b70d, 32'sh3e48fe33, 32'sh3e484533, 32'sh3e478c0b, 32'sh3e46d2be, 32'sh3e46194a, 32'sh3e455fb0, 
               32'sh3e44a5ef, 32'sh3e43ec08, 32'sh3e4331fa, 32'sh3e4277c6, 32'sh3e41bd6c, 32'sh3e4102eb, 32'sh3e404844, 32'sh3e3f8d76, 
               32'sh3e3ed282, 32'sh3e3e1768, 32'sh3e3d5c27, 32'sh3e3ca0c0, 32'sh3e3be532, 32'sh3e3b297e, 32'sh3e3a6da4, 32'sh3e39b1a3, 
               32'sh3e38f57c, 32'sh3e38392f, 32'sh3e377cbb, 32'sh3e36c021, 32'sh3e360360, 32'sh3e354679, 32'sh3e34896c, 32'sh3e33cc38, 
               32'sh3e330ede, 32'sh3e32515d, 32'sh3e3193b7, 32'sh3e30d5e9, 32'sh3e3017f6, 32'sh3e2f59dc, 32'sh3e2e9b9c, 32'sh3e2ddd35, 
               32'sh3e2d1ea8, 32'sh3e2c5ff5, 32'sh3e2ba11b, 32'sh3e2ae21b, 32'sh3e2a22f4, 32'sh3e2963a8, 32'sh3e28a435, 32'sh3e27e49b, 
               32'sh3e2724db, 32'sh3e2664f5, 32'sh3e25a4e9, 32'sh3e24e4b6, 32'sh3e24245d, 32'sh3e2363dd, 32'sh3e22a338, 32'sh3e21e26c, 
               32'sh3e212179, 32'sh3e206060, 32'sh3e1f9f21, 32'sh3e1eddbc, 32'sh3e1e1c30, 32'sh3e1d5a7e, 32'sh3e1c98a6, 32'sh3e1bd6a7, 
               32'sh3e1b1482, 32'sh3e1a5237, 32'sh3e198fc5, 32'sh3e18cd2d, 32'sh3e180a6f, 32'sh3e17478a, 32'sh3e168480, 32'sh3e15c14f, 
               32'sh3e14fdf7, 32'sh3e143a79, 32'sh3e1376d5, 32'sh3e12b30b, 32'sh3e11ef1b, 32'sh3e112b04, 32'sh3e1066c7, 32'sh3e0fa263, 
               32'sh3e0eddd9, 32'sh3e0e1929, 32'sh3e0d5453, 32'sh3e0c8f57, 32'sh3e0bca34, 32'sh3e0b04eb, 32'sh3e0a3f7b, 32'sh3e0979e6, 
               32'sh3e08b42a, 32'sh3e07ee47, 32'sh3e07283f, 32'sh3e066210, 32'sh3e059bbb, 32'sh3e04d540, 32'sh3e040e9f, 32'sh3e0347d7, 
               32'sh3e0280e9, 32'sh3e01b9d5, 32'sh3e00f29a, 32'sh3e002b39, 32'sh3dff63b2, 32'sh3dfe9c05, 32'sh3dfdd432, 32'sh3dfd0c38, 
               32'sh3dfc4418, 32'sh3dfb7bd2, 32'sh3dfab365, 32'sh3df9ead3, 32'sh3df9221a, 32'sh3df8593b, 32'sh3df79036, 32'sh3df6c70a, 
               32'sh3df5fdb8, 32'sh3df53440, 32'sh3df46aa2, 32'sh3df3a0de, 32'sh3df2d6f3, 32'sh3df20ce2, 32'sh3df142ab, 32'sh3df0784e, 
               32'sh3defadca, 32'sh3deee321, 32'sh3dee1851, 32'sh3ded4d5b, 32'sh3dec823e, 32'sh3debb6fc, 32'sh3deaeb93, 32'sh3dea2004, 
               32'sh3de9544f, 32'sh3de88874, 32'sh3de7bc72, 32'sh3de6f04b, 32'sh3de623fd, 32'sh3de55789, 32'sh3de48aef, 32'sh3de3be2e, 
               32'sh3de2f148, 32'sh3de2243b, 32'sh3de15708, 32'sh3de089af, 32'sh3ddfbc30, 32'sh3ddeee8a, 32'sh3dde20bf, 32'sh3ddd52cd, 
               32'sh3ddc84b5, 32'sh3ddbb677, 32'sh3ddae813, 32'sh3dda1989, 32'sh3dd94ad8, 32'sh3dd87c02, 32'sh3dd7ad05, 32'sh3dd6dde2, 
               32'sh3dd60e99, 32'sh3dd53f29, 32'sh3dd46f94, 32'sh3dd39fd8, 32'sh3dd2cff7, 32'sh3dd1ffef, 32'sh3dd12fc1, 32'sh3dd05f6d, 
               32'sh3dcf8ef3, 32'sh3dcebe52, 32'sh3dcded8c, 32'sh3dcd1c9f, 32'sh3dcc4b8d, 32'sh3dcb7a54, 32'sh3dcaa8f5, 32'sh3dc9d770, 
               32'sh3dc905c5, 32'sh3dc833f3, 32'sh3dc761fc, 32'sh3dc68fdf, 32'sh3dc5bd9b, 32'sh3dc4eb31, 32'sh3dc418a1, 32'sh3dc345eb, 
               32'sh3dc2730f, 32'sh3dc1a00d, 32'sh3dc0cce5, 32'sh3dbff997, 32'sh3dbf2622, 32'sh3dbe5288, 32'sh3dbd7ec7, 32'sh3dbcaae1, 
               32'sh3dbbd6d4, 32'sh3dbb02a1, 32'sh3dba2e48, 32'sh3db959c9, 32'sh3db88524, 32'sh3db7b059, 32'sh3db6db68, 32'sh3db60651, 
               32'sh3db53113, 32'sh3db45bb0, 32'sh3db38627, 32'sh3db2b077, 32'sh3db1daa2, 32'sh3db104a6, 32'sh3db02e84, 32'sh3daf583d, 
               32'sh3dae81cf, 32'sh3dadab3b, 32'sh3dacd481, 32'sh3dabfda1, 32'sh3dab269b, 32'sh3daa4f6f, 32'sh3da9781d, 32'sh3da8a0a5, 
               32'sh3da7c907, 32'sh3da6f143, 32'sh3da61959, 32'sh3da54149, 32'sh3da46912, 32'sh3da390b6, 32'sh3da2b834, 32'sh3da1df8c, 
               32'sh3da106bd, 32'sh3da02dc9, 32'sh3d9f54af, 32'sh3d9e7b6e, 32'sh3d9da208, 32'sh3d9cc87b, 32'sh3d9beec9, 32'sh3d9b14f1, 
               32'sh3d9a3af2, 32'sh3d9960ce, 32'sh3d988684, 32'sh3d97ac13, 32'sh3d96d17d, 32'sh3d95f6c1, 32'sh3d951bde, 32'sh3d9440d6, 
               32'sh3d9365a8, 32'sh3d928a53, 32'sh3d91aed9, 32'sh3d90d339, 32'sh3d8ff772, 32'sh3d8f1b86, 32'sh3d8e3f74, 32'sh3d8d633c, 
               32'sh3d8c86de, 32'sh3d8baa5a, 32'sh3d8acdb0, 32'sh3d89f0e0, 32'sh3d8913ea, 32'sh3d8836ce, 32'sh3d87598c, 32'sh3d867c24, 
               32'sh3d859e96, 32'sh3d84c0e2, 32'sh3d83e309, 32'sh3d830509, 32'sh3d8226e4, 32'sh3d814898, 32'sh3d806a27, 32'sh3d7f8b8f, 
               32'sh3d7eacd2, 32'sh3d7dcdef, 32'sh3d7ceee5, 32'sh3d7c0fb6, 32'sh3d7b3061, 32'sh3d7a50e6, 32'sh3d797145, 32'sh3d78917e, 
               32'sh3d77b192, 32'sh3d76d17f, 32'sh3d75f147, 32'sh3d7510e8, 32'sh3d743064, 32'sh3d734fb9, 32'sh3d726ee9, 32'sh3d718df3, 
               32'sh3d70acd7, 32'sh3d6fcb95, 32'sh3d6eea2d, 32'sh3d6e08a0, 32'sh3d6d26ec, 32'sh3d6c4513, 32'sh3d6b6313, 32'sh3d6a80ee, 
               32'sh3d699ea3, 32'sh3d68bc32, 32'sh3d67d99b, 32'sh3d66f6de, 32'sh3d6613fb, 32'sh3d6530f3, 32'sh3d644dc4, 32'sh3d636a70, 
               32'sh3d6286f6, 32'sh3d61a356, 32'sh3d60bf90, 32'sh3d5fdba4, 32'sh3d5ef793, 32'sh3d5e135b, 32'sh3d5d2efe, 32'sh3d5c4a7b, 
               32'sh3d5b65d2, 32'sh3d5a8103, 32'sh3d599c0e, 32'sh3d58b6f4, 32'sh3d57d1b3, 32'sh3d56ec4d, 32'sh3d5606c1, 32'sh3d55210f, 
               32'sh3d543b37, 32'sh3d53553a, 32'sh3d526f16, 32'sh3d5188cd, 32'sh3d50a25e, 32'sh3d4fbbc9, 32'sh3d4ed50f, 32'sh3d4dee2e, 
               32'sh3d4d0728, 32'sh3d4c1ffc, 32'sh3d4b38aa, 32'sh3d4a5132, 32'sh3d496994, 32'sh3d4881d1, 32'sh3d4799e8, 32'sh3d46b1d9, 
               32'sh3d45c9a4, 32'sh3d44e14a, 32'sh3d43f8c9, 32'sh3d431023, 32'sh3d422757, 32'sh3d413e65, 32'sh3d40554e, 32'sh3d3f6c11, 
               32'sh3d3e82ae, 32'sh3d3d9925, 32'sh3d3caf76, 32'sh3d3bc5a2, 32'sh3d3adba7, 32'sh3d39f188, 32'sh3d390742, 32'sh3d381cd6, 
               32'sh3d373245, 32'sh3d36478e, 32'sh3d355cb1, 32'sh3d3471af, 32'sh3d338687, 32'sh3d329b39, 32'sh3d31afc5, 32'sh3d30c42b, 
               32'sh3d2fd86c, 32'sh3d2eec87, 32'sh3d2e007c, 32'sh3d2d144c, 32'sh3d2c27f6, 32'sh3d2b3b7a, 32'sh3d2a4ed8, 32'sh3d296210, 
               32'sh3d287523, 32'sh3d278810, 32'sh3d269ad8, 32'sh3d25ad7a, 32'sh3d24bff6, 32'sh3d23d24c, 32'sh3d22e47c, 32'sh3d21f687, 
               32'sh3d21086c, 32'sh3d201a2c, 32'sh3d1f2bc5, 32'sh3d1e3d39, 32'sh3d1d4e88, 32'sh3d1c5fb0, 32'sh3d1b70b3, 32'sh3d1a8190, 
               32'sh3d199248, 32'sh3d18a2da, 32'sh3d17b346, 32'sh3d16c38c, 32'sh3d15d3ad, 32'sh3d14e3a8, 32'sh3d13f37e, 32'sh3d13032d, 
               32'sh3d1212b7, 32'sh3d11221c, 32'sh3d10315a, 32'sh3d0f4074, 32'sh3d0e4f67, 32'sh3d0d5e35, 32'sh3d0c6cdd, 32'sh3d0b7b5f, 
               32'sh3d0a89bc, 32'sh3d0997f3, 32'sh3d08a604, 32'sh3d07b3f0, 32'sh3d06c1b6, 32'sh3d05cf57, 32'sh3d04dcd2, 32'sh3d03ea27, 
               32'sh3d02f757, 32'sh3d020461, 32'sh3d011145, 32'sh3d001e04, 32'sh3cff2a9d, 32'sh3cfe3710, 32'sh3cfd435e, 32'sh3cfc4f86, 
               32'sh3cfb5b89, 32'sh3cfa6766, 32'sh3cf9731d, 32'sh3cf87eaf, 32'sh3cf78a1b, 32'sh3cf69561, 32'sh3cf5a082, 32'sh3cf4ab7e, 
               32'sh3cf3b653, 32'sh3cf2c103, 32'sh3cf1cb8e, 32'sh3cf0d5f3, 32'sh3cefe032, 32'sh3ceeea4c, 32'sh3cedf440, 32'sh3cecfe0f, 
               32'sh3cec07b8, 32'sh3ceb113b, 32'sh3cea1a99, 32'sh3ce923d1, 32'sh3ce82ce4, 32'sh3ce735d1, 32'sh3ce63e98, 32'sh3ce5473a, 
               32'sh3ce44fb7, 32'sh3ce3580e, 32'sh3ce2603f, 32'sh3ce1684b, 32'sh3ce07031, 32'sh3cdf77f2, 32'sh3cde7f8d, 32'sh3cdd8702, 
               32'sh3cdc8e52, 32'sh3cdb957d, 32'sh3cda9c81, 32'sh3cd9a361, 32'sh3cd8aa1b, 32'sh3cd7b0af, 32'sh3cd6b71e, 32'sh3cd5bd67, 
               32'sh3cd4c38b, 32'sh3cd3c989, 32'sh3cd2cf62, 32'sh3cd1d515, 32'sh3cd0daa2, 32'sh3ccfe00b, 32'sh3ccee54d, 32'sh3ccdea6a, 
               32'sh3cccef62, 32'sh3ccbf434, 32'sh3ccaf8e0, 32'sh3cc9fd68, 32'sh3cc901c9, 32'sh3cc80605, 32'sh3cc70a1c, 32'sh3cc60e0d, 
               32'sh3cc511d9, 32'sh3cc4157f, 32'sh3cc318ff, 32'sh3cc21c5b, 32'sh3cc11f90, 32'sh3cc022a0, 32'sh3cbf258b, 32'sh3cbe2850, 
               32'sh3cbd2af0, 32'sh3cbc2d6b, 32'sh3cbb2fbf, 32'sh3cba31ef, 32'sh3cb933f9, 32'sh3cb835dd, 32'sh3cb7379c, 32'sh3cb63936, 
               32'sh3cb53aaa, 32'sh3cb43bf9, 32'sh3cb33d22, 32'sh3cb23e26, 32'sh3cb13f04, 32'sh3cb03fbd, 32'sh3caf4051, 32'sh3cae40bf, 
               32'sh3cad4107, 32'sh3cac412a, 32'sh3cab4128, 32'sh3caa4100, 32'sh3ca940b3, 32'sh3ca84041, 32'sh3ca73fa9, 32'sh3ca63eec, 
               32'sh3ca53e09, 32'sh3ca43d01, 32'sh3ca33bd3, 32'sh3ca23a80, 32'sh3ca13908, 32'sh3ca0376a, 32'sh3c9f35a7, 32'sh3c9e33be, 
               32'sh3c9d31b0, 32'sh3c9c2f7d, 32'sh3c9b2d24, 32'sh3c9a2aa6, 32'sh3c992803, 32'sh3c98253a, 32'sh3c97224c, 32'sh3c961f38, 
               32'sh3c951bff, 32'sh3c9418a1, 32'sh3c93151d, 32'sh3c921174, 32'sh3c910da5, 32'sh3c9009b2, 32'sh3c8f0598, 32'sh3c8e015a, 
               32'sh3c8cfcf6, 32'sh3c8bf86d, 32'sh3c8af3be, 32'sh3c89eeea, 32'sh3c88e9f1, 32'sh3c87e4d2, 32'sh3c86df8e, 32'sh3c85da25, 
               32'sh3c84d496, 32'sh3c83cee2, 32'sh3c82c909, 32'sh3c81c30a, 32'sh3c80bce7, 32'sh3c7fb69d, 32'sh3c7eb02f, 32'sh3c7da99b, 
               32'sh3c7ca2e2, 32'sh3c7b9c03, 32'sh3c7a94ff, 32'sh3c798dd6, 32'sh3c788688, 32'sh3c777f14, 32'sh3c76777b, 32'sh3c756fbd, 
               32'sh3c7467d9, 32'sh3c735fd0, 32'sh3c7257a2, 32'sh3c714f4e, 32'sh3c7046d6, 32'sh3c6f3e37, 32'sh3c6e3574, 32'sh3c6d2c8b, 
               32'sh3c6c237e, 32'sh3c6b1a4a, 32'sh3c6a10f2, 32'sh3c690774, 32'sh3c67fdd1, 32'sh3c66f409, 32'sh3c65ea1c, 32'sh3c64e009, 
               32'sh3c63d5d1, 32'sh3c62cb74, 32'sh3c61c0f1, 32'sh3c60b649, 32'sh3c5fab7c, 32'sh3c5ea08a, 32'sh3c5d9573, 32'sh3c5c8a36, 
               32'sh3c5b7ed4, 32'sh3c5a734d, 32'sh3c5967a1, 32'sh3c585bcf, 32'sh3c574fd8, 32'sh3c5643bc, 32'sh3c55377b, 32'sh3c542b14, 
               32'sh3c531e88, 32'sh3c5211d8, 32'sh3c510501, 32'sh3c4ff806, 32'sh3c4eeae5, 32'sh3c4ddda0, 32'sh3c4cd035, 32'sh3c4bc2a5, 
               32'sh3c4ab4ef, 32'sh3c49a715, 32'sh3c489915, 32'sh3c478af0, 32'sh3c467ca6, 32'sh3c456e37, 32'sh3c445fa2, 32'sh3c4350e9, 
               32'sh3c42420a, 32'sh3c413306, 32'sh3c4023dd, 32'sh3c3f148f, 32'sh3c3e051b, 32'sh3c3cf582, 32'sh3c3be5c5, 32'sh3c3ad5e2, 
               32'sh3c39c5da, 32'sh3c38b5ac, 32'sh3c37a55a, 32'sh3c3694e2, 32'sh3c358446, 32'sh3c347384, 32'sh3c33629d, 32'sh3c325191, 
               32'sh3c314060, 32'sh3c302f09, 32'sh3c2f1d8e, 32'sh3c2e0bed, 32'sh3c2cfa28, 32'sh3c2be83d, 32'sh3c2ad62d, 32'sh3c29c3f8, 
               32'sh3c28b19e, 32'sh3c279f1e, 32'sh3c268c7a, 32'sh3c2579b0, 32'sh3c2466c2, 32'sh3c2353ae, 32'sh3c224075, 32'sh3c212d17, 
               32'sh3c201994, 32'sh3c1f05ec, 32'sh3c1df21f, 32'sh3c1cde2d, 32'sh3c1bca16, 32'sh3c1ab5d9, 32'sh3c19a178, 32'sh3c188cf1, 
               32'sh3c177845, 32'sh3c166375, 32'sh3c154e7f, 32'sh3c143964, 32'sh3c132424, 32'sh3c120ebf, 32'sh3c10f935, 32'sh3c0fe386, 
               32'sh3c0ecdb2, 32'sh3c0db7b9, 32'sh3c0ca19b, 32'sh3c0b8b58, 32'sh3c0a74f0, 32'sh3c095e62, 32'sh3c0847b0, 32'sh3c0730d9, 
               32'sh3c0619dc, 32'sh3c0502bb, 32'sh3c03eb74, 32'sh3c02d409, 32'sh3c01bc78, 32'sh3c00a4c3, 32'sh3bff8ce8, 32'sh3bfe74e9, 
               32'sh3bfd5cc4, 32'sh3bfc447b, 32'sh3bfb2c0c, 32'sh3bfa1379, 32'sh3bf8fac0, 32'sh3bf7e1e3, 32'sh3bf6c8e0, 32'sh3bf5afb9, 
               32'sh3bf4966c, 32'sh3bf37cfb, 32'sh3bf26364, 32'sh3bf149a9, 32'sh3bf02fc9, 32'sh3bef15c3, 32'sh3bedfb99, 32'sh3bece149, 
               32'sh3bebc6d5, 32'sh3beaac3c, 32'sh3be9917e, 32'sh3be8769b, 32'sh3be75b93, 32'sh3be64065, 32'sh3be52513, 32'sh3be4099c, 
               32'sh3be2ee01, 32'sh3be1d240, 32'sh3be0b65a, 32'sh3bdf9a4f, 32'sh3bde7e20, 32'sh3bdd61cb, 32'sh3bdc4552, 32'sh3bdb28b3, 
               32'sh3bda0bf0, 32'sh3bd8ef07, 32'sh3bd7d1fa, 32'sh3bd6b4c8, 32'sh3bd59771, 32'sh3bd479f5, 32'sh3bd35c54, 32'sh3bd23e8f, 
               32'sh3bd120a4, 32'sh3bd00295, 32'sh3bcee460, 32'sh3bcdc607, 32'sh3bcca789, 32'sh3bcb88e5, 32'sh3bca6a1d, 32'sh3bc94b31, 
               32'sh3bc82c1f, 32'sh3bc70ce8, 32'sh3bc5ed8d, 32'sh3bc4ce0c, 32'sh3bc3ae67, 32'sh3bc28e9d, 32'sh3bc16eae, 32'sh3bc04e9a, 
               32'sh3bbf2e62, 32'sh3bbe0e04, 32'sh3bbced82, 32'sh3bbbccda, 32'sh3bbaac0e, 32'sh3bb98b1d, 32'sh3bb86a08, 32'sh3bb748cd, 
               32'sh3bb6276e, 32'sh3bb505e9, 32'sh3bb3e440, 32'sh3bb2c272, 32'sh3bb1a080, 32'sh3bb07e68, 32'sh3baf5c2c, 32'sh3bae39ca, 
               32'sh3bad1744, 32'sh3babf499, 32'sh3baad1ca, 32'sh3ba9aed5, 32'sh3ba88bbc, 32'sh3ba7687e, 32'sh3ba6451b, 32'sh3ba52194, 
               32'sh3ba3fde7, 32'sh3ba2da16, 32'sh3ba1b620, 32'sh3ba09205, 32'sh3b9f6dc5, 32'sh3b9e4961, 32'sh3b9d24d8, 32'sh3b9c002a, 
               32'sh3b9adb57, 32'sh3b99b660, 32'sh3b989144, 32'sh3b976c03, 32'sh3b96469d, 32'sh3b952112, 32'sh3b93fb63, 32'sh3b92d58f, 
               32'sh3b91af97, 32'sh3b908979, 32'sh3b8f6337, 32'sh3b8e3cd0, 32'sh3b8d1644, 32'sh3b8bef94, 32'sh3b8ac8bf, 32'sh3b89a1c5, 
               32'sh3b887aa6, 32'sh3b875363, 32'sh3b862bfb, 32'sh3b85046e, 32'sh3b83dcbc, 32'sh3b82b4e6, 32'sh3b818ceb, 32'sh3b8064cc, 
               32'sh3b7f3c87, 32'sh3b7e141e, 32'sh3b7ceb90, 32'sh3b7bc2de, 32'sh3b7a9a07, 32'sh3b79710b, 32'sh3b7847eb, 32'sh3b771ea5, 
               32'sh3b75f53c, 32'sh3b74cbad, 32'sh3b73a1fa, 32'sh3b727822, 32'sh3b714e25, 32'sh3b702404, 32'sh3b6ef9be, 32'sh3b6dcf54, 
               32'sh3b6ca4c4, 32'sh3b6b7a11, 32'sh3b6a4f38, 32'sh3b69243b, 32'sh3b67f919, 32'sh3b66cdd3, 32'sh3b65a268, 32'sh3b6476d8, 
               32'sh3b634b23, 32'sh3b621f4a, 32'sh3b60f34d, 32'sh3b5fc72a, 32'sh3b5e9ae4, 32'sh3b5d6e78, 32'sh3b5c41e8, 32'sh3b5b1533, 
               32'sh3b59e85a, 32'sh3b58bb5c, 32'sh3b578e39, 32'sh3b5660f2, 32'sh3b553386, 32'sh3b5405f6, 32'sh3b52d841, 32'sh3b51aa67, 
               32'sh3b507c69, 32'sh3b4f4e46, 32'sh3b4e1fff, 32'sh3b4cf193, 32'sh3b4bc303, 32'sh3b4a944d, 32'sh3b496574, 32'sh3b483676, 
               32'sh3b470753, 32'sh3b45d80b, 32'sh3b44a8a0, 32'sh3b43790f, 32'sh3b42495a, 32'sh3b411980, 32'sh3b3fe982, 32'sh3b3eb960, 
               32'sh3b3d8918, 32'sh3b3c58ad, 32'sh3b3b281c, 32'sh3b39f767, 32'sh3b38c68e, 32'sh3b379590, 32'sh3b36646e, 32'sh3b353327, 
               32'sh3b3401bb, 32'sh3b32d02b, 32'sh3b319e77, 32'sh3b306c9d, 32'sh3b2f3aa0, 32'sh3b2e087e, 32'sh3b2cd637, 32'sh3b2ba3cc, 
               32'sh3b2a713d, 32'sh3b293e89, 32'sh3b280bb0, 32'sh3b26d8b3, 32'sh3b25a591, 32'sh3b24724b, 32'sh3b233ee1, 32'sh3b220b52, 
               32'sh3b20d79e, 32'sh3b1fa3c6, 32'sh3b1e6fca, 32'sh3b1d3ba9, 32'sh3b1c0764, 32'sh3b1ad2fa, 32'sh3b199e6c, 32'sh3b1869b9, 
               32'sh3b1734e2, 32'sh3b15ffe6, 32'sh3b14cac6, 32'sh3b139582, 32'sh3b126019, 32'sh3b112a8b, 32'sh3b0ff4d9, 32'sh3b0ebf03, 
               32'sh3b0d8909, 32'sh3b0c52e9, 32'sh3b0b1ca6, 32'sh3b09e63e, 32'sh3b08afb2, 32'sh3b077901, 32'sh3b06422c, 32'sh3b050b32, 
               32'sh3b03d414, 32'sh3b029cd1, 32'sh3b01656b, 32'sh3b002ddf, 32'sh3afef630, 32'sh3afdbe5c, 32'sh3afc8663, 32'sh3afb4e47, 
               32'sh3afa1605, 32'sh3af8dda0, 32'sh3af7a516, 32'sh3af66c68, 32'sh3af53395, 32'sh3af3fa9e, 32'sh3af2c183, 32'sh3af18843, 
               32'sh3af04edf, 32'sh3aef1556, 32'sh3aeddba9, 32'sh3aeca1d8, 32'sh3aeb67e3, 32'sh3aea2dc9, 32'sh3ae8f38b, 32'sh3ae7b928, 
               32'sh3ae67ea1, 32'sh3ae543f6, 32'sh3ae40926, 32'sh3ae2ce32, 32'sh3ae1931a, 32'sh3ae057de, 32'sh3adf1c7d, 32'sh3adde0f8, 
               32'sh3adca54e, 32'sh3adb6980, 32'sh3ada2d8e, 32'sh3ad8f178, 32'sh3ad7b53d, 32'sh3ad678de, 32'sh3ad53c5b, 32'sh3ad3ffb3, 
               32'sh3ad2c2e8, 32'sh3ad185f7, 32'sh3ad048e3, 32'sh3acf0baa, 32'sh3acdce4d, 32'sh3acc90cc, 32'sh3acb5327, 32'sh3aca155d, 
               32'sh3ac8d76f, 32'sh3ac7995c, 32'sh3ac65b26, 32'sh3ac51ccb, 32'sh3ac3de4c, 32'sh3ac29fa9, 32'sh3ac160e1, 32'sh3ac021f5, 
               32'sh3abee2e5, 32'sh3abda3b1, 32'sh3abc6458, 32'sh3abb24db, 32'sh3ab9e53a, 32'sh3ab8a575, 32'sh3ab7658c, 32'sh3ab6257e, 
               32'sh3ab4e54c, 32'sh3ab3a4f6, 32'sh3ab2647c, 32'sh3ab123dd, 32'sh3aafe31b, 32'sh3aaea234, 32'sh3aad6129, 32'sh3aac1ff9, 
               32'sh3aaadea6, 32'sh3aa99d2e, 32'sh3aa85b92, 32'sh3aa719d2, 32'sh3aa5d7ee, 32'sh3aa495e6, 32'sh3aa353b9, 32'sh3aa21168, 
               32'sh3aa0cef3, 32'sh3a9f8c5a, 32'sh3a9e499d, 32'sh3a9d06bc, 32'sh3a9bc3b6, 32'sh3a9a808c, 32'sh3a993d3e, 32'sh3a97f9cc, 
               32'sh3a96b636, 32'sh3a95727c, 32'sh3a942e9d, 32'sh3a92ea9b, 32'sh3a91a674, 32'sh3a906229, 32'sh3a8f1dba, 32'sh3a8dd927, 
               32'sh3a8c9470, 32'sh3a8b4f95, 32'sh3a8a0a95, 32'sh3a88c572, 32'sh3a87802a, 32'sh3a863abe, 32'sh3a84f52f, 32'sh3a83af7b, 
               32'sh3a8269a3, 32'sh3a8123a6, 32'sh3a7fdd86, 32'sh3a7e9742, 32'sh3a7d50da, 32'sh3a7c0a4d, 32'sh3a7ac39d, 32'sh3a797cc8, 
               32'sh3a7835cf, 32'sh3a76eeb2, 32'sh3a75a772, 32'sh3a74600d, 32'sh3a731884, 32'sh3a71d0d7, 32'sh3a708906, 32'sh3a6f4111, 
               32'sh3a6df8f8, 32'sh3a6cb0ba, 32'sh3a6b6859, 32'sh3a6a1fd4, 32'sh3a68d72b, 32'sh3a678e5d, 32'sh3a66456c, 32'sh3a64fc57, 
               32'sh3a63b31d, 32'sh3a6269c0, 32'sh3a61203e, 32'sh3a5fd699, 32'sh3a5e8cd0, 32'sh3a5d42e2, 32'sh3a5bf8d1, 32'sh3a5aae9b, 
               32'sh3a596442, 32'sh3a5819c4, 32'sh3a56cf23, 32'sh3a55845d, 32'sh3a543974, 32'sh3a52ee67, 32'sh3a51a335, 32'sh3a5057e0, 
               32'sh3a4f0c67, 32'sh3a4dc0c9, 32'sh3a4c7508, 32'sh3a4b2923, 32'sh3a49dd1a, 32'sh3a4890ed, 32'sh3a47449c, 32'sh3a45f827, 
               32'sh3a44ab8e, 32'sh3a435ed1, 32'sh3a4211f0, 32'sh3a40c4eb, 32'sh3a3f77c3, 32'sh3a3e2a76, 32'sh3a3cdd05, 32'sh3a3b8f71, 
               32'sh3a3a41b9, 32'sh3a38f3dc, 32'sh3a37a5dc, 32'sh3a3657b8, 32'sh3a350970, 32'sh3a33bb04, 32'sh3a326c74, 32'sh3a311dc0, 
               32'sh3a2fcee8, 32'sh3a2e7fed, 32'sh3a2d30cd, 32'sh3a2be18a, 32'sh3a2a9223, 32'sh3a294298, 32'sh3a27f2e9, 32'sh3a26a316, 
               32'sh3a25531f, 32'sh3a240305, 32'sh3a22b2c6, 32'sh3a216264, 32'sh3a2011de, 32'sh3a1ec134, 32'sh3a1d7066, 32'sh3a1c1f74, 
               32'sh3a1ace5f, 32'sh3a197d25, 32'sh3a182bc8, 32'sh3a16da47, 32'sh3a1588a2, 32'sh3a1436d9, 32'sh3a12e4ed, 32'sh3a1192dc, 
               32'sh3a1040a8, 32'sh3a0eee50, 32'sh3a0d9bd4, 32'sh3a0c4935, 32'sh3a0af671, 32'sh3a09a38a, 32'sh3a08507f, 32'sh3a06fd50, 
               32'sh3a05a9fd, 32'sh3a045687, 32'sh3a0302ed, 32'sh3a01af2f, 32'sh3a005b4d, 32'sh39ff0747, 32'sh39fdb31e, 32'sh39fc5ed1, 
               32'sh39fb0a60, 32'sh39f9b5cb, 32'sh39f86113, 32'sh39f70c37, 32'sh39f5b737, 32'sh39f46213, 32'sh39f30ccc, 32'sh39f1b761, 
               32'sh39f061d2, 32'sh39ef0c1f, 32'sh39edb649, 32'sh39ec604e, 32'sh39eb0a31, 32'sh39e9b3ef, 32'sh39e85d8a, 32'sh39e70701, 
               32'sh39e5b054, 32'sh39e45983, 32'sh39e3028f, 32'sh39e1ab77, 32'sh39e0543c, 32'sh39defcdd, 32'sh39dda55a, 32'sh39dc4db3, 
               32'sh39daf5e8, 32'sh39d99dfa, 32'sh39d845e9, 32'sh39d6edb3, 32'sh39d5955a, 32'sh39d43cdd, 32'sh39d2e43d, 32'sh39d18b79, 
               32'sh39d03291, 32'sh39ced986, 32'sh39cd8056, 32'sh39cc2704, 32'sh39cacd8d, 32'sh39c973f3, 32'sh39c81a36, 32'sh39c6c054, 
               32'sh39c5664f, 32'sh39c40c27, 32'sh39c2b1da, 32'sh39c1576a, 32'sh39bffcd7, 32'sh39bea220, 32'sh39bd4745, 32'sh39bbec47, 
               32'sh39ba9125, 32'sh39b935df, 32'sh39b7da76, 32'sh39b67ee9, 32'sh39b52339, 32'sh39b3c765, 32'sh39b26b6d, 32'sh39b10f52, 
               32'sh39afb313, 32'sh39ae56b1, 32'sh39acfa2b, 32'sh39ab9d81, 32'sh39aa40b4, 32'sh39a8e3c4, 32'sh39a786af, 32'sh39a62978, 
               32'sh39a4cc1c, 32'sh39a36e9d, 32'sh39a210fb, 32'sh39a0b335, 32'sh399f554b, 32'sh399df73e, 32'sh399c990d, 32'sh399b3ab9, 
               32'sh3999dc42, 32'sh39987da6, 32'sh39971ee7, 32'sh3995c005, 32'sh399460ff, 32'sh399301d6, 32'sh3991a289, 32'sh39904319, 
               32'sh398ee385, 32'sh398d83ce, 32'sh398c23f3, 32'sh398ac3f4, 32'sh398963d2, 32'sh3988038d, 32'sh3986a324, 32'sh39854298, 
               32'sh3983e1e8, 32'sh39828115, 32'sh3981201e, 32'sh397fbf04, 32'sh397e5dc6, 32'sh397cfc65, 32'sh397b9ae0, 32'sh397a3938, 
               32'sh3978d76c, 32'sh3977757d, 32'sh3976136b, 32'sh3974b135, 32'sh39734edc, 32'sh3971ec5f, 32'sh397089bf, 32'sh396f26fb, 
               32'sh396dc414, 32'sh396c610a, 32'sh396afddc, 32'sh39699a8a, 32'sh39683715, 32'sh3966d37d, 32'sh39656fc2, 32'sh39640be3, 
               32'sh3962a7e0, 32'sh396143bb, 32'sh395fdf71, 32'sh395e7b05, 32'sh395d1675, 32'sh395bb1c2, 32'sh395a4ceb, 32'sh3958e7f1, 
               32'sh395782d3, 32'sh39561d92, 32'sh3954b82e, 32'sh395352a7, 32'sh3951ecfc, 32'sh3950872d, 32'sh394f213c, 32'sh394dbb27, 
               32'sh394c54ee, 32'sh394aee93, 32'sh39498814, 32'sh39482171, 32'sh3946baac, 32'sh394553c3, 32'sh3943ecb6, 32'sh39428586, 
               32'sh39411e33, 32'sh393fb6bd, 32'sh393e4f23, 32'sh393ce767, 32'sh393b7f86, 32'sh393a1783, 32'sh3938af5c, 32'sh39374712, 
               32'sh3935dea4, 32'sh39347613, 32'sh39330d5f, 32'sh3931a488, 32'sh39303b8e, 32'sh392ed270, 32'sh392d692f, 32'sh392bffca, 
               32'sh392a9642, 32'sh39292c97, 32'sh3927c2c9, 32'sh392658d8, 32'sh3924eec3, 32'sh3923848b, 32'sh39221a30, 32'sh3920afb1, 
               32'sh391f4510, 32'sh391dda4b, 32'sh391c6f63, 32'sh391b0457, 32'sh39199929, 32'sh39182dd7, 32'sh3916c262, 32'sh391556ca, 
               32'sh3913eb0e, 32'sh39127f2f, 32'sh3911132d, 32'sh390fa708, 32'sh390e3ac0, 32'sh390cce55, 32'sh390b61c6, 32'sh3909f514, 
               32'sh3908883f, 32'sh39071b47, 32'sh3905ae2b, 32'sh390440ed, 32'sh3902d38b, 32'sh39016606, 32'sh38fff85e, 32'sh38fe8a93, 
               32'sh38fd1ca4, 32'sh38fbae93, 32'sh38fa405e, 32'sh38f8d206, 32'sh38f7638b, 32'sh38f5f4ed, 32'sh38f4862c, 32'sh38f31747, 
               32'sh38f1a840, 32'sh38f03915, 32'sh38eec9c7, 32'sh38ed5a56, 32'sh38ebeac2, 32'sh38ea7b0b, 32'sh38e90b31, 32'sh38e79b34, 
               32'sh38e62b13, 32'sh38e4bad0, 32'sh38e34a69, 32'sh38e1d9df, 32'sh38e06932, 32'sh38def863, 32'sh38dd8770, 32'sh38dc165a, 
               32'sh38daa520, 32'sh38d933c4, 32'sh38d7c245, 32'sh38d650a3, 32'sh38d4dedd, 32'sh38d36cf5, 32'sh38d1fae9, 32'sh38d088bb, 
               32'sh38cf1669, 32'sh38cda3f4, 32'sh38cc315d, 32'sh38cabea2, 32'sh38c94bc4, 32'sh38c7d8c3, 32'sh38c665a0, 32'sh38c4f259, 
               32'sh38c37eef, 32'sh38c20b62, 32'sh38c097b2, 32'sh38bf23df, 32'sh38bdafea, 32'sh38bc3bd1, 32'sh38bac795, 32'sh38b95336, 
               32'sh38b7deb4, 32'sh38b66a0f, 32'sh38b4f547, 32'sh38b3805c, 32'sh38b20b4f, 32'sh38b0961e, 32'sh38af20ca, 32'sh38adab54, 
               32'sh38ac35ba, 32'sh38aabffd, 32'sh38a94a1e, 32'sh38a7d41b, 32'sh38a65df6, 32'sh38a4e7ad, 32'sh38a37142, 32'sh38a1fab4, 
               32'sh38a08402, 32'sh389f0d2e, 32'sh389d9637, 32'sh389c1f1d, 32'sh389aa7e0, 32'sh38993080, 32'sh3897b8fe, 32'sh38964158, 
               32'sh3894c98f, 32'sh389351a4, 32'sh3891d995, 32'sh38906164, 32'sh388ee910, 32'sh388d7099, 32'sh388bf7ff, 32'sh388a7f42, 
               32'sh38890663, 32'sh38878d60, 32'sh3886143b, 32'sh38849af2, 32'sh38832187, 32'sh3881a7f9, 32'sh38802e48, 32'sh387eb474, 
               32'sh387d3a7e, 32'sh387bc064, 32'sh387a4628, 32'sh3878cbc9, 32'sh38775147, 32'sh3875d6a2, 32'sh38745bdb, 32'sh3872e0f0, 
               32'sh387165e3, 32'sh386feab3, 32'sh386e6f60, 32'sh386cf3ea, 32'sh386b7852, 32'sh3869fc97, 32'sh386880b8, 32'sh386704b8, 
               32'sh38658894, 32'sh38640c4d, 32'sh38628fe4, 32'sh38611358, 32'sh385f96a9, 32'sh385e19d8, 32'sh385c9ce3, 32'sh385b1fcc, 
               32'sh3859a292, 32'sh38582536, 32'sh3856a7b6, 32'sh38552a14, 32'sh3853ac4f, 32'sh38522e68, 32'sh3850b05d, 32'sh384f3230, 
               32'sh384db3e0, 32'sh384c356e, 32'sh384ab6d8, 32'sh38493820, 32'sh3847b946, 32'sh38463a48, 32'sh3844bb28, 32'sh38433be5, 
               32'sh3841bc7f, 32'sh38403cf7, 32'sh383ebd4c, 32'sh383d3d7e, 32'sh383bbd8e, 32'sh383a3d7b, 32'sh3838bd45, 32'sh38373ced, 
               32'sh3835bc71, 32'sh38343bd4, 32'sh3832bb13, 32'sh38313a30, 32'sh382fb92a, 32'sh382e3802, 32'sh382cb6b7, 32'sh382b3549, 
               32'sh3829b3b9, 32'sh38283205, 32'sh3826b030, 32'sh38252e37, 32'sh3823ac1d, 32'sh382229df, 32'sh3820a77f, 32'sh381f24fc, 
               32'sh381da256, 32'sh381c1f8e, 32'sh381a9ca4, 32'sh38191996, 32'sh38179666, 32'sh38161314, 32'sh38148f9f, 32'sh38130c07, 
               32'sh3811884d, 32'sh38100470, 32'sh380e8071, 32'sh380cfc4f, 32'sh380b780a, 32'sh3809f3a3, 32'sh38086f19, 32'sh3806ea6d, 
               32'sh3805659e, 32'sh3803e0ac, 32'sh38025b98, 32'sh3800d662, 32'sh37ff5109, 32'sh37fdcb8d, 32'sh37fc45ef, 32'sh37fac02e, 
               32'sh37f93a4b, 32'sh37f7b446, 32'sh37f62e1d, 32'sh37f4a7d2, 32'sh37f32165, 32'sh37f19ad5, 32'sh37f01423, 32'sh37ee8d4e, 
               32'sh37ed0657, 32'sh37eb7f3d, 32'sh37e9f801, 32'sh37e870a2, 32'sh37e6e921, 32'sh37e5617d, 32'sh37e3d9b7, 32'sh37e251ce, 
               32'sh37e0c9c3, 32'sh37df4195, 32'sh37ddb945, 32'sh37dc30d2, 32'sh37daa83d, 32'sh37d91f86, 32'sh37d796ac, 32'sh37d60daf, 
               32'sh37d48490, 32'sh37d2fb4f, 32'sh37d171eb, 32'sh37cfe865, 32'sh37ce5ebd, 32'sh37ccd4f2, 32'sh37cb4b04, 32'sh37c9c0f4, 
               32'sh37c836c2, 32'sh37c6ac6d, 32'sh37c521f6, 32'sh37c3975d, 32'sh37c20ca1, 32'sh37c081c3, 32'sh37bef6c2, 32'sh37bd6b9f, 
               32'sh37bbe05a, 32'sh37ba54f2, 32'sh37b8c968, 32'sh37b73dbb, 32'sh37b5b1ec, 32'sh37b425fb, 32'sh37b299e7, 32'sh37b10db1, 
               32'sh37af8159, 32'sh37adf4de, 32'sh37ac6841, 32'sh37aadb82, 32'sh37a94ea0, 32'sh37a7c19c, 32'sh37a63476, 32'sh37a4a72d, 
               32'sh37a319c2, 32'sh37a18c34, 32'sh379ffe85, 32'sh379e70b3, 32'sh379ce2be, 32'sh379b54a8, 32'sh3799c66f, 32'sh37983814, 
               32'sh3796a996, 32'sh37951af6, 32'sh37938c34, 32'sh3791fd50, 32'sh37906e49, 32'sh378edf20, 32'sh378d4fd5, 32'sh378bc068, 
               32'sh378a30d8, 32'sh3788a126, 32'sh37871152, 32'sh3785815b, 32'sh3783f143, 32'sh37826108, 32'sh3780d0aa, 32'sh377f402b, 
               32'sh377daf89, 32'sh377c1ec5, 32'sh377a8ddf, 32'sh3778fcd7, 32'sh37776bac, 32'sh3775da5f, 32'sh377448f0, 32'sh3772b75f, 
               32'sh377125ac, 32'sh376f93d6, 32'sh376e01de, 32'sh376c6fc4, 32'sh376add88, 32'sh37694b2a, 32'sh3767b8a9, 32'sh37662606, 
               32'sh37649341, 32'sh3763005a, 32'sh37616d51, 32'sh375fda26, 32'sh375e46d8, 32'sh375cb368, 32'sh375b1fd7, 32'sh37598c23, 
               32'sh3757f84c, 32'sh37566454, 32'sh3754d03a, 32'sh37533bfd, 32'sh3751a79e, 32'sh3750131e, 32'sh374e7e7b, 32'sh374ce9b6, 
               32'sh374b54ce, 32'sh3749bfc5, 32'sh37482a9a, 32'sh3746954c, 32'sh3744ffdd, 32'sh37436a4b, 32'sh3741d497, 32'sh37403ec1, 
               32'sh373ea8ca, 32'sh373d12b0, 32'sh373b7c73, 32'sh3739e615, 32'sh37384f95, 32'sh3736b8f3, 32'sh3735222f, 32'sh37338b48, 
               32'sh3731f440, 32'sh37305d15, 32'sh372ec5c9, 32'sh372d2e5a, 32'sh372b96ca, 32'sh3729ff17, 32'sh37286742, 32'sh3726cf4c, 
               32'sh37253733, 32'sh37239ef8, 32'sh3722069b, 32'sh37206e1d, 32'sh371ed57c, 32'sh371d3cb9, 32'sh371ba3d4, 32'sh371a0ace, 
               32'sh371871a5, 32'sh3716d85a, 32'sh37153eee, 32'sh3713a55f, 32'sh37120bae, 32'sh371071dc, 32'sh370ed7e7, 32'sh370d3dd0, 
               32'sh370ba398, 32'sh370a093d, 32'sh37086ec1, 32'sh3706d423, 32'sh37053962, 32'sh37039e80, 32'sh3702037c, 32'sh37006856, 
               32'sh36fecd0e, 32'sh36fd31a4, 32'sh36fb9618, 32'sh36f9fa6a, 32'sh36f85e9a, 32'sh36f6c2a9, 32'sh36f52695, 32'sh36f38a60, 
               32'sh36f1ee09, 32'sh36f0518f, 32'sh36eeb4f4, 32'sh36ed1837, 32'sh36eb7b58, 32'sh36e9de58, 32'sh36e84135, 32'sh36e6a3f1, 
               32'sh36e5068a, 32'sh36e36902, 32'sh36e1cb58, 32'sh36e02d8c, 32'sh36de8f9e, 32'sh36dcf18f, 32'sh36db535d, 32'sh36d9b50a, 
               32'sh36d81695, 32'sh36d677fe, 32'sh36d4d945, 32'sh36d33a6a, 32'sh36d19b6e, 32'sh36cffc50, 32'sh36ce5d10, 32'sh36ccbdae, 
               32'sh36cb1e2a, 32'sh36c97e85, 32'sh36c7debd, 32'sh36c63ed4, 32'sh36c49ec9, 32'sh36c2fe9d, 32'sh36c15e4e, 32'sh36bfbdde, 
               32'sh36be1d4c, 32'sh36bc7c98, 32'sh36badbc3, 32'sh36b93acc, 32'sh36b799b3, 32'sh36b5f878, 32'sh36b4571b, 32'sh36b2b59d, 
               32'sh36b113fd, 32'sh36af723b, 32'sh36add058, 32'sh36ac2e53, 32'sh36aa8c2c, 32'sh36a8e9e3, 32'sh36a74779, 32'sh36a5a4ed, 
               32'sh36a4023f, 32'sh36a25f70, 32'sh36a0bc7e, 32'sh369f196b, 32'sh369d7637, 32'sh369bd2e1, 32'sh369a2f69, 32'sh36988bcf, 
               32'sh3696e814, 32'sh36954437, 32'sh3693a038, 32'sh3691fc18, 32'sh369057d6, 32'sh368eb372, 32'sh368d0eed, 32'sh368b6a46, 
               32'sh3689c57d, 32'sh36882093, 32'sh36867b87, 32'sh3684d65a, 32'sh3683310b, 32'sh36818b9a, 32'sh367fe608, 32'sh367e4054, 
               32'sh367c9a7e, 32'sh367af487, 32'sh36794e6e, 32'sh3677a833, 32'sh367601d7, 32'sh36745b5a, 32'sh3672b4bb, 32'sh36710dfa, 
               32'sh366f6717, 32'sh366dc013, 32'sh366c18ee, 32'sh366a71a7, 32'sh3668ca3e, 32'sh366722b4, 32'sh36657b08, 32'sh3663d33b, 
               32'sh36622b4c, 32'sh3660833b, 32'sh365edb09, 32'sh365d32b6, 32'sh365b8a41, 32'sh3659e1aa, 32'sh365838f2, 32'sh36569019, 
               32'sh3654e71d, 32'sh36533e01, 32'sh365194c3, 32'sh364feb63, 32'sh364e41e2, 32'sh364c983f, 32'sh364aee7b, 32'sh36494495, 
               32'sh36479a8e, 32'sh3645f065, 32'sh3644461b, 32'sh36429bb0, 32'sh3640f123, 32'sh363f4674, 32'sh363d9ba4, 32'sh363bf0b3, 
               32'sh363a45a0, 32'sh36389a6b, 32'sh3636ef16, 32'sh3635439e, 32'sh36339806, 32'sh3631ec4c, 32'sh36304070, 32'sh362e9473, 
               32'sh362ce855, 32'sh362b3c15, 32'sh36298fb4, 32'sh3627e331, 32'sh3626368d, 32'sh362489c7, 32'sh3622dce1, 32'sh36212fd8, 
               32'sh361f82af, 32'sh361dd564, 32'sh361c27f7, 32'sh361a7a6a, 32'sh3618ccba, 32'sh36171eea, 32'sh361570f8, 32'sh3613c2e5, 
               32'sh361214b0, 32'sh3610665a, 32'sh360eb7e3, 32'sh360d094a, 32'sh360b5a90, 32'sh3609abb5, 32'sh3607fcb8, 32'sh36064d9a, 
               32'sh36049e5b, 32'sh3602eefa, 32'sh36013f78, 32'sh35ff8fd5, 32'sh35fde011, 32'sh35fc302b, 32'sh35fa8023, 32'sh35f8cffb, 
               32'sh35f71fb1, 32'sh35f56f46, 32'sh35f3beba, 32'sh35f20e0c, 32'sh35f05d3d, 32'sh35eeac4d, 32'sh35ecfb3c, 32'sh35eb4a09, 
               32'sh35e998b5, 32'sh35e7e740, 32'sh35e635a9, 32'sh35e483f2, 32'sh35e2d219, 32'sh35e1201e, 32'sh35df6e03, 32'sh35ddbbc6, 
               32'sh35dc0968, 32'sh35da56e9, 32'sh35d8a449, 32'sh35d6f187, 32'sh35d53ea5, 32'sh35d38ba1, 32'sh35d1d87c, 32'sh35d02535, 
               32'sh35ce71ce, 32'sh35ccbe45, 32'sh35cb0a9b, 32'sh35c956d0, 32'sh35c7a2e3, 32'sh35c5eed6, 32'sh35c43aa7, 32'sh35c28658, 
               32'sh35c0d1e7, 32'sh35bf1d54, 32'sh35bd68a1, 32'sh35bbb3cd, 32'sh35b9fed7, 32'sh35b849c0, 32'sh35b69489, 32'sh35b4df30, 
               32'sh35b329b5, 32'sh35b1741a, 32'sh35afbe5e, 32'sh35ae0880, 32'sh35ac5282, 32'sh35aa9c62, 32'sh35a8e621, 32'sh35a72fbf, 
               32'sh35a5793c, 32'sh35a3c298, 32'sh35a20bd3, 32'sh35a054ed, 32'sh359e9de5, 32'sh359ce6bd, 32'sh359b2f73, 32'sh35997809, 
               32'sh3597c07d, 32'sh359608d1, 32'sh35945103, 32'sh35929914, 32'sh3590e104, 32'sh358f28d3, 32'sh358d7081, 32'sh358bb80e, 
               32'sh3589ff7a, 32'sh358846c5, 32'sh35868def, 32'sh3584d4f8, 32'sh35831be0, 32'sh358162a7, 32'sh357fa94d, 32'sh357defd2, 
               32'sh357c3636, 32'sh357a7c79, 32'sh3578c29b, 32'sh3577089c, 32'sh35754e7c, 32'sh3573943b, 32'sh3571d9d9, 32'sh35701f56, 
               32'sh356e64b2, 32'sh356ca9ed, 32'sh356aef08, 32'sh35693401, 32'sh356778d9, 32'sh3565bd90, 32'sh35640227, 32'sh3562469c, 
               32'sh35608af1, 32'sh355ecf25, 32'sh355d1337, 32'sh355b5729, 32'sh35599afa, 32'sh3557deaa, 32'sh35562239, 32'sh355465a7, 
               32'sh3552a8f4, 32'sh3550ec21, 32'sh354f2f2c, 32'sh354d7217, 32'sh354bb4e1, 32'sh3549f789, 32'sh35483a11, 32'sh35467c78, 
               32'sh3544bebf, 32'sh354300e4, 32'sh354142e9, 32'sh353f84cc, 32'sh353dc68f, 32'sh353c0831, 32'sh353a49b2, 32'sh35388b13, 
               32'sh3536cc52, 32'sh35350d71, 32'sh35334e6f, 32'sh35318f4c, 32'sh352fd008, 32'sh352e10a3, 32'sh352c511e, 32'sh352a9178, 
               32'sh3528d1b1, 32'sh352711c9, 32'sh352551c0, 32'sh35239197, 32'sh3521d14d, 32'sh352010e2, 32'sh351e5056, 32'sh351c8faa, 
               32'sh351acedd, 32'sh35190def, 32'sh35174ce0, 32'sh35158bb1, 32'sh3513ca60, 32'sh351208ef, 32'sh3510475e, 32'sh350e85ab, 
               32'sh350cc3d8, 32'sh350b01e4, 32'sh35093fd0, 32'sh35077d9a, 32'sh3505bb44, 32'sh3503f8ce, 32'sh35023636, 32'sh3500737e, 
               32'sh34feb0a5, 32'sh34fcedac, 32'sh34fb2a92, 32'sh34f96757, 32'sh34f7a3fb, 32'sh34f5e07f, 32'sh34f41ce2, 32'sh34f25924, 
               32'sh34f09546, 32'sh34eed147, 32'sh34ed0d28, 32'sh34eb48e8, 32'sh34e98487, 32'sh34e7c005, 32'sh34e5fb63, 32'sh34e436a1, 
               32'sh34e271bd, 32'sh34e0acb9, 32'sh34dee795, 32'sh34dd224f, 32'sh34db5cea, 32'sh34d99763, 32'sh34d7d1bc, 32'sh34d60bf5, 
               32'sh34d4460c, 32'sh34d28004, 32'sh34d0b9da, 32'sh34cef390, 32'sh34cd2d26, 32'sh34cb669b, 32'sh34c99fef, 32'sh34c7d923, 
               32'sh34c61236, 32'sh34c44b29, 32'sh34c283fb, 32'sh34c0bcac, 32'sh34bef53d, 32'sh34bd2dae, 32'sh34bb65fe, 32'sh34b99e2d, 
               32'sh34b7d63c, 32'sh34b60e2b, 32'sh34b445f8, 32'sh34b27da6, 32'sh34b0b533, 32'sh34aeec9f, 32'sh34ad23eb, 32'sh34ab5b16, 
               32'sh34a99221, 32'sh34a7c90c, 32'sh34a5ffd5, 32'sh34a4367f, 32'sh34a26d08, 32'sh34a0a370, 32'sh349ed9b8, 32'sh349d0fe0, 
               32'sh349b45e7, 32'sh34997bce, 32'sh3497b194, 32'sh3495e73a, 32'sh34941cbf, 32'sh34925224, 32'sh34908768, 32'sh348ebc8d, 
               32'sh348cf190, 32'sh348b2673, 32'sh34895b36, 32'sh34878fd9, 32'sh3485c45b, 32'sh3483f8bc, 32'sh34822cfd, 32'sh3480611e, 
               32'sh347e951f, 32'sh347cc8ff, 32'sh347afcbe, 32'sh3479305e, 32'sh347763dd, 32'sh3475973b, 32'sh3473ca79, 32'sh3471fd97, 
               32'sh34703095, 32'sh346e6372, 32'sh346c962f, 32'sh346ac8cb, 32'sh3468fb47, 32'sh34672da3, 32'sh34655fdf, 32'sh346391fa, 
               32'sh3461c3f5, 32'sh345ff5cf, 32'sh345e2789, 32'sh345c5923, 32'sh345a8a9d, 32'sh3458bbf6, 32'sh3456ed2f, 32'sh34551e48, 
               32'sh34534f41, 32'sh34518019, 32'sh344fb0d1, 32'sh344de168, 32'sh344c11e0, 32'sh344a4237, 32'sh3448726e, 32'sh3446a284, 
               32'sh3444d27b, 32'sh34430251, 32'sh34413207, 32'sh343f619c, 32'sh343d9112, 32'sh343bc067, 32'sh3439ef9c, 32'sh34381eb1, 
               32'sh34364da6, 32'sh34347c7a, 32'sh3432ab2e, 32'sh3430d9c2, 32'sh342f0836, 32'sh342d3689, 32'sh342b64bd, 32'sh342992d0, 
               32'sh3427c0c3, 32'sh3425ee96, 32'sh34241c49, 32'sh342249db, 32'sh3420774d, 32'sh341ea4a0, 32'sh341cd1d2, 32'sh341afee4, 
               32'sh34192bd5, 32'sh341758a7, 32'sh34158559, 32'sh3413b1ea, 32'sh3411de5b, 32'sh34100aac, 32'sh340e36dd, 32'sh340c62ee, 
               32'sh340a8edf, 32'sh3408bab0, 32'sh3406e660, 32'sh340511f1, 32'sh34033d61, 32'sh340168b2, 32'sh33ff93e2, 32'sh33fdbef2, 
               32'sh33fbe9e2, 32'sh33fa14b2, 32'sh33f83f62, 32'sh33f669f2, 32'sh33f49462, 32'sh33f2beb2, 32'sh33f0e8e2, 32'sh33ef12f2, 
               32'sh33ed3ce1, 32'sh33eb66b1, 32'sh33e99061, 32'sh33e7b9f0, 32'sh33e5e360, 32'sh33e40cb0, 32'sh33e235df, 32'sh33e05eef, 
               32'sh33de87de, 32'sh33dcb0ae, 32'sh33dad95e, 32'sh33d901ed, 32'sh33d72a5d, 32'sh33d552ac, 32'sh33d37adc, 32'sh33d1a2ec, 
               32'sh33cfcadc, 32'sh33cdf2ab, 32'sh33cc1a5b, 32'sh33ca41eb, 32'sh33c8695b, 32'sh33c690ab, 32'sh33c4b7db, 32'sh33c2deeb, 
               32'sh33c105db, 32'sh33bf2cac, 32'sh33bd535c, 32'sh33bb79ec, 32'sh33b9a05d, 32'sh33b7c6ae, 32'sh33b5ecde, 32'sh33b412ef, 
               32'sh33b238e0, 32'sh33b05eb1, 32'sh33ae8462, 32'sh33aca9f4, 32'sh33aacf65, 32'sh33a8f4b6, 32'sh33a719e8, 32'sh33a53efa, 
               32'sh33a363ec, 32'sh33a188be, 32'sh339fad70, 32'sh339dd203, 32'sh339bf675, 32'sh339a1ac8, 32'sh33983efb, 32'sh3396630e, 
               32'sh33948701, 32'sh3392aad4, 32'sh3390ce88, 32'sh338ef21c, 32'sh338d1590, 32'sh338b38e4, 32'sh33895c18, 32'sh33877f2d, 
               32'sh3385a222, 32'sh3383c4f7, 32'sh3381e7ac, 32'sh33800a42, 32'sh337e2cb7, 32'sh337c4f0d, 32'sh337a7144, 32'sh3378935a, 
               32'sh3376b551, 32'sh3374d728, 32'sh3372f8df, 32'sh33711a76, 32'sh336f3bee, 32'sh336d5d46, 32'sh336b7e7e, 32'sh33699f97, 
               32'sh3367c090, 32'sh3365e169, 32'sh33640223, 32'sh336222bc, 32'sh33604336, 32'sh335e6391, 32'sh335c83cb, 32'sh335aa3e6, 
               32'sh3358c3e2, 32'sh3356e3bd, 32'sh33550379, 32'sh33532316, 32'sh33514292, 32'sh334f61ef, 32'sh334d812d, 32'sh334ba04a, 
               32'sh3349bf48, 32'sh3347de27, 32'sh3345fce6, 32'sh33441b85, 32'sh33423a04, 32'sh33405864, 32'sh333e76a4, 32'sh333c94c5, 
               32'sh333ab2c6, 32'sh3338d0a8, 32'sh3336ee6a, 32'sh33350c0c, 32'sh3333298f, 32'sh333146f2, 32'sh332f6435, 32'sh332d8159, 
               32'sh332b9e5e, 32'sh3329bb43, 32'sh3327d808, 32'sh3325f4ae, 32'sh33241134, 32'sh33222d9a, 32'sh332049e1, 32'sh331e6609, 
               32'sh331c8211, 32'sh331a9dfa, 32'sh3318b9c2, 32'sh3316d56c, 32'sh3314f0f6, 32'sh33130c60, 32'sh331127ab, 32'sh330f42d7, 
               32'sh330d5de3, 32'sh330b78cf, 32'sh3309939c, 32'sh3307ae49, 32'sh3305c8d7, 32'sh3303e346, 32'sh3301fd95, 32'sh330017c4, 
               32'sh32fe31d5, 32'sh32fc4bc5, 32'sh32fa6596, 32'sh32f87f48, 32'sh32f698db, 32'sh32f4b24d, 32'sh32f2cba1, 32'sh32f0e4d5, 
               32'sh32eefdea, 32'sh32ed16df, 32'sh32eb2fb5, 32'sh32e9486b, 32'sh32e76102, 32'sh32e57979, 32'sh32e391d2, 32'sh32e1aa0a, 
               32'sh32dfc224, 32'sh32ddda1e, 32'sh32dbf1f8, 32'sh32da09b4, 32'sh32d82150, 32'sh32d638cc, 32'sh32d45029, 32'sh32d26767, 
               32'sh32d07e85, 32'sh32ce9585, 32'sh32ccac64, 32'sh32cac325, 32'sh32c8d9c6, 32'sh32c6f048, 32'sh32c506aa, 32'sh32c31ced, 
               32'sh32c13311, 32'sh32bf4916, 32'sh32bd5efb, 32'sh32bb74c1, 32'sh32b98a67, 32'sh32b79fef, 32'sh32b5b557, 32'sh32b3caa0, 
               32'sh32b1dfc9, 32'sh32aff4d3, 32'sh32ae09be, 32'sh32ac1e8a, 32'sh32aa3336, 32'sh32a847c4, 32'sh32a65c32, 32'sh32a47080, 
               32'sh32a284b0, 32'sh32a098c0, 32'sh329eacb1, 32'sh329cc083, 32'sh329ad435, 32'sh3298e7c9, 32'sh3296fb3d, 32'sh32950e92, 
               32'sh329321c7, 32'sh329134de, 32'sh328f47d5, 32'sh328d5aad, 32'sh328b6d66, 32'sh32898000, 32'sh3287927b, 32'sh3285a4d6, 
               32'sh3283b712, 32'sh3281c92f, 32'sh327fdb2d, 32'sh327ded0c, 32'sh327bfecc, 32'sh327a106c, 32'sh327821ee, 32'sh32763350, 
               32'sh32744493, 32'sh327255b7, 32'sh327066bc, 32'sh326e77a2, 32'sh326c8868, 32'sh326a9910, 32'sh3268a998, 32'sh3266ba02, 
               32'sh3264ca4c, 32'sh3262da77, 32'sh3260ea83, 32'sh325efa70, 32'sh325d0a3e, 32'sh325b19ed, 32'sh3259297d, 32'sh325738ee, 
               32'sh32554840, 32'sh32535772, 32'sh32516686, 32'sh324f757a, 32'sh324d8450, 32'sh324b9306, 32'sh3249a19e, 32'sh3247b016, 
               32'sh3245be70, 32'sh3243ccaa, 32'sh3241dac6, 32'sh323fe8c2, 32'sh323df6a0, 32'sh323c045e, 32'sh323a11fe, 32'sh32381f7e, 
               32'sh32362ce0, 32'sh32343a22, 32'sh32324746, 32'sh3230544a, 32'sh322e6130, 32'sh322c6df7, 32'sh322a7a9e, 32'sh32288727, 
               32'sh32269391, 32'sh32249fdc, 32'sh3222ac08, 32'sh3220b815, 32'sh321ec403, 32'sh321ccfd2, 32'sh321adb83, 32'sh3218e714, 
               32'sh3216f287, 32'sh3214fdda, 32'sh3213090f, 32'sh32111425, 32'sh320f1f1c, 32'sh320d29f4, 32'sh320b34ad, 32'sh32093f47, 
               32'sh320749c3, 32'sh3205541f, 32'sh32035e5d, 32'sh3201687c, 32'sh31ff727c, 32'sh31fd7c5d, 32'sh31fb8620, 32'sh31f98fc3, 
               32'sh31f79948, 32'sh31f5a2ae, 32'sh31f3abf5, 32'sh31f1b51d, 32'sh31efbe27, 32'sh31edc711, 32'sh31ebcfdd, 32'sh31e9d88a, 
               32'sh31e7e118, 32'sh31e5e988, 32'sh31e3f1d8, 32'sh31e1fa0a, 32'sh31e0021e, 32'sh31de0a12, 32'sh31dc11e8, 32'sh31da199e, 
               32'sh31d82137, 32'sh31d628b0, 32'sh31d4300b, 32'sh31d23746, 32'sh31d03e64, 32'sh31ce4562, 32'sh31cc4c42, 32'sh31ca5303, 
               32'sh31c859a5, 32'sh31c66029, 32'sh31c4668d, 32'sh31c26cd4, 32'sh31c072fb, 32'sh31be7904, 32'sh31bc7eee, 32'sh31ba84b9, 
               32'sh31b88a66, 32'sh31b68ff4, 32'sh31b49564, 32'sh31b29ab4, 32'sh31b09fe7, 32'sh31aea4fa, 32'sh31aca9ef, 32'sh31aaaec5, 
               32'sh31a8b37c, 32'sh31a6b815, 32'sh31a4bc90, 32'sh31a2c0eb, 32'sh31a0c528, 32'sh319ec947, 32'sh319ccd46, 32'sh319ad128, 
               32'sh3198d4ea, 32'sh3196d88e, 32'sh3194dc14, 32'sh3192df7a, 32'sh3190e2c3, 32'sh318ee5ec, 32'sh318ce8f7, 32'sh318aebe4, 
               32'sh3188eeb2, 32'sh3186f161, 32'sh3184f3f2, 32'sh3182f665, 32'sh3180f8b8, 32'sh317efaee, 32'sh317cfd04, 32'sh317afefc, 
               32'sh317900d6, 32'sh31770291, 32'sh3175042e, 32'sh317305ac, 32'sh3171070c, 32'sh316f084d, 32'sh316d096f, 32'sh316b0a74, 
               32'sh31690b59, 32'sh31670c20, 32'sh31650cc9, 32'sh31630d53, 32'sh31610dbf, 32'sh315f0e0c, 32'sh315d0e3b, 32'sh315b0e4c, 
               32'sh31590e3e, 32'sh31570e11, 32'sh31550dc6, 32'sh31530d5d, 32'sh31510cd5, 32'sh314f0c2f, 32'sh314d0b6a, 32'sh314b0a87, 
               32'sh31490986, 32'sh31470866, 32'sh31450728, 32'sh314305cb, 32'sh31410450, 32'sh313f02b7, 32'sh313d00ff, 32'sh313aff29, 
               32'sh3138fd35, 32'sh3136fb22, 32'sh3134f8f1, 32'sh3132f6a1, 32'sh3130f433, 32'sh312ef1a7, 32'sh312ceefc, 32'sh312aec33, 
               32'sh3128e94c, 32'sh3126e646, 32'sh3124e322, 32'sh3122dfe0, 32'sh3120dc80, 32'sh311ed901, 32'sh311cd564, 32'sh311ad1a8, 
               32'sh3118cdcf, 32'sh3116c9d7, 32'sh3114c5c0, 32'sh3112c18c, 32'sh3110bd39, 32'sh310eb8c8, 32'sh310cb438, 32'sh310aaf8b, 
               32'sh3108aabf, 32'sh3106a5d5, 32'sh3104a0cc, 32'sh31029ba6, 32'sh31009661, 32'sh30fe90fe, 32'sh30fc8b7d, 32'sh30fa85dd, 
               32'sh30f8801f, 32'sh30f67a44, 32'sh30f47449, 32'sh30f26e31, 32'sh30f067fb, 32'sh30ee61a6, 32'sh30ec5b33, 32'sh30ea54a2, 
               32'sh30e84df3, 32'sh30e64725, 32'sh30e4403a, 32'sh30e23930, 32'sh30e03208, 32'sh30de2ac2, 32'sh30dc235e, 32'sh30da1bdc, 
               32'sh30d8143b, 32'sh30d60c7d, 32'sh30d404a0, 32'sh30d1fca5, 32'sh30cff48c, 32'sh30cdec55, 32'sh30cbe400, 32'sh30c9db8d, 
               32'sh30c7d2fb, 32'sh30c5ca4c, 32'sh30c3c17e, 32'sh30c1b893, 32'sh30bfaf89, 32'sh30bda661, 32'sh30bb9d1c, 32'sh30b993b8, 
               32'sh30b78a36, 32'sh30b58096, 32'sh30b376d8, 32'sh30b16cfc, 32'sh30af6302, 32'sh30ad58ea, 32'sh30ab4eb3, 32'sh30a9445f, 
               32'sh30a739ed, 32'sh30a52f5d, 32'sh30a324af, 32'sh30a119e2, 32'sh309f0ef8, 32'sh309d03f0, 32'sh309af8ca, 32'sh3098ed86, 
               32'sh3096e223, 32'sh3094d6a3, 32'sh3092cb05, 32'sh3090bf49, 32'sh308eb36f, 32'sh308ca777, 32'sh308a9b61, 32'sh30888f2d, 
               32'sh308682dc, 32'sh3084766c, 32'sh308269de, 32'sh30805d33, 32'sh307e5069, 32'sh307c4382, 32'sh307a367c, 32'sh30782959, 
               32'sh30761c18, 32'sh30740eb9, 32'sh3072013c, 32'sh306ff3a1, 32'sh306de5e9, 32'sh306bd812, 32'sh3069ca1e, 32'sh3067bc0b, 
               32'sh3065addb, 32'sh30639f8d, 32'sh30619121, 32'sh305f8298, 32'sh305d73f0, 32'sh305b652b, 32'sh30595648, 32'sh30574747, 
               32'sh30553828, 32'sh305328eb, 32'sh30511991, 32'sh304f0a19, 32'sh304cfa83, 32'sh304aeacf, 32'sh3048dafd, 32'sh3046cb0e, 
               32'sh3044bb00, 32'sh3042aad5, 32'sh30409a8d, 32'sh303e8a26, 32'sh303c79a2, 32'sh303a6900, 32'sh30385840, 32'sh30364763, 
               32'sh30343667, 32'sh3032254e, 32'sh30301418, 32'sh302e02c3, 32'sh302bf151, 32'sh3029dfc1, 32'sh3027ce14, 32'sh3025bc48, 
               32'sh3023aa5f, 32'sh30219859, 32'sh301f8634, 32'sh301d73f2, 32'sh301b6193, 32'sh30194f15, 32'sh30173c7a, 32'sh301529c1, 
               32'sh301316eb, 32'sh301103f7, 32'sh300ef0e5, 32'sh300cddb6, 32'sh300aca69, 32'sh3008b6fe, 32'sh3006a376, 32'sh30048fd0, 
               32'sh30027c0c, 32'sh3000682b, 32'sh2ffe542d, 32'sh2ffc4010, 32'sh2ffa2bd6, 32'sh2ff8177f, 32'sh2ff6030a, 32'sh2ff3ee77, 
               32'sh2ff1d9c7, 32'sh2fefc4f9, 32'sh2fedb00d, 32'sh2feb9b04, 32'sh2fe985de, 32'sh2fe7709a, 32'sh2fe55b38, 32'sh2fe345b9, 
               32'sh2fe1301c, 32'sh2fdf1a62, 32'sh2fdd048a, 32'sh2fdaee95, 32'sh2fd8d882, 32'sh2fd6c252, 32'sh2fd4ac04, 32'sh2fd29598, 
               32'sh2fd07f0f, 32'sh2fce6869, 32'sh2fcc51a5, 32'sh2fca3ac4, 32'sh2fc823c5, 32'sh2fc60ca9, 32'sh2fc3f56f, 32'sh2fc1de18, 
               32'sh2fbfc6a3, 32'sh2fbdaf11, 32'sh2fbb9761, 32'sh2fb97f94, 32'sh2fb767aa, 32'sh2fb54fa2, 32'sh2fb3377c, 32'sh2fb11f3a, 
               32'sh2faf06da, 32'sh2facee5c, 32'sh2faad5c1, 32'sh2fa8bd09, 32'sh2fa6a433, 32'sh2fa48b40, 32'sh2fa2722f, 32'sh2fa05901, 
               32'sh2f9e3fb6, 32'sh2f9c264d, 32'sh2f9a0cc7, 32'sh2f97f323, 32'sh2f95d963, 32'sh2f93bf84, 32'sh2f91a589, 32'sh2f8f8b70, 
               32'sh2f8d713a, 32'sh2f8b56e6, 32'sh2f893c75, 32'sh2f8721e7, 32'sh2f85073c, 32'sh2f82ec73, 32'sh2f80d18d, 32'sh2f7eb689, 
               32'sh2f7c9b69, 32'sh2f7a802b, 32'sh2f7864cf, 32'sh2f764957, 32'sh2f742dc1, 32'sh2f72120e, 32'sh2f6ff63d, 32'sh2f6dda50, 
               32'sh2f6bbe45, 32'sh2f69a21d, 32'sh2f6785d7, 32'sh2f656975, 32'sh2f634cf5, 32'sh2f613058, 32'sh2f5f139d, 32'sh2f5cf6c6, 
               32'sh2f5ad9d1, 32'sh2f58bcbf, 32'sh2f569f90, 32'sh2f548243, 32'sh2f5264da, 32'sh2f504753, 32'sh2f4e29af, 32'sh2f4c0bee, 
               32'sh2f49ee0f, 32'sh2f47d014, 32'sh2f45b1fb, 32'sh2f4393c6, 32'sh2f417573, 32'sh2f3f5702, 32'sh2f3d3875, 32'sh2f3b19cb, 
               32'sh2f38fb03, 32'sh2f36dc1f, 32'sh2f34bd1d, 32'sh2f329dfe, 32'sh2f307ec2, 32'sh2f2e5f69, 32'sh2f2c3ff2, 32'sh2f2a205f, 
               32'sh2f2800af, 32'sh2f25e0e1, 32'sh2f23c0f6, 32'sh2f21a0ef, 32'sh2f1f80ca, 32'sh2f1d6088, 32'sh2f1b4029, 32'sh2f191fad, 
               32'sh2f16ff14, 32'sh2f14de5e, 32'sh2f12bd8b, 32'sh2f109c9b, 32'sh2f0e7b8e, 32'sh2f0c5a64, 32'sh2f0a391d, 32'sh2f0817b8, 
               32'sh2f05f637, 32'sh2f03d499, 32'sh2f01b2de, 32'sh2eff9105, 32'sh2efd6f10, 32'sh2efb4cfe, 32'sh2ef92acf, 32'sh2ef70883, 
               32'sh2ef4e619, 32'sh2ef2c393, 32'sh2ef0a0f0, 32'sh2eee7e30, 32'sh2eec5b53, 32'sh2eea3859, 32'sh2ee81543, 32'sh2ee5f20f, 
               32'sh2ee3cebe, 32'sh2ee1ab50, 32'sh2edf87c6, 32'sh2edd641e, 32'sh2edb405a, 32'sh2ed91c79, 32'sh2ed6f87a, 32'sh2ed4d45f, 
               32'sh2ed2b027, 32'sh2ed08bd3, 32'sh2ece6761, 32'sh2ecc42d2, 32'sh2eca1e27, 32'sh2ec7f95e, 32'sh2ec5d479, 32'sh2ec3af77, 
               32'sh2ec18a58, 32'sh2ebf651d, 32'sh2ebd3fc4, 32'sh2ebb1a4f, 32'sh2eb8f4bc, 32'sh2eb6cf0d, 32'sh2eb4a942, 32'sh2eb28359, 
               32'sh2eb05d53, 32'sh2eae3731, 32'sh2eac10f2, 32'sh2ea9ea96, 32'sh2ea7c41e, 32'sh2ea59d88, 32'sh2ea376d6, 32'sh2ea15007, 
               32'sh2e9f291b, 32'sh2e9d0213, 32'sh2e9adaee, 32'sh2e98b3ac, 32'sh2e968c4d, 32'sh2e9464d1, 32'sh2e923d39, 32'sh2e901584, 
               32'sh2e8dedb3, 32'sh2e8bc5c4, 32'sh2e899db9, 32'sh2e877591, 32'sh2e854d4d, 32'sh2e8324ec, 32'sh2e80fc6e, 32'sh2e7ed3d3, 
               32'sh2e7cab1c, 32'sh2e7a8248, 32'sh2e785958, 32'sh2e76304a, 32'sh2e740720, 32'sh2e71ddda, 32'sh2e6fb477, 32'sh2e6d8af7, 
               32'sh2e6b615a, 32'sh2e6937a1, 32'sh2e670dcb, 32'sh2e64e3d9, 32'sh2e62b9ca, 32'sh2e608f9e, 32'sh2e5e6556, 32'sh2e5c3af1, 
               32'sh2e5a1070, 32'sh2e57e5d2, 32'sh2e55bb17, 32'sh2e539040, 32'sh2e51654c, 32'sh2e4f3a3c, 32'sh2e4d0f0f, 32'sh2e4ae3c6, 
               32'sh2e48b860, 32'sh2e468cdd, 32'sh2e44613e, 32'sh2e423582, 32'sh2e4009aa, 32'sh2e3dddb5, 32'sh2e3bb1a4, 32'sh2e398576, 
               32'sh2e37592c, 32'sh2e352cc5, 32'sh2e330042, 32'sh2e30d3a2, 32'sh2e2ea6e6, 32'sh2e2c7a0d, 32'sh2e2a4d18, 32'sh2e282006, 
               32'sh2e25f2d8, 32'sh2e23c58d, 32'sh2e219826, 32'sh2e1f6aa3, 32'sh2e1d3d03, 32'sh2e1b0f46, 32'sh2e18e16d, 32'sh2e16b378, 
               32'sh2e148566, 32'sh2e125738, 32'sh2e1028ed, 32'sh2e0dfa86, 32'sh2e0bcc03, 32'sh2e099d63, 32'sh2e076ea7, 32'sh2e053fce, 
               32'sh2e0310d9, 32'sh2e00e1c8, 32'sh2dfeb29a, 32'sh2dfc8350, 32'sh2dfa53e9, 32'sh2df82466, 32'sh2df5f4c7, 32'sh2df3c50c, 
               32'sh2df19534, 32'sh2def653f, 32'sh2ded352f, 32'sh2deb0502, 32'sh2de8d4b8, 32'sh2de6a453, 32'sh2de473d1, 32'sh2de24333, 
               32'sh2de01278, 32'sh2ddde1a1, 32'sh2ddbb0ae, 32'sh2dd97f9f, 32'sh2dd74e73, 32'sh2dd51d2b, 32'sh2dd2ebc7, 32'sh2dd0ba47, 
               32'sh2dce88aa, 32'sh2dcc56f1, 32'sh2dca251c, 32'sh2dc7f32a, 32'sh2dc5c11c, 32'sh2dc38ef2, 32'sh2dc15cac, 32'sh2dbf2a4a, 
               32'sh2dbcf7cb, 32'sh2dbac530, 32'sh2db89279, 32'sh2db65fa6, 32'sh2db42cb6, 32'sh2db1f9ab, 32'sh2dafc683, 32'sh2dad933f, 
               32'sh2dab5fdf, 32'sh2da92c62, 32'sh2da6f8ca, 32'sh2da4c515, 32'sh2da29144, 32'sh2da05d57, 32'sh2d9e294e, 32'sh2d9bf529, 
               32'sh2d99c0e7, 32'sh2d978c8a, 32'sh2d955810, 32'sh2d93237a, 32'sh2d90eec8, 32'sh2d8eb9fa, 32'sh2d8c8510, 32'sh2d8a500a, 
               32'sh2d881ae8, 32'sh2d85e5a9, 32'sh2d83b04f, 32'sh2d817ad8, 32'sh2d7f4545, 32'sh2d7d0f97, 32'sh2d7ad9cc, 32'sh2d78a3e5, 
               32'sh2d766de2, 32'sh2d7437c3, 32'sh2d720189, 32'sh2d6fcb32, 32'sh2d6d94bf, 32'sh2d6b5e30, 32'sh2d692784, 32'sh2d66f0bd, 
               32'sh2d64b9da, 32'sh2d6282db, 32'sh2d604bc0, 32'sh2d5e1489, 32'sh2d5bdd36, 32'sh2d59a5c7, 32'sh2d576e3c, 32'sh2d553695, 
               32'sh2d52fed2, 32'sh2d50c6f3, 32'sh2d4e8ef9, 32'sh2d4c56e2, 32'sh2d4a1eaf, 32'sh2d47e661, 32'sh2d45adf6, 32'sh2d43756f, 
               32'sh2d413ccd, 32'sh2d3f040f, 32'sh2d3ccb34, 32'sh2d3a923e, 32'sh2d38592c, 32'sh2d361ffe, 32'sh2d33e6b4, 32'sh2d31ad4f, 
               32'sh2d2f73cd, 32'sh2d2d3a30, 32'sh2d2b0076, 32'sh2d28c6a1, 32'sh2d268cb0, 32'sh2d2452a3, 32'sh2d22187a, 32'sh2d1fde36, 
               32'sh2d1da3d5, 32'sh2d1b6959, 32'sh2d192ec1, 32'sh2d16f40d, 32'sh2d14b93d, 32'sh2d127e52, 32'sh2d10434a, 32'sh2d0e0827, 
               32'sh2d0bcce8, 32'sh2d09918e, 32'sh2d075617, 32'sh2d051a85, 32'sh2d02ded7, 32'sh2d00a30d, 32'sh2cfe6728, 32'sh2cfc2b26, 
               32'sh2cf9ef09, 32'sh2cf7b2d0, 32'sh2cf5767c, 32'sh2cf33a0c, 32'sh2cf0fd80, 32'sh2ceec0d8, 32'sh2cec8414, 32'sh2cea4735, 
               32'sh2ce80a3a, 32'sh2ce5cd24, 32'sh2ce38ff1, 32'sh2ce152a4, 32'sh2cdf153a, 32'sh2cdcd7b5, 32'sh2cda9a14, 32'sh2cd85c57, 
               32'sh2cd61e7f, 32'sh2cd3e08b, 32'sh2cd1a27b, 32'sh2ccf6450, 32'sh2ccd2609, 32'sh2ccae7a6, 32'sh2cc8a928, 32'sh2cc66a8e, 
               32'sh2cc42bd9, 32'sh2cc1ed08, 32'sh2cbfae1b, 32'sh2cbd6f13, 32'sh2cbb2fef, 32'sh2cb8f0b0, 32'sh2cb6b155, 32'sh2cb471de, 
               32'sh2cb2324c, 32'sh2caff29e, 32'sh2cadb2d5, 32'sh2cab72f0, 32'sh2ca932ef, 32'sh2ca6f2d4, 32'sh2ca4b29c, 32'sh2ca27249, 
               32'sh2ca031da, 32'sh2c9df150, 32'sh2c9bb0ab, 32'sh2c996fe9, 32'sh2c972f0d, 32'sh2c94ee15, 32'sh2c92ad01, 32'sh2c906bd2, 
               32'sh2c8e2a87, 32'sh2c8be921, 32'sh2c89a79f, 32'sh2c876602, 32'sh2c85244a, 32'sh2c82e276, 32'sh2c80a086, 32'sh2c7e5e7b, 
               32'sh2c7c1c55, 32'sh2c79da13, 32'sh2c7797b6, 32'sh2c75553d, 32'sh2c7312a9, 32'sh2c70cff9, 32'sh2c6e8d2e, 32'sh2c6c4a48, 
               32'sh2c6a0746, 32'sh2c67c429, 32'sh2c6580f1, 32'sh2c633d9d, 32'sh2c60fa2d, 32'sh2c5eb6a3, 32'sh2c5c72fd, 32'sh2c5a2f3b, 
               32'sh2c57eb5e, 32'sh2c55a766, 32'sh2c536353, 32'sh2c511f24, 32'sh2c4edada, 32'sh2c4c9674, 32'sh2c4a51f3, 32'sh2c480d57, 
               32'sh2c45c8a0, 32'sh2c4383cd, 32'sh2c413edf, 32'sh2c3ef9d6, 32'sh2c3cb4b1, 32'sh2c3a6f71, 32'sh2c382a16, 32'sh2c35e49f, 
               32'sh2c339f0e, 32'sh2c315961, 32'sh2c2f1398, 32'sh2c2ccdb5, 32'sh2c2a87b6, 32'sh2c28419c, 32'sh2c25fb66, 32'sh2c23b516, 
               32'sh2c216eaa, 32'sh2c1f2823, 32'sh2c1ce181, 32'sh2c1a9ac4, 32'sh2c1853eb, 32'sh2c160cf7, 32'sh2c13c5e8, 32'sh2c117ebe, 
               32'sh2c0f3779, 32'sh2c0cf018, 32'sh2c0aa89c, 32'sh2c086106, 32'sh2c061953, 32'sh2c03d186, 32'sh2c01899e, 32'sh2bff419a, 
               32'sh2bfcf97c, 32'sh2bfab142, 32'sh2bf868ed, 32'sh2bf6207d, 32'sh2bf3d7f2, 32'sh2bf18f4c, 32'sh2bef468a, 32'sh2becfdae, 
               32'sh2beab4b6, 32'sh2be86ba4, 32'sh2be62276, 32'sh2be3d92d, 32'sh2be18fc9, 32'sh2bdf464a, 32'sh2bdcfcb0, 32'sh2bdab2fb, 
               32'sh2bd8692b, 32'sh2bd61f40, 32'sh2bd3d53a, 32'sh2bd18b18, 32'sh2bcf40dc, 32'sh2bccf685, 32'sh2bcaac12, 32'sh2bc86185, 
               32'sh2bc616dd, 32'sh2bc3cc19, 32'sh2bc1813b, 32'sh2bbf3642, 32'sh2bbceb2d, 32'sh2bba9ffe, 32'sh2bb854b4, 32'sh2bb6094f, 
               32'sh2bb3bdce, 32'sh2bb17233, 32'sh2baf267d, 32'sh2bacdaac, 32'sh2baa8ec0, 32'sh2ba842b9, 32'sh2ba5f697, 32'sh2ba3aa5b, 
               32'sh2ba15e03, 32'sh2b9f1190, 32'sh2b9cc503, 32'sh2b9a785a, 32'sh2b982b97, 32'sh2b95deb9, 32'sh2b9391c0, 32'sh2b9144ac, 
               32'sh2b8ef77d, 32'sh2b8caa33, 32'sh2b8a5cce, 32'sh2b880f4f, 32'sh2b85c1b5, 32'sh2b837400, 32'sh2b812630, 32'sh2b7ed845, 
               32'sh2b7c8a3f, 32'sh2b7a3c1f, 32'sh2b77ede3, 32'sh2b759f8d, 32'sh2b73511c, 32'sh2b710291, 32'sh2b6eb3ea, 32'sh2b6c6529, 
               32'sh2b6a164d, 32'sh2b67c756, 32'sh2b657844, 32'sh2b632918, 32'sh2b60d9d0, 32'sh2b5e8a6f, 32'sh2b5c3af2, 32'sh2b59eb5a, 
               32'sh2b579ba8, 32'sh2b554bdb, 32'sh2b52fbf4, 32'sh2b50abf1, 32'sh2b4e5bd4, 32'sh2b4c0b9c, 32'sh2b49bb4a, 32'sh2b476add, 
               32'sh2b451a55, 32'sh2b42c9b2, 32'sh2b4078f5, 32'sh2b3e281d, 32'sh2b3bd72a, 32'sh2b39861d, 32'sh2b3734f5, 32'sh2b34e3b2, 
               32'sh2b329255, 32'sh2b3040dd, 32'sh2b2def4b, 32'sh2b2b9d9d, 32'sh2b294bd5, 32'sh2b26f9f3, 32'sh2b24a7f6, 32'sh2b2255de, 
               32'sh2b2003ac, 32'sh2b1db15f, 32'sh2b1b5ef8, 32'sh2b190c75, 32'sh2b16b9d9, 32'sh2b146722, 32'sh2b121450, 32'sh2b0fc163, 
               32'sh2b0d6e5c, 32'sh2b0b1b3b, 32'sh2b08c7ff, 32'sh2b0674a8, 32'sh2b042137, 32'sh2b01cdab, 32'sh2aff7a05, 32'sh2afd2644, 
               32'sh2afad269, 32'sh2af87e73, 32'sh2af62a63, 32'sh2af3d638, 32'sh2af181f3, 32'sh2aef2d93, 32'sh2aecd919, 32'sh2aea8484, 
               32'sh2ae82fd5, 32'sh2ae5db0b, 32'sh2ae38627, 32'sh2ae13129, 32'sh2adedc10, 32'sh2adc86dc, 32'sh2ada318e, 32'sh2ad7dc26, 
               32'sh2ad586a3, 32'sh2ad33106, 32'sh2ad0db4e, 32'sh2ace857c, 32'sh2acc2f90, 32'sh2ac9d989, 32'sh2ac78368, 32'sh2ac52d2c, 
               32'sh2ac2d6d6, 32'sh2ac08066, 32'sh2abe29db, 32'sh2abbd336, 32'sh2ab97c77, 32'sh2ab7259d, 32'sh2ab4cea9, 32'sh2ab2779a, 
               32'sh2ab02071, 32'sh2aadc92e, 32'sh2aab71d0, 32'sh2aa91a59, 32'sh2aa6c2c6, 32'sh2aa46b1a, 32'sh2aa21353, 32'sh2a9fbb72, 
               32'sh2a9d6377, 32'sh2a9b0b61, 32'sh2a98b331, 32'sh2a965ae7, 32'sh2a940283, 32'sh2a91aa04, 32'sh2a8f516b, 32'sh2a8cf8b8, 
               32'sh2a8a9fea, 32'sh2a884702, 32'sh2a85ee00, 32'sh2a8394e4, 32'sh2a813bae, 32'sh2a7ee25d, 32'sh2a7c88f2, 32'sh2a7a2f6d, 
               32'sh2a77d5ce, 32'sh2a757c15, 32'sh2a732241, 32'sh2a70c853, 32'sh2a6e6e4b, 32'sh2a6c1429, 32'sh2a69b9ec, 32'sh2a675f96, 
               32'sh2a650525, 32'sh2a62aa9a, 32'sh2a604ff5, 32'sh2a5df536, 32'sh2a5b9a5d, 32'sh2a593f6a, 32'sh2a56e45c, 32'sh2a548935, 
               32'sh2a522df3, 32'sh2a4fd297, 32'sh2a4d7721, 32'sh2a4b1b91, 32'sh2a48bfe7, 32'sh2a466423, 32'sh2a440844, 32'sh2a41ac4c, 
               32'sh2a3f503a, 32'sh2a3cf40d, 32'sh2a3a97c7, 32'sh2a383b66, 32'sh2a35deeb, 32'sh2a338257, 32'sh2a3125a8, 32'sh2a2ec8df, 
               32'sh2a2c6bfd, 32'sh2a2a0f00, 32'sh2a27b1e9, 32'sh2a2554b8, 32'sh2a22f76e, 32'sh2a209a09, 32'sh2a1e3c8a, 32'sh2a1bdef1, 
               32'sh2a19813f, 32'sh2a172372, 32'sh2a14c58b, 32'sh2a12678b, 32'sh2a100970, 32'sh2a0dab3c, 32'sh2a0b4ced, 32'sh2a08ee85, 
               32'sh2a069003, 32'sh2a043166, 32'sh2a01d2b0, 32'sh29ff73e0, 32'sh29fd14f6, 32'sh29fab5f3, 32'sh29f856d5, 32'sh29f5f79d, 
               32'sh29f3984c, 32'sh29f138e0, 32'sh29eed95b, 32'sh29ec79bc, 32'sh29ea1a03, 32'sh29e7ba30, 32'sh29e55a43, 32'sh29e2fa3d, 
               32'sh29e09a1c, 32'sh29de39e2, 32'sh29dbd98e, 32'sh29d97920, 32'sh29d71899, 32'sh29d4b7f7, 32'sh29d2573c, 32'sh29cff667, 
               32'sh29cd9578, 32'sh29cb346f, 32'sh29c8d34d, 32'sh29c67210, 32'sh29c410ba, 32'sh29c1af4b, 32'sh29bf4dc1, 32'sh29bcec1e, 
               32'sh29ba8a61, 32'sh29b8288a, 32'sh29b5c69a, 32'sh29b3648f, 32'sh29b1026c, 32'sh29aea02e, 32'sh29ac3dd7, 32'sh29a9db65, 
               32'sh29a778db, 32'sh29a51636, 32'sh29a2b378, 32'sh29a050a0, 32'sh299dedaf, 32'sh299b8aa4, 32'sh2999277f, 32'sh2996c440, 
               32'sh299460e8, 32'sh2991fd76, 32'sh298f99eb, 32'sh298d3646, 32'sh298ad287, 32'sh29886eaf, 32'sh29860abd, 32'sh2983a6b1, 
               32'sh2981428c, 32'sh297ede4d, 32'sh297c79f5, 32'sh297a1583, 32'sh2977b0f7, 32'sh29754c52, 32'sh2972e793, 32'sh297082bb, 
               32'sh296e1dc9, 32'sh296bb8be, 32'sh29695399, 32'sh2966ee5a, 32'sh29648902, 32'sh29622391, 32'sh295fbe06, 32'sh295d5861, 
               32'sh295af2a3, 32'sh29588ccb, 32'sh295626da, 32'sh2953c0cf, 32'sh29515aab, 32'sh294ef46e, 32'sh294c8e16, 32'sh294a27a6, 
               32'sh2947c11c, 32'sh29455a78, 32'sh2942f3bb, 32'sh29408ce5, 32'sh293e25f5, 32'sh293bbeec, 32'sh293957c9, 32'sh2936f08d, 
               32'sh29348937, 32'sh293221c8, 32'sh292fba40, 32'sh292d529e, 32'sh292aeae3, 32'sh2928830e, 32'sh29261b20, 32'sh2923b319, 
               32'sh29214af8, 32'sh291ee2be, 32'sh291c7a6a, 32'sh291a11fd, 32'sh2917a977, 32'sh291540d8, 32'sh2912d81f, 32'sh29106f4c, 
               32'sh290e0661, 32'sh290b9d5c, 32'sh2909343e, 32'sh2906cb06, 32'sh290461b5, 32'sh2901f84b, 32'sh28ff8ec8, 32'sh28fd252b, 
               32'sh28fabb75, 32'sh28f851a6, 32'sh28f5e7bd, 32'sh28f37dbb, 32'sh28f113a0, 32'sh28eea96c, 32'sh28ec3f1e, 32'sh28e9d4b7, 
               32'sh28e76a37, 32'sh28e4ff9e, 32'sh28e294eb, 32'sh28e02a20, 32'sh28ddbf3b, 32'sh28db543c, 32'sh28d8e925, 32'sh28d67df4, 
               32'sh28d412ab, 32'sh28d1a748, 32'sh28cf3bcc, 32'sh28ccd036, 32'sh28ca6488, 32'sh28c7f8c0, 32'sh28c58cdf, 32'sh28c320e5, 
               32'sh28c0b4d2, 32'sh28be48a6, 32'sh28bbdc61, 32'sh28b97002, 32'sh28b7038b, 32'sh28b496fa, 32'sh28b22a50, 32'sh28afbd8d, 
               32'sh28ad50b1, 32'sh28aae3bc, 32'sh28a876ae, 32'sh28a60987, 32'sh28a39c46, 32'sh28a12eed, 32'sh289ec17a, 32'sh289c53ef, 
               32'sh2899e64a, 32'sh2897788c, 32'sh28950ab6, 32'sh28929cc6, 32'sh28902ebd, 32'sh288dc09c, 32'sh288b5261, 32'sh2888e40d, 
               32'sh288675a0, 32'sh2884071a, 32'sh2881987c, 32'sh287f29c4, 32'sh287cbaf3, 32'sh287a4c09, 32'sh2877dd07, 32'sh28756deb, 
               32'sh2872feb6, 32'sh28708f69, 32'sh286e2002, 32'sh286bb083, 32'sh286940ea, 32'sh2866d139, 32'sh2864616f, 32'sh2861f18c, 
               32'sh285f8190, 32'sh285d117b, 32'sh285aa14d, 32'sh28583106, 32'sh2855c0a6, 32'sh2853502e, 32'sh2850df9d, 32'sh284e6ef2, 
               32'sh284bfe2f, 32'sh28498d53, 32'sh28471c5e, 32'sh2844ab51, 32'sh28423a2a, 32'sh283fc8eb, 32'sh283d5793, 32'sh283ae622, 
               32'sh28387498, 32'sh283602f5, 32'sh2833913a, 32'sh28311f65, 32'sh282ead78, 32'sh282c3b73, 32'sh2829c954, 32'sh2827571d, 
               32'sh2824e4cc, 32'sh28227264, 32'sh281fffe2, 32'sh281d8d48, 32'sh281b1a94, 32'sh2818a7c8, 32'sh281634e4, 32'sh2813c1e6, 
               32'sh28114ed0, 32'sh280edba2, 32'sh280c685a, 32'sh2809f4fa, 32'sh28078181, 32'sh28050def, 32'sh28029a45, 32'sh28002682, 
               32'sh27fdb2a7, 32'sh27fb3eb2, 32'sh27f8caa5, 32'sh27f65680, 32'sh27f3e241, 32'sh27f16dea, 32'sh27eef97b, 32'sh27ec84f3, 
               32'sh27ea1052, 32'sh27e79b98, 32'sh27e526c6, 32'sh27e2b1dc, 32'sh27e03cd8, 32'sh27ddc7bd, 32'sh27db5288, 32'sh27d8dd3b, 
               32'sh27d667d5, 32'sh27d3f257, 32'sh27d17cc1, 32'sh27cf0711, 32'sh27cc9149, 32'sh27ca1b69, 32'sh27c7a570, 32'sh27c52f5e, 
               32'sh27c2b934, 32'sh27c042f2, 32'sh27bdcc97, 32'sh27bb5623, 32'sh27b8df97, 32'sh27b668f2, 32'sh27b3f235, 32'sh27b17b60, 
               32'sh27af0472, 32'sh27ac8d6b, 32'sh27aa164c, 32'sh27a79f14, 32'sh27a527c4, 32'sh27a2b05c, 32'sh27a038db, 32'sh279dc142, 
               32'sh279b4990, 32'sh2798d1c6, 32'sh279659e3, 32'sh2793e1e8, 32'sh279169d5, 32'sh278ef1a9, 32'sh278c7965, 32'sh278a0108, 
               32'sh27878893, 32'sh27851006, 32'sh27829760, 32'sh27801ea2, 32'sh277da5cb, 32'sh277b2cdc, 32'sh2778b3d5, 32'sh27763ab5, 
               32'sh2773c17d, 32'sh2771482d, 32'sh276ecec5, 32'sh276c5544, 32'sh2769dbaa, 32'sh276761f9, 32'sh2764e82f, 32'sh27626e4d, 
               32'sh275ff452, 32'sh275d7a40, 32'sh275b0014, 32'sh275885d1, 32'sh27560b76, 32'sh27539102, 32'sh27511676, 32'sh274e9bd1, 
               32'sh274c2115, 32'sh2749a640, 32'sh27472b53, 32'sh2744b04d, 32'sh27423530, 32'sh273fb9fa, 32'sh273d3eac, 32'sh273ac346, 
               32'sh273847c8, 32'sh2735cc31, 32'sh27335082, 32'sh2730d4bb, 32'sh272e58dc, 32'sh272bdce5, 32'sh272960d6, 32'sh2726e4ae, 
               32'sh2724686e, 32'sh2721ec16, 32'sh271f6fa6, 32'sh271cf31e, 32'sh271a767e, 32'sh2717f9c6, 32'sh27157cf5, 32'sh2713000c, 
               32'sh2710830c, 32'sh270e05f3, 32'sh270b88c2, 32'sh27090b79, 32'sh27068e18, 32'sh2704109f, 32'sh2701930e, 32'sh26ff1564, 
               32'sh26fc97a3, 32'sh26fa19ca, 32'sh26f79bd8, 32'sh26f51dcf, 32'sh26f29fad, 32'sh26f02174, 32'sh26eda322, 32'sh26eb24b9, 
               32'sh26e8a637, 32'sh26e6279d, 32'sh26e3a8ec, 32'sh26e12a22, 32'sh26deab41, 32'sh26dc2c47, 32'sh26d9ad36, 32'sh26d72e0c, 
               32'sh26d4aecb, 32'sh26d22f72, 32'sh26cfb000, 32'sh26cd3077, 32'sh26cab0d6, 32'sh26c8311d, 32'sh26c5b14c, 32'sh26c33163, 
               32'sh26c0b162, 32'sh26be3149, 32'sh26bbb119, 32'sh26b930d0, 32'sh26b6b070, 32'sh26b42ff7, 32'sh26b1af67, 32'sh26af2ebf, 
               32'sh26acadff, 32'sh26aa2d27, 32'sh26a7ac38, 32'sh26a52b30, 32'sh26a2aa11, 32'sh26a028da, 32'sh269da78b, 32'sh269b2624, 
               32'sh2698a4a6, 32'sh2696230f, 32'sh2693a161, 32'sh26911f9b, 32'sh268e9dbd, 32'sh268c1bc8, 32'sh268999ba, 32'sh26871795, 
               32'sh26849558, 32'sh26821303, 32'sh267f9097, 32'sh267d0e13, 32'sh267a8b77, 32'sh267808c3, 32'sh267585f8, 32'sh26730315, 
               32'sh2670801a, 32'sh266dfd08, 32'sh266b79dd, 32'sh2668f69b, 32'sh26667342, 32'sh2663efd1, 32'sh26616c48, 32'sh265ee8a7, 
               32'sh265c64ef, 32'sh2659e11f, 32'sh26575d37, 32'sh2654d938, 32'sh26525521, 32'sh264fd0f2, 32'sh264d4cac, 32'sh264ac84e, 
               32'sh264843d9, 32'sh2645bf4b, 32'sh26433aa7, 32'sh2640b5eb, 32'sh263e3117, 32'sh263bac2b, 32'sh26392728, 32'sh2636a20d, 
               32'sh26341cdb, 32'sh26319792, 32'sh262f1230, 32'sh262c8cb7, 32'sh262a0727, 32'sh2627817f, 32'sh2624fbbf, 32'sh262275e8, 
               32'sh261feffa, 32'sh261d69f4, 32'sh261ae3d6, 32'sh26185da1, 32'sh2615d754, 32'sh261350f0, 32'sh2610ca75, 32'sh260e43e2, 
               32'sh260bbd37, 32'sh26093675, 32'sh2606af9c, 32'sh260428ab, 32'sh2601a1a2, 32'sh25ff1a83, 32'sh25fc934b, 32'sh25fa0bfd, 
               32'sh25f78497, 32'sh25f4fd19, 32'sh25f27584, 32'sh25efedd8, 32'sh25ed6614, 32'sh25eade39, 32'sh25e85646, 32'sh25e5ce3c, 
               32'sh25e3461b, 32'sh25e0bde2, 32'sh25de3592, 32'sh25dbad2b, 32'sh25d924ac, 32'sh25d69c16, 32'sh25d41369, 32'sh25d18aa4, 
               32'sh25cf01c8, 32'sh25cc78d4, 32'sh25c9efca, 32'sh25c766a8, 32'sh25c4dd6e, 32'sh25c2541e, 32'sh25bfcab6, 32'sh25bd4136, 
               32'sh25bab7a0, 32'sh25b82df2, 32'sh25b5a42d, 32'sh25b31a51, 32'sh25b0905d, 32'sh25ae0652, 32'sh25ab7c30, 32'sh25a8f1f7, 
               32'sh25a667a7, 32'sh25a3dd3f, 32'sh25a152c0, 32'sh259ec82a, 32'sh259c3d7c, 32'sh2599b2b8, 32'sh259727dc, 32'sh25949ce9, 
               32'sh259211df, 32'sh258f86be, 32'sh258cfb85, 32'sh258a7035, 32'sh2587e4cf, 32'sh25855951, 32'sh2582cdbc, 32'sh2580420f, 
               32'sh257db64c, 32'sh257b2a71, 32'sh25789e80, 32'sh25761277, 32'sh25738657, 32'sh2570fa20, 32'sh256e6dd2, 32'sh256be16d, 
               32'sh256954f1, 32'sh2566c85e, 32'sh25643bb3, 32'sh2561aef2, 32'sh255f2219, 32'sh255c952a, 32'sh255a0823, 32'sh25577b06, 
               32'sh2554edd1, 32'sh25526085, 32'sh254fd323, 32'sh254d45a9, 32'sh254ab818, 32'sh25482a70, 32'sh25459cb2, 32'sh25430edc, 
               32'sh254080ef, 32'sh253df2eb, 32'sh253b64d1, 32'sh2538d69f, 32'sh25364857, 32'sh2533b9f7, 32'sh25312b81, 32'sh252e9cf3, 
               32'sh252c0e4f, 32'sh25297f93, 32'sh2526f0c1, 32'sh252461d8, 32'sh2521d2d8, 32'sh251f43c1, 32'sh251cb493, 32'sh251a254e, 
               32'sh251795f3, 32'sh25150680, 32'sh251276f7, 32'sh250fe757, 32'sh250d57a0, 32'sh250ac7d2, 32'sh250837ed, 32'sh2505a7f1, 
               32'sh250317df, 32'sh250087b5, 32'sh24fdf775, 32'sh24fb671e, 32'sh24f8d6b0, 32'sh24f6462c, 32'sh24f3b590, 32'sh24f124de, 
               32'sh24ee9415, 32'sh24ec0335, 32'sh24e9723f, 32'sh24e6e132, 32'sh24e4500e, 32'sh24e1bed3, 32'sh24df2d81, 32'sh24dc9c19, 
               32'sh24da0a9a, 32'sh24d77904, 32'sh24d4e757, 32'sh24d25594, 32'sh24cfc3ba, 32'sh24cd31ca, 32'sh24ca9fc2, 32'sh24c80da4, 
               32'sh24c57b6f, 32'sh24c2e924, 32'sh24c056c2, 32'sh24bdc449, 32'sh24bb31ba, 32'sh24b89f14, 32'sh24b60c57, 32'sh24b37983, 
               32'sh24b0e699, 32'sh24ae5399, 32'sh24abc082, 32'sh24a92d54, 32'sh24a69a0f, 32'sh24a406b4, 32'sh24a17342, 32'sh249edfba, 
               32'sh249c4c1b, 32'sh2499b865, 32'sh24972499, 32'sh249490b7, 32'sh2491fcbe, 32'sh248f68ae, 32'sh248cd487, 32'sh248a404b, 
               32'sh2487abf7, 32'sh2485178d, 32'sh2482830d, 32'sh247fee76, 32'sh247d59c8, 32'sh247ac504, 32'sh2478302a, 32'sh24759b39, 
               32'sh24730631, 32'sh24707113, 32'sh246ddbdf, 32'sh246b4694, 32'sh2468b132, 32'sh24661bbb, 32'sh2463862c, 32'sh2460f088, 
               32'sh245e5acc, 32'sh245bc4fb, 32'sh24592f13, 32'sh24569914, 32'sh245402ff, 32'sh24516cd4, 32'sh244ed692, 32'sh244c403a, 
               32'sh2449a9cc, 32'sh24471347, 32'sh24447cac, 32'sh2441e5fa, 32'sh243f4f32, 32'sh243cb854, 32'sh243a215f, 32'sh24378a54, 
               32'sh2434f332, 32'sh24325bfb, 32'sh242fc4ad, 32'sh242d2d48, 32'sh242a95ce, 32'sh2427fe3d, 32'sh24256695, 32'sh2422ced8, 
               32'sh24203704, 32'sh241d9f1a, 32'sh241b0719, 32'sh24186f02, 32'sh2415d6d5, 32'sh24133e92, 32'sh2410a639, 32'sh240e0dc9, 
               32'sh240b7543, 32'sh2408dca7, 32'sh240643f4, 32'sh2403ab2c, 32'sh2401124d, 32'sh23fe7958, 32'sh23fbe04c, 32'sh23f9472b, 
               32'sh23f6adf3, 32'sh23f414a5, 32'sh23f17b41, 32'sh23eee1c7, 32'sh23ec4837, 32'sh23e9ae90, 32'sh23e714d3, 32'sh23e47b00, 
               32'sh23e1e117, 32'sh23df4718, 32'sh23dcad03, 32'sh23da12d8, 32'sh23d77896, 32'sh23d4de3f, 32'sh23d243d1, 32'sh23cfa94d, 
               32'sh23cd0eb3, 32'sh23ca7403, 32'sh23c7d93d, 32'sh23c53e61, 32'sh23c2a36f, 32'sh23c00867, 32'sh23bd6d48, 32'sh23bad214, 
               32'sh23b836ca, 32'sh23b59b69, 32'sh23b2fff3, 32'sh23b06466, 32'sh23adc8c4, 32'sh23ab2d0b, 32'sh23a8913d, 32'sh23a5f558, 
               32'sh23a3595e, 32'sh23a0bd4e, 32'sh239e2127, 32'sh239b84eb, 32'sh2398e898, 32'sh23964c30, 32'sh2393afb2, 32'sh2391131e, 
               32'sh238e7673, 32'sh238bd9b3, 32'sh23893cdd, 32'sh23869ff1, 32'sh238402ef, 32'sh238165d8, 32'sh237ec8aa, 32'sh237c2b66, 
               32'sh23798e0d, 32'sh2376f09e, 32'sh23745318, 32'sh2371b57d, 32'sh236f17cc, 32'sh236c7a06, 32'sh2369dc29, 32'sh23673e36, 
               32'sh2364a02e, 32'sh23620210, 32'sh235f63dc, 32'sh235cc592, 32'sh235a2733, 32'sh235788bd, 32'sh2354ea32, 32'sh23524b91, 
               32'sh234facda, 32'sh234d0e0d, 32'sh234a6f2b, 32'sh2347d033, 32'sh23453125, 32'sh23429201, 32'sh233ff2c8, 32'sh233d5379, 
               32'sh233ab414, 32'sh23381499, 32'sh23357509, 32'sh2332d563, 32'sh233035a7, 32'sh232d95d6, 32'sh232af5ee, 32'sh232855f2, 
               32'sh2325b5df, 32'sh232315b7, 32'sh23207579, 32'sh231dd525, 32'sh231b34bc, 32'sh2318943d, 32'sh2315f3a8, 32'sh231352fe, 
               32'sh2310b23e, 32'sh230e1169, 32'sh230b707e, 32'sh2308cf7d, 32'sh23062e67, 32'sh23038d3b, 32'sh2300ebf9, 32'sh22fe4aa2, 
               32'sh22fba936, 32'sh22f907b3, 32'sh22f6661c, 32'sh22f3c46e, 32'sh22f122ab, 32'sh22ee80d3, 32'sh22ebdee5, 32'sh22e93ce1, 
               32'sh22e69ac8, 32'sh22e3f899, 32'sh22e15655, 32'sh22deb3fb, 32'sh22dc118c, 32'sh22d96f07, 32'sh22d6cc6d, 32'sh22d429bd, 
               32'sh22d186f8, 32'sh22cee41d, 32'sh22cc412d, 32'sh22c99e28, 32'sh22c6fb0c, 32'sh22c457dc, 32'sh22c1b496, 32'sh22bf113b, 
               32'sh22bc6dca, 32'sh22b9ca43, 32'sh22b726a8, 32'sh22b482f7, 32'sh22b1df30, 32'sh22af3b54, 32'sh22ac9763, 32'sh22a9f35c, 
               32'sh22a74f40, 32'sh22a4ab0f, 32'sh22a206c8, 32'sh229f626c, 32'sh229cbdfa, 32'sh229a1973, 32'sh229774d7, 32'sh2294d025, 
               32'sh22922b5e, 32'sh228f8682, 32'sh228ce191, 32'sh228a3c8a, 32'sh2287976e, 32'sh2284f23c, 32'sh22824cf5, 32'sh227fa799, 
               32'sh227d0228, 32'sh227a5ca1, 32'sh2277b705, 32'sh22751154, 32'sh22726b8e, 32'sh226fc5b2, 32'sh226d1fc1, 32'sh226a79bb, 
               32'sh2267d3a0, 32'sh22652d6f, 32'sh22628729, 32'sh225fe0ce, 32'sh225d3a5e, 32'sh225a93d9, 32'sh2257ed3e, 32'sh2255468e, 
               32'sh22529fca, 32'sh224ff8ef, 32'sh224d5200, 32'sh224aaafc, 32'sh224803e2, 32'sh22455cb3, 32'sh2242b56f, 32'sh22400e16, 
               32'sh223d66a8, 32'sh223abf25, 32'sh2238178d, 32'sh22356fdf, 32'sh2232c81c, 32'sh22302045, 32'sh222d7858, 32'sh222ad056, 
               32'sh2228283f, 32'sh22258013, 32'sh2222d7d2, 32'sh22202f7c, 32'sh221d8711, 32'sh221ade91, 32'sh221835fb, 32'sh22158d51, 
               32'sh2212e492, 32'sh22103bbd, 32'sh220d92d4, 32'sh220ae9d6, 32'sh220840c2, 32'sh2205979a, 32'sh2202ee5d, 32'sh2200450a, 
               32'sh21fd9ba3, 32'sh21faf227, 32'sh21f84895, 32'sh21f59eef, 32'sh21f2f534, 32'sh21f04b64, 32'sh21eda17f, 32'sh21eaf785, 
               32'sh21e84d76, 32'sh21e5a353, 32'sh21e2f91a, 32'sh21e04ecc, 32'sh21dda46a, 32'sh21daf9f2, 32'sh21d84f66, 32'sh21d5a4c5, 
               32'sh21d2fa0f, 32'sh21d04f44, 32'sh21cda465, 32'sh21caf970, 32'sh21c84e67, 32'sh21c5a348, 32'sh21c2f815, 32'sh21c04ccd, 
               32'sh21bda171, 32'sh21baf5ff, 32'sh21b84a79, 32'sh21b59ede, 32'sh21b2f32e, 32'sh21b04769, 32'sh21ad9b8f, 32'sh21aaefa1, 
               32'sh21a8439e, 32'sh21a59786, 32'sh21a2eb5a, 32'sh21a03f18, 32'sh219d92c2, 32'sh219ae657, 32'sh219839d8, 32'sh21958d44, 
               32'sh2192e09b, 32'sh219033dd, 32'sh218d870b, 32'sh218ada24, 32'sh21882d28, 32'sh21858017, 32'sh2182d2f2, 32'sh218025b8, 
               32'sh217d786a, 32'sh217acb07, 32'sh21781d8f, 32'sh21757003, 32'sh2172c262, 32'sh217014ac, 32'sh216d66e2, 32'sh216ab903, 
               32'sh21680b0f, 32'sh21655d07, 32'sh2162aeea, 32'sh216000b9, 32'sh215d5273, 32'sh215aa418, 32'sh2157f5a9, 32'sh21554726, 
               32'sh2152988d, 32'sh214fe9e1, 32'sh214d3b1f, 32'sh214a8c49, 32'sh2147dd5f, 32'sh21452e60, 32'sh21427f4d, 32'sh213fd025, 
               32'sh213d20e8, 32'sh213a7197, 32'sh2137c232, 32'sh213512b8, 32'sh21326329, 32'sh212fb386, 32'sh212d03cf, 32'sh212a5403, 
               32'sh2127a423, 32'sh2124f42e, 32'sh21224425, 32'sh211f9407, 32'sh211ce3d5, 32'sh211a338e, 32'sh21178334, 32'sh2114d2c4, 
               32'sh21122240, 32'sh210f71a8, 32'sh210cc0fc, 32'sh210a103b, 32'sh21075f65, 32'sh2104ae7c, 32'sh2101fd7e, 32'sh20ff4c6b, 
               32'sh20fc9b44, 32'sh20f9ea09, 32'sh20f738ba, 32'sh20f48756, 32'sh20f1d5de, 32'sh20ef2451, 32'sh20ec72b1, 32'sh20e9c0fc, 
               32'sh20e70f32, 32'sh20e45d55, 32'sh20e1ab63, 32'sh20def95c, 32'sh20dc4742, 32'sh20d99513, 32'sh20d6e2d0, 32'sh20d43079, 
               32'sh20d17e0d, 32'sh20cecb8d, 32'sh20cc18f9, 32'sh20c96651, 32'sh20c6b395, 32'sh20c400c4, 32'sh20c14ddf, 32'sh20be9ae6, 
               32'sh20bbe7d8, 32'sh20b934b7, 32'sh20b68181, 32'sh20b3ce37, 32'sh20b11ad9, 32'sh20ae6767, 32'sh20abb3e1, 32'sh20a90046, 
               32'sh20a64c97, 32'sh20a398d5, 32'sh20a0e4fe, 32'sh209e3112, 32'sh209b7d13, 32'sh2098c900, 32'sh209614d9, 32'sh2093609d, 
               32'sh2090ac4d, 32'sh208df7ea, 32'sh208b4372, 32'sh20888ee6, 32'sh2085da46, 32'sh20832592, 32'sh208070ca, 32'sh207dbbee, 
               32'sh207b06fe, 32'sh207851fa, 32'sh20759ce1, 32'sh2072e7b5, 32'sh20703275, 32'sh206d7d21, 32'sh206ac7b8, 32'sh2068123c, 
               32'sh20655cac, 32'sh2062a708, 32'sh205ff14f, 32'sh205d3b83, 32'sh205a85a3, 32'sh2057cfaf, 32'sh205519a7, 32'sh2052638b, 
               32'sh204fad5b, 32'sh204cf717, 32'sh204a40bf, 32'sh20478a54, 32'sh2044d3d4, 32'sh20421d41, 32'sh203f6699, 32'sh203cafde, 
               32'sh2039f90f, 32'sh2037422c, 32'sh20348b35, 32'sh2031d42a, 32'sh202f1d0b, 32'sh202c65d9, 32'sh2029ae92, 32'sh2026f738, 
               32'sh20243fca, 32'sh20218848, 32'sh201ed0b2, 32'sh201c1909, 32'sh2019614c, 32'sh2016a97a, 32'sh2013f196, 32'sh2011399d, 
               32'sh200e8190, 32'sh200bc970, 32'sh2009113c, 32'sh200658f4, 32'sh2003a099, 32'sh2000e829, 32'sh1ffe2fa6, 32'sh1ffb7710, 
               32'sh1ff8be65, 32'sh1ff605a7, 32'sh1ff34cd5, 32'sh1ff093ef, 32'sh1feddaf6, 32'sh1feb21e9, 32'sh1fe868c8, 32'sh1fe5af94, 
               32'sh1fe2f64c, 32'sh1fe03cf0, 32'sh1fdd8381, 32'sh1fdac9fe, 32'sh1fd81067, 32'sh1fd556bd, 32'sh1fd29cff, 32'sh1fcfe32d, 
               32'sh1fcd2948, 32'sh1fca6f4f, 32'sh1fc7b542, 32'sh1fc4fb22, 32'sh1fc240ef, 32'sh1fbf86a7, 32'sh1fbccc4d, 32'sh1fba11de, 
               32'sh1fb7575c, 32'sh1fb49cc7, 32'sh1fb1e21d, 32'sh1faf2761, 32'sh1fac6c91, 32'sh1fa9b1ad, 32'sh1fa6f6b6, 32'sh1fa43bab, 
               32'sh1fa1808c, 32'sh1f9ec55b, 32'sh1f9c0a15, 32'sh1f994ebc, 32'sh1f969350, 32'sh1f93d7d0, 32'sh1f911c3d, 32'sh1f8e6096, 
               32'sh1f8ba4dc, 32'sh1f88e90e, 32'sh1f862d2d, 32'sh1f837139, 32'sh1f80b531, 32'sh1f7df915, 32'sh1f7b3ce6, 32'sh1f7880a4, 
               32'sh1f75c44e, 32'sh1f7307e5, 32'sh1f704b69, 32'sh1f6d8ed9, 32'sh1f6ad235, 32'sh1f68157f, 32'sh1f6558b5, 32'sh1f629bd7, 
               32'sh1f5fdee6, 32'sh1f5d21e2, 32'sh1f5a64cb, 32'sh1f57a7a0, 32'sh1f54ea62, 32'sh1f522d10, 32'sh1f4f6fab, 32'sh1f4cb233, 
               32'sh1f49f4a8, 32'sh1f473709, 32'sh1f447957, 32'sh1f41bb92, 32'sh1f3efdb9, 32'sh1f3c3fcd, 32'sh1f3981ce, 32'sh1f36c3bc, 
               32'sh1f340596, 32'sh1f31475d, 32'sh1f2e8911, 32'sh1f2bcab2, 32'sh1f290c3f, 32'sh1f264db9, 32'sh1f238f20, 32'sh1f20d074, 
               32'sh1f1e11b5, 32'sh1f1b52e2, 32'sh1f1893fc, 32'sh1f15d503, 32'sh1f1315f7, 32'sh1f1056d8, 32'sh1f0d97a5, 32'sh1f0ad860, 
               32'sh1f081907, 32'sh1f05599b, 32'sh1f029a1c, 32'sh1effda89, 32'sh1efd1ae4, 32'sh1efa5b2c, 32'sh1ef79b60, 32'sh1ef4db81, 
               32'sh1ef21b90, 32'sh1eef5b8b, 32'sh1eec9b73, 32'sh1ee9db48, 32'sh1ee71b0a, 32'sh1ee45ab9, 32'sh1ee19a54, 32'sh1eded9dd, 
               32'sh1edc1953, 32'sh1ed958b6, 32'sh1ed69805, 32'sh1ed3d742, 32'sh1ed1166b, 32'sh1ece5582, 32'sh1ecb9486, 32'sh1ec8d376, 
               32'sh1ec61254, 32'sh1ec3511f, 32'sh1ec08fd6, 32'sh1ebdce7b, 32'sh1ebb0d0d, 32'sh1eb84b8b, 32'sh1eb589f7, 32'sh1eb2c850, 
               32'sh1eb00696, 32'sh1ead44c9, 32'sh1eaa82e9, 32'sh1ea7c0f6, 32'sh1ea4fef0, 32'sh1ea23cd8, 32'sh1e9f7aac, 32'sh1e9cb86e, 
               32'sh1e99f61d, 32'sh1e9733b8, 32'sh1e947141, 32'sh1e91aeb7, 32'sh1e8eec1b, 32'sh1e8c296b, 32'sh1e8966a8, 32'sh1e86a3d3, 
               32'sh1e83e0eb, 32'sh1e811df0, 32'sh1e7e5ae2, 32'sh1e7b97c2, 32'sh1e78d48e, 32'sh1e761148, 32'sh1e734def, 32'sh1e708a83, 
               32'sh1e6dc705, 32'sh1e6b0373, 32'sh1e683fcf, 32'sh1e657c19, 32'sh1e62b84f, 32'sh1e5ff473, 32'sh1e5d3084, 32'sh1e5a6c82, 
               32'sh1e57a86d, 32'sh1e54e446, 32'sh1e52200c, 32'sh1e4f5bbf, 32'sh1e4c9760, 32'sh1e49d2ee, 32'sh1e470e69, 32'sh1e4449d2, 
               32'sh1e418528, 32'sh1e3ec06b, 32'sh1e3bfb9c, 32'sh1e3936ba, 32'sh1e3671c5, 32'sh1e33acbe, 32'sh1e30e7a4, 32'sh1e2e2277, 
               32'sh1e2b5d38, 32'sh1e2897e6, 32'sh1e25d282, 32'sh1e230d0b, 32'sh1e204781, 32'sh1e1d81e5, 32'sh1e1abc36, 32'sh1e17f675, 
               32'sh1e1530a1, 32'sh1e126abb, 32'sh1e0fa4c2, 32'sh1e0cdeb6, 32'sh1e0a1898, 32'sh1e075268, 32'sh1e048c24, 32'sh1e01c5cf, 
               32'sh1dfeff67, 32'sh1dfc38ec, 32'sh1df9725f, 32'sh1df6abbf, 32'sh1df3e50d, 32'sh1df11e49, 32'sh1dee5771, 32'sh1deb9088, 
               32'sh1de8c98c, 32'sh1de6027e, 32'sh1de33b5d, 32'sh1de07429, 32'sh1dddace4, 32'sh1ddae58b, 32'sh1dd81e21, 32'sh1dd556a4, 
               32'sh1dd28f15, 32'sh1dcfc773, 32'sh1dccffbf, 32'sh1dca37f8, 32'sh1dc7701f, 32'sh1dc4a834, 32'sh1dc1e036, 32'sh1dbf1826, 
               32'sh1dbc5004, 32'sh1db987cf, 32'sh1db6bf88, 32'sh1db3f72f, 32'sh1db12ec3, 32'sh1dae6645, 32'sh1dab9db5, 32'sh1da8d512, 
               32'sh1da60c5d, 32'sh1da34396, 32'sh1da07abc, 32'sh1d9db1d1, 32'sh1d9ae8d2, 32'sh1d981fc2, 32'sh1d9556a0, 32'sh1d928d6b, 
               32'sh1d8fc424, 32'sh1d8cfaca, 32'sh1d8a315f, 32'sh1d8767e1, 32'sh1d849e51, 32'sh1d81d4af, 32'sh1d7f0afb, 32'sh1d7c4134, 
               32'sh1d79775c, 32'sh1d76ad71, 32'sh1d73e374, 32'sh1d711964, 32'sh1d6e4f43, 32'sh1d6b850f, 32'sh1d68baca, 32'sh1d65f072, 
               32'sh1d632608, 32'sh1d605b8c, 32'sh1d5d90fd, 32'sh1d5ac65d, 32'sh1d57fbaa, 32'sh1d5530e6, 32'sh1d52660f, 32'sh1d4f9b26, 
               32'sh1d4cd02c, 32'sh1d4a051f, 32'sh1d473a00, 32'sh1d446ecf, 32'sh1d41a38c, 32'sh1d3ed837, 32'sh1d3c0ccf, 32'sh1d394156, 
               32'sh1d3675cb, 32'sh1d33aa2e, 32'sh1d30de7e, 32'sh1d2e12bd, 32'sh1d2b46ea, 32'sh1d287b05, 32'sh1d25af0d, 32'sh1d22e304, 
               32'sh1d2016e9, 32'sh1d1d4abc, 32'sh1d1a7e7d, 32'sh1d17b22c, 32'sh1d14e5c9, 32'sh1d121954, 32'sh1d0f4ccd, 32'sh1d0c8034, 
               32'sh1d09b389, 32'sh1d06e6cc, 32'sh1d0419fe, 32'sh1d014d1d, 32'sh1cfe802b, 32'sh1cfbb327, 32'sh1cf8e611, 32'sh1cf618e9, 
               32'sh1cf34baf, 32'sh1cf07e63, 32'sh1cedb106, 32'sh1ceae396, 32'sh1ce81615, 32'sh1ce54882, 32'sh1ce27add, 32'sh1cdfad26, 
               32'sh1cdcdf5e, 32'sh1cda1183, 32'sh1cd74397, 32'sh1cd47599, 32'sh1cd1a78a, 32'sh1cced968, 32'sh1ccc0b35, 32'sh1cc93cf0, 
               32'sh1cc66e99, 32'sh1cc3a031, 32'sh1cc0d1b6, 32'sh1cbe032a, 32'sh1cbb348d, 32'sh1cb865dd, 32'sh1cb5971c, 32'sh1cb2c849, 
               32'sh1caff965, 32'sh1cad2a6e, 32'sh1caa5b66, 32'sh1ca78c4d, 32'sh1ca4bd21, 32'sh1ca1ede4, 32'sh1c9f1e96, 32'sh1c9c4f35, 
               32'sh1c997fc4, 32'sh1c96b040, 32'sh1c93e0ab, 32'sh1c911104, 32'sh1c8e414b, 32'sh1c8b7181, 32'sh1c88a1a6, 32'sh1c85d1b8, 
               32'sh1c8301b9, 32'sh1c8031a9, 32'sh1c7d6187, 32'sh1c7a9153, 32'sh1c77c10e, 32'sh1c74f0b7, 32'sh1c72204f, 32'sh1c6f4fd5, 
               32'sh1c6c7f4a, 32'sh1c69aead, 32'sh1c66ddfe, 32'sh1c640d3e, 32'sh1c613c6d, 32'sh1c5e6b8a, 32'sh1c5b9a95, 32'sh1c58c98f, 
               32'sh1c55f878, 32'sh1c53274f, 32'sh1c505614, 32'sh1c4d84c8, 32'sh1c4ab36b, 32'sh1c47e1fc, 32'sh1c45107c, 32'sh1c423eea, 
               32'sh1c3f6d47, 32'sh1c3c9b93, 32'sh1c39c9cd, 32'sh1c36f7f5, 32'sh1c34260c, 32'sh1c315412, 32'sh1c2e8207, 32'sh1c2bafea, 
               32'sh1c28ddbb, 32'sh1c260b7c, 32'sh1c23392b, 32'sh1c2066c8, 32'sh1c1d9454, 32'sh1c1ac1cf, 32'sh1c17ef39, 32'sh1c151c91, 
               32'sh1c1249d8, 32'sh1c0f770e, 32'sh1c0ca432, 32'sh1c09d145, 32'sh1c06fe46, 32'sh1c042b37, 32'sh1c015816, 32'sh1bfe84e4, 
               32'sh1bfbb1a0, 32'sh1bf8de4c, 32'sh1bf60ae6, 32'sh1bf3376f, 32'sh1bf063e6, 32'sh1bed904c, 32'sh1beabca1, 32'sh1be7e8e5, 
               32'sh1be51518, 32'sh1be24139, 32'sh1bdf6d4a, 32'sh1bdc9949, 32'sh1bd9c537, 32'sh1bd6f113, 32'sh1bd41cdf, 32'sh1bd14899, 
               32'sh1bce7442, 32'sh1bcb9fda, 32'sh1bc8cb61, 32'sh1bc5f6d7, 32'sh1bc3223c, 32'sh1bc04d8f, 32'sh1bbd78d2, 32'sh1bbaa403, 
               32'sh1bb7cf23, 32'sh1bb4fa32, 32'sh1bb22530, 32'sh1baf501d, 32'sh1bac7af9, 32'sh1ba9a5c4, 32'sh1ba6d07d, 32'sh1ba3fb26, 
               32'sh1ba125bd, 32'sh1b9e5044, 32'sh1b9b7ab9, 32'sh1b98a51e, 32'sh1b95cf71, 32'sh1b92f9b4, 32'sh1b9023e5, 32'sh1b8d4e06, 
               32'sh1b8a7815, 32'sh1b87a213, 32'sh1b84cc01, 32'sh1b81f5dd, 32'sh1b7f1fa9, 32'sh1b7c4963, 32'sh1b79730d, 32'sh1b769ca6, 
               32'sh1b73c62d, 32'sh1b70efa4, 32'sh1b6e190a, 32'sh1b6b425f, 32'sh1b686ba3, 32'sh1b6594d6, 32'sh1b62bdf8, 32'sh1b5fe709, 
               32'sh1b5d100a, 32'sh1b5a38f9, 32'sh1b5761d8, 32'sh1b548aa6, 32'sh1b51b363, 32'sh1b4edc0f, 32'sh1b4c04aa, 32'sh1b492d35, 
               32'sh1b4655ae, 32'sh1b437e17, 32'sh1b40a66f, 32'sh1b3dceb6, 32'sh1b3af6ec, 32'sh1b381f12, 32'sh1b354727, 32'sh1b326f2b, 
               32'sh1b2f971e, 32'sh1b2cbf00, 32'sh1b29e6d2, 32'sh1b270e93, 32'sh1b243643, 32'sh1b215de2, 32'sh1b1e8571, 32'sh1b1bacef, 
               32'sh1b18d45c, 32'sh1b15fbb8, 32'sh1b132304, 32'sh1b104a3f, 32'sh1b0d716a, 32'sh1b0a9883, 32'sh1b07bf8c, 32'sh1b04e685, 
               32'sh1b020d6c, 32'sh1aff3444, 32'sh1afc5b0a, 32'sh1af981c0, 32'sh1af6a865, 32'sh1af3cef9, 32'sh1af0f57d, 32'sh1aee1bf0, 
               32'sh1aeb4253, 32'sh1ae868a5, 32'sh1ae58ee6, 32'sh1ae2b517, 32'sh1adfdb37, 32'sh1add0147, 32'sh1ada2746, 32'sh1ad74d34, 
               32'sh1ad47312, 32'sh1ad198e0, 32'sh1acebe9d, 32'sh1acbe449, 32'sh1ac909e5, 32'sh1ac62f70, 32'sh1ac354eb, 32'sh1ac07a55, 
               32'sh1abd9faf, 32'sh1abac4f8, 32'sh1ab7ea31, 32'sh1ab50f59, 32'sh1ab23471, 32'sh1aaf5978, 32'sh1aac7e6f, 32'sh1aa9a355, 
               32'sh1aa6c82b, 32'sh1aa3ecf1, 32'sh1aa111a6, 32'sh1a9e364b, 32'sh1a9b5adf, 32'sh1a987f63, 32'sh1a95a3d6, 32'sh1a92c839, 
               32'sh1a8fec8c, 32'sh1a8d10ce, 32'sh1a8a3500, 32'sh1a875922, 32'sh1a847d33, 32'sh1a81a134, 32'sh1a7ec524, 32'sh1a7be904, 
               32'sh1a790cd4, 32'sh1a763093, 32'sh1a735442, 32'sh1a7077e1, 32'sh1a6d9b70, 32'sh1a6abeee, 32'sh1a67e25c, 32'sh1a6505b9, 
               32'sh1a622907, 32'sh1a5f4c44, 32'sh1a5c6f70, 32'sh1a59928d, 32'sh1a56b599, 32'sh1a53d895, 32'sh1a50fb81, 32'sh1a4e1e5d, 
               32'sh1a4b4128, 32'sh1a4863e3, 32'sh1a45868e, 32'sh1a42a929, 32'sh1a3fcbb3, 32'sh1a3cee2d, 32'sh1a3a1097, 32'sh1a3732f1, 
               32'sh1a34553b, 32'sh1a317775, 32'sh1a2e999e, 32'sh1a2bbbb7, 32'sh1a28ddc0, 32'sh1a25ffb9, 32'sh1a2321a2, 32'sh1a20437b, 
               32'sh1a1d6544, 32'sh1a1a86fc, 32'sh1a17a8a5, 32'sh1a14ca3d, 32'sh1a11ebc5, 32'sh1a0f0d3d, 32'sh1a0c2ea5, 32'sh1a094ffd, 
               32'sh1a067145, 32'sh1a03927d, 32'sh1a00b3a5, 32'sh19fdd4bd, 32'sh19faf5c5, 32'sh19f816bc, 32'sh19f537a4, 32'sh19f2587c, 
               32'sh19ef7944, 32'sh19ec99fb, 32'sh19e9baa3, 32'sh19e6db3b, 32'sh19e3fbc3, 32'sh19e11c3a, 32'sh19de3ca2, 32'sh19db5cfa, 
               32'sh19d87d42, 32'sh19d59d7a, 32'sh19d2bda2, 32'sh19cfddba, 32'sh19ccfdc2, 32'sh19ca1dbb, 32'sh19c73da3, 32'sh19c45d7b, 
               32'sh19c17d44, 32'sh19be9cfd, 32'sh19bbbca6, 32'sh19b8dc3e, 32'sh19b5fbc8, 32'sh19b31b41, 32'sh19b03aaa, 32'sh19ad5a04, 
               32'sh19aa794d, 32'sh19a79887, 32'sh19a4b7b1, 32'sh19a1d6cb, 32'sh199ef5d6, 32'sh199c14d0, 32'sh199933bb, 32'sh19965296, 
               32'sh19937161, 32'sh1990901d, 32'sh198daec8, 32'sh198acd64, 32'sh1987ebf0, 32'sh19850a6d, 32'sh198228d9, 32'sh197f4736, 
               32'sh197c6584, 32'sh197983c1, 32'sh1976a1ef, 32'sh1973c00d, 32'sh1970de1b, 32'sh196dfc1a, 32'sh196b1a09, 32'sh196837e8, 
               32'sh196555b8, 32'sh19627378, 32'sh195f9128, 32'sh195caec9, 32'sh1959cc5a, 32'sh1956e9db, 32'sh1954074d, 32'sh195124af, 
               32'sh194e4201, 32'sh194b5f44, 32'sh19487c77, 32'sh1945999b, 32'sh1942b6af, 32'sh193fd3b4, 32'sh193cf0a9, 32'sh193a0d8e, 
               32'sh19372a64, 32'sh1934472a, 32'sh193163e1, 32'sh192e8088, 32'sh192b9d1f, 32'sh1928b9a8, 32'sh1925d620, 32'sh1922f289, 
               32'sh19200ee3, 32'sh191d2b2d, 32'sh191a4767, 32'sh19176393, 32'sh19147fae, 32'sh19119bba, 32'sh190eb7b7, 32'sh190bd3a4, 
               32'sh1908ef82, 32'sh19060b50, 32'sh1903270f, 32'sh190042bf, 32'sh18fd5e5f, 32'sh18fa79ef, 32'sh18f79571, 32'sh18f4b0e2, 
               32'sh18f1cc45, 32'sh18eee798, 32'sh18ec02db, 32'sh18e91e10, 32'sh18e63935, 32'sh18e3544a, 32'sh18e06f50, 32'sh18dd8a47, 
               32'sh18daa52f, 32'sh18d7c007, 32'sh18d4dad0, 32'sh18d1f589, 32'sh18cf1034, 32'sh18cc2acf, 32'sh18c9455a, 32'sh18c65fd7, 
               32'sh18c37a44, 32'sh18c094a1, 32'sh18bdaef0, 32'sh18bac92f, 32'sh18b7e35f, 32'sh18b4fd80, 32'sh18b21791, 32'sh18af3194, 
               32'sh18ac4b87, 32'sh18a9656b, 32'sh18a67f3f, 32'sh18a39905, 32'sh18a0b2bb, 32'sh189dcc62, 32'sh189ae5fa, 32'sh1897ff82, 
               32'sh189518fc, 32'sh18923266, 32'sh188f4bc2, 32'sh188c650e, 32'sh18897e4a, 32'sh18869778, 32'sh1883b097, 32'sh1880c9a6, 
               32'sh187de2a7, 32'sh187afb98, 32'sh1878147a, 32'sh18752d4d, 32'sh18724611, 32'sh186f5ec6, 32'sh186c776c, 32'sh18699003, 
               32'sh1866a88a, 32'sh1863c103, 32'sh1860d96d, 32'sh185df1c7, 32'sh185b0a13, 32'sh1858224f, 32'sh18553a7d, 32'sh1852529b, 
               32'sh184f6aab, 32'sh184c82ab, 32'sh18499a9d, 32'sh1846b280, 32'sh1843ca53, 32'sh1840e218, 32'sh183df9cd, 32'sh183b1174, 
               32'sh1838290c, 32'sh18354094, 32'sh1832580e, 32'sh182f6f79, 32'sh182c86d5, 32'sh18299e22, 32'sh1826b561, 32'sh1823cc90, 
               32'sh1820e3b0, 32'sh181dfac2, 32'sh181b11c4, 32'sh181828b8, 32'sh18153f9d, 32'sh18125673, 32'sh180f6d3a, 32'sh180c83f3, 
               32'sh18099a9c, 32'sh1806b137, 32'sh1803c7c3, 32'sh1800de40, 32'sh17fdf4ae, 32'sh17fb0b0e, 32'sh17f8215e, 32'sh17f537a0, 
               32'sh17f24dd3, 32'sh17ef63f8, 32'sh17ec7a0d, 32'sh17e99014, 32'sh17e6a60c, 32'sh17e3bbf6, 32'sh17e0d1d0, 32'sh17dde79c, 
               32'sh17dafd59, 32'sh17d81308, 32'sh17d528a7, 32'sh17d23e38, 32'sh17cf53bb, 32'sh17cc692e, 32'sh17c97e93, 32'sh17c693ea, 
               32'sh17c3a931, 32'sh17c0be6a, 32'sh17bdd394, 32'sh17bae8b0, 32'sh17b7fdbd, 32'sh17b512bb, 32'sh17b227ab, 32'sh17af3c8c, 
               32'sh17ac515f, 32'sh17a96623, 32'sh17a67ad8, 32'sh17a38f7f, 32'sh17a0a417, 32'sh179db8a1, 32'sh179acd1c, 32'sh1797e188, 
               32'sh1794f5e6, 32'sh17920a35, 32'sh178f1e76, 32'sh178c32a9, 32'sh178946cc, 32'sh17865ae2, 32'sh17836ee8, 32'sh178082e1, 
               32'sh177d96ca, 32'sh177aaaa6, 32'sh1777be72, 32'sh1774d231, 32'sh1771e5e0, 32'sh176ef982, 32'sh176c0d15, 32'sh17692099, 
               32'sh1766340f, 32'sh17634777, 32'sh17605ad0, 32'sh175d6e1b, 32'sh175a8157, 32'sh17579485, 32'sh1754a7a4, 32'sh1751bab5, 
               32'sh174ecdb8, 32'sh174be0ad, 32'sh1748f393, 32'sh1746066a, 32'sh17431933, 32'sh17402bee, 32'sh173d3e9b, 32'sh173a5139, 
               32'sh173763c9, 32'sh1734764b, 32'sh173188be, 32'sh172e9b23, 32'sh172bad7a, 32'sh1728bfc2, 32'sh1725d1fc, 32'sh1722e428, 
               32'sh171ff646, 32'sh171d0855, 32'sh171a1a56, 32'sh17172c49, 32'sh17143e2d, 32'sh17115003, 32'sh170e61cc, 32'sh170b7385, 
               32'sh17088531, 32'sh170596ce, 32'sh1702a85e, 32'sh16ffb9df, 32'sh16fccb51, 32'sh16f9dcb6, 32'sh16f6ee0d, 32'sh16f3ff55, 
               32'sh16f1108f, 32'sh16ee21bb, 32'sh16eb32d9, 32'sh16e843e9, 32'sh16e554ea, 32'sh16e265de, 32'sh16df76c3, 32'sh16dc879a, 
               32'sh16d99864, 32'sh16d6a91f, 32'sh16d3b9cc, 32'sh16d0ca6a, 32'sh16cddafb, 32'sh16caeb7e, 32'sh16c7fbf3, 32'sh16c50c59, 
               32'sh16c21cb2, 32'sh16bf2cfc, 32'sh16bc3d39, 32'sh16b94d67, 32'sh16b65d88, 32'sh16b36d9a, 32'sh16b07d9f, 32'sh16ad8d95, 
               32'sh16aa9d7e, 32'sh16a7ad58, 32'sh16a4bd25, 32'sh16a1cce3, 32'sh169edc94, 32'sh169bec37, 32'sh1698fbcb, 32'sh16960b52, 
               32'sh16931acb, 32'sh16902a36, 32'sh168d3993, 32'sh168a48e2, 32'sh16875823, 32'sh16846756, 32'sh1681767c, 32'sh167e8593, 
               32'sh167b949d, 32'sh1678a398, 32'sh1675b286, 32'sh1672c166, 32'sh166fd039, 32'sh166cdefd, 32'sh1669edb3, 32'sh1666fc5c, 
               32'sh16640af7, 32'sh16611984, 32'sh165e2803, 32'sh165b3675, 32'sh165844d8, 32'sh1655532e, 32'sh16526176, 32'sh164f6fb1, 
               32'sh164c7ddd, 32'sh16498bfc, 32'sh16469a0d, 32'sh1643a810, 32'sh1640b606, 32'sh163dc3ee, 32'sh163ad1c8, 32'sh1637df95, 
               32'sh1634ed53, 32'sh1631fb04, 32'sh162f08a8, 32'sh162c163d, 32'sh162923c5, 32'sh16263140, 32'sh16233eac, 32'sh16204c0b, 
               32'sh161d595d, 32'sh161a66a0, 32'sh161773d6, 32'sh161480ff, 32'sh16118e1a, 32'sh160e9b27, 32'sh160ba826, 32'sh1608b518, 
               32'sh1605c1fd, 32'sh1602ced4, 32'sh15ffdb9d, 32'sh15fce859, 32'sh15f9f507, 32'sh15f701a7, 32'sh15f40e3a, 32'sh15f11ac0, 
               32'sh15ee2738, 32'sh15eb33a2, 32'sh15e83fff, 32'sh15e54c4e, 32'sh15e25890, 32'sh15df64c5, 32'sh15dc70eb, 32'sh15d97d05, 
               32'sh15d68911, 32'sh15d3950f, 32'sh15d0a100, 32'sh15cdace4, 32'sh15cab8ba, 32'sh15c7c482, 32'sh15c4d03e, 32'sh15c1dbeb, 
               32'sh15bee78c, 32'sh15bbf31f, 32'sh15b8fea4, 32'sh15b60a1c, 32'sh15b31587, 32'sh15b020e4, 32'sh15ad2c34, 32'sh15aa3777, 
               32'sh15a742ac, 32'sh15a44dd4, 32'sh15a158ee, 32'sh159e63fc, 32'sh159b6efb, 32'sh159879ee, 32'sh159584d3, 32'sh15928fab, 
               32'sh158f9a76, 32'sh158ca533, 32'sh1589afe3, 32'sh1586ba86, 32'sh1583c51b, 32'sh1580cfa3, 32'sh157dda1e, 32'sh157ae48c, 
               32'sh1577eeec, 32'sh1574f93f, 32'sh15720385, 32'sh156f0dbe, 32'sh156c17e9, 32'sh15692207, 32'sh15662c18, 32'sh1563361c, 
               32'sh15604013, 32'sh155d49fc, 32'sh155a53d9, 32'sh15575da8, 32'sh1554676a, 32'sh1551711e, 32'sh154e7ac6, 32'sh154b8461, 
               32'sh15488dee, 32'sh1545976e, 32'sh1542a0e1, 32'sh153faa47, 32'sh153cb3a0, 32'sh1539bcec, 32'sh1536c62b, 32'sh1533cf5c, 
               32'sh1530d881, 32'sh152de198, 32'sh152aeaa3, 32'sh1527f3a0, 32'sh1524fc90, 32'sh15220573, 32'sh151f0e4a, 32'sh151c1713, 
               32'sh15191fcf, 32'sh1516287e, 32'sh15133120, 32'sh151039b5, 32'sh150d423d, 32'sh150a4ab9, 32'sh15075327, 32'sh15045b88, 
               32'sh150163dc, 32'sh14fe6c23, 32'sh14fb745e, 32'sh14f87c8b, 32'sh14f584ac, 32'sh14f28cbf, 32'sh14ef94c6, 32'sh14ec9cbf, 
               32'sh14e9a4ac, 32'sh14e6ac8c, 32'sh14e3b45f, 32'sh14e0bc25, 32'sh14ddc3de, 32'sh14dacb8b, 32'sh14d7d32a, 32'sh14d4dabd, 
               32'sh14d1e242, 32'sh14cee9bb, 32'sh14cbf127, 32'sh14c8f887, 32'sh14c5ffd9, 32'sh14c3071f, 32'sh14c00e58, 32'sh14bd1584, 
               32'sh14ba1ca3, 32'sh14b723b5, 32'sh14b42abb, 32'sh14b131b4, 32'sh14ae38a0, 32'sh14ab3f7f, 32'sh14a84652, 32'sh14a54d18, 
               32'sh14a253d1, 32'sh149f5a7e, 32'sh149c611d, 32'sh149967b0, 32'sh14966e36, 32'sh149374b0, 32'sh14907b1d, 32'sh148d817d, 
               32'sh148a87d1, 32'sh14878e18, 32'sh14849452, 32'sh14819a7f, 32'sh147ea0a0, 32'sh147ba6b4, 32'sh1478acbc, 32'sh1475b2b7, 
               32'sh1472b8a5, 32'sh146fbe87, 32'sh146cc45c, 32'sh1469ca25, 32'sh1466cfe1, 32'sh1463d590, 32'sh1460db33, 32'sh145de0c9, 
               32'sh145ae653, 32'sh1457ebd0, 32'sh1454f140, 32'sh1451f6a4, 32'sh144efbfc, 32'sh144c0147, 32'sh14490685, 32'sh14460bb7, 
               32'sh144310dd, 32'sh144015f5, 32'sh143d1b02, 32'sh143a2002, 32'sh143724f5, 32'sh143429dc, 32'sh14312eb7, 32'sh142e3385, 
               32'sh142b3846, 32'sh14283cfc, 32'sh142541a4, 32'sh14224641, 32'sh141f4ad1, 32'sh141c4f54, 32'sh141953cb, 32'sh14165836, 
               32'sh14135c94, 32'sh141060e6, 32'sh140d652c, 32'sh140a6965, 32'sh14076d91, 32'sh140471b2, 32'sh140175c6, 32'sh13fe79ce, 
               32'sh13fb7dc9, 32'sh13f881b8, 32'sh13f5859b, 32'sh13f28972, 32'sh13ef8d3c, 32'sh13ec90fa, 32'sh13e994ab, 32'sh13e69850, 
               32'sh13e39be9, 32'sh13e09f76, 32'sh13dda2f7, 32'sh13daa66b, 32'sh13d7a9d3, 32'sh13d4ad2f, 32'sh13d1b07e, 32'sh13ceb3c1, 
               32'sh13cbb6f8, 32'sh13c8ba23, 32'sh13c5bd42, 32'sh13c2c054, 32'sh13bfc35b, 32'sh13bcc655, 32'sh13b9c943, 32'sh13b6cc24, 
               32'sh13b3cefa, 32'sh13b0d1c3, 32'sh13add481, 32'sh13aad732, 32'sh13a7d9d7, 32'sh13a4dc70, 32'sh13a1defd, 32'sh139ee17d, 
               32'sh139be3f2, 32'sh1398e65a, 32'sh1395e8b7, 32'sh1392eb07, 32'sh138fed4b, 32'sh138cef83, 32'sh1389f1af, 32'sh1386f3cf, 
               32'sh1383f5e3, 32'sh1380f7eb, 32'sh137df9e7, 32'sh137afbd7, 32'sh1377fdbb, 32'sh1374ff93, 32'sh1372015f, 32'sh136f031f, 
               32'sh136c04d2, 32'sh1369067a, 32'sh13660816, 32'sh136309a6, 32'sh13600b2a, 32'sh135d0ca2, 32'sh135a0e0e, 32'sh13570f6f, 
               32'sh135410c3, 32'sh1351120b, 32'sh134e1348, 32'sh134b1478, 32'sh1348159d, 32'sh134516b5, 32'sh134217c2, 32'sh133f18c3, 
               32'sh133c19b8, 32'sh13391aa1, 32'sh13361b7f, 32'sh13331c50, 32'sh13301d16, 32'sh132d1dd0, 32'sh132a1e7e, 32'sh13271f20, 
               32'sh13241fb6, 32'sh13212041, 32'sh131e20c0, 32'sh131b2132, 32'sh1318219a, 32'sh131521f5, 32'sh13122245, 32'sh130f2288, 
               32'sh130c22c1, 32'sh130922ed, 32'sh1306230d, 32'sh13032322, 32'sh1300232c, 32'sh12fd2329, 32'sh12fa231b, 32'sh12f72301, 
               32'sh12f422db, 32'sh12f122aa, 32'sh12ee226c, 32'sh12eb2224, 32'sh12e821cf, 32'sh12e5216f, 32'sh12e22103, 32'sh12df208c, 
               32'sh12dc2009, 32'sh12d91f7a, 32'sh12d61ee0, 32'sh12d31e3a, 32'sh12d01d89, 32'sh12cd1ccc, 32'sh12ca1c03, 32'sh12c71b2e, 
               32'sh12c41a4f, 32'sh12c11963, 32'sh12be186c, 32'sh12bb1769, 32'sh12b8165b, 32'sh12b51542, 32'sh12b2141c, 32'sh12af12ec, 
               32'sh12ac11af, 32'sh12a91067, 32'sh12a60f14, 32'sh12a30db5, 32'sh12a00c4b, 32'sh129d0ad5, 32'sh129a0954, 32'sh129707c7, 
               32'sh1294062f, 32'sh1291048b, 32'sh128e02dc, 32'sh128b0121, 32'sh1287ff5b, 32'sh1284fd8a, 32'sh1281fbad, 32'sh127ef9c5, 
               32'sh127bf7d1, 32'sh1278f5d2, 32'sh1275f3c7, 32'sh1272f1b1, 32'sh126fef90, 32'sh126ced63, 32'sh1269eb2b, 32'sh1266e8e8, 
               32'sh1263e699, 32'sh1260e43f, 32'sh125de1da, 32'sh125adf69, 32'sh1257dced, 32'sh1254da66, 32'sh1251d7d3, 32'sh124ed535, 
               32'sh124bd28c, 32'sh1248cfd7, 32'sh1245cd17, 32'sh1242ca4c, 32'sh123fc776, 32'sh123cc494, 32'sh1239c1a7, 32'sh1236beaf, 
               32'sh1233bbac, 32'sh1230b89d, 32'sh122db583, 32'sh122ab25e, 32'sh1227af2e, 32'sh1224abf3, 32'sh1221a8ac, 32'sh121ea55a, 
               32'sh121ba1fd, 32'sh12189e95, 32'sh12159b22, 32'sh121297a3, 32'sh120f941a, 32'sh120c9085, 32'sh12098ce5, 32'sh1206893a, 
               32'sh12038584, 32'sh120081c3, 32'sh11fd7df6, 32'sh11fa7a1f, 32'sh11f7763c, 32'sh11f4724f, 32'sh11f16e56, 32'sh11ee6a52, 
               32'sh11eb6643, 32'sh11e86229, 32'sh11e55e04, 32'sh11e259d4, 32'sh11df5599, 32'sh11dc5153, 32'sh11d94d02, 32'sh11d648a6, 
               32'sh11d3443f, 32'sh11d03fcd, 32'sh11cd3b50, 32'sh11ca36c8, 32'sh11c73235, 32'sh11c42d97, 32'sh11c128ee, 32'sh11be243a, 
               32'sh11bb1f7c, 32'sh11b81ab2, 32'sh11b515dd, 32'sh11b210fe, 32'sh11af0c13, 32'sh11ac071e, 32'sh11a9021d, 32'sh11a5fd12, 
               32'sh11a2f7fc, 32'sh119ff2db, 32'sh119cedaf, 32'sh1199e878, 32'sh1196e337, 32'sh1193ddea, 32'sh1190d893, 32'sh118dd331, 
               32'sh118acdc4, 32'sh1187c84c, 32'sh1184c2ca, 32'sh1181bd3c, 32'sh117eb7a4, 32'sh117bb201, 32'sh1178ac53, 32'sh1175a69b, 
               32'sh1172a0d7, 32'sh116f9b09, 32'sh116c9531, 32'sh11698f4d, 32'sh1166895f, 32'sh11638366, 32'sh11607d62, 32'sh115d7753, 
               32'sh115a713a, 32'sh11576b16, 32'sh115464e8, 32'sh11515eae, 32'sh114e586a, 32'sh114b521c, 32'sh11484bc2, 32'sh1145455e, 
               32'sh11423ef0, 32'sh113f3876, 32'sh113c31f3, 32'sh11392b64, 32'sh113624cb, 32'sh11331e27, 32'sh11301779, 32'sh112d10c0, 
               32'sh112a09fc, 32'sh1127032e, 32'sh1123fc55, 32'sh1120f572, 32'sh111dee84, 32'sh111ae78b, 32'sh1117e088, 32'sh1114d97b, 
               32'sh1111d263, 32'sh110ecb40, 32'sh110bc413, 32'sh1108bcdb, 32'sh1105b599, 32'sh1102ae4c, 32'sh10ffa6f5, 32'sh10fc9f94, 
               32'sh10f99827, 32'sh10f690b1, 32'sh10f38930, 32'sh10f081a4, 32'sh10ed7a0e, 32'sh10ea726e, 32'sh10e76ac3, 32'sh10e4630e, 
               32'sh10e15b4e, 32'sh10de5384, 32'sh10db4baf, 32'sh10d843d1, 32'sh10d53be7, 32'sh10d233f4, 32'sh10cf2bf6, 32'sh10cc23ed, 
               32'sh10c91bda, 32'sh10c613bd, 32'sh10c30b96, 32'sh10c00364, 32'sh10bcfb28, 32'sh10b9f2e1, 32'sh10b6ea90, 32'sh10b3e235, 
               32'sh10b0d9d0, 32'sh10add160, 32'sh10aac8e6, 32'sh10a7c062, 32'sh10a4b7d3, 32'sh10a1af3a, 32'sh109ea697, 32'sh109b9dea, 
               32'sh10989532, 32'sh10958c71, 32'sh109283a5, 32'sh108f7ace, 32'sh108c71ee, 32'sh10896903, 32'sh1086600e, 32'sh1083570f, 
               32'sh10804e06, 32'sh107d44f2, 32'sh107a3bd5, 32'sh107732ad, 32'sh1074297b, 32'sh1071203f, 32'sh106e16f9, 32'sh106b0da8, 
               32'sh1068044e, 32'sh1064fae9, 32'sh1061f17b, 32'sh105ee802, 32'sh105bde7f, 32'sh1058d4f2, 32'sh1055cb5b, 32'sh1052c1b9, 
               32'sh104fb80e, 32'sh104cae59, 32'sh1049a49a, 32'sh10469ad0, 32'sh104390fd, 32'sh1040871f, 32'sh103d7d38, 32'sh103a7346, 
               32'sh1037694b, 32'sh10345f45, 32'sh10315535, 32'sh102e4b1c, 32'sh102b40f8, 32'sh102836cb, 32'sh10252c94, 32'sh10222252, 
               32'sh101f1807, 32'sh101c0db1, 32'sh10190352, 32'sh1015f8e9, 32'sh1012ee76, 32'sh100fe3f9, 32'sh100cd972, 32'sh1009cee1, 
               32'sh1006c446, 32'sh1003b9a2, 32'sh1000aef3, 32'sh0ffda43b, 32'sh0ffa9979, 32'sh0ff78ead, 32'sh0ff483d7, 32'sh0ff178f7, 
               32'sh0fee6e0d, 32'sh0feb631a, 32'sh0fe8581d, 32'sh0fe54d16, 32'sh0fe24205, 32'sh0fdf36ea, 32'sh0fdc2bc6, 32'sh0fd92098, 
               32'sh0fd6155f, 32'sh0fd30a1e, 32'sh0fcffed2, 32'sh0fccf37d, 32'sh0fc9e81e, 32'sh0fc6dcb5, 32'sh0fc3d143, 32'sh0fc0c5c6, 
               32'sh0fbdba40, 32'sh0fbaaeb1, 32'sh0fb7a317, 32'sh0fb49774, 32'sh0fb18bc8, 32'sh0fae8011, 32'sh0fab7451, 32'sh0fa86887, 
               32'sh0fa55cb4, 32'sh0fa250d7, 32'sh0f9f44f0, 32'sh0f9c3900, 32'sh0f992d06, 32'sh0f962102, 32'sh0f9314f5, 32'sh0f9008de, 
               32'sh0f8cfcbe, 32'sh0f89f094, 32'sh0f86e460, 32'sh0f83d823, 32'sh0f80cbdc, 32'sh0f7dbf8c, 32'sh0f7ab332, 32'sh0f77a6ce, 
               32'sh0f749a61, 32'sh0f718deb, 32'sh0f6e816b, 32'sh0f6b74e1, 32'sh0f68684e, 32'sh0f655bb2, 32'sh0f624f0c, 32'sh0f5f425c, 
               32'sh0f5c35a3, 32'sh0f5928e1, 32'sh0f561c15, 32'sh0f530f3f, 32'sh0f500260, 32'sh0f4cf578, 32'sh0f49e886, 32'sh0f46db8b, 
               32'sh0f43ce86, 32'sh0f40c178, 32'sh0f3db461, 32'sh0f3aa740, 32'sh0f379a16, 32'sh0f348ce2, 32'sh0f317fa5, 32'sh0f2e725f, 
               32'sh0f2b650f, 32'sh0f2857b6, 32'sh0f254a53, 32'sh0f223ce8, 32'sh0f1f2f73, 32'sh0f1c21f4, 32'sh0f19146c, 32'sh0f1606db, 
               32'sh0f12f941, 32'sh0f0feb9d, 32'sh0f0cddf0, 32'sh0f09d03a, 32'sh0f06c27a, 32'sh0f03b4b1, 32'sh0f00a6df, 32'sh0efd9904, 
               32'sh0efa8b20, 32'sh0ef77d32, 32'sh0ef46f3b, 32'sh0ef1613a, 32'sh0eee5331, 32'sh0eeb451e, 32'sh0ee83702, 32'sh0ee528dd, 
               32'sh0ee21aaf, 32'sh0edf0c77, 32'sh0edbfe37, 32'sh0ed8efed, 32'sh0ed5e19a, 32'sh0ed2d33e, 32'sh0ecfc4d9, 32'sh0eccb66a, 
               32'sh0ec9a7f3, 32'sh0ec69972, 32'sh0ec38ae8, 32'sh0ec07c55, 32'sh0ebd6db9, 32'sh0eba5f14, 32'sh0eb75066, 32'sh0eb441af, 
               32'sh0eb132ef, 32'sh0eae2425, 32'sh0eab1553, 32'sh0ea80677, 32'sh0ea4f793, 32'sh0ea1e8a5, 32'sh0e9ed9af, 32'sh0e9bcaaf, 
               32'sh0e98bba7, 32'sh0e95ac95, 32'sh0e929d7a, 32'sh0e8f8e57, 32'sh0e8c7f2a, 32'sh0e896ff5, 32'sh0e8660b6, 32'sh0e83516f, 
               32'sh0e80421e, 32'sh0e7d32c5, 32'sh0e7a2363, 32'sh0e7713f7, 32'sh0e740483, 32'sh0e70f506, 32'sh0e6de580, 32'sh0e6ad5f1, 
               32'sh0e67c65a, 32'sh0e64b6b9, 32'sh0e61a70f, 32'sh0e5e975d, 32'sh0e5b87a2, 32'sh0e5877de, 32'sh0e556811, 32'sh0e52583b, 
               32'sh0e4f485c, 32'sh0e4c3875, 32'sh0e492884, 32'sh0e46188b, 32'sh0e430889, 32'sh0e3ff87f, 32'sh0e3ce86b, 32'sh0e39d84f, 
               32'sh0e36c82a, 32'sh0e33b7fc, 32'sh0e30a7c5, 32'sh0e2d9786, 32'sh0e2a873e, 32'sh0e2776ed, 32'sh0e246693, 32'sh0e215631, 
               32'sh0e1e45c6, 32'sh0e1b3552, 32'sh0e1824d6, 32'sh0e151451, 32'sh0e1203c3, 32'sh0e0ef32d, 32'sh0e0be28e, 32'sh0e08d1e6, 
               32'sh0e05c135, 32'sh0e02b07c, 32'sh0dff9fba, 32'sh0dfc8ef0, 32'sh0df97e1d, 32'sh0df66d41, 32'sh0df35c5d, 32'sh0df04b70, 
               32'sh0ded3a7b, 32'sh0dea297d, 32'sh0de71876, 32'sh0de40767, 32'sh0de0f64f, 32'sh0ddde52f, 32'sh0ddad406, 32'sh0dd7c2d4, 
               32'sh0dd4b19a, 32'sh0dd1a058, 32'sh0dce8f0d, 32'sh0dcb7db9, 32'sh0dc86c5d, 32'sh0dc55af9, 32'sh0dc2498c, 32'sh0dbf3816, 
               32'sh0dbc2698, 32'sh0db91512, 32'sh0db60383, 32'sh0db2f1eb, 32'sh0dafe04b, 32'sh0daccea3, 32'sh0da9bcf2, 32'sh0da6ab39, 
               32'sh0da39978, 32'sh0da087ae, 32'sh0d9d75db, 32'sh0d9a6400, 32'sh0d97521d, 32'sh0d944032, 32'sh0d912e3e, 32'sh0d8e1c41, 
               32'sh0d8b0a3d, 32'sh0d87f830, 32'sh0d84e61a, 32'sh0d81d3fc, 32'sh0d7ec1d6, 32'sh0d7bafa8, 32'sh0d789d71, 32'sh0d758b32, 
               32'sh0d7278eb, 32'sh0d6f669b, 32'sh0d6c5443, 32'sh0d6941e3, 32'sh0d662f7b, 32'sh0d631d0a, 32'sh0d600a91, 32'sh0d5cf810, 
               32'sh0d59e586, 32'sh0d56d2f5, 32'sh0d53c05b, 32'sh0d50adb9, 32'sh0d4d9b0e, 32'sh0d4a885c, 32'sh0d4775a1, 32'sh0d4462de, 
               32'sh0d415013, 32'sh0d3e3d40, 32'sh0d3b2a64, 32'sh0d381780, 32'sh0d350495, 32'sh0d31f1a1, 32'sh0d2edea5, 32'sh0d2bcba0, 
               32'sh0d28b894, 32'sh0d25a57f, 32'sh0d229263, 32'sh0d1f7f3e, 32'sh0d1c6c11, 32'sh0d1958dd, 32'sh0d1645a0, 32'sh0d13325b, 
               32'sh0d101f0e, 32'sh0d0d0bb8, 32'sh0d09f85b, 32'sh0d06e4f6, 32'sh0d03d189, 32'sh0d00be13, 32'sh0cfdaa96, 32'sh0cfa9711, 
               32'sh0cf78383, 32'sh0cf46fee, 32'sh0cf15c51, 32'sh0cee48ab, 32'sh0ceb34fe, 32'sh0ce82149, 32'sh0ce50d8c, 32'sh0ce1f9c7, 
               32'sh0cdee5f9, 32'sh0cdbd224, 32'sh0cd8be47, 32'sh0cd5aa62, 32'sh0cd29676, 32'sh0ccf8281, 32'sh0ccc6e84, 32'sh0cc95a80, 
               32'sh0cc64673, 32'sh0cc3325f, 32'sh0cc01e43, 32'sh0cbd0a1f, 32'sh0cb9f5f3, 32'sh0cb6e1bf, 32'sh0cb3cd84, 32'sh0cb0b940, 
               32'sh0cada4f5, 32'sh0caa90a2, 32'sh0ca77c47, 32'sh0ca467e4, 32'sh0ca1537a, 32'sh0c9e3f07, 32'sh0c9b2a8d, 32'sh0c98160c, 
               32'sh0c950182, 32'sh0c91ecf1, 32'sh0c8ed857, 32'sh0c8bc3b7, 32'sh0c88af0e, 32'sh0c859a5e, 32'sh0c8285a5, 32'sh0c7f70e6, 
               32'sh0c7c5c1e, 32'sh0c79474f, 32'sh0c763278, 32'sh0c731d9a, 32'sh0c7008b3, 32'sh0c6cf3c5, 32'sh0c69ded0, 32'sh0c66c9d3, 
               32'sh0c63b4ce, 32'sh0c609fc1, 32'sh0c5d8aad, 32'sh0c5a7591, 32'sh0c57606e, 32'sh0c544b43, 32'sh0c513610, 32'sh0c4e20d6, 
               32'sh0c4b0b94, 32'sh0c47f64a, 32'sh0c44e0f9, 32'sh0c41cba1, 32'sh0c3eb641, 32'sh0c3ba0d9, 32'sh0c388b6a, 32'sh0c3575f3, 
               32'sh0c326075, 32'sh0c2f4aef, 32'sh0c2c3562, 32'sh0c291fcd, 32'sh0c260a31, 32'sh0c22f48d, 32'sh0c1fdee1, 32'sh0c1cc92f, 
               32'sh0c19b374, 32'sh0c169db3, 32'sh0c1387e9, 32'sh0c107219, 32'sh0c0d5c41, 32'sh0c0a4661, 32'sh0c07307a, 32'sh0c041a8c, 
               32'sh0c010496, 32'sh0bfdee99, 32'sh0bfad894, 32'sh0bf7c288, 32'sh0bf4ac75, 32'sh0bf1965a, 32'sh0bee8038, 32'sh0beb6a0f, 
               32'sh0be853de, 32'sh0be53da6, 32'sh0be22766, 32'sh0bdf111f, 32'sh0bdbfad1, 32'sh0bd8e47c, 32'sh0bd5ce1f, 32'sh0bd2b7bb, 
               32'sh0bcfa150, 32'sh0bcc8add, 32'sh0bc97463, 32'sh0bc65de2, 32'sh0bc34759, 32'sh0bc030ca, 32'sh0bbd1a33, 32'sh0bba0395, 
               32'sh0bb6ecef, 32'sh0bb3d642, 32'sh0bb0bf8f, 32'sh0bada8d4, 32'sh0baa9211, 32'sh0ba77b48, 32'sh0ba46477, 32'sh0ba14d9f, 
               32'sh0b9e36c0, 32'sh0b9b1fda, 32'sh0b9808ed, 32'sh0b94f1f8, 32'sh0b91dafc, 32'sh0b8ec3fa, 32'sh0b8bacf0, 32'sh0b8895df, 
               32'sh0b857ec7, 32'sh0b8267a7, 32'sh0b7f5081, 32'sh0b7c3953, 32'sh0b79221f, 32'sh0b760ae3, 32'sh0b72f3a1, 32'sh0b6fdc57, 
               32'sh0b6cc506, 32'sh0b69adae, 32'sh0b66964f, 32'sh0b637ee9, 32'sh0b60677c, 32'sh0b5d5008, 32'sh0b5a388d, 32'sh0b57210b, 
               32'sh0b540982, 32'sh0b50f1f3, 32'sh0b4dda5c, 32'sh0b4ac2be, 32'sh0b47ab19, 32'sh0b44936d, 32'sh0b417bba, 32'sh0b3e6400, 
               32'sh0b3b4c40, 32'sh0b383478, 32'sh0b351caa, 32'sh0b3204d4, 32'sh0b2eecf8, 32'sh0b2bd515, 32'sh0b28bd2a, 32'sh0b25a539, 
               32'sh0b228d42, 32'sh0b1f7543, 32'sh0b1c5d3d, 32'sh0b194531, 32'sh0b162d1d, 32'sh0b131503, 32'sh0b0ffce2, 32'sh0b0ce4ba, 
               32'sh0b09cc8c, 32'sh0b06b456, 32'sh0b039c1a, 32'sh0b0083d7, 32'sh0afd6b8d, 32'sh0afa533d, 32'sh0af73ae5, 32'sh0af42287, 
               32'sh0af10a22, 32'sh0aedf1b7, 32'sh0aead944, 32'sh0ae7c0cb, 32'sh0ae4a84b, 32'sh0ae18fc5, 32'sh0ade7737, 32'sh0adb5ea3, 
               32'sh0ad84609, 32'sh0ad52d67, 32'sh0ad214bf, 32'sh0acefc11, 32'sh0acbe35b, 32'sh0ac8ca9f, 32'sh0ac5b1dc, 32'sh0ac29913, 
               32'sh0abf8043, 32'sh0abc676d, 32'sh0ab94e8f, 32'sh0ab635ab, 32'sh0ab31cc1, 32'sh0ab003d0, 32'sh0aacead8, 32'sh0aa9d1da, 
               32'sh0aa6b8d5, 32'sh0aa39fca, 32'sh0aa086b8, 32'sh0a9d6d9f, 32'sh0a9a5480, 32'sh0a973b5b, 32'sh0a94222f, 32'sh0a9108fc, 
               32'sh0a8defc3, 32'sh0a8ad683, 32'sh0a87bd3d, 32'sh0a84a3f0, 32'sh0a818a9d, 32'sh0a7e7143, 32'sh0a7b57e3, 32'sh0a783e7d, 
               32'sh0a752510, 32'sh0a720b9c, 32'sh0a6ef222, 32'sh0a6bd8a2, 32'sh0a68bf1b, 32'sh0a65a58e, 32'sh0a628bfa, 32'sh0a5f7260, 
               32'sh0a5c58c0, 32'sh0a593f19, 32'sh0a56256c, 32'sh0a530bb8, 32'sh0a4ff1fe, 32'sh0a4cd83e, 32'sh0a49be77, 32'sh0a46a4aa, 
               32'sh0a438ad7, 32'sh0a4070fd, 32'sh0a3d571d, 32'sh0a3a3d37, 32'sh0a37234a, 32'sh0a340957, 32'sh0a30ef5e, 32'sh0a2dd55e, 
               32'sh0a2abb59, 32'sh0a27a14d, 32'sh0a24873a, 32'sh0a216d22, 32'sh0a1e5303, 32'sh0a1b38de, 32'sh0a181eb2, 32'sh0a150481, 
               32'sh0a11ea49, 32'sh0a0ed00b, 32'sh0a0bb5c7, 32'sh0a089b7c, 32'sh0a05812c, 32'sh0a0266d5, 32'sh09ff4c78, 32'sh09fc3215, 
               32'sh09f917ac, 32'sh09f5fd3d, 32'sh09f2e2c7, 32'sh09efc84b, 32'sh09ecadc9, 32'sh09e99342, 32'sh09e678b4, 32'sh09e35e1f, 
               32'sh09e04385, 32'sh09dd28e5, 32'sh09da0e3e, 32'sh09d6f392, 32'sh09d3d8df, 32'sh09d0be27, 32'sh09cda368, 32'sh09ca88a3, 
               32'sh09c76dd8, 32'sh09c45308, 32'sh09c13831, 32'sh09be1d54, 32'sh09bb0271, 32'sh09b7e788, 32'sh09b4cc99, 32'sh09b1b1a4, 
               32'sh09ae96aa, 32'sh09ab7ba9, 32'sh09a860a2, 32'sh09a54595, 32'sh09a22a83, 32'sh099f0f6a, 32'sh099bf44c, 32'sh0998d927, 
               32'sh0995bdfd, 32'sh0992a2cc, 32'sh098f8796, 32'sh098c6c5a, 32'sh09895118, 32'sh098635d0, 32'sh09831a82, 32'sh097fff2f, 
               32'sh097ce3d5, 32'sh0979c876, 32'sh0976ad11, 32'sh097391a6, 32'sh09707635, 32'sh096d5abe, 32'sh096a3f42, 32'sh096723bf, 
               32'sh09640837, 32'sh0960eca9, 32'sh095dd116, 32'sh095ab57c, 32'sh095799dd, 32'sh09547e38, 32'sh0951628d, 32'sh094e46dd, 
               32'sh094b2b27, 32'sh09480f6b, 32'sh0944f3a9, 32'sh0941d7e2, 32'sh093ebc14, 32'sh093ba042, 32'sh09388469, 32'sh0935688b, 
               32'sh09324ca7, 32'sh092f30bd, 32'sh092c14ce, 32'sh0928f8d9, 32'sh0925dcdf, 32'sh0922c0df, 32'sh091fa4d9, 32'sh091c88cd, 
               32'sh09196cbc, 32'sh091650a6, 32'sh09133489, 32'sh09101868, 32'sh090cfc40, 32'sh0909e013, 32'sh0906c3e0, 32'sh0903a7a8, 
               32'sh09008b6a, 32'sh08fd6f27, 32'sh08fa52de, 32'sh08f73690, 32'sh08f41a3c, 32'sh08f0fde3, 32'sh08ede184, 32'sh08eac51f, 
               32'sh08e7a8b5, 32'sh08e48c46, 32'sh08e16fd1, 32'sh08de5356, 32'sh08db36d6, 32'sh08d81a51, 32'sh08d4fdc6, 32'sh08d1e136, 
               32'sh08cec4a0, 32'sh08cba805, 32'sh08c88b65, 32'sh08c56ebf, 32'sh08c25213, 32'sh08bf3563, 32'sh08bc18ac, 32'sh08b8fbf1, 
               32'sh08b5df30, 32'sh08b2c26a, 32'sh08afa59e, 32'sh08ac88cd, 32'sh08a96bf6, 32'sh08a64f1b, 32'sh08a3323a, 32'sh08a01553, 
               32'sh089cf867, 32'sh0899db76, 32'sh0896be80, 32'sh0893a184, 32'sh08908483, 32'sh088d677d, 32'sh088a4a72, 32'sh08872d61, 
               32'sh0884104b, 32'sh0880f330, 32'sh087dd60f, 32'sh087ab8e9, 32'sh08779bbe, 32'sh08747e8e, 32'sh08716159, 32'sh086e441e, 
               32'sh086b26de, 32'sh08680999, 32'sh0864ec4f, 32'sh0861cf00, 32'sh085eb1ab, 32'sh085b9451, 32'sh085876f3, 32'sh0855598f, 
               32'sh08523c25, 32'sh084f1eb7, 32'sh084c0144, 32'sh0848e3cb, 32'sh0845c64d, 32'sh0842a8cb, 32'sh083f8b43, 32'sh083c6db6, 
               32'sh08395024, 32'sh0836328d, 32'sh083314f1, 32'sh082ff74f, 32'sh082cd9a9, 32'sh0829bbfe, 32'sh08269e4d, 32'sh08238098, 
               32'sh082062de, 32'sh081d451e, 32'sh081a275a, 32'sh08170990, 32'sh0813ebc2, 32'sh0810cdef, 32'sh080db016, 32'sh080a9239, 
               32'sh08077457, 32'sh0804566f, 32'sh08013883, 32'sh07fe1a92, 32'sh07fafc9c, 32'sh07f7dea1, 32'sh07f4c0a1, 32'sh07f1a29c, 
               32'sh07ee8493, 32'sh07eb6684, 32'sh07e84871, 32'sh07e52a58, 32'sh07e20c3b, 32'sh07deee19, 32'sh07dbcff2, 32'sh07d8b1c6, 
               32'sh07d59396, 32'sh07d27560, 32'sh07cf5726, 32'sh07cc38e7, 32'sh07c91aa3, 32'sh07c5fc5a, 32'sh07c2de0d, 32'sh07bfbfba, 
               32'sh07bca163, 32'sh07b98307, 32'sh07b664a7, 32'sh07b34641, 32'sh07b027d7, 32'sh07ad0968, 32'sh07a9eaf5, 32'sh07a6cc7d, 
               32'sh07a3adff, 32'sh07a08f7e, 32'sh079d70f7, 32'sh079a526c, 32'sh079733dc, 32'sh07941548, 32'sh0790f6ae, 32'sh078dd811, 
               32'sh078ab96e, 32'sh07879ac7, 32'sh07847c1b, 32'sh07815d6b, 32'sh077e3eb5, 32'sh077b1ffc, 32'sh0778013d, 32'sh0774e27a, 
               32'sh0771c3b3, 32'sh076ea4e7, 32'sh076b8616, 32'sh07686741, 32'sh07654867, 32'sh07622988, 32'sh075f0aa5, 32'sh075bebbe, 
               32'sh0758ccd2, 32'sh0755ade1, 32'sh07528eec, 32'sh074f6ff3, 32'sh074c50f4, 32'sh074931f2, 32'sh074612eb, 32'sh0742f3df, 
               32'sh073fd4cf, 32'sh073cb5ba, 32'sh073996a1, 32'sh07367784, 32'sh07335862, 32'sh0730393b, 32'sh072d1a10, 32'sh0729fae1, 
               32'sh0726dbae, 32'sh0723bc75, 32'sh07209d39, 32'sh071d7df8, 32'sh071a5eb3, 32'sh07173f69, 32'sh0714201b, 32'sh071100c9, 
               32'sh070de172, 32'sh070ac217, 32'sh0707a2b7, 32'sh07048354, 32'sh070163eb, 32'sh06fe447f, 32'sh06fb250e, 32'sh06f80599, 
               32'sh06f4e620, 32'sh06f1c6a2, 32'sh06eea720, 32'sh06eb879a, 32'sh06e86810, 32'sh06e54881, 32'sh06e228ee, 32'sh06df0957, 
               32'sh06dbe9bb, 32'sh06d8ca1b, 32'sh06d5aa77, 32'sh06d28acf, 32'sh06cf6b23, 32'sh06cc4b72, 32'sh06c92bbe, 32'sh06c60c05, 
               32'sh06c2ec48, 32'sh06bfcc86, 32'sh06bcacc1, 32'sh06b98cf7, 32'sh06b66d29, 32'sh06b34d58, 32'sh06b02d81, 32'sh06ad0da7, 
               32'sh06a9edc9, 32'sh06a6cde7, 32'sh06a3ae00, 32'sh06a08e16, 32'sh069d6e27, 32'sh069a4e34, 32'sh06972e3d, 32'sh06940e42, 
               32'sh0690ee44, 32'sh068dce41, 32'sh068aae3a, 32'sh06878e2e, 32'sh06846e1f, 32'sh06814e0c, 32'sh067e2df5, 32'sh067b0dda, 
               32'sh0677edbb, 32'sh0674cd98, 32'sh0671ad71, 32'sh066e8d45, 32'sh066b6d16, 32'sh06684ce3, 32'sh06652cac, 32'sh06620c72, 
               32'sh065eec33, 32'sh065bcbf0, 32'sh0658aba9, 32'sh06558b5f, 32'sh06526b10, 32'sh064f4abe, 32'sh064c2a67, 32'sh06490a0d, 
               32'sh0645e9af, 32'sh0642c94d, 32'sh063fa8e7, 32'sh063c887e, 32'sh06396810, 32'sh0636479f, 32'sh0633272a, 32'sh063006b1, 
               32'sh062ce634, 32'sh0629c5b3, 32'sh0626a52f, 32'sh062384a6, 32'sh0620641a, 32'sh061d438b, 32'sh061a22f7, 32'sh06170260, 
               32'sh0613e1c5, 32'sh0610c126, 32'sh060da083, 32'sh060a7fdd, 32'sh06075f33, 32'sh06043e85, 32'sh06011dd4, 32'sh05fdfd1f, 
               32'sh05fadc66, 32'sh05f7bba9, 32'sh05f49ae9, 32'sh05f17a25, 32'sh05ee595d, 32'sh05eb3892, 32'sh05e817c3, 32'sh05e4f6f1, 
               32'sh05e1d61b, 32'sh05deb541, 32'sh05db9463, 32'sh05d87382, 32'sh05d5529e, 32'sh05d231b5, 32'sh05cf10ca, 32'sh05cbefda, 
               32'sh05c8cee7, 32'sh05c5adf1, 32'sh05c28cf7, 32'sh05bf6bf9, 32'sh05bc4af8, 32'sh05b929f3, 32'sh05b608eb, 32'sh05b2e7df, 
               32'sh05afc6d0, 32'sh05aca5bd, 32'sh05a984a6, 32'sh05a6638d, 32'sh05a3426f, 32'sh05a0214f, 32'sh059d002a, 32'sh0599df03, 
               32'sh0596bdd7, 32'sh05939ca9, 32'sh05907b77, 32'sh058d5a41, 32'sh058a3908, 32'sh058717cc, 32'sh0583f68c, 32'sh0580d549, 
               32'sh057db403, 32'sh057a92b9, 32'sh0577716b, 32'sh0574501b, 32'sh05712ec7, 32'sh056e0d6f, 32'sh056aec15, 32'sh0567cab6, 
               32'sh0564a955, 32'sh056187f0, 32'sh055e6688, 32'sh055b451d, 32'sh055823ae, 32'sh0555023c, 32'sh0551e0c7, 32'sh054ebf4e, 
               32'sh054b9dd3, 32'sh05487c53, 32'sh05455ad1, 32'sh0542394c, 32'sh053f17c3, 32'sh053bf637, 32'sh0538d4a7, 32'sh0535b315, 
               32'sh0532917f, 32'sh052f6fe6, 32'sh052c4e4a, 32'sh05292cab, 32'sh05260b08, 32'sh0522e962, 32'sh051fc7b9, 32'sh051ca60d, 
               32'sh0519845e, 32'sh051662ac, 32'sh051340f6, 32'sh05101f3e, 32'sh050cfd82, 32'sh0509dbc3, 32'sh0506ba01, 32'sh0503983c, 
               32'sh05007674, 32'sh04fd54a9, 32'sh04fa32db, 32'sh04f71109, 32'sh04f3ef35, 32'sh04f0cd5d, 32'sh04edab83, 32'sh04ea89a5, 
               32'sh04e767c5, 32'sh04e445e1, 32'sh04e123fa, 32'sh04de0211, 32'sh04dae024, 32'sh04d7be34, 32'sh04d49c42, 32'sh04d17a4c, 
               32'sh04ce5854, 32'sh04cb3658, 32'sh04c81459, 32'sh04c4f258, 32'sh04c1d054, 32'sh04beae4c, 32'sh04bb8c42, 32'sh04b86a35, 
               32'sh04b54825, 32'sh04b22612, 32'sh04af03fc, 32'sh04abe1e3, 32'sh04a8bfc7, 32'sh04a59da9, 32'sh04a27b87, 32'sh049f5963, 
               32'sh049c373c, 32'sh04991512, 32'sh0495f2e5, 32'sh0492d0b6, 32'sh048fae83, 32'sh048c8c4e, 32'sh04896a16, 32'sh048647db, 
               32'sh0483259d, 32'sh0480035d, 32'sh047ce11a, 32'sh0479bed4, 32'sh04769c8b, 32'sh04737a3f, 32'sh047057f1, 32'sh046d35a0, 
               32'sh046a134c, 32'sh0466f0f6, 32'sh0463ce9d, 32'sh0460ac41, 32'sh045d89e2, 32'sh045a6781, 32'sh0457451d, 32'sh045422b7, 
               32'sh0451004d, 32'sh044ddde1, 32'sh044abb73, 32'sh04479901, 32'sh0444768d, 32'sh04415417, 32'sh043e319e, 32'sh043b0f22, 
               32'sh0437eca4, 32'sh0434ca23, 32'sh0431a79f, 32'sh042e8519, 32'sh042b6290, 32'sh04284005, 32'sh04251d77, 32'sh0421fae7, 
               32'sh041ed854, 32'sh041bb5be, 32'sh04189326, 32'sh0415708b, 32'sh04124dee, 32'sh040f2b4f, 32'sh040c08ad, 32'sh0408e608, 
               32'sh0405c361, 32'sh0402a0b7, 32'sh03ff7e0b, 32'sh03fc5b5d, 32'sh03f938ac, 32'sh03f615f8, 32'sh03f2f342, 32'sh03efd08a, 
               32'sh03ecadcf, 32'sh03e98b12, 32'sh03e66852, 32'sh03e34591, 32'sh03e022cc, 32'sh03dd0005, 32'sh03d9dd3c, 32'sh03d6ba71, 
               32'sh03d397a3, 32'sh03d074d2, 32'sh03cd5200, 32'sh03ca2f2b, 32'sh03c70c54, 32'sh03c3e97a, 32'sh03c0c69e, 32'sh03bda3c0, 
               32'sh03ba80df, 32'sh03b75dfc, 32'sh03b43b17, 32'sh03b11830, 32'sh03adf546, 32'sh03aad25a, 32'sh03a7af6c, 32'sh03a48c7b, 
               32'sh03a16988, 32'sh039e4693, 32'sh039b239c, 32'sh039800a3, 32'sh0394dda7, 32'sh0391baa9, 32'sh038e97a9, 32'sh038b74a7, 
               32'sh038851a2, 32'sh03852e9c, 32'sh03820b93, 32'sh037ee888, 32'sh037bc57b, 32'sh0378a26b, 32'sh03757f5a, 32'sh03725c46, 
               32'sh036f3931, 32'sh036c1619, 32'sh0368f2ff, 32'sh0365cfe3, 32'sh0362acc5, 32'sh035f89a5, 32'sh035c6682, 32'sh0359435e, 
               32'sh03562038, 32'sh0352fd0f, 32'sh034fd9e5, 32'sh034cb6b8, 32'sh03499389, 32'sh03467059, 32'sh03434d26, 32'sh034029f2, 
               32'sh033d06bb, 32'sh0339e382, 32'sh0336c047, 32'sh03339d0b, 32'sh033079cc, 32'sh032d568c, 32'sh032a3349, 32'sh03271005, 
               32'sh0323ecbe, 32'sh0320c976, 32'sh031da62b, 32'sh031a82df, 32'sh03175f91, 32'sh03143c41, 32'sh031118ef, 32'sh030df59b, 
               32'sh030ad245, 32'sh0307aeee, 32'sh03048b94, 32'sh03016839, 32'sh02fe44dc, 32'sh02fb217d, 32'sh02f7fe1c, 32'sh02f4dab9, 
               32'sh02f1b755, 32'sh02ee93ee, 32'sh02eb7086, 32'sh02e84d1c, 32'sh02e529b0, 32'sh02e20643, 32'sh02dee2d4, 32'sh02dbbf63, 
               32'sh02d89bf0, 32'sh02d5787b, 32'sh02d25505, 32'sh02cf318d, 32'sh02cc0e13, 32'sh02c8ea97, 32'sh02c5c71a, 32'sh02c2a39b, 
               32'sh02bf801a, 32'sh02bc5c98, 32'sh02b93914, 32'sh02b6158e, 32'sh02b2f207, 32'sh02afce7e, 32'sh02acaaf3, 32'sh02a98766, 
               32'sh02a663d8, 32'sh02a34049, 32'sh02a01cb8, 32'sh029cf925, 32'sh0299d590, 32'sh0296b1fa, 32'sh02938e62, 32'sh02906ac9, 
               32'sh028d472e, 32'sh028a2392, 32'sh0286fff3, 32'sh0283dc54, 32'sh0280b8b3, 32'sh027d9510, 32'sh027a716c, 32'sh02774dc6, 
               32'sh02742a1f, 32'sh02710676, 32'sh026de2cc, 32'sh026abf20, 32'sh02679b73, 32'sh026477c4, 32'sh02615414, 32'sh025e3062, 
               32'sh025b0caf, 32'sh0257e8fa, 32'sh0254c544, 32'sh0251a18c, 32'sh024e7dd4, 32'sh024b5a19, 32'sh0248365d, 32'sh024512a0, 
               32'sh0241eee2, 32'sh023ecb22, 32'sh023ba760, 32'sh0238839e, 32'sh02355fd9, 32'sh02323c14, 32'sh022f184d, 32'sh022bf485, 
               32'sh0228d0bb, 32'sh0225acf1, 32'sh02228924, 32'sh021f6557, 32'sh021c4188, 32'sh02191db8, 32'sh0215f9e7, 32'sh0212d614, 
               32'sh020fb240, 32'sh020c8e6b, 32'sh02096a94, 32'sh020646bc, 32'sh020322e3, 32'sh01ffff09, 32'sh01fcdb2e, 32'sh01f9b751, 
               32'sh01f69373, 32'sh01f36f94, 32'sh01f04bb4, 32'sh01ed27d2, 32'sh01ea03ef, 32'sh01e6e00b, 32'sh01e3bc26, 32'sh01e09840, 
               32'sh01dd7459, 32'sh01da5070, 32'sh01d72c87, 32'sh01d4089c, 32'sh01d0e4b0, 32'sh01cdc0c3, 32'sh01ca9cd4, 32'sh01c778e5, 
               32'sh01c454f5, 32'sh01c13103, 32'sh01be0d11, 32'sh01bae91d, 32'sh01b7c528, 32'sh01b4a133, 32'sh01b17d3c, 32'sh01ae5944, 
               32'sh01ab354b, 32'sh01a81151, 32'sh01a4ed56, 32'sh01a1c95a, 32'sh019ea55d, 32'sh019b815f, 32'sh01985d60, 32'sh01953960, 
               32'sh0192155f, 32'sh018ef15e, 32'sh018bcd5b, 32'sh0188a957, 32'sh01858552, 32'sh0182614c, 32'sh017f3d46, 32'sh017c193e, 
               32'sh0178f536, 32'sh0175d12c, 32'sh0172ad22, 32'sh016f8917, 32'sh016c650b, 32'sh016940fe, 32'sh01661cf0, 32'sh0162f8e2, 
               32'sh015fd4d2, 32'sh015cb0c2, 32'sh01598cb1, 32'sh0156689f, 32'sh0153448c, 32'sh01502078, 32'sh014cfc63, 32'sh0149d84e, 
               32'sh0146b438, 32'sh01439021, 32'sh01406c0a, 32'sh013d47f1, 32'sh013a23d8, 32'sh0136ffbe, 32'sh0133dba3, 32'sh0130b788, 
               32'sh012d936c, 32'sh012a6f4f, 32'sh01274b31, 32'sh01242713, 32'sh012102f4, 32'sh011dded4, 32'sh011abab4, 32'sh01179693, 
               32'sh01147271, 32'sh01114e4e, 32'sh010e2a2b, 32'sh010b0608, 32'sh0107e1e3, 32'sh0104bdbe, 32'sh01019998, 32'sh00fe7572, 
               32'sh00fb514b, 32'sh00f82d24, 32'sh00f508fc, 32'sh00f1e4d3, 32'sh00eec0aa, 32'sh00eb9c80, 32'sh00e87856, 32'sh00e5542b, 
               32'sh00e22fff, 32'sh00df0bd3, 32'sh00dbe7a6, 32'sh00d8c379, 32'sh00d59f4c, 32'sh00d27b1d, 32'sh00cf56ef, 32'sh00cc32c0, 
               32'sh00c90e90, 32'sh00c5ea60, 32'sh00c2c62f, 32'sh00bfa1fe, 32'sh00bc7dcc, 32'sh00b9599a, 32'sh00b63568, 32'sh00b31135, 
               32'sh00afed02, 32'sh00acc8ce, 32'sh00a9a49a, 32'sh00a68065, 32'sh00a35c30, 32'sh00a037fb, 32'sh009d13c5, 32'sh0099ef8f, 
               32'sh0096cb58, 32'sh0093a722, 32'sh009082ea, 32'sh008d5eb3, 32'sh008a3a7b, 32'sh00871643, 32'sh0083f20a, 32'sh0080cdd1, 
               32'sh007da998, 32'sh007a855e, 32'sh00776125, 32'sh00743cea, 32'sh007118b0, 32'sh006df475, 32'sh006ad03b, 32'sh0067abff, 
               32'sh006487c4, 32'sh00616388, 32'sh005e3f4c, 32'sh005b1b10, 32'sh0057f6d4, 32'sh0054d297, 32'sh0051ae5b, 32'sh004e8a1e, 
               32'sh004b65e1, 32'sh004841a3, 32'sh00451d66, 32'sh0041f928, 32'sh003ed4ea, 32'sh003bb0ac, 32'sh00388c6e, 32'sh00356830, 
               32'sh003243f1, 32'sh002f1fb3, 32'sh002bfb74, 32'sh0028d736, 32'sh0025b2f7, 32'sh00228eb8, 32'sh001f6a79, 32'sh001c463a, 
               32'sh001921fb, 32'sh0015fdbb, 32'sh0012d97c, 32'sh000fb53d, 32'sh000c90fe, 32'sh00096cbe, 32'sh0006487f, 32'sh0003243f, 
               32'sh00000000, 32'shfffcdbc1, 32'shfff9b781, 32'shfff69342, 32'shfff36f02, 32'shfff04ac3, 32'shffed2684, 32'shffea0245, 
               32'shffe6de05, 32'shffe3b9c6, 32'shffe09587, 32'shffdd7148, 32'shffda4d09, 32'shffd728ca, 32'shffd4048c, 32'shffd0e04d, 
               32'shffcdbc0f, 32'shffca97d0, 32'shffc77392, 32'shffc44f54, 32'shffc12b16, 32'shffbe06d8, 32'shffbae29a, 32'shffb7be5d, 
               32'shffb49a1f, 32'shffb175e2, 32'shffae51a5, 32'shffab2d69, 32'shffa8092c, 32'shffa4e4f0, 32'shffa1c0b4, 32'shff9e9c78, 
               32'shff9b783c, 32'shff985401, 32'shff952fc5, 32'shff920b8b, 32'shff8ee750, 32'shff8bc316, 32'shff889edb, 32'shff857aa2, 
               32'shff825668, 32'shff7f322f, 32'shff7c0df6, 32'shff78e9bd, 32'shff75c585, 32'shff72a14d, 32'shff6f7d16, 32'shff6c58de, 
               32'shff6934a8, 32'shff661071, 32'shff62ec3b, 32'shff5fc805, 32'shff5ca3d0, 32'shff597f9b, 32'shff565b66, 32'shff533732, 
               32'shff5012fe, 32'shff4ceecb, 32'shff49ca98, 32'shff46a666, 32'shff438234, 32'shff405e02, 32'shff3d39d1, 32'shff3a15a0, 
               32'shff36f170, 32'shff33cd40, 32'shff30a911, 32'shff2d84e3, 32'shff2a60b4, 32'shff273c87, 32'shff24185a, 32'shff20f42d, 
               32'shff1dd001, 32'shff1aabd5, 32'shff1787aa, 32'shff146380, 32'shff113f56, 32'shff0e1b2d, 32'shff0af704, 32'shff07d2dc, 
               32'shff04aeb5, 32'shff018a8e, 32'shfefe6668, 32'shfefb4242, 32'shfef81e1d, 32'shfef4f9f8, 32'shfef1d5d5, 32'shfeeeb1b2, 
               32'shfeeb8d8f, 32'shfee8696d, 32'shfee5454c, 32'shfee2212c, 32'shfedefd0c, 32'shfedbd8ed, 32'shfed8b4cf, 32'shfed590b1, 
               32'shfed26c94, 32'shfecf4878, 32'shfecc245d, 32'shfec90042, 32'shfec5dc28, 32'shfec2b80f, 32'shfebf93f6, 32'shfebc6fdf, 
               32'shfeb94bc8, 32'shfeb627b2, 32'shfeb3039d, 32'shfeafdf88, 32'shfeacbb74, 32'shfea99761, 32'shfea6734f, 32'shfea34f3e, 
               32'shfea02b2e, 32'shfe9d071e, 32'shfe99e310, 32'shfe96bf02, 32'shfe939af5, 32'shfe9076e9, 32'shfe8d52de, 32'shfe8a2ed4, 
               32'shfe870aca, 32'shfe83e6c2, 32'shfe80c2ba, 32'shfe7d9eb4, 32'shfe7a7aae, 32'shfe7756a9, 32'shfe7432a5, 32'shfe710ea2, 
               32'shfe6deaa1, 32'shfe6ac6a0, 32'shfe67a2a0, 32'shfe647ea1, 32'shfe615aa3, 32'shfe5e36a6, 32'shfe5b12aa, 32'shfe57eeaf, 
               32'shfe54cab5, 32'shfe51a6bc, 32'shfe4e82c4, 32'shfe4b5ecd, 32'shfe483ad8, 32'shfe4516e3, 32'shfe41f2ef, 32'shfe3ecefd, 
               32'shfe3bab0b, 32'shfe38871b, 32'shfe35632c, 32'shfe323f3d, 32'shfe2f1b50, 32'shfe2bf764, 32'shfe28d379, 32'shfe25af90, 
               32'shfe228ba7, 32'shfe1f67c0, 32'shfe1c43da, 32'shfe191ff5, 32'shfe15fc11, 32'shfe12d82e, 32'shfe0fb44c, 32'shfe0c906c, 
               32'shfe096c8d, 32'shfe0648af, 32'shfe0324d2, 32'shfe0000f7, 32'shfdfcdd1d, 32'shfdf9b944, 32'shfdf6956c, 32'shfdf37195, 
               32'shfdf04dc0, 32'shfded29ec, 32'shfdea0619, 32'shfde6e248, 32'shfde3be78, 32'shfde09aa9, 32'shfddd76dc, 32'shfdda530f, 
               32'shfdd72f45, 32'shfdd40b7b, 32'shfdd0e7b3, 32'shfdcdc3ec, 32'shfdcaa027, 32'shfdc77c62, 32'shfdc458a0, 32'shfdc134de, 
               32'shfdbe111e, 32'shfdbaed60, 32'shfdb7c9a3, 32'shfdb4a5e7, 32'shfdb1822c, 32'shfdae5e74, 32'shfdab3abc, 32'shfda81706, 
               32'shfda4f351, 32'shfda1cf9e, 32'shfd9eabec, 32'shfd9b883c, 32'shfd98648d, 32'shfd9540e0, 32'shfd921d34, 32'shfd8ef98a, 
               32'shfd8bd5e1, 32'shfd88b23a, 32'shfd858e94, 32'shfd826af0, 32'shfd7f474d, 32'shfd7c23ac, 32'shfd79000d, 32'shfd75dc6e, 
               32'shfd72b8d2, 32'shfd6f9537, 32'shfd6c719e, 32'shfd694e06, 32'shfd662a70, 32'shfd6306db, 32'shfd5fe348, 32'shfd5cbfb7, 
               32'shfd599c28, 32'shfd56789a, 32'shfd53550d, 32'shfd503182, 32'shfd4d0df9, 32'shfd49ea72, 32'shfd46c6ec, 32'shfd43a368, 
               32'shfd407fe6, 32'shfd3d5c65, 32'shfd3a38e6, 32'shfd371569, 32'shfd33f1ed, 32'shfd30ce73, 32'shfd2daafb, 32'shfd2a8785, 
               32'shfd276410, 32'shfd24409d, 32'shfd211d2c, 32'shfd1df9bd, 32'shfd1ad650, 32'shfd17b2e4, 32'shfd148f7a, 32'shfd116c12, 
               32'shfd0e48ab, 32'shfd0b2547, 32'shfd0801e4, 32'shfd04de83, 32'shfd01bb24, 32'shfcfe97c7, 32'shfcfb746c, 32'shfcf85112, 
               32'shfcf52dbb, 32'shfcf20a65, 32'shfceee711, 32'shfcebc3bf, 32'shfce8a06f, 32'shfce57d21, 32'shfce259d5, 32'shfcdf368a, 
               32'shfcdc1342, 32'shfcd8effb, 32'shfcd5ccb7, 32'shfcd2a974, 32'shfccf8634, 32'shfccc62f5, 32'shfcc93fb9, 32'shfcc61c7e, 
               32'shfcc2f945, 32'shfcbfd60e, 32'shfcbcb2da, 32'shfcb98fa7, 32'shfcb66c77, 32'shfcb34948, 32'shfcb0261b, 32'shfcad02f1, 
               32'shfca9dfc8, 32'shfca6bca2, 32'shfca3997e, 32'shfca0765b, 32'shfc9d533b, 32'shfc9a301d, 32'shfc970d01, 32'shfc93e9e7, 
               32'shfc90c6cf, 32'shfc8da3ba, 32'shfc8a80a6, 32'shfc875d95, 32'shfc843a85, 32'shfc811778, 32'shfc7df46d, 32'shfc7ad164, 
               32'shfc77ae5e, 32'shfc748b59, 32'shfc716857, 32'shfc6e4557, 32'shfc6b2259, 32'shfc67ff5d, 32'shfc64dc64, 32'shfc61b96d, 
               32'shfc5e9678, 32'shfc5b7385, 32'shfc585094, 32'shfc552da6, 32'shfc520aba, 32'shfc4ee7d0, 32'shfc4bc4e9, 32'shfc48a204, 
               32'shfc457f21, 32'shfc425c40, 32'shfc3f3962, 32'shfc3c1686, 32'shfc38f3ac, 32'shfc35d0d5, 32'shfc32ae00, 32'shfc2f8b2e, 
               32'shfc2c685d, 32'shfc29458f, 32'shfc2622c4, 32'shfc22fffb, 32'shfc1fdd34, 32'shfc1cba6f, 32'shfc1997ae, 32'shfc1674ee, 
               32'shfc135231, 32'shfc102f76, 32'shfc0d0cbe, 32'shfc09ea08, 32'shfc06c754, 32'shfc03a4a3, 32'shfc0081f5, 32'shfbfd5f49, 
               32'shfbfa3c9f, 32'shfbf719f8, 32'shfbf3f753, 32'shfbf0d4b1, 32'shfbedb212, 32'shfbea8f75, 32'shfbe76cda, 32'shfbe44a42, 
               32'shfbe127ac, 32'shfbde0519, 32'shfbdae289, 32'shfbd7bffb, 32'shfbd49d70, 32'shfbd17ae7, 32'shfbce5861, 32'shfbcb35dd, 
               32'shfbc8135c, 32'shfbc4f0de, 32'shfbc1ce62, 32'shfbbeabe9, 32'shfbbb8973, 32'shfbb866ff, 32'shfbb5448d, 32'shfbb2221f, 
               32'shfbaeffb3, 32'shfbabdd49, 32'shfba8bae3, 32'shfba5987f, 32'shfba2761e, 32'shfb9f53bf, 32'shfb9c3163, 32'shfb990f0a, 
               32'shfb95ecb4, 32'shfb92ca60, 32'shfb8fa80f, 32'shfb8c85c1, 32'shfb896375, 32'shfb86412c, 32'shfb831ee6, 32'shfb7ffca3, 
               32'shfb7cda63, 32'shfb79b825, 32'shfb7695ea, 32'shfb7373b2, 32'shfb70517d, 32'shfb6d2f4a, 32'shfb6a0d1b, 32'shfb66eaee, 
               32'shfb63c8c4, 32'shfb60a69d, 32'shfb5d8479, 32'shfb5a6257, 32'shfb574039, 32'shfb541e1d, 32'shfb50fc04, 32'shfb4dd9ee, 
               32'shfb4ab7db, 32'shfb4795cb, 32'shfb4473be, 32'shfb4151b4, 32'shfb3e2fac, 32'shfb3b0da8, 32'shfb37eba7, 32'shfb34c9a8, 
               32'shfb31a7ac, 32'shfb2e85b4, 32'shfb2b63be, 32'shfb2841cc, 32'shfb251fdc, 32'shfb21fdef, 32'shfb1edc06, 32'shfb1bba1f, 
               32'shfb18983b, 32'shfb15765b, 32'shfb12547d, 32'shfb0f32a3, 32'shfb0c10cb, 32'shfb08eef7, 32'shfb05cd25, 32'shfb02ab57, 
               32'shfaff898c, 32'shfafc67c4, 32'shfaf945ff, 32'shfaf6243d, 32'shfaf3027e, 32'shfaefe0c2, 32'shfaecbf0a, 32'shfae99d54, 
               32'shfae67ba2, 32'shfae359f3, 32'shfae03847, 32'shfadd169e, 32'shfad9f4f8, 32'shfad6d355, 32'shfad3b1b6, 32'shfad0901a, 
               32'shfacd6e81, 32'shfaca4ceb, 32'shfac72b59, 32'shfac409c9, 32'shfac0e83d, 32'shfabdc6b4, 32'shfabaa52f, 32'shfab783ad, 
               32'shfab4622d, 32'shfab140b2, 32'shfaae1f39, 32'shfaaafdc4, 32'shfaa7dc52, 32'shfaa4bae3, 32'shfaa19978, 32'shfa9e7810, 
               32'shfa9b56ab, 32'shfa98354a, 32'shfa9513eb, 32'shfa91f291, 32'shfa8ed139, 32'shfa8bafe5, 32'shfa888e95, 32'shfa856d47, 
               32'shfa824bfd, 32'shfa7f2ab7, 32'shfa7c0974, 32'shfa78e834, 32'shfa75c6f8, 32'shfa72a5bf, 32'shfa6f8489, 32'shfa6c6357, 
               32'shfa694229, 32'shfa6620fd, 32'shfa62ffd6, 32'shfa5fdeb1, 32'shfa5cbd91, 32'shfa599c73, 32'shfa567b5a, 32'shfa535a43, 
               32'shfa503930, 32'shfa4d1821, 32'shfa49f715, 32'shfa46d60d, 32'shfa43b508, 32'shfa409407, 32'shfa3d7309, 32'shfa3a520f, 
               32'shfa373119, 32'shfa341026, 32'shfa30ef36, 32'shfa2dce4b, 32'shfa2aad62, 32'shfa278c7e, 32'shfa246b9d, 32'shfa214abf, 
               32'shfa1e29e5, 32'shfa1b090f, 32'shfa17e83d, 32'shfa14c76e, 32'shfa11a6a3, 32'shfa0e85db, 32'shfa0b6517, 32'shfa084457, 
               32'shfa05239a, 32'shfa0202e1, 32'shf9fee22c, 32'shf9fbc17b, 32'shf9f8a0cd, 32'shf9f58023, 32'shf9f25f7d, 32'shf9ef3eda, 
               32'shf9ec1e3b, 32'shf9e8fda0, 32'shf9e5dd09, 32'shf9e2bc75, 32'shf9df9be6, 32'shf9dc7b5a, 32'shf9d95ad1, 32'shf9d63a4d, 
               32'shf9d319cc, 32'shf9cff94f, 32'shf9ccd8d6, 32'shf9c9b861, 32'shf9c697f0, 32'shf9c37782, 32'shf9c05719, 32'shf9bd36b3, 
               32'shf9ba1651, 32'shf9b6f5f3, 32'shf9b3d599, 32'shf9b0b542, 32'shf9ad94f0, 32'shf9aa74a1, 32'shf9a75457, 32'shf9a43410, 
               32'shf9a113cd, 32'shf99df38e, 32'shf99ad354, 32'shf997b31d, 32'shf99492ea, 32'shf99172bb, 32'shf98e528f, 32'shf98b3268, 
               32'shf9881245, 32'shf984f226, 32'shf981d20b, 32'shf97eb1f4, 32'shf97b91e1, 32'shf97871d2, 32'shf97551c6, 32'shf97231bf, 
               32'shf96f11bc, 32'shf96bf1be, 32'shf968d1c3, 32'shf965b1cc, 32'shf96291d9, 32'shf95f71ea, 32'shf95c5200, 32'shf9593219, 
               32'shf9561237, 32'shf952f259, 32'shf94fd27f, 32'shf94cb2a8, 32'shf94992d7, 32'shf9467309, 32'shf943533f, 32'shf940337a, 
               32'shf93d13b8, 32'shf939f3fb, 32'shf936d442, 32'shf933b48e, 32'shf93094dd, 32'shf92d7531, 32'shf92a5589, 32'shf92735e5, 
               32'shf9241645, 32'shf920f6a9, 32'shf91dd712, 32'shf91ab77f, 32'shf91797f0, 32'shf9147866, 32'shf91158e0, 32'shf90e395e, 
               32'shf90b19e0, 32'shf907fa67, 32'shf904daf2, 32'shf901bb81, 32'shf8fe9c15, 32'shf8fb7cac, 32'shf8f85d49, 32'shf8f53de9, 
               32'shf8f21e8e, 32'shf8eeff37, 32'shf8ebdfe5, 32'shf8e8c097, 32'shf8e5a14d, 32'shf8e28208, 32'shf8df62c7, 32'shf8dc438b, 
               32'shf8d92452, 32'shf8d6051f, 32'shf8d2e5f0, 32'shf8cfc6c5, 32'shf8cca79e, 32'shf8c9887c, 32'shf8c6695f, 32'shf8c34a46, 
               32'shf8c02b31, 32'shf8bd0c21, 32'shf8b9ed15, 32'shf8b6ce0e, 32'shf8b3af0c, 32'shf8b0900d, 32'shf8ad7114, 32'shf8aa521f, 
               32'shf8a7332e, 32'shf8a41442, 32'shf8a0f55b, 32'shf89dd678, 32'shf89ab799, 32'shf89798bf, 32'shf89479ea, 32'shf8915b19, 
               32'shf88e3c4d, 32'shf88b1d86, 32'shf887fec3, 32'shf884e004, 32'shf881c14b, 32'shf87ea295, 32'shf87b83e5, 32'shf8786539, 
               32'shf8754692, 32'shf87227ef, 32'shf86f0952, 32'shf86beab8, 32'shf868cc24, 32'shf865ad94, 32'shf8628f09, 32'shf85f7082, 
               32'shf85c5201, 32'shf8593383, 32'shf856150b, 32'shf852f698, 32'shf84fd829, 32'shf84cb9bf, 32'shf8499b59, 32'shf8467cf9, 
               32'shf8435e9d, 32'shf8404046, 32'shf83d21f3, 32'shf83a03a6, 32'shf836e55d, 32'shf833c719, 32'shf830a8da, 32'shf82d8aa0, 
               32'shf82a6c6a, 32'shf8274e3a, 32'shf824300e, 32'shf82111e7, 32'shf81df3c5, 32'shf81ad5a8, 32'shf817b78f, 32'shf814997c, 
               32'shf8117b6d, 32'shf80e5d64, 32'shf80b3f5f, 32'shf808215f, 32'shf8050364, 32'shf801e56e, 32'shf7fec77d, 32'shf7fba991, 
               32'shf7f88ba9, 32'shf7f56dc7, 32'shf7f24fea, 32'shf7ef3211, 32'shf7ec143e, 32'shf7e8f670, 32'shf7e5d8a6, 32'shf7e2bae2, 
               32'shf7df9d22, 32'shf7dc7f68, 32'shf7d961b3, 32'shf7d64402, 32'shf7d32657, 32'shf7d008b1, 32'shf7cceb0f, 32'shf7c9cd73, 
               32'shf7c6afdc, 32'shf7c3924a, 32'shf7c074bd, 32'shf7bd5735, 32'shf7ba39b3, 32'shf7b71c35, 32'shf7b3febc, 32'shf7b0e149, 
               32'shf7adc3db, 32'shf7aaa671, 32'shf7a7890d, 32'shf7a46baf, 32'shf7a14e55, 32'shf79e3100, 32'shf79b13b1, 32'shf797f667, 
               32'shf794d922, 32'shf791bbe2, 32'shf78e9ea7, 32'shf78b8172, 32'shf7886442, 32'shf7854717, 32'shf78229f1, 32'shf77f0cd0, 
               32'shf77befb5, 32'shf778d29f, 32'shf775b58e, 32'shf7729883, 32'shf76f7b7d, 32'shf76c5e7c, 32'shf7694180, 32'shf766248a, 
               32'shf7630799, 32'shf75feaad, 32'shf75ccdc6, 32'shf759b0e5, 32'shf756940a, 32'shf7537733, 32'shf7505a62, 32'shf74d3d96, 
               32'shf74a20d0, 32'shf747040f, 32'shf743e754, 32'shf740ca9d, 32'shf73daded, 32'shf73a9141, 32'shf737749b, 32'shf73457fb, 
               32'shf7313b60, 32'shf72e1eca, 32'shf72b023a, 32'shf727e5af, 32'shf724c92a, 32'shf721acaa, 32'shf71e902f, 32'shf71b73ba, 
               32'shf718574b, 32'shf7153ae1, 32'shf7121e7c, 32'shf70f021d, 32'shf70be5c4, 32'shf708c970, 32'shf705ad22, 32'shf70290d9, 
               32'shf6ff7496, 32'shf6fc5858, 32'shf6f93c20, 32'shf6f61fed, 32'shf6f303c0, 32'shf6efe798, 32'shf6eccb77, 32'shf6e9af5a, 
               32'shf6e69344, 32'shf6e37733, 32'shf6e05b27, 32'shf6dd3f21, 32'shf6da2321, 32'shf6d70727, 32'shf6d3eb32, 32'shf6d0cf43, 
               32'shf6cdb359, 32'shf6ca9775, 32'shf6c77b97, 32'shf6c45fbe, 32'shf6c143ec, 32'shf6be281e, 32'shf6bb0c57, 32'shf6b7f095, 
               32'shf6b4d4d9, 32'shf6b1b923, 32'shf6ae9d73, 32'shf6ab81c8, 32'shf6a86623, 32'shf6a54a84, 32'shf6a22eea, 32'shf69f1357, 
               32'shf69bf7c9, 32'shf698dc41, 32'shf695c0be, 32'shf692a542, 32'shf68f89cb, 32'shf68c6e5a, 32'shf68952ef, 32'shf686378a, 
               32'shf6831c2b, 32'shf68000d1, 32'shf67ce57e, 32'shf679ca30, 32'shf676aee8, 32'shf67393a6, 32'shf670786a, 32'shf66d5d34, 
               32'shf66a4203, 32'shf66726d9, 32'shf6640bb4, 32'shf660f096, 32'shf65dd57d, 32'shf65aba6b, 32'shf6579f5e, 32'shf6548457, 
               32'shf6516956, 32'shf64e4e5c, 32'shf64b3367, 32'shf6481878, 32'shf644fd8f, 32'shf641e2ac, 32'shf63ec7cf, 32'shf63bacf8, 
               32'shf6389228, 32'shf635775d, 32'shf6325c98, 32'shf62f41d9, 32'shf62c2721, 32'shf6290c6e, 32'shf625f1c2, 32'shf622d71b, 
               32'shf61fbc7b, 32'shf61ca1e1, 32'shf619874c, 32'shf6166cbe, 32'shf6135237, 32'shf61037b5, 32'shf60d1d39, 32'shf60a02c3, 
               32'shf606e854, 32'shf603cdeb, 32'shf600b388, 32'shf5fd992b, 32'shf5fa7ed4, 32'shf5f76484, 32'shf5f44a39, 32'shf5f12ff5, 
               32'shf5ee15b7, 32'shf5eafb7f, 32'shf5e7e14e, 32'shf5e4c722, 32'shf5e1acfd, 32'shf5de92de, 32'shf5db78c6, 32'shf5d85eb3, 
               32'shf5d544a7, 32'shf5d22aa2, 32'shf5cf10a2, 32'shf5cbf6a9, 32'shf5c8dcb6, 32'shf5c5c2c9, 32'shf5c2a8e3, 32'shf5bf8f03, 
               32'shf5bc7529, 32'shf5b95b56, 32'shf5b64189, 32'shf5b327c2, 32'shf5b00e02, 32'shf5acf448, 32'shf5a9da94, 32'shf5a6c0e7, 
               32'shf5a3a740, 32'shf5a08da0, 32'shf59d7406, 32'shf59a5a72, 32'shf59740e5, 32'shf594275e, 32'shf5910dde, 32'shf58df464, 
               32'shf58adaf0, 32'shf587c183, 32'shf584a81d, 32'shf5818ebd, 32'shf57e7563, 32'shf57b5c10, 32'shf57842c3, 32'shf575297d, 
               32'shf572103d, 32'shf56ef704, 32'shf56bddd1, 32'shf568c4a5, 32'shf565ab80, 32'shf5629261, 32'shf55f7948, 32'shf55c6036, 
               32'shf559472b, 32'shf5562e26, 32'shf5531528, 32'shf54ffc30, 32'shf54ce33f, 32'shf549ca55, 32'shf546b171, 32'shf5439893, 
               32'shf5407fbd, 32'shf53d66ed, 32'shf53a4e24, 32'shf5373561, 32'shf5341ca5, 32'shf53103ef, 32'shf52deb41, 32'shf52ad299, 
               32'shf527b9f7, 32'shf524a15d, 32'shf52188c9, 32'shf51e703b, 32'shf51b57b5, 32'shf5183f35, 32'shf51526bc, 32'shf5120e49, 
               32'shf50ef5de, 32'shf50bdd79, 32'shf508c51b, 32'shf505acc3, 32'shf5029473, 32'shf4ff7c29, 32'shf4fc63e6, 32'shf4f94baa, 
               32'shf4f63374, 32'shf4f31b46, 32'shf4f0031e, 32'shf4eceafd, 32'shf4e9d2e3, 32'shf4e6bacf, 32'shf4e3a2c3, 32'shf4e08abd, 
               32'shf4dd72be, 32'shf4da5ac7, 32'shf4d742d6, 32'shf4d42aeb, 32'shf4d11308, 32'shf4cdfb2c, 32'shf4cae356, 32'shf4c7cb88, 
               32'shf4c4b3c0, 32'shf4c19c00, 32'shf4be8446, 32'shf4bb6c93, 32'shf4b854e7, 32'shf4b53d42, 32'shf4b225a4, 32'shf4af0e0d, 
               32'shf4abf67e, 32'shf4a8def5, 32'shf4a5c773, 32'shf4a2aff8, 32'shf49f9884, 32'shf49c8117, 32'shf49969b1, 32'shf4965252, 
               32'shf4933afa, 32'shf49023a9, 32'shf48d0c5f, 32'shf489f51d, 32'shf486dde1, 32'shf483c6ad, 32'shf480af7f, 32'shf47d9859, 
               32'shf47a8139, 32'shf4776a21, 32'shf4745310, 32'shf4713c06, 32'shf46e2504, 32'shf46b0e08, 32'shf467f713, 32'shf464e026, 
               32'shf461c940, 32'shf45eb261, 32'shf45b9b89, 32'shf45884b8, 32'shf4556def, 32'shf452572c, 32'shf44f4071, 32'shf44c29be, 
               32'shf4491311, 32'shf445fc6b, 32'shf442e5cd, 32'shf43fcf36, 32'shf43cb8a7, 32'shf439a21e, 32'shf4368b9d, 32'shf4337523, 
               32'shf4305eb0, 32'shf42d4845, 32'shf42a31e1, 32'shf4271b84, 32'shf424052f, 32'shf420eee1, 32'shf41dd89a, 32'shf41ac25a, 
               32'shf417ac22, 32'shf41495f1, 32'shf4117fc8, 32'shf40e69a6, 32'shf40b538b, 32'shf4083d78, 32'shf405276c, 32'shf4021167, 
               32'shf3fefb6a, 32'shf3fbe574, 32'shf3f8cf86, 32'shf3f5b99f, 32'shf3f2a3bf, 32'shf3ef8de7, 32'shf3ec7817, 32'shf3e9624d, 
               32'shf3e64c8c, 32'shf3e336d1, 32'shf3e0211f, 32'shf3dd0b73, 32'shf3d9f5cf, 32'shf3d6e033, 32'shf3d3ca9e, 32'shf3d0b511, 
               32'shf3cd9f8b, 32'shf3ca8a0d, 32'shf3c77496, 32'shf3c45f27, 32'shf3c149bf, 32'shf3be345f, 32'shf3bb1f07, 32'shf3b809b6, 
               32'shf3b4f46c, 32'shf3b1df2a, 32'shf3aec9f0, 32'shf3abb4bd, 32'shf3a89f92, 32'shf3a58a6f, 32'shf3a27553, 32'shf39f603f, 
               32'shf39c4b32, 32'shf399362d, 32'shf3962130, 32'shf3930c3b, 32'shf38ff74d, 32'shf38ce266, 32'shf389cd88, 32'shf386b8b1, 
               32'shf383a3e2, 32'shf3808f1a, 32'shf37d7a5b, 32'shf37a65a2, 32'shf37750f2, 32'shf3743c49, 32'shf37127a9, 32'shf36e130f, 
               32'shf36afe7e, 32'shf367e9f4, 32'shf364d573, 32'shf361c0f9, 32'shf35eac86, 32'shf35b981c, 32'shf35883b9, 32'shf3556f5e, 
               32'shf3525b0b, 32'shf34f46c0, 32'shf34c327c, 32'shf3491e41, 32'shf3460a0d, 32'shf342f5e1, 32'shf33fe1bd, 32'shf33ccda1, 
               32'shf339b98d, 32'shf336a580, 32'shf333917c, 32'shf3307d7f, 32'shf32d698a, 32'shf32a559e, 32'shf32741b9, 32'shf3242ddc, 
               32'shf3211a07, 32'shf31e0639, 32'shf31af274, 32'shf317deb7, 32'shf314cb02, 32'shf311b755, 32'shf30ea3af, 32'shf30b9012, 
               32'shf3087c7d, 32'shf30568ef, 32'shf302556a, 32'shf2ff41ed, 32'shf2fc2e77, 32'shf2f91b0a, 32'shf2f607a5, 32'shf2f2f448, 
               32'shf2efe0f2, 32'shf2eccda5, 32'shf2e9ba60, 32'shf2e6a723, 32'shf2e393ef, 32'shf2e080c2, 32'shf2dd6d9d, 32'shf2da5a81, 
               32'shf2d7476c, 32'shf2d43460, 32'shf2d1215b, 32'shf2ce0e5f, 32'shf2cafb6b, 32'shf2c7e880, 32'shf2c4d59c, 32'shf2c1c2c0, 
               32'shf2beafed, 32'shf2bb9d22, 32'shf2b88a5f, 32'shf2b577a4, 32'shf2b264f2, 32'shf2af5247, 32'shf2ac3fa5, 32'shf2a92d0b, 
               32'shf2a61a7a, 32'shf2a307f0, 32'shf29ff56f, 32'shf29ce2f6, 32'shf299d085, 32'shf296be1d, 32'shf293abbd, 32'shf2909965, 
               32'shf28d8715, 32'shf28a74ce, 32'shf287628f, 32'shf2845058, 32'shf2813e2a, 32'shf27e2c04, 32'shf27b19e6, 32'shf27807d0, 
               32'shf274f5c3, 32'shf271e3bf, 32'shf26ed1c2, 32'shf26bbfce, 32'shf268ade3, 32'shf2659c00, 32'shf2628a25, 32'shf25f7852, 
               32'shf25c6688, 32'shf25954c7, 32'shf256430e, 32'shf253315d, 32'shf2501fb5, 32'shf24d0e15, 32'shf249fc7d, 32'shf246eaee, 
               32'shf243d968, 32'shf240c7ea, 32'shf23db674, 32'shf23aa507, 32'shf23793a3, 32'shf2348247, 32'shf23170f3, 32'shf22e5fa8, 
               32'shf22b4e66, 32'shf2283d2c, 32'shf2252bfa, 32'shf2221ad1, 32'shf21f09b1, 32'shf21bf899, 32'shf218e78a, 32'shf215d683, 
               32'shf212c585, 32'shf20fb490, 32'shf20ca3a3, 32'shf20992bf, 32'shf20681e3, 32'shf2037110, 32'shf2006046, 32'shf1fd4f84, 
               32'shf1fa3ecb, 32'shf1f72e1a, 32'shf1f41d72, 32'shf1f10cd3, 32'shf1edfc3d, 32'shf1eaebaf, 32'shf1e7db2a, 32'shf1e4caae, 
               32'shf1e1ba3a, 32'shf1dea9cf, 32'shf1db996d, 32'shf1d88913, 32'shf1d578c2, 32'shf1d2687a, 32'shf1cf583b, 32'shf1cc4804, 
               32'shf1c937d6, 32'shf1c627b1, 32'shf1c31795, 32'shf1c00781, 32'shf1bcf777, 32'shf1b9e775, 32'shf1b6d77c, 32'shf1b3c78b, 
               32'shf1b0b7a4, 32'shf1ada7c5, 32'shf1aa97ef, 32'shf1a78822, 32'shf1a4785e, 32'shf1a168a3, 32'shf19e58f1, 32'shf19b4947, 
               32'shf19839a6, 32'shf1952a0f, 32'shf1921a80, 32'shf18f0afa, 32'shf18bfb7d, 32'shf188ec09, 32'shf185dc9d, 32'shf182cd3b, 
               32'shf17fbde2, 32'shf17cae91, 32'shf1799f4a, 32'shf176900b, 32'shf17380d6, 32'shf17071a9, 32'shf16d6286, 32'shf16a536b, 
               32'shf1674459, 32'shf1643551, 32'shf1612651, 32'shf15e175b, 32'shf15b086d, 32'shf157f989, 32'shf154eaad, 32'shf151dbdb, 
               32'shf14ecd11, 32'shf14bbe51, 32'shf148af9a, 32'shf145a0ec, 32'shf1429247, 32'shf13f83ab, 32'shf13c7518, 32'shf139668e, 
               32'shf136580d, 32'shf1334996, 32'shf1303b27, 32'shf12d2cc2, 32'shf12a1e66, 32'shf1271013, 32'shf12401c9, 32'shf120f389, 
               32'shf11de551, 32'shf11ad723, 32'shf117c8fe, 32'shf114bae2, 32'shf111accf, 32'shf10e9ec6, 32'shf10b90c5, 32'shf10882ce, 
               32'shf10574e0, 32'shf10266fc, 32'shf0ff5921, 32'shf0fc4b4f, 32'shf0f93d86, 32'shf0f62fc6, 32'shf0f32210, 32'shf0f01463, 
               32'shf0ed06bf, 32'shf0e9f925, 32'shf0e6eb94, 32'shf0e3de0c, 32'shf0e0d08d, 32'shf0ddc318, 32'shf0dab5ad, 32'shf0d7a84a, 
               32'shf0d49af1, 32'shf0d18da1, 32'shf0ce805b, 32'shf0cb731e, 32'shf0c865ea, 32'shf0c558c0, 32'shf0c24b9f, 32'shf0bf3e88, 
               32'shf0bc317a, 32'shf0b92475, 32'shf0b6177a, 32'shf0b30a88, 32'shf0affda0, 32'shf0acf0c1, 32'shf0a9e3eb, 32'shf0a6d71f, 
               32'shf0a3ca5d, 32'shf0a0bda4, 32'shf09db0f4, 32'shf09aa44e, 32'shf09797b2, 32'shf0948b1f, 32'shf0917e95, 32'shf08e7215, 
               32'shf08b659f, 32'shf0885932, 32'shf0854cce, 32'shf0824074, 32'shf07f3424, 32'shf07c27dd, 32'shf0791ba0, 32'shf0760f6c, 
               32'shf0730342, 32'shf06ff722, 32'shf06ceb0b, 32'shf069defe, 32'shf066d2fa, 32'shf063c700, 32'shf060bb10, 32'shf05daf29, 
               32'shf05aa34c, 32'shf0579779, 32'shf0548baf, 32'shf0517fef, 32'shf04e7438, 32'shf04b688c, 32'shf0485ce9, 32'shf045514f, 
               32'shf04245c0, 32'shf03f3a3a, 32'shf03c2ebd, 32'shf039234b, 32'shf03617e2, 32'shf0330c83, 32'shf030012e, 32'shf02cf5e2, 
               32'shf029eaa1, 32'shf026df68, 32'shf023d43a, 32'shf020c916, 32'shf01dbdfb, 32'shf01ab2ea, 32'shf017a7e3, 32'shf0149ce6, 
               32'shf01191f3, 32'shf00e8709, 32'shf00b7c29, 32'shf0087153, 32'shf0056687, 32'shf0025bc5, 32'shefff510d, 32'sheffc465e, 
               32'sheff93bba, 32'sheff6311f, 32'sheff3268e, 32'sheff01c07, 32'shefed118a, 32'shefea0717, 32'shefe6fcae, 32'shefe3f24f, 
               32'shefe0e7f9, 32'shefddddae, 32'shefdad36c, 32'shefd7c935, 32'shefd4bf08, 32'shefd1b4e4, 32'shefceaacb, 32'shefcba0bb, 
               32'shefc896b5, 32'shefc58cba, 32'shefc282c8, 32'shefbf78e1, 32'shefbc6f03, 32'shefb96530, 32'shefb65b66, 32'shefb351a7, 
               32'shefb047f2, 32'shefad3e47, 32'shefaa34a5, 32'shefa72b0e, 32'shefa42181, 32'shefa117fe, 32'shef9e0e85, 32'shef9b0517, 
               32'shef97fbb2, 32'shef94f258, 32'shef91e907, 32'shef8edfc1, 32'shef8bd685, 32'shef88cd53, 32'shef85c42b, 32'shef82bb0e, 
               32'shef7fb1fa, 32'shef7ca8f1, 32'shef799ff2, 32'shef7696fd, 32'shef738e12, 32'shef708532, 32'shef6d7c5b, 32'shef6a738f, 
               32'shef676ace, 32'shef646216, 32'shef615969, 32'shef5e50c6, 32'shef5b482d, 32'shef583f9e, 32'shef55371a, 32'shef522ea0, 
               32'shef4f2630, 32'shef4c1dcb, 32'shef491570, 32'shef460d1f, 32'shef4304d8, 32'shef3ffc9c, 32'shef3cf46a, 32'shef39ec43, 
               32'shef36e426, 32'shef33dc13, 32'shef30d40a, 32'shef2dcc0c, 32'shef2ac419, 32'shef27bc2f, 32'shef24b451, 32'shef21ac7c, 
               32'shef1ea4b2, 32'shef1b9cf2, 32'shef18953d, 32'shef158d92, 32'shef1285f2, 32'shef0f7e5c, 32'shef0c76d0, 32'shef096f4f, 
               32'shef0667d9, 32'shef03606c, 32'shef00590b, 32'sheefd51b4, 32'sheefa4a67, 32'sheef74325, 32'sheef43bed, 32'sheef134c0, 
               32'sheeee2d9d, 32'sheeeb2685, 32'sheee81f78, 32'sheee51875, 32'sheee2117c, 32'sheedf0a8e, 32'sheedc03ab, 32'sheed8fcd2, 
               32'sheed5f604, 32'sheed2ef40, 32'sheecfe887, 32'sheecce1d9, 32'sheec9db35, 32'sheec6d49c, 32'sheec3ce0d, 32'sheec0c78a, 
               32'sheebdc110, 32'sheebabaa2, 32'sheeb7b43e, 32'sheeb4ade4, 32'sheeb1a796, 32'sheeaea152, 32'sheeab9b18, 32'sheea894ea, 
               32'sheea58ec6, 32'sheea288ad, 32'shee9f829e, 32'shee9c7c9a, 32'shee9976a1, 32'shee9670b3, 32'shee936acf, 32'shee9064f7, 
               32'shee8d5f29, 32'shee8a5965, 32'shee8753ad, 32'shee844dff, 32'shee81485c, 32'shee7e42c4, 32'shee7b3d36, 32'shee7837b4, 
               32'shee75323c, 32'shee722ccf, 32'shee6f276d, 32'shee6c2216, 32'shee691cc9, 32'shee661788, 32'shee631251, 32'shee600d25, 
               32'shee5d0804, 32'shee5a02ee, 32'shee56fde3, 32'shee53f8e2, 32'shee50f3ed, 32'shee4def02, 32'shee4aea23, 32'shee47e54e, 
               32'shee44e084, 32'shee41dbc6, 32'shee3ed712, 32'shee3bd269, 32'shee38cdcb, 32'shee35c938, 32'shee32c4b0, 32'shee2fc033, 
               32'shee2cbbc1, 32'shee29b75a, 32'shee26b2fe, 32'shee23aead, 32'shee20aa67, 32'shee1da62c, 32'shee1aa1fc, 32'shee179dd7, 
               32'shee1499bd, 32'shee1195ae, 32'shee0e91aa, 32'shee0b8db1, 32'shee0889c4, 32'shee0585e1, 32'shee02820a, 32'shedff7e3d, 
               32'shedfc7a7c, 32'shedf976c6, 32'shedf6731b, 32'shedf36f7b, 32'shedf06be6, 32'sheded685d, 32'shedea64de, 32'shede7616b, 
               32'shede45e03, 32'shede15aa6, 32'shedde5754, 32'sheddb540d, 32'shedd850d2, 32'shedd54da2, 32'shedd24a7d, 32'shedcf4763, 
               32'shedcc4454, 32'shedc94151, 32'shedc63e59, 32'shedc33b6c, 32'shedc0388a, 32'shedbd35b4, 32'shedba32e9, 32'shedb73029, 
               32'shedb42d74, 32'shedb12acb, 32'shedae282d, 32'shedab259a, 32'sheda82313, 32'sheda52097, 32'sheda21e26, 32'shed9f1bc1, 
               32'shed9c1967, 32'shed991718, 32'shed9614d5, 32'shed93129d, 32'shed901070, 32'shed8d0e4f, 32'shed8a0c39, 32'shed870a2e, 
               32'shed84082f, 32'shed81063b, 32'shed7e0453, 32'shed7b0276, 32'shed7800a5, 32'shed74fedf, 32'shed71fd24, 32'shed6efb75, 
               32'shed6bf9d1, 32'shed68f839, 32'shed65f6ac, 32'shed62f52b, 32'shed5ff3b5, 32'shed5cf24b, 32'shed59f0ec, 32'shed56ef99, 
               32'shed53ee51, 32'shed50ed14, 32'shed4debe4, 32'shed4aeabe, 32'shed47e9a5, 32'shed44e897, 32'shed41e794, 32'shed3ee69d, 
               32'shed3be5b1, 32'shed38e4d2, 32'shed35e3fd, 32'shed32e334, 32'shed2fe277, 32'shed2ce1c6, 32'shed29e120, 32'shed26e086, 
               32'shed23dff7, 32'shed20df74, 32'shed1ddefd, 32'shed1ade91, 32'shed17de31, 32'shed14dddc, 32'shed11dd94, 32'shed0edd56, 
               32'shed0bdd25, 32'shed08dcff, 32'shed05dce5, 32'shed02dcd7, 32'shecffdcd4, 32'shecfcdcde, 32'shecf9dcf3, 32'shecf6dd13, 
               32'shecf3dd3f, 32'shecf0dd78, 32'shecedddbb, 32'sheceade0b, 32'shece7de66, 32'shece4dece, 32'shece1df40, 32'shecdedfbf, 
               32'shecdbe04a, 32'shecd8e0e0, 32'shecd5e182, 32'shecd2e230, 32'sheccfe2ea, 32'sheccce3b0, 32'shecc9e481, 32'shecc6e55f, 
               32'shecc3e648, 32'shecc0e73d, 32'shecbde83e, 32'shecbae94b, 32'shecb7ea63, 32'shecb4eb88, 32'shecb1ecb8, 32'shecaeedf5, 
               32'shecabef3d, 32'sheca8f091, 32'sheca5f1f2, 32'sheca2f35e, 32'shec9ff4d6, 32'shec9cf65a, 32'shec99f7ea, 32'shec96f986, 
               32'shec93fb2e, 32'shec90fce1, 32'shec8dfea1, 32'shec8b006d, 32'shec880245, 32'shec850429, 32'shec820619, 32'shec7f0815, 
               32'shec7c0a1d, 32'shec790c31, 32'shec760e51, 32'shec73107d, 32'shec7012b5, 32'shec6d14f9, 32'shec6a1749, 32'shec6719a6, 
               32'shec641c0e, 32'shec611e83, 32'shec5e2103, 32'shec5b2390, 32'shec582629, 32'shec5528ce, 32'shec522b7f, 32'shec4f2e3d, 
               32'shec4c3106, 32'shec4933dc, 32'shec4636bd, 32'shec4339ab, 32'shec403ca5, 32'shec3d3fac, 32'shec3a42be, 32'shec3745dd, 
               32'shec344908, 32'shec314c3f, 32'shec2e4f82, 32'shec2b52d1, 32'shec28562d, 32'shec255995, 32'shec225d09, 32'shec1f608a, 
               32'shec1c6417, 32'shec1967b0, 32'shec166b55, 32'shec136f06, 32'shec1072c4, 32'shec0d768e, 32'shec0a7a65, 32'shec077e48, 
               32'shec048237, 32'shec018632, 32'shebfe8a3a, 32'shebfb8e4e, 32'shebf8926f, 32'shebf5969b, 32'shebf29ad4, 32'shebef9f1a, 
               32'shebeca36c, 32'shebe9a7ca, 32'shebe6ac35, 32'shebe3b0ac, 32'shebe0b52f, 32'shebddb9bf, 32'shebdabe5c, 32'shebd7c304, 
               32'shebd4c7ba, 32'shebd1cc7b, 32'shebced149, 32'shebcbd624, 32'shebc8db0b, 32'shebc5dffe, 32'shebc2e4fe, 32'shebbfea0b, 
               32'shebbcef23, 32'shebb9f449, 32'shebb6f97b, 32'shebb3feb9, 32'shebb10404, 32'shebae095c, 32'shebab0ec0, 32'sheba81430, 
               32'sheba519ad, 32'sheba21f37, 32'sheb9f24cd, 32'sheb9c2a70, 32'sheb99301f, 32'sheb9635db, 32'sheb933ba4, 32'sheb904179, 
               32'sheb8d475b, 32'sheb8a4d49, 32'sheb875344, 32'sheb84594c, 32'sheb815f60, 32'sheb7e6581, 32'sheb7b6bae, 32'sheb7871e8, 
               32'sheb75782f, 32'sheb727e83, 32'sheb6f84e3, 32'sheb6c8b50, 32'sheb6991ca, 32'sheb669850, 32'sheb639ee3, 32'sheb60a582, 
               32'sheb5dac2f, 32'sheb5ab2e8, 32'sheb57b9ae, 32'sheb54c081, 32'sheb51c760, 32'sheb4ece4c, 32'sheb4bd545, 32'sheb48dc4b, 
               32'sheb45e35d, 32'sheb42ea7c, 32'sheb3ff1a8, 32'sheb3cf8e1, 32'sheb3a0027, 32'sheb370779, 32'sheb340ed9, 32'sheb311645, 
               32'sheb2e1dbe, 32'sheb2b2543, 32'sheb282cd6, 32'sheb253475, 32'sheb223c22, 32'sheb1f43db, 32'sheb1c4ba1, 32'sheb195374, 
               32'sheb165b54, 32'sheb136341, 32'sheb106b3a, 32'sheb0d7341, 32'sheb0a7b54, 32'sheb078375, 32'sheb048ba2, 32'sheb0193dd, 
               32'sheafe9c24, 32'sheafba478, 32'sheaf8acd9, 32'sheaf5b547, 32'sheaf2bdc3, 32'sheaefc64b, 32'sheaeccee0, 32'sheae9d782, 
               32'sheae6e031, 32'sheae3e8ed, 32'sheae0f1b6, 32'sheaddfa8d, 32'sheadb0370, 32'shead80c60, 32'shead5155d, 32'shead21e68, 
               32'sheacf277f, 32'sheacc30a4, 32'sheac939d5, 32'sheac64314, 32'sheac34c60, 32'sheac055b9, 32'sheabd5f1f, 32'sheaba6892, 
               32'sheab77212, 32'sheab47b9f, 32'sheab1853a, 32'sheaae8ee2, 32'sheaab9896, 32'sheaa8a258, 32'sheaa5ac27, 32'sheaa2b604, 
               32'shea9fbfed, 32'shea9cc9e4, 32'shea99d3e8, 32'shea96ddf9, 32'shea93e817, 32'shea90f242, 32'shea8dfc7b, 32'shea8b06c1, 
               32'shea881114, 32'shea851b74, 32'shea8225e2, 32'shea7f305d, 32'shea7c3ae5, 32'shea79457a, 32'shea76501d, 32'shea735acd, 
               32'shea70658a, 32'shea6d7055, 32'shea6a7b2d, 32'shea678612, 32'shea649105, 32'shea619c04, 32'shea5ea712, 32'shea5bb22c, 
               32'shea58bd54, 32'shea55c889, 32'shea52d3cc, 32'shea4fdf1c, 32'shea4cea79, 32'shea49f5e4, 32'shea47015c, 32'shea440ce1, 
               32'shea411874, 32'shea3e2415, 32'shea3b2fc2, 32'shea383b7e, 32'shea354746, 32'shea32531c, 32'shea2f5f00, 32'shea2c6af1, 
               32'shea2976ef, 32'shea2682fb, 32'shea238f15, 32'shea209b3b, 32'shea1da770, 32'shea1ab3b2, 32'shea17c001, 32'shea14cc5e, 
               32'shea11d8c8, 32'shea0ee540, 32'shea0bf1c6, 32'shea08fe59, 32'shea060af9, 32'shea0317a7, 32'shea002463, 32'she9fd312c, 
               32'she9fa3e03, 32'she9f74ae8, 32'she9f457da, 32'she9f164d9, 32'she9ee71e6, 32'she9eb7f01, 32'she9e88c2a, 32'she9e59960, 
               32'she9e2a6a3, 32'she9dfb3f5, 32'she9dcc154, 32'she9d9cec0, 32'she9d6dc3b, 32'she9d3e9c3, 32'she9d0f758, 32'she9ce04fc, 
               32'she9cb12ad, 32'she9c8206b, 32'she9c52e38, 32'she9c23c12, 32'she9bf49fa, 32'she9bc57f0, 32'she9b965f3, 32'she9b67404, 
               32'she9b38223, 32'she9b0904f, 32'she9ad9e8a, 32'she9aaacd2, 32'she9a7bb28, 32'she9a4c98b, 32'she9a1d7fd, 32'she99ee67c, 
               32'she99bf509, 32'she99903a4, 32'she996124d, 32'she9932103, 32'she9902fc7, 32'she98d3e9a, 32'she98a4d7a, 32'she9875c68, 
               32'she9846b63, 32'she9817a6d, 32'she97e8984, 32'she97b98aa, 32'she978a7dd, 32'she975b71e, 32'she972c66d, 32'she96fd5ca, 
               32'she96ce535, 32'she969f4ae, 32'she9670435, 32'she96413c9, 32'she961236c, 32'she95e331d, 32'she95b42db, 32'she95852a8, 
               32'she9556282, 32'she952726b, 32'she94f8261, 32'she94c9266, 32'she949a278, 32'she946b299, 32'she943c2c7, 32'she940d304, 
               32'she93de34e, 32'she93af3a7, 32'she938040d, 32'she9351482, 32'she9322505, 32'she92f3596, 32'she92c4634, 32'she92956e1, 
               32'she926679c, 32'she9237866, 32'she920893d, 32'she91d9a22, 32'she91aab16, 32'she917bc17, 32'she914cd27, 32'she911de45, 
               32'she90eef71, 32'she90c00ab, 32'she90911f3, 32'she906234a, 32'she90334af, 32'she9004621, 32'she8fd57a2, 32'she8fa6932, 
               32'she8f77acf, 32'she8f48c7b, 32'she8f19e34, 32'she8eeaffd, 32'she8ebc1d3, 32'she8e8d3b7, 32'she8e5e5aa, 32'she8e2f7ab, 
               32'she8e009ba, 32'she8dd1bd8, 32'she8da2e04, 32'she8d7403e, 32'she8d45286, 32'she8d164dd, 32'she8ce7742, 32'she8cb89b5, 
               32'she8c89c37, 32'she8c5aec7, 32'she8c2c165, 32'she8bfd412, 32'she8bce6cd, 32'she8b9f996, 32'she8b70c6d, 32'she8b41f53, 
               32'she8b13248, 32'she8ae454b, 32'she8ab585c, 32'she8a86b7b, 32'she8a57ea9, 32'she8a291e5, 32'she89fa530, 32'she89cb889, 
               32'she899cbf1, 32'she896df67, 32'she893f2eb, 32'she891067e, 32'she88e1a20, 32'she88b2dcf, 32'she888418e, 32'she885555a, 
               32'she8826936, 32'she87f7d1f, 32'she87c9118, 32'she879a51e, 32'she876b934, 32'she873cd57, 32'she870e18a, 32'she86df5cb, 
               32'she86b0a1a, 32'she8681e78, 32'she86532e4, 32'she862475f, 32'she85f5be9, 32'she85c7081, 32'she8598528, 32'she85699dd, 
               32'she853aea1, 32'she850c374, 32'she84dd855, 32'she84aed45, 32'she8480243, 32'she8451750, 32'she8422c6c, 32'she83f4196, 
               32'she83c56cf, 32'she8396c16, 32'she836816d, 32'she83396d2, 32'she830ac45, 32'she82dc1c8, 32'she82ad759, 32'she827ecf8, 
               32'she82502a7, 32'she8221864, 32'she81f2e30, 32'she81c440a, 32'she81959f4, 32'she8166fec, 32'she81385f3, 32'she8109c08, 
               32'she80db22d, 32'she80ac860, 32'she807dea2, 32'she804f4f2, 32'she8020b52, 32'she7ff21c0, 32'she7fc383d, 32'she7f94ec9, 
               32'she7f66564, 32'she7f37c0d, 32'she7f092c6, 32'she7eda98d, 32'she7eac063, 32'she7e7d748, 32'she7e4ee3c, 32'she7e2053e, 
               32'she7df1c50, 32'she7dc3370, 32'she7d94a9f, 32'she7d661de, 32'she7d3792b, 32'she7d09087, 32'she7cda7f2, 32'she7cabf6c, 
               32'she7c7d6f4, 32'she7c4ee8c, 32'she7c20633, 32'she7bf1de8, 32'she7bc35ad, 32'she7b94d80, 32'she7b66563, 32'she7b37d55, 
               32'she7b09555, 32'she7adad65, 32'she7aac583, 32'she7a7ddb1, 32'she7a4f5ed, 32'she7a20e39, 32'she79f2693, 32'she79c3efd, 
               32'she7995776, 32'she7966ffd, 32'she7938894, 32'she790a13a, 32'she78db9ef, 32'she78ad2b3, 32'she787eb86, 32'she7850468, 
               32'she7821d59, 32'she77f365a, 32'she77c4f69, 32'she7796888, 32'she77681b6, 32'she7739af2, 32'she770b43e, 32'she76dcd9a, 
               32'she76ae704, 32'she768007e, 32'she7651a06, 32'she762339e, 32'she75f4d45, 32'she75c66fb, 32'she75980c1, 32'she7569a95, 
               32'she753b479, 32'she750ce6c, 32'she74de86f, 32'she74b0280, 32'she7481ca1, 32'she74536d1, 32'she7425110, 32'she73f6b5f, 
               32'she73c85bc, 32'she739a029, 32'she736baa6, 32'she733d531, 32'she730efcc, 32'she72e0a77, 32'she72b2530, 32'she7283ff9, 
               32'she7255ad1, 32'she72275b9, 32'she71f90b0, 32'she71cabb6, 32'she719c6cb, 32'she716e1f0, 32'she713fd25, 32'she7111868, 
               32'she70e33bb, 32'she70b4f1e, 32'she7086a8f, 32'she7058611, 32'she702a1a1, 32'she6ffbd41, 32'she6fcd8f1, 32'she6f9f4b0, 
               32'she6f7107e, 32'she6f42c5c, 32'she6f14849, 32'she6ee6446, 32'she6eb8052, 32'she6e89c6d, 32'she6e5b899, 32'she6e2d4d3, 
               32'she6dff11d, 32'she6dd0d77, 32'she6da29e0, 32'she6d74658, 32'she6d462e1, 32'she6d17f78, 32'she6ce9c1f, 32'she6cbb8d6, 
               32'she6c8d59c, 32'she6c5f272, 32'she6c30f57, 32'she6c02c4c, 32'she6bd4951, 32'she6ba6665, 32'she6b78389, 32'she6b4a0bc, 
               32'she6b1bdff, 32'she6aedb51, 32'she6abf8b3, 32'she6a91625, 32'she6a633a6, 32'she6a35137, 32'she6a06ed8, 32'she69d8c88, 
               32'she69aaa48, 32'she697c818, 32'she694e5f7, 32'she69203e6, 32'she68f21e5, 32'she68c3ff3, 32'she6895e11, 32'she6867c3f, 
               32'she6839a7c, 32'she680b8ca, 32'she67dd727, 32'she67af593, 32'she6781410, 32'she675329c, 32'she6725138, 32'she66f6fe3, 
               32'she66c8e9f, 32'she669ad6a, 32'she666cc45, 32'she663eb30, 32'she6610a2a, 32'she65e2935, 32'she65b484f, 32'she6586779, 
               32'she65586b3, 32'she652a5fc, 32'she64fc556, 32'she64ce4bf, 32'she64a0438, 32'she64723c2, 32'she644435a, 32'she6416303, 
               32'she63e82bc, 32'she63ba285, 32'she638c25d, 32'she635e245, 32'she633023e, 32'she6302246, 32'she62d425e, 32'she62a6286, 
               32'she62782be, 32'she624a306, 32'she621c35e, 32'she61ee3c6, 32'she61c043d, 32'she61924c5, 32'she616455d, 32'she6136605, 
               32'she61086bc, 32'she60da784, 32'she60ac85c, 32'she607e944, 32'she6050a3b, 32'she6022b43, 32'she5ff4c5b, 32'she5fc6d83, 
               32'she5f98ebb, 32'she5f6b003, 32'she5f3d15b, 32'she5f0f2c3, 32'she5ee143b, 32'she5eb35c3, 32'she5e8575b, 32'she5e57904, 
               32'she5e29abc, 32'she5dfbc85, 32'she5dcde5e, 32'she5da0047, 32'she5d72240, 32'she5d44449, 32'she5d16662, 32'she5ce888b, 
               32'she5cbaac5, 32'she5c8cd0f, 32'she5c5ef69, 32'she5c311d3, 32'she5c0344d, 32'she5bd56d7, 32'she5ba7972, 32'she5b79c1d, 
               32'she5b4bed8, 32'she5b1e1a3, 32'she5af047f, 32'she5ac276b, 32'she5a94a67, 32'she5a66d73, 32'she5a39090, 32'she5a0b3bc, 
               32'she59dd6f9, 32'she59afa47, 32'she5981da4, 32'she5954112, 32'she5926490, 32'she58f881f, 32'she58cabbe, 32'she589cf6d, 
               32'she586f32c, 32'she58416fc, 32'she5813adc, 32'she57e5ecc, 32'she57b82cd, 32'she578a6de, 32'she575cb00, 32'she572ef32, 
               32'she5701374, 32'she56d37c7, 32'she56a5c2a, 32'she567809d, 32'she564a521, 32'she561c9b5, 32'she55eee5a, 32'she55c130f, 
               32'she55937d5, 32'she5565cab, 32'she5538191, 32'she550a688, 32'she54dcb8f, 32'she54af0a7, 32'she54815cf, 32'she5453b08, 
               32'she5426051, 32'she53f85ab, 32'she53cab15, 32'she539d090, 32'she536f61b, 32'she5341bb7, 32'she5314163, 32'she52e6720, 
               32'she52b8cee, 32'she528b2cc, 32'she525d8ba, 32'she522feb9, 32'she52024c9, 32'she51d4ae9, 32'she51a711a, 32'she517975b, 
               32'she514bdad, 32'she511e410, 32'she50f0a83, 32'she50c3107, 32'she509579b, 32'she5067e40, 32'she503a4f6, 32'she500cbbc, 
               32'she4fdf294, 32'she4fb197b, 32'she4f84074, 32'she4f5677d, 32'she4f28e96, 32'she4efb5c1, 32'she4ecdcfc, 32'she4ea0448, 
               32'she4e72ba4, 32'she4e45311, 32'she4e17a8f, 32'she4dea21e, 32'she4dbc9bd, 32'she4d8f16d, 32'she4d6192e, 32'she4d34100, 
               32'she4d068e2, 32'she4cd90d5, 32'she4cab8d9, 32'she4c7e0ee, 32'she4c50914, 32'she4c2314a, 32'she4bf5991, 32'she4bc81e9, 
               32'she4b9aa52, 32'she4b6d2cb, 32'she4b3fb56, 32'she4b123f1, 32'she4ae4c9d, 32'she4ab755a, 32'she4a89e28, 32'she4a5c707, 
               32'she4a2eff6, 32'she4a018f7, 32'she49d4208, 32'she49a6b2a, 32'she497945d, 32'she494bda1, 32'she491e6f6, 32'she48f105c, 
               32'she48c39d3, 32'she489635a, 32'she4868cf3, 32'she483b69d, 32'she480e057, 32'she47e0a23, 32'she47b33ff, 32'she4785ded, 
               32'she47587eb, 32'she472b1fa, 32'she46fdc1b, 32'she46d064c, 32'she46a308f, 32'she4675ae2, 32'she4648547, 32'she461afbc, 
               32'she45eda43, 32'she45c04da, 32'she4592f83, 32'she4565a3c, 32'she4538507, 32'she450afe3, 32'she44ddad0, 32'she44b05ce, 
               32'she44830dd, 32'she4455bfd, 32'she442872e, 32'she43fb271, 32'she43cddc4, 32'she43a0929, 32'she437349f, 32'she4346026, 
               32'she4318bbe, 32'she42eb767, 32'she42be321, 32'she4290eed, 32'she4263ac9, 32'she42366b7, 32'she42092b6, 32'she41dbec7, 
               32'she41aeae8, 32'she418171b, 32'she415435f, 32'she4126fb4, 32'she40f9c1a, 32'she40cc891, 32'she409f51a, 32'she40721b4, 
               32'she4044e60, 32'she4017b1c, 32'she3fea7ea, 32'she3fbd4c9, 32'she3f901ba, 32'she3f62ebb, 32'she3f35bce, 32'she3f088f2, 
               32'she3edb628, 32'she3eae36f, 32'she3e810c7, 32'she3e53e31, 32'she3e26bac, 32'she3df9938, 32'she3dcc6d5, 32'she3d9f484, 
               32'she3d72245, 32'she3d45016, 32'she3d17df9, 32'she3ceabee, 32'she3cbd9f4, 32'she3c9080b, 32'she3c63633, 32'she3c3646d, 
               32'she3c092b9, 32'she3bdc116, 32'she3baef84, 32'she3b81e04, 32'she3b54c95, 32'she3b27b38, 32'she3afa9ec, 32'she3acd8b1, 
               32'she3aa0788, 32'she3a73671, 32'she3a4656b, 32'she3a19476, 32'she39ec393, 32'she39bf2c2, 32'she3992202, 32'she3965153, 
               32'she39380b6, 32'she390b02b, 32'she38ddfb1, 32'she38b0f49, 32'she3883ef2, 32'she3856ead, 32'she3829e79, 32'she37fce57, 
               32'she37cfe47, 32'she37a2e48, 32'she3775e5a, 32'she3748e7f, 32'she371beb5, 32'she36eeefc, 32'she36c1f55, 32'she3694fc0, 
               32'she366803c, 32'she363b0cb, 32'she360e16a, 32'she35e121c, 32'she35b42df, 32'she35873b3, 32'she355a49a, 32'she352d592, 
               32'she350069b, 32'she34d37b7, 32'she34a68e4, 32'she3479a23, 32'she344cb73, 32'she341fcd6, 32'she33f2e4a, 32'she33c5fcf, 
               32'she3399167, 32'she336c310, 32'she333f4cb, 32'she3312698, 32'she32e5876, 32'she32b8a67, 32'she328bc69, 32'she325ee7d, 
               32'she32320a2, 32'she32052da, 32'she31d8523, 32'she31ab77e, 32'she317e9eb, 32'she3151c6a, 32'she3124efa, 32'she30f819d, 
               32'she30cb451, 32'she309e717, 32'she30719ef, 32'she3044cd9, 32'she3017fd5, 32'she2feb2e3, 32'she2fbe602, 32'she2f91934, 
               32'she2f64c77, 32'she2f37fcc, 32'she2f0b333, 32'she2ede6ac, 32'she2eb1a37, 32'she2e84dd4, 32'she2e58183, 32'she2e2b544, 
               32'she2dfe917, 32'she2dd1cfc, 32'she2da50f3, 32'she2d784fb, 32'she2d4b916, 32'she2d1ed43, 32'she2cf2182, 32'she2cc55d2, 
               32'she2c98a35, 32'she2c6beaa, 32'she2c3f331, 32'she2c127c9, 32'she2be5c74, 32'she2bb9131, 32'she2b8c600, 32'she2b5fae1, 
               32'she2b32fd4, 32'she2b064da, 32'she2ad99f1, 32'she2aacf1a, 32'she2a80456, 32'she2a539a3, 32'she2a26f03, 32'she29fa474, 
               32'she29cd9f8, 32'she29a0f8e, 32'she2974536, 32'she2947af1, 32'she291b0bd, 32'she28ee69c, 32'she28c1c8c, 32'she289528f, 
               32'she28688a4, 32'she283becc, 32'she280f505, 32'she27e2b51, 32'she27b61af, 32'she278981f, 32'she275cea1, 32'she2730536, 
               32'she2703bdc, 32'she26d7295, 32'she26aa960, 32'she267e03e, 32'she265172e, 32'she2624e2f, 32'she25f8544, 32'she25cbc6a, 
               32'she259f3a3, 32'she2572aee, 32'she254624b, 32'she25199bb, 32'she24ed13d, 32'she24c08d1, 32'she2494078, 32'she2467831, 
               32'she243affc, 32'she240e7da, 32'she23e1fca, 32'she23b57cc, 32'she2388fe1, 32'she235c808, 32'she2330041, 32'she230388d, 
               32'she22d70eb, 32'she22aa95c, 32'she227e1df, 32'she2251a75, 32'she222531c, 32'she21f8bd7, 32'she21cc4a3, 32'she219fd82, 
               32'she2173674, 32'she2146f78, 32'she211a88f, 32'she20ee1b7, 32'she20c1af3, 32'she2095441, 32'she2068da1, 32'she203c714, 
               32'she2010099, 32'she1fe3a31, 32'she1fb73dc, 32'she1f8ad98, 32'she1f5e768, 32'she1f3214a, 32'she1f05b3e, 32'she1ed9545, 
               32'she1eacf5f, 32'she1e8098b, 32'she1e543ca, 32'she1e27e1b, 32'she1dfb87f, 32'she1dcf2f5, 32'she1da2d7e, 32'she1d7681a, 
               32'she1d4a2c8, 32'she1d1dd89, 32'she1cf185c, 32'she1cc5342, 32'she1c98e3b, 32'she1c6c946, 32'she1c40464, 32'she1c13f95, 
               32'she1be7ad8, 32'she1bbb62e, 32'she1b8f197, 32'she1b62d12, 32'she1b368a0, 32'she1b0a441, 32'she1addff4, 32'she1ab1bba, 
               32'she1a85793, 32'she1a5937e, 32'she1a2cf7c, 32'she1a00b8d, 32'she19d47b1, 32'she19a83e7, 32'she197c031, 32'she194fc8d, 
               32'she19238fb, 32'she18f757d, 32'she18cb211, 32'she189eeb8, 32'she1872b72, 32'she184683e, 32'she181a51e, 32'she17ee210, 
               32'she17c1f15, 32'she1795c2d, 32'she1769958, 32'she173d695, 32'she17113e5, 32'she16e5149, 32'she16b8ebf, 32'she168cc48, 
               32'she16609e3, 32'she1634792, 32'she1608554, 32'she15dc328, 32'she15b0110, 32'she1583f0a, 32'she1557d17, 32'she152bb37, 
               32'she14ff96a, 32'she14d37b0, 32'she14a7609, 32'she147b475, 32'she144f2f3, 32'she1423185, 32'she13f702a, 32'she13caee1, 
               32'she139edac, 32'she1372c8a, 32'she1346b7a, 32'she131aa7e, 32'she12ee995, 32'she12c28be, 32'she12967fb, 32'she126a74a, 
               32'she123e6ad, 32'she1212623, 32'she11e65ac, 32'she11ba547, 32'she118e4f6, 32'she11624b8, 32'she113648d, 32'she110a475, 
               32'she10de470, 32'she10b247f, 32'she10864a0, 32'she105a4d4, 32'she102e51c, 32'she1002577, 32'she0fd65e4, 32'she0faa665, 
               32'she0f7e6f9, 32'she0f527a0, 32'she0f2685b, 32'she0efa928, 32'she0ecea09, 32'she0ea2afd, 32'she0e76c04, 32'she0e4ad1e, 
               32'she0e1ee4b, 32'she0df2f8c, 32'she0dc70e0, 32'she0d9b247, 32'she0d6f3c1, 32'she0d4354e, 32'she0d176ef, 32'she0ceb8a3, 
               32'she0cbfa6a, 32'she0c93c44, 32'she0c67e32, 32'she0c3c033, 32'she0c10247, 32'she0be446e, 32'she0bb86a9, 32'she0b8c8f7, 
               32'she0b60b58, 32'she0b34dcd, 32'she0b09055, 32'she0add2f0, 32'she0ab159e, 32'she0a85860, 32'she0a59b35, 32'she0a2de1e, 
               32'she0a0211a, 32'she09d6429, 32'she09aa74b, 32'she097ea81, 32'she0952dcb, 32'she0927127, 32'she08fb497, 32'she08cf81b, 
               32'she08a3bb2, 32'she0877f5c, 32'she084c31a, 32'she08206eb, 32'she07f4acf, 32'she07c8ec7, 32'she079d2d3, 32'she07716f2, 
               32'she0745b24, 32'she0719f6a, 32'she06ee3c3, 32'she06c2830, 32'she0696cb0, 32'she066b144, 32'she063f5eb, 32'she0613aa5, 
               32'she05e7f74, 32'she05bc455, 32'she059094a, 32'she0564e53, 32'she053936f, 32'she050d89f, 32'she04e1de3, 32'she04b6339, 
               32'she048a8a4, 32'she045ee22, 32'she04333b3, 32'she0407959, 32'she03dbf11, 32'she03b04de, 32'she0384abe, 32'she03590b1, 
               32'she032d6b8, 32'she0301cd3, 32'she02d6301, 32'she02aa943, 32'she027ef99, 32'she0253602, 32'she0227c7f, 32'she01fc310, 
               32'she01d09b4, 32'she01a506c, 32'she0179738, 32'she014de17, 32'she012250a, 32'she00f6c11, 32'she00cb32b, 32'she009fa59, 
               32'she007419b, 32'she00488f0, 32'she001d05a, 32'shdfff17d7, 32'shdffc5f67, 32'shdff9a70c, 32'shdff6eec4, 32'shdff43690, 
               32'shdff17e70, 32'shdfeec663, 32'shdfec0e6a, 32'shdfe95686, 32'shdfe69eb4, 32'shdfe3e6f7, 32'shdfe12f4e, 32'shdfde77b8, 
               32'shdfdbc036, 32'shdfd908c8, 32'shdfd6516e, 32'shdfd39a27, 32'shdfd0e2f5, 32'shdfce2bd6, 32'shdfcb74cb, 32'shdfc8bdd4, 
               32'shdfc606f1, 32'shdfc35022, 32'shdfc09967, 32'shdfbde2bf, 32'shdfbb2c2c, 32'shdfb875ac, 32'shdfb5bf41, 32'shdfb308e9, 
               32'shdfb052a5, 32'shdfad9c75, 32'shdfaae659, 32'shdfa83051, 32'shdfa57a5d, 32'shdfa2c47d, 32'shdfa00eb1, 32'shdf9d58f8, 
               32'shdf9aa354, 32'shdf97edc4, 32'shdf953848, 32'shdf9282df, 32'shdf8fcd8b, 32'shdf8d184b, 32'shdf8a631f, 32'shdf87ae06, 
               32'shdf84f902, 32'shdf824412, 32'shdf7f8f36, 32'shdf7cda6e, 32'shdf7a25ba, 32'shdf77711a, 32'shdf74bc8e, 32'shdf720816, 
               32'shdf6f53b3, 32'shdf6c9f63, 32'shdf69eb27, 32'shdf673700, 32'shdf6482ed, 32'shdf61ceee, 32'shdf5f1b02, 32'shdf5c672b, 
               32'shdf59b369, 32'shdf56ffba, 32'shdf544c1f, 32'shdf519899, 32'shdf4ee527, 32'shdf4c31c9, 32'shdf497e7f, 32'shdf46cb49, 
               32'shdf441828, 32'shdf41651a, 32'shdf3eb221, 32'shdf3bff3c, 32'shdf394c6b, 32'shdf3699af, 32'shdf33e707, 32'shdf313473, 
               32'shdf2e81f3, 32'shdf2bcf87, 32'shdf291d30, 32'shdf266aed, 32'shdf23b8be, 32'shdf2106a4, 32'shdf1e549d, 32'shdf1ba2ab, 
               32'shdf18f0ce, 32'shdf163f04, 32'shdf138d4f, 32'shdf10dbaf, 32'shdf0e2a22, 32'shdf0b78aa, 32'shdf08c746, 32'shdf0615f7, 
               32'shdf0364bc, 32'shdf00b395, 32'shdefe0282, 32'shdefb5184, 32'shdef8a09b, 32'shdef5efc5, 32'shdef33f04, 32'shdef08e58, 
               32'shdeedddc0, 32'shdeeb2d3c, 32'shdee87ccc, 32'shdee5cc72, 32'shdee31c2b, 32'shdee06bf9, 32'shdeddbbdb, 32'shdedb0bd2, 
               32'shded85bdd, 32'shded5abfd, 32'shded2fc31, 32'shded04c7a, 32'shdecd9cd7, 32'shdecaed48, 32'shdec83dce, 32'shdec58e69, 
               32'shdec2df18, 32'shdec02fdb, 32'shdebd80b3, 32'shdebad1a0, 32'shdeb822a1, 32'shdeb573b7, 32'shdeb2c4e1, 32'shdeb0161f, 
               32'shdead6773, 32'shdeaab8da, 32'shdea80a57, 32'shdea55be8, 32'shdea2ad8d, 32'shde9fff47, 32'shde9d5116, 32'shde9aa2f9, 
               32'shde97f4f1, 32'shde9546fd, 32'shde92991e, 32'shde8feb54, 32'shde8d3d9e, 32'shde8a8ffd, 32'shde87e271, 32'shde8534f9, 
               32'shde828796, 32'shde7fda48, 32'shde7d2d0e, 32'shde7a7fe9, 32'shde77d2d8, 32'shde7525dc, 32'shde7278f5, 32'shde6fcc23, 
               32'shde6d1f65, 32'shde6a72bc, 32'shde67c628, 32'shde6519a9, 32'shde626d3e, 32'shde5fc0e8, 32'shde5d14a6, 32'shde5a687a, 
               32'shde57bc62, 32'shde55105f, 32'shde526471, 32'shde4fb897, 32'shde4d0cd2, 32'shde4a6122, 32'shde47b587, 32'shde450a01, 
               32'shde425e8f, 32'shde3fb333, 32'shde3d07eb, 32'shde3a5cb8, 32'shde37b199, 32'shde350690, 32'shde325b9b, 32'shde2fb0bc, 
               32'shde2d05f1, 32'shde2a5b3b, 32'shde27b09a, 32'shde25060e, 32'shde225b96, 32'shde1fb134, 32'shde1d06e6, 32'shde1a5cad, 
               32'shde17b28a, 32'shde15087b, 32'shde125e81, 32'shde0fb49c, 32'shde0d0acc, 32'shde0a6111, 32'shde07b76b, 32'shde050dd9, 
               32'shde02645d, 32'shddffbaf6, 32'shddfd11a3, 32'shddfa6866, 32'shddf7bf3e, 32'shddf5162a, 32'shddf26d2c, 32'shddefc443, 
               32'shdded1b6e, 32'shddea72af, 32'shdde7ca05, 32'shdde5216f, 32'shdde278ef, 32'shdddfd084, 32'shdddd282e, 32'shddda7fed, 
               32'shddd7d7c1, 32'shddd52faa, 32'shddd287a8, 32'shddcfdfbb, 32'shddcd37e4, 32'shddca9021, 32'shddc7e873, 32'shddc540db, 
               32'shddc29958, 32'shddbff1ea, 32'shddbd4a91, 32'shddbaa34d, 32'shddb7fc1e, 32'shddb55504, 32'shddb2ae00, 32'shddb00711, 
               32'shddad6036, 32'shddaab972, 32'shdda812c2, 32'shdda56c27, 32'shdda2c5a2, 32'shdda01f32, 32'shdd9d78d7, 32'shdd9ad291, 
               32'shdd982c60, 32'shdd958645, 32'shdd92e03f, 32'shdd903a4e, 32'shdd8d9472, 32'shdd8aeeac, 32'shdd8848fb, 32'shdd85a35f, 
               32'shdd82fdd8, 32'shdd805867, 32'shdd7db30b, 32'shdd7b0dc4, 32'shdd786892, 32'shdd75c376, 32'shdd731e6f, 32'shdd70797e, 
               32'shdd6dd4a2, 32'shdd6b2fdb, 32'shdd688b29, 32'shdd65e68d, 32'shdd634206, 32'shdd609d94, 32'shdd5df938, 32'shdd5b54f1, 
               32'shdd58b0c0, 32'shdd560ca4, 32'shdd53689d, 32'shdd50c4ac, 32'shdd4e20d0, 32'shdd4b7d09, 32'shdd48d958, 32'shdd4635bd, 
               32'shdd439236, 32'shdd40eec5, 32'shdd3e4b6a, 32'shdd3ba824, 32'shdd3904f4, 32'shdd3661d8, 32'shdd33bed3, 32'shdd311be3, 
               32'shdd2e7908, 32'shdd2bd643, 32'shdd293393, 32'shdd2690f9, 32'shdd23ee74, 32'shdd214c05, 32'shdd1ea9ab, 32'shdd1c0767, 
               32'shdd196538, 32'shdd16c31f, 32'shdd14211b, 32'shdd117f2d, 32'shdd0edd55, 32'shdd0c3b92, 32'shdd0999e4, 32'shdd06f84d, 
               32'shdd0456ca, 32'shdd01b55e, 32'shdcff1407, 32'shdcfc72c5, 32'shdcf9d199, 32'shdcf73083, 32'shdcf48f82, 32'shdcf1ee97, 
               32'shdcef4dc2, 32'shdcecad02, 32'shdcea0c58, 32'shdce76bc3, 32'shdce4cb44, 32'shdce22adb, 32'shdcdf8a87, 32'shdcdcea49, 
               32'shdcda4a21, 32'shdcd7aa0e, 32'shdcd50a12, 32'shdcd26a2a, 32'shdccfca59, 32'shdccd2a9d, 32'shdcca8af7, 32'shdcc7eb67, 
               32'shdcc54bec, 32'shdcc2ac87, 32'shdcc00d38, 32'shdcbd6dff, 32'shdcbacedb, 32'shdcb82fcd, 32'shdcb590d5, 32'shdcb2f1f3, 
               32'shdcb05326, 32'shdcadb46f, 32'shdcab15ce, 32'shdca87743, 32'shdca5d8cd, 32'shdca33a6e, 32'shdca09c24, 32'shdc9dfdf0, 
               32'shdc9b5fd2, 32'shdc98c1ca, 32'shdc9623d7, 32'shdc9385fa, 32'shdc90e834, 32'shdc8e4a83, 32'shdc8bace8, 32'shdc890f62, 
               32'shdc8671f3, 32'shdc83d49a, 32'shdc813756, 32'shdc7e9a28, 32'shdc7bfd11, 32'shdc79600f, 32'shdc76c323, 32'shdc74264d, 
               32'shdc71898d, 32'shdc6eece2, 32'shdc6c504e, 32'shdc69b3d0, 32'shdc671768, 32'shdc647b15, 32'shdc61ded9, 32'shdc5f42b2, 
               32'shdc5ca6a2, 32'shdc5a0aa8, 32'shdc576ec3, 32'shdc54d2f5, 32'shdc52373c, 32'shdc4f9b9a, 32'shdc4d000d, 32'shdc4a6497, 
               32'shdc47c936, 32'shdc452dec, 32'shdc4292b8, 32'shdc3ff799, 32'shdc3d5c91, 32'shdc3ac19f, 32'shdc3826c3, 32'shdc358bfd, 
               32'shdc32f14d, 32'shdc3056b3, 32'shdc2dbc2f, 32'shdc2b21c1, 32'shdc28876a, 32'shdc25ed28, 32'shdc2352fd, 32'shdc20b8e8, 
               32'shdc1e1ee9, 32'shdc1b8500, 32'shdc18eb2d, 32'shdc165170, 32'shdc13b7c9, 32'shdc111e39, 32'shdc0e84bf, 32'shdc0beb5b, 
               32'shdc09520d, 32'shdc06b8d5, 32'shdc041fb4, 32'shdc0186a8, 32'shdbfeedb3, 32'shdbfc54d4, 32'shdbf9bc0c, 32'shdbf72359, 
               32'shdbf48abd, 32'shdbf1f237, 32'shdbef59c7, 32'shdbecc16e, 32'shdbea292b, 32'shdbe790fe, 32'shdbe4f8e7, 32'shdbe260e6, 
               32'shdbdfc8fc, 32'shdbdd3128, 32'shdbda996b, 32'shdbd801c3, 32'shdbd56a32, 32'shdbd2d2b8, 32'shdbd03b53, 32'shdbcda405, 
               32'shdbcb0cce, 32'shdbc875ac, 32'shdbc5dea1, 32'shdbc347ac, 32'shdbc0b0ce, 32'shdbbe1a06, 32'shdbbb8354, 32'shdbb8ecb9, 
               32'shdbb65634, 32'shdbb3bfc6, 32'shdbb1296e, 32'shdbae932c, 32'shdbabfd01, 32'shdba966ec, 32'shdba6d0ed, 32'shdba43b05, 
               32'shdba1a534, 32'shdb9f0f78, 32'shdb9c79d4, 32'shdb99e445, 32'shdb974ece, 32'shdb94b96c, 32'shdb922421, 32'shdb8f8eed, 
               32'shdb8cf9cf, 32'shdb8a64c7, 32'shdb87cfd6, 32'shdb853afc, 32'shdb82a638, 32'shdb80118a, 32'shdb7d7cf3, 32'shdb7ae873, 
               32'shdb785409, 32'shdb75bfb5, 32'shdb732b79, 32'shdb709752, 32'shdb6e0342, 32'shdb6b6f49, 32'shdb68db67, 32'shdb66479b, 
               32'shdb63b3e5, 32'shdb612046, 32'shdb5e8cbe, 32'shdb5bf94c, 32'shdb5965f1, 32'shdb56d2ac, 32'shdb543f7e, 32'shdb51ac67, 
               32'shdb4f1967, 32'shdb4c867d, 32'shdb49f3a9, 32'shdb4760ec, 32'shdb44ce46, 32'shdb423bb7, 32'shdb3fa93e, 32'shdb3d16dc, 
               32'shdb3a8491, 32'shdb37f25c, 32'shdb35603e, 32'shdb32ce36, 32'shdb303c46, 32'shdb2daa6c, 32'shdb2b18a9, 32'shdb2886fc, 
               32'shdb25f566, 32'shdb2363e7, 32'shdb20d27f, 32'shdb1e412d, 32'shdb1baff2, 32'shdb191ece, 32'shdb168dc1, 32'shdb13fccb, 
               32'shdb116beb, 32'shdb0edb22, 32'shdb0c4a70, 32'shdb09b9d4, 32'shdb072950, 32'shdb0498e2, 32'shdb02088b, 32'shdaff784b, 
               32'shdafce821, 32'shdafa580f, 32'shdaf7c813, 32'shdaf5382e, 32'shdaf2a860, 32'shdaf018a9, 32'shdaed8909, 32'shdaeaf980, 
               32'shdae86a0d, 32'shdae5dab2, 32'shdae34b6d, 32'shdae0bc3f, 32'shdade2d28, 32'shdadb9e28, 32'shdad90f3f, 32'shdad6806d, 
               32'shdad3f1b1, 32'shdad1630d, 32'shdaced47f, 32'shdacc4609, 32'shdac9b7a9, 32'shdac72961, 32'shdac49b2f, 32'shdac20d15, 
               32'shdabf7f11, 32'shdabcf124, 32'shdaba634e, 32'shdab7d590, 32'shdab547e8, 32'shdab2ba57, 32'shdab02cdd, 32'shdaad9f7b, 
               32'shdaab122f, 32'shdaa884fa, 32'shdaa5f7dd, 32'shdaa36ad6, 32'shdaa0dde7, 32'shda9e510e, 32'shda9bc44d, 32'shda9937a2, 
               32'shda96ab0f, 32'shda941e93, 32'shda91922e, 32'shda8f05e0, 32'shda8c79a9, 32'shda89ed89, 32'shda876180, 32'shda84d58f, 
               32'shda8249b4, 32'shda7fbdf1, 32'shda7d3244, 32'shda7aa6af, 32'shda781b31, 32'shda758fcb, 32'shda73047b, 32'shda707942, 
               32'shda6dee21, 32'shda6b6317, 32'shda68d824, 32'shda664d48, 32'shda63c284, 32'shda6137d6, 32'shda5ead40, 32'shda5c22c1, 
               32'shda599859, 32'shda570e09, 32'shda5483d0, 32'shda51f9ae, 32'shda4f6fa3, 32'shda4ce5af, 32'shda4a5bd3, 32'shda47d20e, 
               32'shda454860, 32'shda42beca, 32'shda40354a, 32'shda3dabe2, 32'shda3b2292, 32'shda389958, 32'shda361036, 32'shda33872c, 
               32'shda30fe38, 32'shda2e755c, 32'shda2bec97, 32'shda2963ea, 32'shda26db54, 32'shda2452d5, 32'shda21ca6e, 32'shda1f421e, 
               32'shda1cb9e5, 32'shda1a31c4, 32'shda17a9ba, 32'shda1521c7, 32'shda1299ec, 32'shda101228, 32'shda0d8a7c, 32'shda0b02e7, 
               32'shda087b69, 32'shda05f403, 32'shda036cb5, 32'shda00e57d, 32'shd9fe5e5e, 32'shd9fbd755, 32'shd9f95064, 32'shd9f6c98b, 
               32'shd9f442c9, 32'shd9f1bc1e, 32'shd9ef358b, 32'shd9ecaf10, 32'shd9ea28ac, 32'shd9e7a25f, 32'shd9e51c2a, 32'shd9e2960c, 
               32'shd9e01006, 32'shd9dd8a18, 32'shd9db0441, 32'shd9d87e81, 32'shd9d5f8d9, 32'shd9d37349, 32'shd9d0edd0, 32'shd9ce686e, 
               32'shd9cbe325, 32'shd9c95df3, 32'shd9c6d8d8, 32'shd9c453d5, 32'shd9c1cee9, 32'shd9bf4a15, 32'shd9bcc559, 32'shd9ba40b5, 
               32'shd9b7bc27, 32'shd9b537b2, 32'shd9b2b354, 32'shd9b02f0e, 32'shd9adaadf, 32'shd9ab26c8, 32'shd9a8a2c9, 32'shd9a61ee1, 
               32'shd9a39b11, 32'shd9a11759, 32'shd99e93b8, 32'shd99c102f, 32'shd9998cbe, 32'shd9970965, 32'shd9948623, 32'shd99202f8, 
               32'shd98f7fe6, 32'shd98cfceb, 32'shd98a7a08, 32'shd987f73d, 32'shd9857489, 32'shd982f1ed, 32'shd9806f69, 32'shd97decfd, 
               32'shd97b6aa8, 32'shd978e86b, 32'shd9766646, 32'shd973e438, 32'shd9716243, 32'shd96ee065, 32'shd96c5e9f, 32'shd969dcf1, 
               32'shd9675b5a, 32'shd964d9dc, 32'shd9625875, 32'shd95fd726, 32'shd95d55ef, 32'shd95ad4d0, 32'shd95853c8, 32'shd955d2d9, 
               32'shd9535201, 32'shd950d141, 32'shd94e5099, 32'shd94bd009, 32'shd9494f90, 32'shd946cf30, 32'shd9444ee7, 32'shd941ceb7, 
               32'shd93f4e9e, 32'shd93cce9d, 32'shd93a4eb4, 32'shd937cee3, 32'shd9354f2a, 32'shd932cf89, 32'shd9305000, 32'shd92dd08e, 
               32'shd92b5135, 32'shd928d1f4, 32'shd92652ca, 32'shd923d3b9, 32'shd92154bf, 32'shd91ed5de, 32'shd91c5714, 32'shd919d863, 
               32'shd91759c9, 32'shd914db47, 32'shd9125cde, 32'shd90fde8c, 32'shd90d6053, 32'shd90ae231, 32'shd9086428, 32'shd905e636, 
               32'shd903685d, 32'shd900ea9c, 32'shd8fe6cf2, 32'shd8fbef61, 32'shd8f971e8, 32'shd8f6f487, 32'shd8f4773e, 32'shd8f1fa0d, 
               32'shd8ef7cf4, 32'shd8ecfff4, 32'shd8ea830b, 32'shd8e8063a, 32'shd8e58982, 32'shd8e30ce2, 32'shd8e0905a, 32'shd8de13ea, 
               32'shd8db9792, 32'shd8d91b52, 32'shd8d69f2a, 32'shd8d4231b, 32'shd8d1a724, 32'shd8cf2b45, 32'shd8ccaf7e, 32'shd8ca33cf, 
               32'shd8c7b838, 32'shd8c53cba, 32'shd8c2c154, 32'shd8c04606, 32'shd8bdcad0, 32'shd8bb4fb3, 32'shd8b8d4ad, 32'shd8b659c0, 
               32'shd8b3deeb, 32'shd8b1642f, 32'shd8aee98a, 32'shd8ac6efe, 32'shd8a9f48a, 32'shd8a77a2f, 32'shd8a4ffec, 32'shd8a285c0, 
               32'shd8a00bae, 32'shd89d91b3, 32'shd89b17d1, 32'shd8989e07, 32'shd8962456, 32'shd893aabc, 32'shd891313b, 32'shd88eb7d3, 
               32'shd88c3e83, 32'shd889c54b, 32'shd8874c2b, 32'shd884d324, 32'shd8825a35, 32'shd87fe15e, 32'shd87d68a0, 32'shd87aeffa, 
               32'shd878776d, 32'shd875fef8, 32'shd873869b, 32'shd8710e57, 32'shd86e962b, 32'shd86c1e18, 32'shd869a61d, 32'shd8672e3a, 
               32'shd864b670, 32'shd8623ebe, 32'shd85fc725, 32'shd85d4fa4, 32'shd85ad83c, 32'shd85860ec, 32'shd855e9b4, 32'shd8537295, 
               32'shd850fb8e, 32'shd84e84a0, 32'shd84c0dcb, 32'shd849970e, 32'shd8472069, 32'shd844a9dd, 32'shd8423369, 32'shd83fbd0e, 
               32'shd83d46cc, 32'shd83ad0a2, 32'shd8385a90, 32'shd835e497, 32'shd8336eb7, 32'shd830f8ef, 32'shd82e833f, 32'shd82c0da9, 
               32'shd829982b, 32'shd82722c5, 32'shd824ad78, 32'shd8223843, 32'shd81fc328, 32'shd81d4e24, 32'shd81ad93a, 32'shd8186468, 
               32'shd815efae, 32'shd8137b0d, 32'shd8110685, 32'shd80e9216, 32'shd80c1dbf, 32'shd809a980, 32'shd807355b, 32'shd804c14e, 
               32'shd8024d59, 32'shd7ffd97e, 32'shd7fd65bb, 32'shd7faf211, 32'shd7f87e7f, 32'shd7f60b06, 32'shd7f397a6, 32'shd7f1245e, 
               32'shd7eeb130, 32'shd7ec3e1a, 32'shd7e9cb1c, 32'shd7e75838, 32'shd7e4e56c, 32'shd7e272b8, 32'shd7e0001e, 32'shd7dd8d9c, 
               32'shd7db1b34, 32'shd7d8a8e3, 32'shd7d636ac, 32'shd7d3c48d, 32'shd7d15288, 32'shd7cee09b, 32'shd7cc6ec6, 32'shd7c9fd0b, 
               32'shd7c78b68, 32'shd7c519de, 32'shd7c2a86d, 32'shd7c03715, 32'shd7bdc5d6, 32'shd7bb54af, 32'shd7b8e3a2, 32'shd7b672ad, 
               32'shd7b401d1, 32'shd7b1910e, 32'shd7af2063, 32'shd7acafd2, 32'shd7aa3f5a, 32'shd7a7cefa, 32'shd7a55eb3, 32'shd7a2ee85, 
               32'shd7a07e70, 32'shd79e0e74, 32'shd79b9e91, 32'shd7992ec7, 32'shd796bf16, 32'shd7944f7d, 32'shd791dffe, 32'shd78f7097, 
               32'shd78d014a, 32'shd78a9215, 32'shd78822f9, 32'shd785b3f7, 32'shd783450d, 32'shd780d63c, 32'shd77e6784, 32'shd77bf8e6, 
               32'shd7798a60, 32'shd7771bf3, 32'shd774ad9f, 32'shd7723f64, 32'shd76fd143, 32'shd76d633a, 32'shd76af54a, 32'shd7688774, 
               32'shd76619b6, 32'shd763ac11, 32'shd7613e86, 32'shd75ed113, 32'shd75c63ba, 32'shd759f679, 32'shd7578952, 32'shd7551c44, 
               32'shd752af4f, 32'shd7504273, 32'shd74dd5b0, 32'shd74b6906, 32'shd748fc75, 32'shd7468ffe, 32'shd744239f, 32'shd741b75a, 
               32'shd73f4b2e, 32'shd73cdf1b, 32'shd73a7321, 32'shd7380740, 32'shd7359b78, 32'shd7332fca, 32'shd730c434, 32'shd72e58b8, 
               32'shd72bed55, 32'shd729820c, 32'shd72716db, 32'shd724abc4, 32'shd72240c5, 32'shd71fd5e0, 32'shd71d6b15, 32'shd71b0062, 
               32'shd71895c9, 32'shd7162b49, 32'shd713c0e2, 32'shd7115694, 32'shd70eec60, 32'shd70c8245, 32'shd70a1843, 32'shd707ae5a, 
               32'shd705448b, 32'shd702dad5, 32'shd7007138, 32'shd6fe07b5, 32'shd6fb9e4b, 32'shd6f934fa, 32'shd6f6cbc2, 32'shd6f462a4, 
               32'shd6f1f99f, 32'shd6ef90b4, 32'shd6ed27e1, 32'shd6eabf28, 32'shd6e85689, 32'shd6e5ee03, 32'shd6e38596, 32'shd6e11d42, 
               32'shd6deb508, 32'shd6dc4ce7, 32'shd6d9e4e0, 32'shd6d77cf2, 32'shd6d5151d, 32'shd6d2ad62, 32'shd6d045c0, 32'shd6cdde38, 
               32'shd6cb76c9, 32'shd6c90f73, 32'shd6c6a837, 32'shd6c44114, 32'shd6c1da0b, 32'shd6bf731b, 32'shd6bd0c45, 32'shd6baa588, 
               32'shd6b83ee4, 32'shd6b5d85a, 32'shd6b371ea, 32'shd6b10b92, 32'shd6aea555, 32'shd6ac3f31, 32'shd6a9d926, 32'shd6a77335, 
               32'shd6a50d5d, 32'shd6a2a79f, 32'shd6a041fa, 32'shd69ddc6f, 32'shd69b76fe, 32'shd69911a6, 32'shd696ac67, 32'shd6944742, 
               32'shd691e237, 32'shd68f7d45, 32'shd68d186d, 32'shd68ab3ae, 32'shd6884f09, 32'shd685ea7d, 32'shd683860b, 32'shd68121b3, 
               32'shd67ebd74, 32'shd67c594f, 32'shd679f543, 32'shd6779151, 32'shd6752d79, 32'shd672c9ba, 32'shd6706615, 32'shd66e028a, 
               32'shd66b9f18, 32'shd6693bc0, 32'shd666d881, 32'shd664755c, 32'shd6621251, 32'shd65faf60, 32'shd65d4c88, 32'shd65ae9ca, 
               32'shd6588725, 32'shd656249b, 32'shd653c229, 32'shd6515fd2, 32'shd64efd94, 32'shd64c9b71, 32'shd64a3966, 32'shd647d776, 
               32'shd645759f, 32'shd64313e2, 32'shd640b23f, 32'shd63e50b5, 32'shd63bef46, 32'shd6398df0, 32'shd6372cb3, 32'shd634cb91, 
               32'shd6326a88, 32'shd6300999, 32'shd62da8c4, 32'shd62b4809, 32'shd628e767, 32'shd62686e0, 32'shd6242672, 32'shd621c61e, 
               32'shd61f65e4, 32'shd61d05c3, 32'shd61aa5bd, 32'shd61845d0, 32'shd615e5fd, 32'shd6138644, 32'shd61126a5, 32'shd60ec720, 
               32'shd60c67b4, 32'shd60a0863, 32'shd607a92b, 32'shd6054a0d, 32'shd602eb0a, 32'shd6008c20, 32'shd5fe2d50, 32'shd5fbce9a, 
               32'shd5f96ffd, 32'shd5f7117b, 32'shd5f4b313, 32'shd5f254c4, 32'shd5eff690, 32'shd5ed9875, 32'shd5eb3a75, 32'shd5e8dc8e, 
               32'shd5e67ec1, 32'shd5e4210f, 32'shd5e1c376, 32'shd5df65f7, 32'shd5dd0892, 32'shd5daab48, 32'shd5d84e17, 32'shd5d5f100, 
               32'shd5d39403, 32'shd5d13721, 32'shd5ceda58, 32'shd5cc7da9, 32'shd5ca2115, 32'shd5c7c49a, 32'shd5c56839, 32'shd5c30bf3, 
               32'shd5c0afc6, 32'shd5be53b4, 32'shd5bbf7bc, 32'shd5b99bdd, 32'shd5b74019, 32'shd5b4e46f, 32'shd5b288df, 32'shd5b02d69, 
               32'shd5add20d, 32'shd5ab76cb, 32'shd5a91ba4, 32'shd5a6c096, 32'shd5a465a3, 32'shd5a20aca, 32'shd59fb00b, 32'shd59d5566, 
               32'shd59afadb, 32'shd598a06a, 32'shd5964614, 32'shd593ebd7, 32'shd59191b5, 32'shd58f37ad, 32'shd58cddbf, 32'shd58a83eb, 
               32'shd5882a32, 32'shd585d093, 32'shd583770e, 32'shd5811da3, 32'shd57ec452, 32'shd57c6b1c, 32'shd57a1200, 32'shd577b8fe, 
               32'shd5756016, 32'shd5730748, 32'shd570ae95, 32'shd56e55fc, 32'shd56bfd7d, 32'shd569a519, 32'shd5674ccf, 32'shd564f49f, 
               32'shd5629c89, 32'shd560448e, 32'shd55decad, 32'shd55b94e6, 32'shd5593d3a, 32'shd556e5a7, 32'shd5548e30, 32'shd55236d2, 
               32'shd54fdf8f, 32'shd54d8866, 32'shd54b3157, 32'shd548da63, 32'shd5468389, 32'shd5442cca, 32'shd541d625, 32'shd53f7f9a, 
               32'shd53d292a, 32'shd53ad2d4, 32'shd5387c98, 32'shd5362677, 32'shd533d070, 32'shd5317a84, 32'shd52f24b2, 32'shd52ccefa, 
               32'shd52a795d, 32'shd52823da, 32'shd525ce72, 32'shd5237924, 32'shd52123f0, 32'shd51eced7, 32'shd51c79d9, 32'shd51a24f5, 
               32'shd517d02b, 32'shd5157b7c, 32'shd51326e7, 32'shd510d26d, 32'shd50e7e0d, 32'shd50c29c8, 32'shd509d59d, 32'shd507818d, 
               32'shd5052d97, 32'shd502d9bc, 32'shd50085fb, 32'shd4fe3255, 32'shd4fbdec9, 32'shd4f98b58, 32'shd4f73801, 32'shd4f4e4c5, 
               32'shd4f291a4, 32'shd4f03e9d, 32'shd4edebb0, 32'shd4eb98de, 32'shd4e94627, 32'shd4e6f38b, 32'shd4e4a108, 32'shd4e24ea1, 
               32'shd4dffc54, 32'shd4ddaa22, 32'shd4db580a, 32'shd4d9060d, 32'shd4d6b42b, 32'shd4d46263, 32'shd4d210b5, 32'shd4cfbf23, 
               32'shd4cd6dab, 32'shd4cb1c4e, 32'shd4c8cb0b, 32'shd4c679e3, 32'shd4c428d6, 32'shd4c1d7e3, 32'shd4bf870b, 32'shd4bd364e, 
               32'shd4bae5ab, 32'shd4b89523, 32'shd4b644b6, 32'shd4b3f464, 32'shd4b1a42c, 32'shd4af540f, 32'shd4ad040c, 32'shd4aab425, 
               32'shd4a86458, 32'shd4a614a6, 32'shd4a3c50e, 32'shd4a17591, 32'shd49f2630, 32'shd49cd6e8, 32'shd49a87bc, 32'shd49838aa, 
               32'shd495e9b3, 32'shd4939ad7, 32'shd4914c16, 32'shd48efd6f, 32'shd48caee4, 32'shd48a6073, 32'shd488121d, 32'shd485c3e1, 
               32'shd48375c1, 32'shd48127bb, 32'shd47ed9d0, 32'shd47c8c00, 32'shd47a3e4b, 32'shd477f0b1, 32'shd475a332, 32'shd47355cd, 
               32'shd4710883, 32'shd46ebb54, 32'shd46c6e40, 32'shd46a2147, 32'shd467d469, 32'shd46587a6, 32'shd4633afd, 32'shd460ee70, 
               32'shd45ea1fd, 32'shd45c55a5, 32'shd45a0969, 32'shd457bd47, 32'shd4557140, 32'shd4532554, 32'shd450d983, 32'shd44e8dcd, 
               32'shd44c4232, 32'shd449f6b1, 32'shd447ab4c, 32'shd4456002, 32'shd44314d3, 32'shd440c9be, 32'shd43e7ec5, 32'shd43c33e7, 
               32'shd439e923, 32'shd4379e7b, 32'shd43553ee, 32'shd433097b, 32'shd430bf24, 32'shd42e74e8, 32'shd42c2ac6, 32'shd429e0c0, 
               32'shd42796d5, 32'shd4254d05, 32'shd4230350, 32'shd420b9b6, 32'shd41e7037, 32'shd41c26d3, 32'shd419dd8a, 32'shd417945c, 
               32'shd4154b4a, 32'shd4130252, 32'shd410b976, 32'shd40e70b4, 32'shd40c280e, 32'shd409df83, 32'shd4079713, 32'shd4054ebe, 
               32'shd4030684, 32'shd400be66, 32'shd3fe7662, 32'shd3fc2e7a, 32'shd3f9e6ad, 32'shd3f79efa, 32'shd3f55764, 32'shd3f30fe8, 
               32'shd3f0c887, 32'shd3ee8142, 32'shd3ec3a18, 32'shd3e9f309, 32'shd3e7ac15, 32'shd3e5653c, 32'shd3e31e7f, 32'shd3e0d7dd, 
               32'shd3de9156, 32'shd3dc4aea, 32'shd3da049a, 32'shd3d7be64, 32'shd3d5784a, 32'shd3d3324b, 32'shd3d0ec68, 32'shd3cea69f, 
               32'shd3cc60f2, 32'shd3ca1b61, 32'shd3c7d5ea, 32'shd3c5908f, 32'shd3c34b4f, 32'shd3c1062a, 32'shd3bec121, 32'shd3bc7c33, 
               32'shd3ba3760, 32'shd3b7f2a9, 32'shd3b5ae0d, 32'shd3b3698c, 32'shd3b12526, 32'shd3aee0dc, 32'shd3ac9cad, 32'shd3aa589a, 
               32'shd3a814a2, 32'shd3a5d0c5, 32'shd3a38d03, 32'shd3a1495d, 32'shd39f05d3, 32'shd39cc263, 32'shd39a7f0f, 32'shd3983bd7, 
               32'shd395f8ba, 32'shd393b5b8, 32'shd39172d2, 32'shd38f3007, 32'shd38ced57, 32'shd38aaac3, 32'shd388684a, 32'shd38625ed, 
               32'shd383e3ab, 32'shd381a185, 32'shd37f5f7a, 32'shd37d1d8a, 32'shd37adbb6, 32'shd37899fe, 32'shd3765861, 32'shd37416df, 
               32'shd371d579, 32'shd36f942e, 32'shd36d52ff, 32'shd36b11eb, 32'shd368d0f3, 32'shd3669017, 32'shd3644f55, 32'shd3620eb0, 
               32'shd35fce26, 32'shd35d8db7, 32'shd35b4d64, 32'shd3590d2c, 32'shd356cd11, 32'shd3548d10, 32'shd3524d2b, 32'shd3500d62, 
               32'shd34dcdb4, 32'shd34b8e22, 32'shd3494eab, 32'shd3470f50, 32'shd344d011, 32'shd34290ed, 32'shd34051e5, 32'shd33e12f8, 
               32'shd33bd427, 32'shd3399572, 32'shd33756d8, 32'shd335185a, 32'shd332d9f7, 32'shd3309bb0, 32'shd32e5d85, 32'shd32c1f75, 
               32'shd329e181, 32'shd327a3a9, 32'shd32565ec, 32'shd323284b, 32'shd320eac6, 32'shd31ead5c, 32'shd31c700f, 32'shd31a32dc, 
               32'shd317f5c6, 32'shd315b8cb, 32'shd3137bec, 32'shd3113f28, 32'shd30f0280, 32'shd30cc5f4, 32'shd30a8984, 32'shd3084d30, 
               32'shd30610f7, 32'shd303d4da, 32'shd30198d8, 32'shd2ff5cf3, 32'shd2fd2129, 32'shd2fae57b, 32'shd2f8a9e9, 32'shd2f66e72, 
               32'shd2f43318, 32'shd2f1f7d9, 32'shd2efbcb6, 32'shd2ed81ae, 32'shd2eb46c3, 32'shd2e90bf3, 32'shd2e6d13f, 32'shd2e496a7, 
               32'shd2e25c2b, 32'shd2e021ca, 32'shd2dde786, 32'shd2dbad5d, 32'shd2d97350, 32'shd2d7395f, 32'shd2d4ff8a, 32'shd2d2c5d0, 
               32'shd2d08c33, 32'shd2ce52b1, 32'shd2cc194c, 32'shd2c9e002, 32'shd2c7a6d4, 32'shd2c56dc2, 32'shd2c334cc, 32'shd2c0fbf1, 
               32'shd2bec333, 32'shd2bc8a91, 32'shd2ba520a, 32'shd2b8199f, 32'shd2b5e151, 32'shd2b3a91e, 32'shd2b17107, 32'shd2af390d, 
               32'shd2ad012e, 32'shd2aac96b, 32'shd2a891c4, 32'shd2a65a39, 32'shd2a422ca, 32'shd2a1eb77, 32'shd29fb440, 32'shd29d7d25, 
               32'shd29b4626, 32'shd2990f43, 32'shd296d87c, 32'shd294a1d0, 32'shd2926b41, 32'shd29034ce, 32'shd28dfe77, 32'shd28bc83d, 
               32'shd289921e, 32'shd2875c1b, 32'shd2852634, 32'shd282f069, 32'shd280babb, 32'shd27e8528, 32'shd27c4fb1, 32'shd27a1a57, 
               32'shd277e518, 32'shd275aff6, 32'shd2737af0, 32'shd2714606, 32'shd26f1138, 32'shd26cdc86, 32'shd26aa7f0, 32'shd2687376, 
               32'shd2663f19, 32'shd2640ad7, 32'shd261d6b2, 32'shd25fa2a9, 32'shd25d6ebc, 32'shd25b3aeb, 32'shd2590736, 32'shd256d39e, 
               32'shd254a021, 32'shd2526cc1, 32'shd250397d, 32'shd24e0655, 32'shd24bd34a, 32'shd249a05a, 32'shd2476d87, 32'shd2453ad0, 
               32'shd2430835, 32'shd240d5b6, 32'shd23ea354, 32'shd23c710e, 32'shd23a3ee4, 32'shd2380cd6, 32'shd235dae4, 32'shd233a90f, 
               32'shd2317756, 32'shd22f45b9, 32'shd22d1439, 32'shd22ae2d5, 32'shd228b18d, 32'shd2268061, 32'shd2244f52, 32'shd2221e5f, 
               32'shd21fed88, 32'shd21dbccd, 32'shd21b8c2f, 32'shd2195bad, 32'shd2172b48, 32'shd214fafe, 32'shd212cad1, 32'shd2109ac1, 
               32'shd20e6acc, 32'shd20c3af4, 32'shd20a0b39, 32'shd207db9a, 32'shd205ac17, 32'shd2037cb0, 32'shd2014d66, 32'shd1ff1e38, 
               32'shd1fcef27, 32'shd1fac032, 32'shd1f89159, 32'shd1f6629d, 32'shd1f433fd, 32'shd1f2057a, 32'shd1efd713, 32'shd1eda8c8, 
               32'shd1eb7a9a, 32'shd1e94c88, 32'shd1e71e93, 32'shd1e4f0ba, 32'shd1e2c2fd, 32'shd1e0955d, 32'shd1de67da, 32'shd1dc3a73, 
               32'shd1da0d28, 32'shd1d7dffa, 32'shd1d5b2e8, 32'shd1d385f3, 32'shd1d1591a, 32'shd1cf2c5e, 32'shd1ccffbe, 32'shd1cad33b, 
               32'shd1c8a6d4, 32'shd1c67a8a, 32'shd1c44e5c, 32'shd1c2224b, 32'shd1bff656, 32'shd1bdca7e, 32'shd1bb9ec2, 32'shd1b97323, 
               32'shd1b747a0, 32'shd1b51c3a, 32'shd1b2f0f1, 32'shd1b0c5c4, 32'shd1ae9ab4, 32'shd1ac6fc0, 32'shd1aa44e9, 32'shd1a81a2e, 
               32'shd1a5ef90, 32'shd1a3c50f, 32'shd1a19aaa, 32'shd19f7062, 32'shd19d4636, 32'shd19b1c27, 32'shd198f235, 32'shd196c85f, 
               32'shd1949ea6, 32'shd1927509, 32'shd1904b89, 32'shd18e2226, 32'shd18bf8e0, 32'shd189cfb6, 32'shd187a6a8, 32'shd1857db8, 
               32'shd18354e4, 32'shd1812c2d, 32'shd17f0392, 32'shd17cdb14, 32'shd17ab2b3, 32'shd1788a6f, 32'shd1766247, 32'shd1743a3c, 
               32'shd172124d, 32'shd16fea7c, 32'shd16dc2c7, 32'shd16b9b2f, 32'shd16973b3, 32'shd1674c54, 32'shd1652512, 32'shd162fded, 
               32'shd160d6e5, 32'shd15eaff9, 32'shd15c892a, 32'shd15a6278, 32'shd1583be2, 32'shd156156a, 32'shd153ef0e, 32'shd151c8cf, 
               32'shd14fa2ad, 32'shd14d7ca7, 32'shd14b56be, 32'shd14930f3, 32'shd1470b44, 32'shd144e5b1, 32'shd142c03c, 32'shd1409ae3, 
               32'shd13e75a8, 32'shd13c5089, 32'shd13a2b87, 32'shd13806a2, 32'shd135e1d9, 32'shd133bd2e, 32'shd131989f, 32'shd12f742d, 
               32'shd12d4fd9, 32'shd12b2ba1, 32'shd1290786, 32'shd126e387, 32'shd124bfa6, 32'shd1229be2, 32'shd120783a, 32'shd11e54b0, 
               32'shd11c3142, 32'shd11a0df1, 32'shd117eabd, 32'shd115c7a7, 32'shd113a4ad, 32'shd11181d0, 32'shd10f5f10, 32'shd10d3c6d, 
               32'shd10b19e7, 32'shd108f77d, 32'shd106d531, 32'shd104b302, 32'shd10290f0, 32'shd1006efb, 32'shd0fe4d22, 32'shd0fc2b67, 
               32'shd0fa09c9, 32'shd0f7e848, 32'shd0f5c6e3, 32'shd0f3a59c, 32'shd0f18472, 32'shd0ef6365, 32'shd0ed4275, 32'shd0eb21a2, 
               32'shd0e900ec, 32'shd0e6e053, 32'shd0e4bfd7, 32'shd0e29f78, 32'shd0e07f36, 32'shd0de5f11, 32'shd0dc3f0a, 32'shd0da1f1f, 
               32'shd0d7ff51, 32'shd0d5dfa1, 32'shd0d3c00e, 32'shd0d1a097, 32'shd0cf813e, 32'shd0cd6202, 32'shd0cb42e3, 32'shd0c923e1, 
               32'shd0c704fd, 32'shd0c4e635, 32'shd0c2c78b, 32'shd0c0a8fe, 32'shd0be8a8d, 32'shd0bc6c3a, 32'shd0ba4e05, 32'shd0b82fec, 
               32'shd0b611f1, 32'shd0b3f412, 32'shd0b1d651, 32'shd0afb8ad, 32'shd0ad9b26, 32'shd0ab7dbd, 32'shd0a96070, 32'shd0a74341, 
               32'shd0a5262f, 32'shd0a3093a, 32'shd0a0ec63, 32'shd09ecfa8, 32'shd09cb30b, 32'shd09a968b, 32'shd0987a29, 32'shd0965de3, 
               32'shd09441bb, 32'shd09225b0, 32'shd09009c3, 32'shd08dedf2, 32'shd08bd23f, 32'shd089b6a9, 32'shd0879b31, 32'shd0857fd5, 
               32'shd0836497, 32'shd0814977, 32'shd07f2e73, 32'shd07d138d, 32'shd07af8c4, 32'shd078de19, 32'shd076c38b, 32'shd074a91a, 
               32'shd0728ec6, 32'shd0707490, 32'shd06e5a77, 32'shd06c407c, 32'shd06a269d, 32'shd0680cdd, 32'shd065f339, 32'shd063d9b3, 
               32'shd061c04a, 32'shd05fa6ff, 32'shd05d8dd1, 32'shd05b74c0, 32'shd0595bcd, 32'shd05742f7, 32'shd0552a3f, 32'shd05311a4, 
               32'shd050f926, 32'shd04ee0c6, 32'shd04cc884, 32'shd04ab05e, 32'shd0489856, 32'shd046806c, 32'shd044689f, 32'shd04250ef, 
               32'shd040395d, 32'shd03e21e8, 32'shd03c0a91, 32'shd039f357, 32'shd037dc3b, 32'shd035c53c, 32'shd033ae5b, 32'shd0319797, 
               32'shd02f80f1, 32'shd02d6a68, 32'shd02b53fc, 32'shd0293dae, 32'shd027277e, 32'shd025116b, 32'shd022fb76, 32'shd020e59e, 
               32'shd01ecfe4, 32'shd01cba47, 32'shd01aa4c8, 32'shd0188f66, 32'shd0167a22, 32'shd01464fc, 32'shd0124ff3, 32'shd0103b07, 
               32'shd00e2639, 32'shd00c1189, 32'shd009fcf6, 32'shd007e881, 32'shd005d42a, 32'shd003bff0, 32'shd001abd3, 32'shcfff97d5, 
               32'shcffd83f4, 32'shcffb7030, 32'shcff95c8a, 32'shcff74902, 32'shcff53597, 32'shcff3224a, 32'shcff10f1b, 32'shcfeefc09, 
               32'shcfece915, 32'shcfead63f, 32'shcfe8c386, 32'shcfe6b0eb, 32'shcfe49e6d, 32'shcfe28c0e, 32'shcfe079cc, 32'shcfde67a7, 
               32'shcfdc55a1, 32'shcfda43b8, 32'shcfd831ec, 32'shcfd6203f, 32'shcfd40eaf, 32'shcfd1fd3d, 32'shcfcfebe8, 32'shcfcddab2, 
               32'shcfcbc999, 32'shcfc9b89d, 32'shcfc7a7c0, 32'shcfc59700, 32'shcfc3865e, 32'shcfc175da, 32'shcfbf6573, 32'shcfbd552b, 
               32'shcfbb4500, 32'shcfb934f2, 32'shcfb72503, 32'shcfb51531, 32'shcfb3057d, 32'shcfb0f5e7, 32'shcfaee66f, 32'shcfacd715, 
               32'shcfaac7d8, 32'shcfa8b8b9, 32'shcfa6a9b8, 32'shcfa49ad5, 32'shcfa28c10, 32'shcfa07d68, 32'shcf9e6edf, 32'shcf9c6073, 
               32'shcf9a5225, 32'shcf9843f5, 32'shcf9635e2, 32'shcf9427ee, 32'shcf921a17, 32'shcf900c5f, 32'shcf8dfec4, 32'shcf8bf147, 
               32'shcf89e3e8, 32'shcf87d6a7, 32'shcf85c984, 32'shcf83bc7e, 32'shcf81af97, 32'shcf7fa2cd, 32'shcf7d9622, 32'shcf7b8994, 
               32'shcf797d24, 32'shcf7770d3, 32'shcf75649f, 32'shcf735889, 32'shcf714c91, 32'shcf6f40b7, 32'shcf6d34fb, 32'shcf6b295d, 
               32'shcf691ddd, 32'shcf67127a, 32'shcf650736, 32'shcf62fc10, 32'shcf60f108, 32'shcf5ee61e, 32'shcf5cdb51, 32'shcf5ad0a3, 
               32'shcf58c613, 32'shcf56bba1, 32'shcf54b14d, 32'shcf52a716, 32'shcf509cfe, 32'shcf4e9304, 32'shcf4c8928, 32'shcf4a7f6a, 
               32'shcf4875ca, 32'shcf466c48, 32'shcf4462e4, 32'shcf42599f, 32'shcf405077, 32'shcf3e476d, 32'shcf3c3e82, 32'shcf3a35b4, 
               32'shcf382d05, 32'shcf362473, 32'shcf341c00, 32'shcf3213ab, 32'shcf300b74, 32'shcf2e035b, 32'shcf2bfb60, 32'shcf29f383, 
               32'shcf27ebc5, 32'shcf25e424, 32'shcf23dca2, 32'shcf21d53e, 32'shcf1fcdf8, 32'shcf1dc6d0, 32'shcf1bbfc6, 32'shcf19b8db, 
               32'shcf17b20d, 32'shcf15ab5e, 32'shcf13a4cd, 32'shcf119e5a, 32'shcf0f9805, 32'shcf0d91cf, 32'shcf0b8bb7, 32'shcf0985bc, 
               32'shcf077fe1, 32'shcf057a23, 32'shcf037483, 32'shcf016f02, 32'shceff699f, 32'shcefd645a, 32'shcefb5f34, 32'shcef95a2b, 
               32'shcef75541, 32'shcef55075, 32'shcef34bc8, 32'shcef14738, 32'shceef42c7, 32'shceed3e74, 32'shceeb3a40, 32'shcee93629, 
               32'shcee73231, 32'shcee52e58, 32'shcee32a9c, 32'shcee126ff, 32'shcedf2380, 32'shcedd2020, 32'shcedb1cde, 32'shced919ba, 
               32'shced716b4, 32'shced513cd, 32'shced31104, 32'shced10e59, 32'shcecf0bcd, 32'shcecd095f, 32'shcecb070f, 32'shcec904de, 
               32'shcec702cb, 32'shcec500d7, 32'shcec2ff01, 32'shcec0fd49, 32'shcebefbb0, 32'shcebcfa35, 32'shcebaf8d8, 32'shceb8f79a, 
               32'shceb6f67a, 32'shceb4f579, 32'shceb2f496, 32'shceb0f3d1, 32'shceaef32b, 32'shceacf2a3, 32'shceaaf23a, 32'shcea8f1ef, 
               32'shcea6f1c2, 32'shcea4f1b4, 32'shcea2f1c5, 32'shcea0f1f4, 32'shce9ef241, 32'shce9cf2ad, 32'shce9af337, 32'shce98f3e0, 
               32'shce96f4a7, 32'shce94f58c, 32'shce92f691, 32'shce90f7b3, 32'shce8ef8f4, 32'shce8cfa54, 32'shce8afbd2, 32'shce88fd6f, 
               32'shce86ff2a, 32'shce850104, 32'shce8302fc, 32'shce810512, 32'shce7f0748, 32'shce7d099b, 32'shce7b0c0e, 32'shce790e9f, 
               32'shce77114e, 32'shce75141c, 32'shce731709, 32'shce711a14, 32'shce6f1d3d, 32'shce6d2086, 32'shce6b23ec, 32'shce692772, 
               32'shce672b16, 32'shce652ed8, 32'shce6332ba, 32'shce6136b9, 32'shce5f3ad8, 32'shce5d3f15, 32'shce5b4370, 32'shce5947eb, 
               32'shce574c84, 32'shce55513b, 32'shce535611, 32'shce515b06, 32'shce4f6019, 32'shce4d654c, 32'shce4b6a9c, 32'shce49700c, 
               32'shce47759a, 32'shce457b47, 32'shce438112, 32'shce4186fc, 32'shce3f8d05, 32'shce3d932c, 32'shce3b9973, 32'shce399fd7, 
               32'shce37a65b, 32'shce35acfd, 32'shce33b3be, 32'shce31ba9e, 32'shce2fc19c, 32'shce2dc8ba, 32'shce2bcff5, 32'shce29d750, 
               32'shce27dec9, 32'shce25e662, 32'shce23ee18, 32'shce21f5ee, 32'shce1ffde2, 32'shce1e05f6, 32'shce1c0e28, 32'shce1a1678, 
               32'shce181ee8, 32'shce162776, 32'shce143023, 32'shce1238ef, 32'shce1041d9, 32'shce0e4ae3, 32'shce0c540b, 32'shce0a5d52, 
               32'shce0866b8, 32'shce06703d, 32'shce0479e0, 32'shce0283a3, 32'shce008d84, 32'shcdfe9784, 32'shcdfca1a3, 32'shcdfaabe1, 
               32'shcdf8b63d, 32'shcdf6c0b9, 32'shcdf4cb53, 32'shcdf2d60c, 32'shcdf0e0e4, 32'shcdeeebdb, 32'shcdecf6f1, 32'shcdeb0226, 
               32'shcde90d79, 32'shcde718ec, 32'shcde5247d, 32'shcde3302e, 32'shcde13bfd, 32'shcddf47eb, 32'shcddd53f8, 32'shcddb6024, 
               32'shcdd96c6f, 32'shcdd778d9, 32'shcdd58562, 32'shcdd39209, 32'shcdd19ed0, 32'shcdcfabb6, 32'shcdcdb8ba, 32'shcdcbc5de, 
               32'shcdc9d320, 32'shcdc7e082, 32'shcdc5ee02, 32'shcdc3fba2, 32'shcdc20960, 32'shcdc0173e, 32'shcdbe253a, 32'shcdbc3356, 
               32'shcdba4190, 32'shcdb84fea, 32'shcdb65e62, 32'shcdb46cfa, 32'shcdb27bb0, 32'shcdb08a86, 32'shcdae997a, 32'shcdaca88e, 
               32'shcdaab7c0, 32'shcda8c712, 32'shcda6d683, 32'shcda4e613, 32'shcda2f5c2, 32'shcda10590, 32'shcd9f157d, 32'shcd9d2589, 
               32'shcd9b35b4, 32'shcd9945fe, 32'shcd975668, 32'shcd9566f0, 32'shcd937798, 32'shcd91885e, 32'shcd8f9944, 32'shcd8daa49, 
               32'shcd8bbb6d, 32'shcd89ccb0, 32'shcd87de12, 32'shcd85ef94, 32'shcd840134, 32'shcd8212f4, 32'shcd8024d3, 32'shcd7e36d1, 
               32'shcd7c48ee, 32'shcd7a5b2a, 32'shcd786d85, 32'shcd768000, 32'shcd74929a, 32'shcd72a553, 32'shcd70b82b, 32'shcd6ecb22, 
               32'shcd6cde39, 32'shcd6af16e, 32'shcd6904c3, 32'shcd671837, 32'shcd652bcb, 32'shcd633f7d, 32'shcd61534f, 32'shcd5f6740, 
               32'shcd5d7b50, 32'shcd5b8f80, 32'shcd59a3ce, 32'shcd57b83c, 32'shcd55ccca, 32'shcd53e176, 32'shcd51f642, 32'shcd500b2d, 
               32'shcd4e2037, 32'shcd4c3560, 32'shcd4a4aa9, 32'shcd486011, 32'shcd467599, 32'shcd448b3f, 32'shcd42a105, 32'shcd40b6ea, 
               32'shcd3eccef, 32'shcd3ce313, 32'shcd3af956, 32'shcd390fb8, 32'shcd37263a, 32'shcd353cdb, 32'shcd33539c, 32'shcd316a7b, 
               32'shcd2f817b, 32'shcd2d9899, 32'shcd2bafd7, 32'shcd29c734, 32'shcd27deb0, 32'shcd25f64c, 32'shcd240e08, 32'shcd2225e2, 
               32'shcd203ddc, 32'shcd1e55f6, 32'shcd1c6e2e, 32'shcd1a8687, 32'shcd189efe, 32'shcd16b795, 32'shcd14d04b, 32'shcd12e921, 
               32'shcd110216, 32'shcd0f1b2b, 32'shcd0d345f, 32'shcd0b4db3, 32'shcd096725, 32'shcd0780b8, 32'shcd059a6a, 32'shcd03b43b, 
               32'shcd01ce2b, 32'shccffe83c, 32'shccfe026b, 32'shccfc1cba, 32'shccfa3729, 32'shccf851b7, 32'shccf66c64, 32'shccf48731, 
               32'shccf2a21d, 32'shccf0bd29, 32'shcceed855, 32'shccecf3a0, 32'shcceb0f0a, 32'shcce92a94, 32'shcce7463e, 32'shcce56206, 
               32'shcce37def, 32'shcce199f7, 32'shccdfb61f, 32'shccddd266, 32'shccdbeecc, 32'shccda0b52, 32'shccd827f8, 32'shccd644bd, 
               32'shccd461a2, 32'shccd27ea7, 32'shccd09bcb, 32'shccceb90e, 32'shccccd671, 32'shcccaf3f4, 32'shccc91196, 32'shccc72f58, 
               32'shccc54d3a, 32'shccc36b3b, 32'shccc1895c, 32'shccbfa79c, 32'shccbdc5fc, 32'shccbbe47b, 32'shccba031a, 32'shccb821d9, 
               32'shccb640b8, 32'shccb45fb6, 32'shccb27ed3, 32'shccb09e11, 32'shccaebd6e, 32'shccacdcea, 32'shccaafc87, 32'shcca91c43, 
               32'shcca73c1e, 32'shcca55c1a, 32'shcca37c35, 32'shcca19c6f, 32'shcc9fbcca, 32'shcc9ddd44, 32'shcc9bfddd, 32'shcc9a1e97, 
               32'shcc983f70, 32'shcc966069, 32'shcc948182, 32'shcc92a2ba, 32'shcc90c412, 32'shcc8ee58a, 32'shcc8d0721, 32'shcc8b28d8, 
               32'shcc894aaf, 32'shcc876ca6, 32'shcc858ebc, 32'shcc83b0f3, 32'shcc81d349, 32'shcc7ff5be, 32'shcc7e1854, 32'shcc7c3b09, 
               32'shcc7a5dde, 32'shcc7880d3, 32'shcc76a3e8, 32'shcc74c71c, 32'shcc72ea70, 32'shcc710de4, 32'shcc6f3178, 32'shcc6d552c, 
               32'shcc6b78ff, 32'shcc699cf2, 32'shcc67c105, 32'shcc65e538, 32'shcc64098b, 32'shcc622dfd, 32'shcc605290, 32'shcc5e7742, 
               32'shcc5c9c14, 32'shcc5ac106, 32'shcc58e618, 32'shcc570b4a, 32'shcc55309b, 32'shcc53560c, 32'shcc517b9e, 32'shcc4fa14f, 
               32'shcc4dc720, 32'shcc4bed11, 32'shcc4a1322, 32'shcc483952, 32'shcc465fa3, 32'shcc448614, 32'shcc42aca4, 32'shcc40d354, 
               32'shcc3efa25, 32'shcc3d2115, 32'shcc3b4825, 32'shcc396f55, 32'shcc3796a5, 32'shcc35be15, 32'shcc33e5a5, 32'shcc320d55, 
               32'shcc303524, 32'shcc2e5d14, 32'shcc2c8524, 32'shcc2aad54, 32'shcc28d5a3, 32'shcc26fe13, 32'shcc2526a2, 32'shcc234f52, 
               32'shcc217822, 32'shcc1fa111, 32'shcc1dca21, 32'shcc1bf350, 32'shcc1a1ca0, 32'shcc184610, 32'shcc166f9f, 32'shcc14994f, 
               32'shcc12c31f, 32'shcc10ed0e, 32'shcc0f171e, 32'shcc0d414e, 32'shcc0b6b9e, 32'shcc09960e, 32'shcc07c09e, 32'shcc05eb4e, 
               32'shcc04161e, 32'shcc02410e, 32'shcc006c1e, 32'shcbfe974e, 32'shcbfcc29f, 32'shcbfaee0f, 32'shcbf919a0, 32'shcbf74550, 
               32'shcbf57121, 32'shcbf39d12, 32'shcbf1c923, 32'shcbeff554, 32'shcbee21a5, 32'shcbec4e16, 32'shcbea7aa7, 32'shcbe8a759, 
               32'shcbe6d42b, 32'shcbe5011c, 32'shcbe32e2e, 32'shcbe15b60, 32'shcbdf88b3, 32'shcbddb625, 32'shcbdbe3b7, 32'shcbda116a, 
               32'shcbd83f3d, 32'shcbd66d30, 32'shcbd49b43, 32'shcbd2c977, 32'shcbd0f7ca, 32'shcbcf263e, 32'shcbcd54d2, 32'shcbcb8386, 
               32'shcbc9b25a, 32'shcbc7e14f, 32'shcbc61064, 32'shcbc43f99, 32'shcbc26eee, 32'shcbc09e64, 32'shcbbecdf9, 32'shcbbcfdaf, 
               32'shcbbb2d85, 32'shcbb95d7c, 32'shcbb78d92, 32'shcbb5bdc9, 32'shcbb3ee20, 32'shcbb21e98, 32'shcbb04f2f, 32'shcbae7fe7, 
               32'shcbacb0bf, 32'shcbaae1b8, 32'shcba912d1, 32'shcba7440a, 32'shcba57563, 32'shcba3a6dd, 32'shcba1d877, 32'shcba00a31, 
               32'shcb9e3c0b, 32'shcb9c6e06, 32'shcb9aa021, 32'shcb98d25d, 32'shcb9704b9, 32'shcb953735, 32'shcb9369d1, 32'shcb919c8e, 
               32'shcb8fcf6b, 32'shcb8e0269, 32'shcb8c3587, 32'shcb8a68c5, 32'shcb889c23, 32'shcb86cfa2, 32'shcb850342, 32'shcb833701, 
               32'shcb816ae1, 32'shcb7f9ee2, 32'shcb7dd303, 32'shcb7c0744, 32'shcb7a3ba5, 32'shcb787027, 32'shcb76a4ca, 32'shcb74d98d, 
               32'shcb730e70, 32'shcb714373, 32'shcb6f7898, 32'shcb6daddc, 32'shcb6be341, 32'shcb6a18c6, 32'shcb684e6c, 32'shcb668432, 
               32'shcb64ba19, 32'shcb62f020, 32'shcb612648, 32'shcb5f5c90, 32'shcb5d92f8, 32'shcb5bc981, 32'shcb5a002b, 32'shcb5836f4, 
               32'shcb566ddf, 32'shcb54a4ea, 32'shcb52dc15, 32'shcb511361, 32'shcb4f4acd, 32'shcb4d825a, 32'shcb4bba08, 32'shcb49f1d5, 
               32'shcb4829c4, 32'shcb4661d3, 32'shcb449a02, 32'shcb42d252, 32'shcb410ac3, 32'shcb3f4354, 32'shcb3d7c05, 32'shcb3bb4d7, 
               32'shcb39edca, 32'shcb3826dd, 32'shcb366011, 32'shcb349965, 32'shcb32d2da, 32'shcb310c70, 32'shcb2f4626, 32'shcb2d7ffc, 
               32'shcb2bb9f4, 32'shcb29f40b, 32'shcb282e44, 32'shcb26689d, 32'shcb24a316, 32'shcb22ddb1, 32'shcb21186b, 32'shcb1f5347, 
               32'shcb1d8e43, 32'shcb1bc95f, 32'shcb1a049d, 32'shcb183ffb, 32'shcb167b79, 32'shcb14b718, 32'shcb12f2d8, 32'shcb112eb9, 
               32'shcb0f6aba, 32'shcb0da6dc, 32'shcb0be31e, 32'shcb0a1f81, 32'shcb085c05, 32'shcb0698a9, 32'shcb04d56e, 32'shcb031254, 
               32'shcb014f5b, 32'shcaff8c82, 32'shcafdc9ca, 32'shcafc0732, 32'shcafa44bc, 32'shcaf88266, 32'shcaf6c030, 32'shcaf4fe1c, 
               32'shcaf33c28, 32'shcaf17a55, 32'shcaefb8a2, 32'shcaedf711, 32'shcaec35a0, 32'shcaea744f, 32'shcae8b320, 32'shcae6f211, 
               32'shcae53123, 32'shcae37056, 32'shcae1afaa, 32'shcadfef1e, 32'shcade2eb3, 32'shcadc6e69, 32'shcadaae40, 32'shcad8ee37, 
               32'shcad72e4f, 32'shcad56e88, 32'shcad3aee2, 32'shcad1ef5d, 32'shcad02ff8, 32'shcace70b4, 32'shcaccb191, 32'shcacaf28f, 
               32'shcac933ae, 32'shcac774ed, 32'shcac5b64e, 32'shcac3f7cf, 32'shcac23971, 32'shcac07b34, 32'shcabebd17, 32'shcabcff1c, 
               32'shcabb4141, 32'shcab98388, 32'shcab7c5ef, 32'shcab60877, 32'shcab44b1f, 32'shcab28de9, 32'shcab0d0d4, 32'shcaaf13df, 
               32'shcaad570c, 32'shcaab9a59, 32'shcaa9ddc7, 32'shcaa82156, 32'shcaa66506, 32'shcaa4a8d7, 32'shcaa2ecc9, 32'shcaa130db, 
               32'shca9f750f, 32'shca9db964, 32'shca9bfdd9, 32'shca9a4270, 32'shca988727, 32'shca96cbff, 32'shca9510f8, 32'shca935613, 
               32'shca919b4e, 32'shca8fe0aa, 32'shca8e2627, 32'shca8c6bc5, 32'shca8ab184, 32'shca88f764, 32'shca873d65, 32'shca858387, 
               32'shca83c9ca, 32'shca82102e, 32'shca8056b3, 32'shca7e9d59, 32'shca7ce420, 32'shca7b2b08, 32'shca797211, 32'shca77b93b, 
               32'shca760086, 32'shca7447f2, 32'shca728f7f, 32'shca70d72d, 32'shca6f1efc, 32'shca6d66ec, 32'shca6baefd, 32'shca69f72f, 
               32'shca683f83, 32'shca6687f7, 32'shca64d08d, 32'shca631943, 32'shca61621b, 32'shca5fab13, 32'shca5df42d, 32'shca5c3d68, 
               32'shca5a86c4, 32'shca58d041, 32'shca5719df, 32'shca55639e, 32'shca53ad7e, 32'shca51f780, 32'shca5041a2, 32'shca4e8be6, 
               32'shca4cd64b, 32'shca4b20d0, 32'shca496b77, 32'shca47b640, 32'shca460129, 32'shca444c33, 32'shca42975f, 32'shca40e2ac, 
               32'shca3f2e19, 32'shca3d79a8, 32'shca3bc559, 32'shca3a112a, 32'shca385d1d, 32'shca36a930, 32'shca34f565, 32'shca3341bb, 
               32'shca318e32, 32'shca2fdacb, 32'shca2e2784, 32'shca2c745f, 32'shca2ac15b, 32'shca290e79, 32'shca275bb7, 32'shca25a917, 
               32'shca23f698, 32'shca22443a, 32'shca2091fd, 32'shca1edfe2, 32'shca1d2de7, 32'shca1b7c0e, 32'shca19ca57, 32'shca1818c0, 
               32'shca16674b, 32'shca14b5f7, 32'shca1304c4, 32'shca1153b3, 32'shca0fa2c3, 32'shca0df1f4, 32'shca0c4146, 32'shca0a90ba, 
               32'shca08e04f, 32'shca073005, 32'shca057fdd, 32'shca03cfd5, 32'shca021fef, 32'shca00702b, 32'shc9fec088, 32'shc9fd1106, 
               32'shc9fb61a5, 32'shc9f9b266, 32'shc9f80348, 32'shc9f6544b, 32'shc9f4a570, 32'shc9f2f6b6, 32'shc9f1481d, 32'shc9ef99a6, 
               32'shc9edeb50, 32'shc9ec3d1b, 32'shc9ea8f08, 32'shc9e8e116, 32'shc9e73346, 32'shc9e58596, 32'shc9e3d809, 32'shc9e22a9c, 
               32'shc9e07d51, 32'shc9ded028, 32'shc9dd231f, 32'shc9db7639, 32'shc9d9c973, 32'shc9d81ccf, 32'shc9d6704c, 32'shc9d4c3eb, 
               32'shc9d317ab, 32'shc9d16b8d, 32'shc9cfbf90, 32'shc9ce13b4, 32'shc9cc67fa, 32'shc9cabc62, 32'shc9c910ea, 32'shc9c76595, 
               32'shc9c5ba60, 32'shc9c40f4d, 32'shc9c2645c, 32'shc9c0b98c, 32'shc9bf0edd, 32'shc9bd6450, 32'shc9bbb9e5, 32'shc9ba0f9b, 
               32'shc9b86572, 32'shc9b6bb6b, 32'shc9b51185, 32'shc9b367c1, 32'shc9b1be1e, 32'shc9b0149d, 32'shc9ae6b3d, 32'shc9acc1ff, 
               32'shc9ab18e3, 32'shc9a96fe7, 32'shc9a7c70e, 32'shc9a61e56, 32'shc9a475bf, 32'shc9a2cd4a, 32'shc9a124f7, 32'shc99f7cc5, 
               32'shc99dd4b4, 32'shc99c2cc5, 32'shc99a84f8, 32'shc998dd4c, 32'shc99735c2, 32'shc9958e59, 32'shc993e712, 32'shc9923fed, 
               32'shc99098e9, 32'shc98ef206, 32'shc98d4b45, 32'shc98ba4a6, 32'shc989fe29, 32'shc98857cd, 32'shc986b192, 32'shc9850b79, 
               32'shc9836582, 32'shc981bfac, 32'shc98019f8, 32'shc97e7466, 32'shc97ccef5, 32'shc97b29a6, 32'shc9798479, 32'shc977df6d, 
               32'shc9763a83, 32'shc97495ba, 32'shc972f113, 32'shc9714c8e, 32'shc96fa82a, 32'shc96e03e8, 32'shc96c5fc8, 32'shc96abbc9, 
               32'shc96917ec, 32'shc9677431, 32'shc965d097, 32'shc9642d1f, 32'shc96289c9, 32'shc960e695, 32'shc95f4382, 32'shc95da090, 
               32'shc95bfdc1, 32'shc95a5b13, 32'shc958b887, 32'shc957161d, 32'shc95573d4, 32'shc953d1ad, 32'shc9522fa8, 32'shc9508dc5, 
               32'shc94eec03, 32'shc94d4a63, 32'shc94ba8e5, 32'shc94a0788, 32'shc948664d, 32'shc946c534, 32'shc945243d, 32'shc9438368, 
               32'shc941e2b4, 32'shc9404222, 32'shc93ea1b2, 32'shc93d0163, 32'shc93b6137, 32'shc939c12c, 32'shc9382143, 32'shc936817b, 
               32'shc934e1d6, 32'shc9334252, 32'shc931a2f0, 32'shc93003b0, 32'shc92e6492, 32'shc92cc596, 32'shc92b26bb, 32'shc9298802, 
               32'shc927e96b, 32'shc9264af6, 32'shc924aca3, 32'shc9230e71, 32'shc9217062, 32'shc91fd274, 32'shc91e34a8, 32'shc91c96fe, 
               32'shc91af976, 32'shc9195c0f, 32'shc917becb, 32'shc91621a8, 32'shc91484a8, 32'shc912e7c9, 32'shc9114b0c, 32'shc90fae71, 
               32'shc90e11f7, 32'shc90c75a0, 32'shc90ad96b, 32'shc9093d57, 32'shc907a166, 32'shc9060596, 32'shc90469e8, 32'shc902ce5c, 
               32'shc90132f2, 32'shc8ff97aa, 32'shc8fdfc84, 32'shc8fc6180, 32'shc8fac69e, 32'shc8f92bdd, 32'shc8f7913f, 32'shc8f5f6c3, 
               32'shc8f45c68, 32'shc8f2c230, 32'shc8f12819, 32'shc8ef8e24, 32'shc8edf452, 32'shc8ec5aa1, 32'shc8eac112, 32'shc8e927a6, 
               32'shc8e78e5b, 32'shc8e5f532, 32'shc8e45c2c, 32'shc8e2c347, 32'shc8e12a84, 32'shc8df91e3, 32'shc8ddf965, 32'shc8dc6108, 
               32'shc8dac8cd, 32'shc8d930b4, 32'shc8d798be, 32'shc8d600e9, 32'shc8d46936, 32'shc8d2d1a6, 32'shc8d13a37, 32'shc8cfa2eb, 
               32'shc8ce0bc0, 32'shc8cc74b8, 32'shc8caddd1, 32'shc8c9470d, 32'shc8c7b06b, 32'shc8c619eb, 32'shc8c4838d, 32'shc8c2ed50, 
               32'shc8c15736, 32'shc8bfc13f, 32'shc8be2b69, 32'shc8bc95b5, 32'shc8bb0023, 32'shc8b96ab4, 32'shc8b7d566, 32'shc8b6403b, 
               32'shc8b4ab32, 32'shc8b3164a, 32'shc8b18185, 32'shc8afece2, 32'shc8ae5862, 32'shc8acc403, 32'shc8ab2fc6, 32'shc8a99bac, 
               32'shc8a807b4, 32'shc8a673dd, 32'shc8a4e029, 32'shc8a34c98, 32'shc8a1b928, 32'shc8a025da, 32'shc89e92af, 32'shc89cffa6, 
               32'shc89b6cbf, 32'shc899d9fa, 32'shc8984757, 32'shc896b4d6, 32'shc8952278, 32'shc893903c, 32'shc891fe22, 32'shc8906c2a, 
               32'shc88eda54, 32'shc88d48a1, 32'shc88bb710, 32'shc88a25a1, 32'shc8889454, 32'shc8870329, 32'shc8857221, 32'shc883e13b, 
               32'shc8825077, 32'shc880bfd5, 32'shc87f2f56, 32'shc87d9ef8, 32'shc87c0ebd, 32'shc87a7ea5, 32'shc878eeae, 32'shc8775eda, 
               32'shc875cf28, 32'shc8743f98, 32'shc872b02b, 32'shc87120e0, 32'shc86f91b7, 32'shc86e02b0, 32'shc86c73cc, 32'shc86ae50a, 
               32'shc869566a, 32'shc867c7ec, 32'shc8663991, 32'shc864ab58, 32'shc8631d42, 32'shc8618f4d, 32'shc860017b, 32'shc85e73cc, 
               32'shc85ce63e, 32'shc85b58d3, 32'shc859cb8a, 32'shc8583e64, 32'shc856b160, 32'shc855247e, 32'shc85397bf, 32'shc8520b22, 
               32'shc8507ea7, 32'shc84ef24f, 32'shc84d6619, 32'shc84bda05, 32'shc84a4e14, 32'shc848c245, 32'shc8473698, 32'shc845ab0e, 
               32'shc8441fa6, 32'shc8429461, 32'shc841093e, 32'shc83f7e3d, 32'shc83df35f, 32'shc83c68a3, 32'shc83ade0a, 32'shc8395393, 
               32'shc837c93e, 32'shc8363f0c, 32'shc834b4fc, 32'shc8332b0e, 32'shc831a143, 32'shc830179b, 32'shc82e8e15, 32'shc82d04b1, 
               32'shc82b7b70, 32'shc829f251, 32'shc8286954, 32'shc826e07a, 32'shc82557c3, 32'shc823cf2e, 32'shc82246bb, 32'shc820be6b, 
               32'shc81f363d, 32'shc81dae32, 32'shc81c2649, 32'shc81a9e83, 32'shc81916df, 32'shc8178f5e, 32'shc81607ff, 32'shc81480c3, 
               32'shc812f9a9, 32'shc81172b2, 32'shc80febdd, 32'shc80e652b, 32'shc80cde9b, 32'shc80b582e, 32'shc809d1e3, 32'shc8084bba, 
               32'shc806c5b5, 32'shc8053fd2, 32'shc803ba11, 32'shc8023473, 32'shc800aef7, 32'shc7ff299e, 32'shc7fda468, 32'shc7fc1f54, 
               32'shc7fa9a62, 32'shc7f91593, 32'shc7f790e7, 32'shc7f60c5d, 32'shc7f487f6, 32'shc7f303b1, 32'shc7f17f8f, 32'shc7effb90, 
               32'shc7ee77b3, 32'shc7ecf3f9, 32'shc7eb7061, 32'shc7e9ecec, 32'shc7e8699a, 32'shc7e6e66a, 32'shc7e5635c, 32'shc7e3e072, 
               32'shc7e25daa, 32'shc7e0db04, 32'shc7df5881, 32'shc7ddd621, 32'shc7dc53e3, 32'shc7dad1c9, 32'shc7d94fd0, 32'shc7d7cdfb, 
               32'shc7d64c47, 32'shc7d4cab7, 32'shc7d34949, 32'shc7d1c7fe, 32'shc7d046d6, 32'shc7cec5d0, 32'shc7cd44ed, 32'shc7cbc42c, 
               32'shc7ca438f, 32'shc7c8c313, 32'shc7c742bb, 32'shc7c5c285, 32'shc7c44272, 32'shc7c2c282, 32'shc7c142b4, 32'shc7bfc309, 
               32'shc7be4381, 32'shc7bcc41b, 32'shc7bb44d8, 32'shc7b9c5b8, 32'shc7b846ba, 32'shc7b6c7e0, 32'shc7b54928, 32'shc7b3ca92, 
               32'shc7b24c20, 32'shc7b0cdd0, 32'shc7af4fa3, 32'shc7add198, 32'shc7ac53b1, 32'shc7aad5ec, 32'shc7a9584a, 32'shc7a7daca, 
               32'shc7a65d6e, 32'shc7a4e034, 32'shc7a3631d, 32'shc7a1e628, 32'shc7a06957, 32'shc79eeca8, 32'shc79d701c, 32'shc79bf3b3, 
               32'shc79a776c, 32'shc798fb48, 32'shc7977f48, 32'shc7960369, 32'shc79487ae, 32'shc7930c16, 32'shc79190a0, 32'shc790154d, 
               32'shc78e9a1d, 32'shc78d1f10, 32'shc78ba425, 32'shc78a295e, 32'shc788aeb9, 32'shc7873437, 32'shc785b9d8, 32'shc7843f9c, 
               32'shc782c582, 32'shc7814b8c, 32'shc77fd1b8, 32'shc77e5807, 32'shc77cde79, 32'shc77b650e, 32'shc779ebc5, 32'shc77872a0, 
               32'shc776f99d, 32'shc77580be, 32'shc7740801, 32'shc7728f67, 32'shc77116f0, 32'shc76f9e9c, 32'shc76e266b, 32'shc76cae5c, 
               32'shc76b3671, 32'shc769bea8, 32'shc7684702, 32'shc766cf80, 32'shc7655820, 32'shc763e0e3, 32'shc76269c9, 32'shc760f2d2, 
               32'shc75f7bfe, 32'shc75e054c, 32'shc75c8ebe, 32'shc75b1853, 32'shc759a20a, 32'shc7582be5, 32'shc756b5e2, 32'shc7554003, 
               32'shc753ca46, 32'shc75254ac, 32'shc750df36, 32'shc74f69e2, 32'shc74df4b1, 32'shc74c7fa4, 32'shc74b0ab9, 32'shc74995f1, 
               32'shc748214c, 32'shc746acca, 32'shc745386b, 32'shc743c42f, 32'shc7425016, 32'shc740dc21, 32'shc73f684e, 32'shc73df49e, 
               32'shc73c8111, 32'shc73b0da7, 32'shc7399a60, 32'shc738273d, 32'shc736b43c, 32'shc735415e, 32'shc733cea3, 32'shc7325c0c, 
               32'shc730e997, 32'shc72f7745, 32'shc72e0517, 32'shc72c930b, 32'shc72b2123, 32'shc729af5d, 32'shc7283dbb, 32'shc726cc3c, 
               32'shc7255ae0, 32'shc723e9a6, 32'shc7227890, 32'shc721079d, 32'shc71f96ce, 32'shc71e2621, 32'shc71cb597, 32'shc71b4530, 
               32'shc719d4ed, 32'shc71864cc, 32'shc716f4cf, 32'shc71584f5, 32'shc714153e, 32'shc712a5aa, 32'shc7113639, 32'shc70fc6eb, 
               32'shc70e57c0, 32'shc70ce8b9, 32'shc70b79d4, 32'shc70a0b13, 32'shc7089c75, 32'shc7072dfa, 32'shc705bfa2, 32'shc704516d, 
               32'shc702e35c, 32'shc701756d, 32'shc70007a2, 32'shc6fe99fa, 32'shc6fd2c75, 32'shc6fbbf13, 32'shc6fa51d5, 32'shc6f8e4b9, 
               32'shc6f777c1, 32'shc6f60aec, 32'shc6f49e3a, 32'shc6f331ab, 32'shc6f1c540, 32'shc6f058f8, 32'shc6eeecd3, 32'shc6ed80d1, 
               32'shc6ec14f2, 32'shc6eaa936, 32'shc6e93d9e, 32'shc6e7d229, 32'shc6e666d7, 32'shc6e4fba9, 32'shc6e3909d, 32'shc6e225b5, 
               32'shc6e0baf0, 32'shc6df504f, 32'shc6dde5d0, 32'shc6dc7b75, 32'shc6db113d, 32'shc6d9a728, 32'shc6d83d37, 32'shc6d6d369, 
               32'shc6d569be, 32'shc6d40036, 32'shc6d296d1, 32'shc6d12d90, 32'shc6cfc472, 32'shc6ce5b78, 32'shc6ccf2a1, 32'shc6cb89ed, 
               32'shc6ca215c, 32'shc6c8b8ee, 32'shc6c750a4, 32'shc6c5e87d, 32'shc6c4807a, 32'shc6c31899, 32'shc6c1b0dd, 32'shc6c04943, 
               32'shc6bee1cd, 32'shc6bd7a7a, 32'shc6bc134a, 32'shc6baac3d, 32'shc6b94554, 32'shc6b7de8f, 32'shc6b677ec, 32'shc6b5116d, 
               32'shc6b3ab12, 32'shc6b244d9, 32'shc6b0dec4, 32'shc6af78d3, 32'shc6ae1304, 32'shc6acad59, 32'shc6ab47d2, 32'shc6a9e26e, 
               32'shc6a87d2d, 32'shc6a7180f, 32'shc6a5b315, 32'shc6a44e3e, 32'shc6a2e98b, 32'shc6a184fb, 32'shc6a0208f, 32'shc69ebc45, 
               32'shc69d5820, 32'shc69bf41d, 32'shc69a903e, 32'shc6992c83, 32'shc697c8eb, 32'shc6966576, 32'shc6950224, 32'shc6939ef6, 
               32'shc6923bec, 32'shc690d905, 32'shc68f7641, 32'shc68e13a1, 32'shc68cb124, 32'shc68b4ecb, 32'shc689ec95, 32'shc6888a83, 
               32'shc6872894, 32'shc685c6c8, 32'shc6846520, 32'shc683039b, 32'shc681a23a, 32'shc68040fc, 32'shc67edfe2, 32'shc67d7eeb, 
               32'shc67c1e18, 32'shc67abd68, 32'shc6795cdc, 32'shc677fc73, 32'shc6769c2e, 32'shc6753c0c, 32'shc673dc0d, 32'shc6727c32, 
               32'shc6711c7b, 32'shc66fbce7, 32'shc66e5d77, 32'shc66cfe2a, 32'shc66b9f01, 32'shc66a3ffb, 32'shc668e119, 32'shc667825a, 
               32'shc66623be, 32'shc664c547, 32'shc66366f3, 32'shc66208c2, 32'shc660aab5, 32'shc65f4ccb, 32'shc65def05, 32'shc65c9163, 
               32'shc65b33e4, 32'shc659d688, 32'shc6587951, 32'shc6571c3c, 32'shc655bf4c, 32'shc654627f, 32'shc65305d5, 32'shc651a94f, 
               32'shc6504ced, 32'shc64ef0ae, 32'shc64d9493, 32'shc64c389b, 32'shc64adcc7, 32'shc6498117, 32'shc648258a, 32'shc646ca21, 
               32'shc6456edb, 32'shc64413b9, 32'shc642b8bb, 32'shc6415de0, 32'shc6400329, 32'shc63ea896, 32'shc63d4e26, 32'shc63bf3d9, 
               32'shc63a99b1, 32'shc6393fac, 32'shc637e5ca, 32'shc6368c0d, 32'shc6353273, 32'shc633d8fc, 32'shc6327faa, 32'shc631267a, 
               32'shc62fcd6f, 32'shc62e7487, 32'shc62d1bc3, 32'shc62bc323, 32'shc62a6aa6, 32'shc629124d, 32'shc627ba17, 32'shc6266206, 
               32'shc6250a18, 32'shc623b24d, 32'shc6225aa6, 32'shc6210323, 32'shc61fabc4, 32'shc61e5489, 32'shc61cfd71, 32'shc61ba67d, 
               32'shc61a4fac, 32'shc618f8ff, 32'shc617a276, 32'shc6164c11, 32'shc614f5cf, 32'shc6139fb2, 32'shc61249b7, 32'shc610f3e1, 
               32'shc60f9e2e, 32'shc60e489f, 32'shc60cf334, 32'shc60b9ded, 32'shc60a48c9, 32'shc608f3c9, 32'shc6079eed, 32'shc6064a35, 
               32'shc604f5a0, 32'shc603a12f, 32'shc6024ce2, 32'shc600f8b9, 32'shc5ffa4b3, 32'shc5fe50d1, 32'shc5fcfd13, 32'shc5fba979, 
               32'shc5fa5603, 32'shc5f902b0, 32'shc5f7af81, 32'shc5f65c76, 32'shc5f5098f, 32'shc5f3b6cb, 32'shc5f2642c, 32'shc5f111b0, 
               32'shc5efbf58, 32'shc5ee6d24, 32'shc5ed1b13, 32'shc5ebc927, 32'shc5ea775e, 32'shc5e925b9, 32'shc5e7d438, 32'shc5e682db, 
               32'shc5e531a1, 32'shc5e3e08c, 32'shc5e28f9a, 32'shc5e13ecc, 32'shc5dfee22, 32'shc5de9d9c, 32'shc5dd4d3a, 32'shc5dbfcfb, 
               32'shc5daace1, 32'shc5d95cea, 32'shc5d80d17, 32'shc5d6bd68, 32'shc5d56ddd, 32'shc5d41e76, 32'shc5d2cf33, 32'shc5d18013, 
               32'shc5d03118, 32'shc5cee240, 32'shc5cd938c, 32'shc5cc44fc, 32'shc5caf690, 32'shc5c9a848, 32'shc5c85a24, 32'shc5c70c24, 
               32'shc5c5be47, 32'shc5c4708f, 32'shc5c322fb, 32'shc5c1d58a, 32'shc5c0883d, 32'shc5bf3b15, 32'shc5bdee10, 32'shc5bca12f, 
               32'shc5bb5472, 32'shc5ba07d9, 32'shc5b8bb64, 32'shc5b76f13, 32'shc5b622e6, 32'shc5b4d6dd, 32'shc5b38af8, 32'shc5b23f37, 
               32'shc5b0f399, 32'shc5afa820, 32'shc5ae5ccb, 32'shc5ad1199, 32'shc5abc68c, 32'shc5aa7ba3, 32'shc5a930dd, 32'shc5a7e63c, 
               32'shc5a69bbe, 32'shc5a55165, 32'shc5a4072f, 32'shc5a2bd1e, 32'shc5a17330, 32'shc5a02967, 32'shc59edfc2, 32'shc59d9640, 
               32'shc59c4ce3, 32'shc59b03a9, 32'shc599ba94, 32'shc59871a3, 32'shc59728d5, 32'shc595e02c, 32'shc59497a7, 32'shc5934f46, 
               32'shc5920708, 32'shc590beef, 32'shc58f76fa, 32'shc58e2f29, 32'shc58ce77c, 32'shc58b9ff3, 32'shc58a588e, 32'shc589114e, 
               32'shc587ca31, 32'shc5868338, 32'shc5853c63, 32'shc583f5b3, 32'shc582af26, 32'shc58168be, 32'shc580227a, 32'shc57edc5a, 
               32'shc57d965d, 32'shc57c5085, 32'shc57b0ad1, 32'shc579c542, 32'shc5787fd6, 32'shc5773a8e, 32'shc575f56b, 32'shc574b06b, 
               32'shc5736b90, 32'shc57226d9, 32'shc570e246, 32'shc56f9dd7, 32'shc56e598c, 32'shc56d1565, 32'shc56bd163, 32'shc56a8d84, 
               32'shc56949ca, 32'shc5680634, 32'shc566c2c2, 32'shc5657f74, 32'shc5643c4a, 32'shc562f944, 32'shc561b663, 32'shc56073a6, 
               32'shc55f310d, 32'shc55dee98, 32'shc55cac47, 32'shc55b6a1a, 32'shc55a2812, 32'shc558e62e, 32'shc557a46e, 32'shc55662d2, 
               32'shc555215a, 32'shc553e007, 32'shc5529ed7, 32'shc5515dcc, 32'shc5501ce5, 32'shc54edc23, 32'shc54d9b84, 32'shc54c5b0a, 
               32'shc54b1ab4, 32'shc549da82, 32'shc5489a74, 32'shc5475a8b, 32'shc5461ac6, 32'shc544db25, 32'shc5439ba8, 32'shc5425c4f, 
               32'shc5411d1b, 32'shc53fde0b, 32'shc53e9f1f, 32'shc53d6057, 32'shc53c21b4, 32'shc53ae335, 32'shc539a4da, 32'shc53866a4, 
               32'shc5372891, 32'shc535eaa3, 32'shc534acd9, 32'shc5336f34, 32'shc53231b3, 32'shc530f456, 32'shc52fb71d, 32'shc52e7a09, 
               32'shc52d3d18, 32'shc52c004d, 32'shc52ac3a5, 32'shc5298722, 32'shc5284ac3, 32'shc5270e88, 32'shc525d272, 32'shc5249680, 
               32'shc5235ab2, 32'shc5221f08, 32'shc520e383, 32'shc51fa822, 32'shc51e6ce6, 32'shc51d31ce, 32'shc51bf6da, 32'shc51abc0a, 
               32'shc519815f, 32'shc51846d8, 32'shc5170c75, 32'shc515d237, 32'shc514981d, 32'shc5135e28, 32'shc5122457, 32'shc510eaaa, 
               32'shc50fb121, 32'shc50e77bd, 32'shc50d3e7d, 32'shc50c0562, 32'shc50acc6b, 32'shc5099398, 32'shc5085aea, 32'shc5072260, 
               32'shc505e9fb, 32'shc504b1b9, 32'shc503799d, 32'shc50241a4, 32'shc50109d0, 32'shc4ffd221, 32'shc4fe9a95, 32'shc4fd632f, 
               32'shc4fc2bec, 32'shc4faf4ce, 32'shc4f9bdd4, 32'shc4f886ff, 32'shc4f7504e, 32'shc4f619c2, 32'shc4f4e35a, 32'shc4f3ad17, 
               32'shc4f276f7, 32'shc4f140fd, 32'shc4f00b27, 32'shc4eed575, 32'shc4ed9fe7, 32'shc4ec6a7e, 32'shc4eb353a, 32'shc4ea001a, 
               32'shc4e8cb1e, 32'shc4e79647, 32'shc4e66194, 32'shc4e52d06, 32'shc4e3f89c, 32'shc4e2c457, 32'shc4e19036, 32'shc4e05c3a, 
               32'shc4df2862, 32'shc4ddf4ae, 32'shc4dcc11f, 32'shc4db8db5, 32'shc4da5a6f, 32'shc4d9274d, 32'shc4d7f450, 32'shc4d6c177, 
               32'shc4d58ec3, 32'shc4d45c34, 32'shc4d329c9, 32'shc4d1f782, 32'shc4d0c560, 32'shc4cf9363, 32'shc4ce6189, 32'shc4cd2fd5, 
               32'shc4cbfe45, 32'shc4caccd9, 32'shc4c99b92, 32'shc4c86a70, 32'shc4c73972, 32'shc4c60899, 32'shc4c4d7e4, 32'shc4c3a753, 
               32'shc4c276e8, 32'shc4c146a0, 32'shc4c0167e, 32'shc4bee680, 32'shc4bdb6a6, 32'shc4bc86f1, 32'shc4bb5760, 32'shc4ba27f5, 
               32'shc4b8f8ad, 32'shc4b7c98a, 32'shc4b69a8c, 32'shc4b56bb3, 32'shc4b43cfd, 32'shc4b30e6d, 32'shc4b1e001, 32'shc4b0b1ba, 
               32'shc4af8397, 32'shc4ae5599, 32'shc4ad27bf, 32'shc4abfa0a, 32'shc4aacc7a, 32'shc4a99f0e, 32'shc4a871c7, 32'shc4a744a4, 
               32'shc4a617a6, 32'shc4a4eacd, 32'shc4a3be18, 32'shc4a29188, 32'shc4a1651c, 32'shc4a038d6, 32'shc49f0cb3, 32'shc49de0b6, 
               32'shc49cb4dd, 32'shc49b8928, 32'shc49a5d98, 32'shc499322d, 32'shc49806e7, 32'shc496dbc5, 32'shc495b0c8, 32'shc49485ef, 
               32'shc4935b3c, 32'shc49230ac, 32'shc4910642, 32'shc48fdbfc, 32'shc48eb1db, 32'shc48d87de, 32'shc48c5e06, 32'shc48b3453, 
               32'shc48a0ac4, 32'shc488e15b, 32'shc487b815, 32'shc4868ef5, 32'shc48565f9, 32'shc4843d22, 32'shc4831470, 32'shc481ebe2, 
               32'shc480c379, 32'shc47f9b34, 32'shc47e7315, 32'shc47d4b1a, 32'shc47c2344, 32'shc47afb92, 32'shc479d405, 32'shc478ac9d, 
               32'shc477855a, 32'shc4765e3b, 32'shc4753741, 32'shc474106c, 32'shc472e9bc, 32'shc471c330, 32'shc4709cc9, 32'shc46f7687, 
               32'shc46e5069, 32'shc46d2a71, 32'shc46c049d, 32'shc46adeee, 32'shc469b963, 32'shc46893fd, 32'shc4676ebc, 32'shc46649a0, 
               32'shc46524a9, 32'shc463ffd6, 32'shc462db28, 32'shc461b69f, 32'shc460923b, 32'shc45f6dfb, 32'shc45e49e0, 32'shc45d25ea, 
               32'shc45c0219, 32'shc45ade6c, 32'shc459bae5, 32'shc4589782, 32'shc4577444, 32'shc456512b, 32'shc4552e36, 32'shc4540b67, 
               32'shc452e8bc, 32'shc451c636, 32'shc450a3d4, 32'shc44f8198, 32'shc44e5f80, 32'shc44d3d8e, 32'shc44c1bc0, 32'shc44afa17, 
               32'shc449d892, 32'shc448b733, 32'shc44795f8, 32'shc44674e3, 32'shc44553f2, 32'shc4443326, 32'shc443127e, 32'shc441f1fc, 
               32'shc440d19e, 32'shc43fb166, 32'shc43e9152, 32'shc43d7163, 32'shc43c5199, 32'shc43b31f4, 32'shc43a1273, 32'shc438f318, 
               32'shc437d3e1, 32'shc436b4cf, 32'shc43595e3, 32'shc434771b, 32'shc4335877, 32'shc43239f9, 32'shc4311ba0, 32'shc42ffd6b, 
               32'shc42edf5c, 32'shc42dc171, 32'shc42ca3ac, 32'shc42b860b, 32'shc42a688f, 32'shc4294b38, 32'shc4282e06, 32'shc42710f9, 
               32'shc425f410, 32'shc424d74d, 32'shc423baae, 32'shc4229e35, 32'shc42181e0, 32'shc42065b1, 32'shc41f49a6, 32'shc41e2dc0, 
               32'shc41d11ff, 32'shc41bf664, 32'shc41adaed, 32'shc419bf9b, 32'shc418a46d, 32'shc4178965, 32'shc4166e82, 32'shc41553c4, 
               32'shc414392b, 32'shc4131eb7, 32'shc4120467, 32'shc410ea3d, 32'shc40fd037, 32'shc40eb657, 32'shc40d9c9c, 32'shc40c8305, 
               32'shc40b6994, 32'shc40a5047, 32'shc4093720, 32'shc4081e1d, 32'shc4070540, 32'shc405ec87, 32'shc404d3f4, 32'shc403bb85, 
               32'shc402a33c, 32'shc4018b17, 32'shc4007318, 32'shc3ff5b3d, 32'shc3fe4388, 32'shc3fd2bf7, 32'shc3fc148c, 32'shc3fafd45, 
               32'shc3f9e624, 32'shc3f8cf27, 32'shc3f7b850, 32'shc3f6a19e, 32'shc3f58b10, 32'shc3f474a8, 32'shc3f35e65, 32'shc3f24847, 
               32'shc3f1324e, 32'shc3f01c7a, 32'shc3ef06cb, 32'shc3edf141, 32'shc3ecdbdc, 32'shc3ebc69c, 32'shc3eab181, 32'shc3e99c8b, 
               32'shc3e887bb, 32'shc3e7730f, 32'shc3e65e88, 32'shc3e54a27, 32'shc3e435ea, 32'shc3e321d3, 32'shc3e20de1, 32'shc3e0fa14, 
               32'shc3dfe66c, 32'shc3ded2e9, 32'shc3ddbf8b, 32'shc3dcac52, 32'shc3db993e, 32'shc3da8650, 32'shc3d97386, 32'shc3d860e2, 
               32'shc3d74e62, 32'shc3d63c08, 32'shc3d529d3, 32'shc3d417c3, 32'shc3d305d8, 32'shc3d1f413, 32'shc3d0e272, 32'shc3cfd0f7, 
               32'shc3cebfa0, 32'shc3cdae6f, 32'shc3cc9d63, 32'shc3cb8c7c, 32'shc3ca7bba, 32'shc3c96b1e, 32'shc3c85aa6, 32'shc3c74a54, 
               32'shc3c63a26, 32'shc3c52a1e, 32'shc3c41a3b, 32'shc3c30a7e, 32'shc3c1fae5, 32'shc3c0eb71, 32'shc3bfdc23, 32'shc3beccfa, 
               32'shc3bdbdf6, 32'shc3bcaf17, 32'shc3bba05e, 32'shc3ba91c9, 32'shc3b9835a, 32'shc3b87510, 32'shc3b766eb, 32'shc3b658eb, 
               32'shc3b54b11, 32'shc3b43d5b, 32'shc3b32fcb, 32'shc3b22260, 32'shc3b1151b, 32'shc3b007fa, 32'shc3aefaff, 32'shc3adee28, 
               32'shc3ace178, 32'shc3abd4ec, 32'shc3aac885, 32'shc3a9bc44, 32'shc3a8b028, 32'shc3a7a431, 32'shc3a6985f, 32'shc3a58cb3, 
               32'shc3a4812c, 32'shc3a375ca, 32'shc3a26a8d, 32'shc3a15f76, 32'shc3a05484, 32'shc39f49b7, 32'shc39e3f0f, 32'shc39d348c, 
               32'shc39c2a2f, 32'shc39b1ff7, 32'shc39a15e4, 32'shc3990bf7, 32'shc398022f, 32'shc396f88c, 32'shc395ef0e, 32'shc394e5b6, 
               32'shc393dc82, 32'shc392d375, 32'shc391ca8c, 32'shc390c1c9, 32'shc38fb92a, 32'shc38eb0b2, 32'shc38da85e, 32'shc38ca030, 
               32'shc38b9827, 32'shc38a9043, 32'shc3898885, 32'shc38880ec, 32'shc3877978, 32'shc386722a, 32'shc3856b01, 32'shc38463fd, 
               32'shc3835d1e, 32'shc3825665, 32'shc3814fd1, 32'shc3804963, 32'shc37f4319, 32'shc37e3cf6, 32'shc37d36f7, 32'shc37c311e, 
               32'shc37b2b6a, 32'shc37a25db, 32'shc3792072, 32'shc3781b2e, 32'shc377160f, 32'shc3761116, 32'shc3750c42, 32'shc3740793, 
               32'shc373030a, 32'shc371fea6, 32'shc370fa68, 32'shc36ff64e, 32'shc36ef25b, 32'shc36dee8c, 32'shc36ceae3, 32'shc36be75f, 
               32'shc36ae401, 32'shc369e0c8, 32'shc368ddb4, 32'shc367dac6, 32'shc366d7fd, 32'shc365d55a, 32'shc364d2dc, 32'shc363d083, 
               32'shc362ce50, 32'shc361cc42, 32'shc360ca59, 32'shc35fc896, 32'shc35ec6f8, 32'shc35dc580, 32'shc35cc42d, 32'shc35bc2ff, 
               32'shc35ac1f7, 32'shc359c114, 32'shc358c057, 32'shc357bfbf, 32'shc356bf4d, 32'shc355bf00, 32'shc354bed8, 32'shc353bed6, 
               32'shc352bef9, 32'shc351bf41, 32'shc350bfaf, 32'shc34fc043, 32'shc34ec0fc, 32'shc34dc1da, 32'shc34cc2de, 32'shc34bc407, 
               32'shc34ac556, 32'shc349c6ca, 32'shc348c864, 32'shc347ca23, 32'shc346cc07, 32'shc345ce11, 32'shc344d041, 32'shc343d295, 
               32'shc342d510, 32'shc341d7b0, 32'shc340da75, 32'shc33fdd60, 32'shc33ee070, 32'shc33de3a5, 32'shc33ce701, 32'shc33bea81, 
               32'shc33aee27, 32'shc339f1f3, 32'shc338f5e4, 32'shc337f9fb, 32'shc336fe37, 32'shc3360298, 32'shc3350720, 32'shc3340bcc, 
               32'shc333109e, 32'shc3321596, 32'shc3311ab3, 32'shc3301ff5, 32'shc32f255e, 32'shc32e2aeb, 32'shc32d309e, 32'shc32c3677, 
               32'shc32b3c75, 32'shc32a4299, 32'shc32948e2, 32'shc3284f51, 32'shc32755e5, 32'shc3265c9f, 32'shc325637f, 32'shc3246a83, 
               32'shc32371ae, 32'shc32278fe, 32'shc3218073, 32'shc320880e, 32'shc31f8fcf, 32'shc31e97b5, 32'shc31d9fc1, 32'shc31ca7f2, 
               32'shc31bb049, 32'shc31ab8c6, 32'shc319c168, 32'shc318ca2f, 32'shc317d31c, 32'shc316dc2f, 32'shc315e567, 32'shc314eec5, 
               32'shc313f848, 32'shc31301f1, 32'shc3120bc0, 32'shc31115b4, 32'shc3101fce, 32'shc30f2a0d, 32'shc30e3472, 32'shc30d3efd, 
               32'shc30c49ad, 32'shc30b5482, 32'shc30a5f7e, 32'shc3096a9f, 32'shc30875e5, 32'shc3078151, 32'shc3068ce3, 32'shc305989a, 
               32'shc304a477, 32'shc303b07a, 32'shc302bca2, 32'shc301c8f0, 32'shc300d563, 32'shc2ffe1fc, 32'shc2feeebb, 32'shc2fdfb9f, 
               32'shc2fd08a9, 32'shc2fc15d9, 32'shc2fb232e, 32'shc2fa30a9, 32'shc2f93e4a, 32'shc2f84c10, 32'shc2f759fc, 32'shc2f6680d, 
               32'shc2f57644, 32'shc2f484a1, 32'shc2f39323, 32'shc2f2a1cb, 32'shc2f1b099, 32'shc2f0bf8c, 32'shc2efcea6, 32'shc2eedde4, 
               32'shc2eded49, 32'shc2ecfcd3, 32'shc2ec0c82, 32'shc2eb1c58, 32'shc2ea2c53, 32'shc2e93c74, 32'shc2e84cba, 32'shc2e75d26, 
               32'shc2e66db8, 32'shc2e57e70, 32'shc2e48f4d, 32'shc2e3a050, 32'shc2e2b178, 32'shc2e1c2c7, 32'shc2e0d43b, 32'shc2dfe5d4, 
               32'shc2def794, 32'shc2de0979, 32'shc2dd1b84, 32'shc2dc2db4, 32'shc2db400a, 32'shc2da5286, 32'shc2d96528, 32'shc2d877f0, 
               32'shc2d78add, 32'shc2d69df0, 32'shc2d5b128, 32'shc2d4c486, 32'shc2d3d80a, 32'shc2d2ebb4, 32'shc2d1ff84, 32'shc2d11379, 
               32'shc2d02794, 32'shc2cf3bd5, 32'shc2ce503b, 32'shc2cd64c7, 32'shc2cc7979, 32'shc2cb8e51, 32'shc2caa34f, 32'shc2c9b872, 
               32'shc2c8cdbb, 32'shc2c7e32a, 32'shc2c6f8be, 32'shc2c60e78, 32'shc2c52459, 32'shc2c43a5e, 32'shc2c3508a, 32'shc2c266db, 
               32'shc2c17d52, 32'shc2c093ef, 32'shc2bfaab2, 32'shc2bec19b, 32'shc2bdd8a9, 32'shc2bcefdd, 32'shc2bc0737, 32'shc2bb1eb6, 
               32'shc2ba365c, 32'shc2b94e27, 32'shc2b86618, 32'shc2b77e2f, 32'shc2b6966c, 32'shc2b5aece, 32'shc2b4c756, 32'shc2b3e004, 
               32'shc2b2f8d8, 32'shc2b211d2, 32'shc2b12af1, 32'shc2b04437, 32'shc2af5da2, 32'shc2ae7733, 32'shc2ad90ea, 32'shc2acaac6, 
               32'shc2abc4c9, 32'shc2aadef1, 32'shc2a9f93f, 32'shc2a913b3, 32'shc2a82e4d, 32'shc2a7490c, 32'shc2a663f2, 32'shc2a57efd, 
               32'shc2a49a2e, 32'shc2a3b585, 32'shc2a2d102, 32'shc2a1eca5, 32'shc2a1086d, 32'shc2a0245c, 32'shc29f4070, 32'shc29e5caa, 
               32'shc29d790a, 32'shc29c9590, 32'shc29bb23c, 32'shc29acf0d, 32'shc299ec05, 32'shc2990922, 32'shc2982665, 32'shc29743ce, 
               32'shc296615d, 32'shc2957f12, 32'shc2949ced, 32'shc293baed, 32'shc292d914, 32'shc291f760, 32'shc29115d3, 32'shc290346b, 
               32'shc28f5329, 32'shc28e720d, 32'shc28d9117, 32'shc28cb047, 32'shc28bcf9c, 32'shc28aef18, 32'shc28a0eb9, 32'shc2892e81, 
               32'shc2884e6e, 32'shc2876e82, 32'shc2868ebb, 32'shc285af1a, 32'shc284cf9f, 32'shc283f04a, 32'shc283111b, 32'shc2823211, 
               32'shc281532e, 32'shc2807471, 32'shc27f95d9, 32'shc27eb768, 32'shc27dd91c, 32'shc27cfaf7, 32'shc27c1cf7, 32'shc27b3f1e, 
               32'shc27a616a, 32'shc27983dc, 32'shc278a674, 32'shc277c932, 32'shc276ec16, 32'shc2760f20, 32'shc2753250, 32'shc27455a6, 
               32'shc2737922, 32'shc2729cc4, 32'shc271c08c, 32'shc270e47a, 32'shc270088e, 32'shc26f2cc7, 32'shc26e5127, 32'shc26d75ad, 
               32'shc26c9a58, 32'shc26bbf2a, 32'shc26ae422, 32'shc26a093f, 32'shc2692e83, 32'shc26853ed, 32'shc267797c, 32'shc2669f32, 
               32'shc265c50e, 32'shc264eb0f, 32'shc2641137, 32'shc2633785, 32'shc2625df8, 32'shc2618492, 32'shc260ab51, 32'shc25fd237, 
               32'shc25ef943, 32'shc25e2074, 32'shc25d47cc, 32'shc25c6f4a, 32'shc25b96ee, 32'shc25abeb7, 32'shc259e6a7, 32'shc2590ebd, 
               32'shc25836f9, 32'shc2575f5b, 32'shc25687e3, 32'shc255b091, 32'shc254d965, 32'shc254025f, 32'shc2532b7f, 32'shc25254c5, 
               32'shc2517e31, 32'shc250a7c3, 32'shc24fd17c, 32'shc24efb5a, 32'shc24e255e, 32'shc24d4f89, 32'shc24c79d9, 32'shc24ba450, 
               32'shc24aceed, 32'shc249f9af, 32'shc2492498, 32'shc2484fa7, 32'shc2477adc, 32'shc246a637, 32'shc245d1b8, 32'shc244fd5f, 
               32'shc244292c, 32'shc243551f, 32'shc2428139, 32'shc241ad78, 32'shc240d9de, 32'shc2400669, 32'shc23f331b, 32'shc23e5ff3, 
               32'shc23d8cf1, 32'shc23cba15, 32'shc23be75f, 32'shc23b14cf, 32'shc23a4265, 32'shc2397021, 32'shc2389e04, 32'shc237cc0d, 
               32'shc236fa3b, 32'shc2362890, 32'shc235570b, 32'shc23485ac, 32'shc233b473, 32'shc232e361, 32'shc2321274, 32'shc23141ae, 
               32'shc230710d, 32'shc22fa093, 32'shc22ed03f, 32'shc22e0011, 32'shc22d3009, 32'shc22c6028, 32'shc22b906c, 32'shc22ac0d7, 
               32'shc229f167, 32'shc229221e, 32'shc22852fb, 32'shc22783fe, 32'shc226b528, 32'shc225e677, 32'shc22517ed, 32'shc2244989, 
               32'shc2237b4b, 32'shc222ad33, 32'shc221df41, 32'shc2211176, 32'shc22043d0, 32'shc21f7651, 32'shc21ea8f8, 32'shc21ddbc5, 
               32'shc21d0eb8, 32'shc21c41d2, 32'shc21b7511, 32'shc21aa877, 32'shc219dc03, 32'shc2190fb5, 32'shc218438e, 32'shc217778c, 
               32'shc216abb1, 32'shc215dffc, 32'shc215146d, 32'shc2144904, 32'shc2137dc2, 32'shc212b2a5, 32'shc211e7af, 32'shc2111cdf, 
               32'shc2105236, 32'shc20f87b2, 32'shc20ebd55, 32'shc20df31e, 32'shc20d290d, 32'shc20c5f22, 32'shc20b955e, 32'shc20acbc0, 
               32'shc20a0248, 32'shc20938f6, 32'shc2086fca, 32'shc207a6c5, 32'shc206dde6, 32'shc206152d, 32'shc2054c9b, 32'shc204842e, 
               32'shc203bbe8, 32'shc202f3c8, 32'shc2022bce, 32'shc20163fb, 32'shc2009c4e, 32'shc1ffd4c7, 32'shc1ff0d66, 32'shc1fe462b, 
               32'shc1fd7f17, 32'shc1fcb829, 32'shc1fbf161, 32'shc1fb2ac0, 32'shc1fa6445, 32'shc1f99df0, 32'shc1f8d7c1, 32'shc1f811b9, 
               32'shc1f74bd6, 32'shc1f6861a, 32'shc1f5c085, 32'shc1f4fb15, 32'shc1f435cc, 32'shc1f370a9, 32'shc1f2abad, 32'shc1f1e6d7, 
               32'shc1f12227, 32'shc1f05d9d, 32'shc1ef9939, 32'shc1eed4fc, 32'shc1ee10e5, 32'shc1ed4cf5, 32'shc1ec892b, 32'shc1ebc587, 
               32'shc1eb0209, 32'shc1ea3eb1, 32'shc1e97b80, 32'shc1e8b876, 32'shc1e7f591, 32'shc1e732d3, 32'shc1e6703b, 32'shc1e5adc9, 
               32'shc1e4eb7e, 32'shc1e42959, 32'shc1e3675a, 32'shc1e2a582, 32'shc1e1e3d0, 32'shc1e12244, 32'shc1e060df, 32'shc1df9fa0, 
               32'shc1dede87, 32'shc1de1d94, 32'shc1dd5cc8, 32'shc1dc9c23, 32'shc1dbdba3, 32'shc1db1b4a, 32'shc1da5b17, 32'shc1d99b0b, 
               32'shc1d8db25, 32'shc1d81b65, 32'shc1d75bcb, 32'shc1d69c58, 32'shc1d5dd0c, 32'shc1d51de5, 32'shc1d45ee5, 32'shc1d3a00b, 
               32'shc1d2e158, 32'shc1d222cb, 32'shc1d16464, 32'shc1d0a624, 32'shc1cfe80a, 32'shc1cf2a17, 32'shc1ce6c49, 32'shc1cdaea3, 
               32'shc1ccf122, 32'shc1cc33c8, 32'shc1cb7694, 32'shc1cab987, 32'shc1c9fca0, 32'shc1c93fdf, 32'shc1c88345, 32'shc1c7c6d1, 
               32'shc1c70a84, 32'shc1c64e5d, 32'shc1c5925c, 32'shc1c4d682, 32'shc1c41ace, 32'shc1c35f40, 32'shc1c2a3d9, 32'shc1c1e898, 
               32'shc1c12d7e, 32'shc1c0728a, 32'shc1bfb7bc, 32'shc1befd15, 32'shc1be4294, 32'shc1bd883a, 32'shc1bcce06, 32'shc1bc13f8, 
               32'shc1bb5a11, 32'shc1baa050, 32'shc1b9e6b6, 32'shc1b92d42, 32'shc1b873f5, 32'shc1b7bacd, 32'shc1b701cd, 32'shc1b648f3, 
               32'shc1b5903f, 32'shc1b4d7b1, 32'shc1b41f4a, 32'shc1b3670a, 32'shc1b2aef0, 32'shc1b1f6fc, 32'shc1b13f2f, 32'shc1b08788, 
               32'shc1afd007, 32'shc1af18ae, 32'shc1ae617a, 32'shc1adaa6d, 32'shc1acf386, 32'shc1ac3cc6, 32'shc1ab862c, 32'shc1aacfb9, 
               32'shc1aa196c, 32'shc1a96346, 32'shc1a8ad46, 32'shc1a7f76c, 32'shc1a741b9, 32'shc1a68c2d, 32'shc1a5d6c7, 32'shc1a52187, 
               32'shc1a46c6e, 32'shc1a3b77b, 32'shc1a302af, 32'shc1a24e09, 32'shc1a1998a, 32'shc1a0e531, 32'shc1a030ff, 32'shc19f7cf3, 
               32'shc19ec90d, 32'shc19e154e, 32'shc19d61b6, 32'shc19cae44, 32'shc19bfaf9, 32'shc19b47d4, 32'shc19a94d5, 32'shc199e1fd, 
               32'shc1992f4c, 32'shc1987cc1, 32'shc197ca5c, 32'shc197181e, 32'shc1966606, 32'shc195b415, 32'shc195024b, 32'shc19450a7, 
               32'shc1939f29, 32'shc192edd2, 32'shc1923ca2, 32'shc1918b98, 32'shc190dab4, 32'shc19029f7, 32'shc18f7961, 32'shc18ec8f1, 
               32'shc18e18a7, 32'shc18d6884, 32'shc18cb888, 32'shc18c08b2, 32'shc18b5903, 32'shc18aa97a, 32'shc189fa17, 32'shc1894adc, 
               32'shc1889bc6, 32'shc187ecd8, 32'shc1873e10, 32'shc1868f6e, 32'shc185e0f3, 32'shc185329e, 32'shc1848470, 32'shc183d669, 
               32'shc1832888, 32'shc1827acd, 32'shc181cd3a, 32'shc1811fcc, 32'shc1807285, 32'shc17fc565, 32'shc17f186c, 32'shc17e6b99, 
               32'shc17dbeec, 32'shc17d1266, 32'shc17c6607, 32'shc17bb9ce, 32'shc17b0dbb, 32'shc17a61d0, 32'shc179b60b, 32'shc1790a6c, 
               32'shc1785ef4, 32'shc177b3a3, 32'shc1770878, 32'shc1765d73, 32'shc175b296, 32'shc17507df, 32'shc1745d4e, 32'shc173b2e4, 
               32'shc17308a1, 32'shc1725e84, 32'shc171b48e, 32'shc1710abe, 32'shc1706115, 32'shc16fb792, 32'shc16f0e36, 32'shc16e6501, 
               32'shc16dbbf3, 32'shc16d130a, 32'shc16c6a49, 32'shc16bc1ae, 32'shc16b193a, 32'shc16a70ec, 32'shc169c8c5, 32'shc16920c5, 
               32'shc16878eb, 32'shc167d137, 32'shc16729ab, 32'shc1668245, 32'shc165db05, 32'shc16533ed, 32'shc1648cfa, 32'shc163e62f, 
               32'shc1633f8a, 32'shc162990c, 32'shc161f2b4, 32'shc1614c83, 32'shc160a678, 32'shc1600095, 32'shc15f5ad7, 32'shc15eb541, 
               32'shc15e0fd1, 32'shc15d6a88, 32'shc15cc565, 32'shc15c2069, 32'shc15b7b94, 32'shc15ad6e5, 32'shc15a325d, 32'shc1598dfb, 
               32'shc158e9c1, 32'shc15845ac, 32'shc157a1bf, 32'shc156fdf8, 32'shc1565a58, 32'shc155b6de, 32'shc155138c, 32'shc154705f, 
               32'shc153cd5a, 32'shc1532a7b, 32'shc15287c3, 32'shc151e531, 32'shc15142c6, 32'shc150a082, 32'shc14ffe64, 32'shc14f5c6d, 
               32'shc14eba9d, 32'shc14e18f3, 32'shc14d7771, 32'shc14cd614, 32'shc14c34df, 32'shc14b93d0, 32'shc14af2e8, 32'shc14a5226, 
               32'shc149b18b, 32'shc1491117, 32'shc14870ca, 32'shc147d0a3, 32'shc14730a3, 32'shc14690ca, 32'shc145f117, 32'shc145518b, 
               32'shc144b225, 32'shc14412e7, 32'shc14373cf, 32'shc142d4de, 32'shc1423613, 32'shc141976f, 32'shc140f8f2, 32'shc1405a9c, 
               32'shc13fbc6c, 32'shc13f1e63, 32'shc13e8081, 32'shc13de2c5, 32'shc13d4530, 32'shc13ca7c2, 32'shc13c0a7b, 32'shc13b6d5a, 
               32'shc13ad060, 32'shc13a338d, 32'shc13996e0, 32'shc138fa5a, 32'shc1385dfb, 32'shc137c1c3, 32'shc13725b1, 32'shc13689c6, 
               32'shc135ee02, 32'shc1355265, 32'shc134b6ee, 32'shc1341b9e, 32'shc1338075, 32'shc132e572, 32'shc1324a96, 32'shc131afe1, 
               32'shc1311553, 32'shc1307aeb, 32'shc12fe0ab, 32'shc12f4690, 32'shc12eac9d, 32'shc12e12d1, 32'shc12d792b, 32'shc12cdfac, 
               32'shc12c4653, 32'shc12bad22, 32'shc12b1417, 32'shc12a7b33, 32'shc129e276, 32'shc12949df, 32'shc128b16f, 32'shc1281926, 
               32'shc1278104, 32'shc126e909, 32'shc1265134, 32'shc125b986, 32'shc12521ff, 32'shc1248a9e, 32'shc123f365, 32'shc1235c52, 
               32'shc122c566, 32'shc1222ea1, 32'shc1219802, 32'shc121018a, 32'shc1206b39, 32'shc11fd50f, 32'shc11f3f0c, 32'shc11ea92f, 
               32'shc11e1379, 32'shc11d7dea, 32'shc11ce882, 32'shc11c5341, 32'shc11bbe26, 32'shc11b2932, 32'shc11a9465, 32'shc119ffbf, 
               32'shc1196b3f, 32'shc118d6e7, 32'shc11842b5, 32'shc117aeaa, 32'shc1171ac6, 32'shc1168708, 32'shc115f372, 32'shc1156002, 
               32'shc114ccb9, 32'shc1143997, 32'shc113a69b, 32'shc11313c7, 32'shc1128119, 32'shc111ee92, 32'shc1115c32, 32'shc110c9f8, 
               32'shc11037e6, 32'shc10fa5fa, 32'shc10f1435, 32'shc10e8297, 32'shc10df120, 32'shc10d5fd0, 32'shc10ccea6, 32'shc10c3da4, 
               32'shc10bacc8, 32'shc10b1c13, 32'shc10a8b85, 32'shc109fb1d, 32'shc1096add, 32'shc108dac3, 32'shc1084ad0, 32'shc107bb04, 
               32'shc1072b5f, 32'shc1069be1, 32'shc1060c89, 32'shc1057d59, 32'shc104ee4f, 32'shc1045f6c, 32'shc103d0b0, 32'shc103421b, 
               32'shc102b3ac, 32'shc1022565, 32'shc1019744, 32'shc101094a, 32'shc1007b77, 32'shc0ffedcb, 32'shc0ff6046, 32'shc0fed2e8, 
               32'shc0fe45b0, 32'shc0fdb8a0, 32'shc0fd2bb6, 32'shc0fc9ef3, 32'shc0fc1257, 32'shc0fb85e2, 32'shc0faf993, 32'shc0fa6d6c, 
               32'shc0f9e16b, 32'shc0f95592, 32'shc0f8c9df, 32'shc0f83e53, 32'shc0f7b2ee, 32'shc0f727b0, 32'shc0f69c99, 32'shc0f611a8, 
               32'shc0f586df, 32'shc0f4fc3c, 32'shc0f471c1, 32'shc0f3e76c, 32'shc0f35d3e, 32'shc0f2d337, 32'shc0f24957, 32'shc0f1bf9d, 
               32'shc0f1360b, 32'shc0f0aca0, 32'shc0f0235b, 32'shc0ef9a3d, 32'shc0ef1147, 32'shc0ee8877, 32'shc0edffce, 32'shc0ed774c, 
               32'shc0eceef1, 32'shc0ec66bc, 32'shc0ebdeaf, 32'shc0eb56c9, 32'shc0eacf09, 32'shc0ea4771, 32'shc0e9bfff, 32'shc0e938b4, 
               32'shc0e8b190, 32'shc0e82a93, 32'shc0e7a3bd, 32'shc0e71d0e, 32'shc0e69686, 32'shc0e61025, 32'shc0e589eb, 32'shc0e503d7, 
               32'shc0e47deb, 32'shc0e3f825, 32'shc0e37287, 32'shc0e2ed0f, 32'shc0e267be, 32'shc0e1e294, 32'shc0e15d92, 32'shc0e0d8b6, 
               32'shc0e05401, 32'shc0dfcf73, 32'shc0df4b0b, 32'shc0dec6cb, 32'shc0de42b2, 32'shc0ddbec0, 32'shc0dd3af4, 32'shc0dcb750, 
               32'shc0dc33d2, 32'shc0dbb07c, 32'shc0db2d4c, 32'shc0daaa44, 32'shc0da2762, 32'shc0d9a4a7, 32'shc0d92214, 32'shc0d89fa7, 
               32'shc0d81d61, 32'shc0d79b42, 32'shc0d7194a, 32'shc0d69779, 32'shc0d615cf, 32'shc0d5944c, 32'shc0d512f0, 32'shc0d491bb, 
               32'shc0d410ad, 32'shc0d38fc6, 32'shc0d30f05, 32'shc0d28e6c, 32'shc0d20dfa, 32'shc0d18dae, 32'shc0d10d8a, 32'shc0d08d8d, 
               32'shc0d00db6, 32'shc0cf8e07, 32'shc0cf0e7f, 32'shc0ce8f1d, 32'shc0ce0fe3, 32'shc0cd90cf, 32'shc0cd11e3, 32'shc0cc931d, 
               32'shc0cc147f, 32'shc0cb9607, 32'shc0cb17b7, 32'shc0ca998d, 32'shc0ca1b8a, 32'shc0c99daf, 32'shc0c91ffa, 32'shc0c8a26d, 
               32'shc0c82506, 32'shc0c7a7c6, 32'shc0c72aae, 32'shc0c6adbc, 32'shc0c630f2, 32'shc0c5b44e, 32'shc0c537d1, 32'shc0c4bb7c, 
               32'shc0c43f4d, 32'shc0c3c346, 32'shc0c34765, 32'shc0c2cbab, 32'shc0c25019, 32'shc0c1d4ad, 32'shc0c15969, 32'shc0c0de4b, 
               32'shc0c06355, 32'shc0bfe885, 32'shc0bf6ddd, 32'shc0bef35b, 32'shc0be7901, 32'shc0bdfecd, 32'shc0bd84c1, 32'shc0bd0adb, 
               32'shc0bc911d, 32'shc0bc1786, 32'shc0bb9e15, 32'shc0bb24cc, 32'shc0baabaa, 32'shc0ba32af, 32'shc0b9b9da, 32'shc0b9412d, 
               32'shc0b8c8a7, 32'shc0b85048, 32'shc0b7d810, 32'shc0b75fff, 32'shc0b6e815, 32'shc0b67052, 32'shc0b5f8b6, 32'shc0b58141, 
               32'shc0b509f3, 32'shc0b492cc, 32'shc0b41bcd, 32'shc0b3a4f4, 32'shc0b32e42, 32'shc0b2b7b8, 32'shc0b24154, 32'shc0b1cb17, 
               32'shc0b15502, 32'shc0b0df13, 32'shc0b0694c, 32'shc0aff3ac, 32'shc0af7e33, 32'shc0af08e0, 32'shc0ae93b5, 32'shc0ae1eb1, 
               32'shc0ada9d4, 32'shc0ad351e, 32'shc0acc08f, 32'shc0ac4c27, 32'shc0abd7e6, 32'shc0ab63cd, 32'shc0aaefda, 32'shc0aa7c0e, 
               32'shc0aa086a, 32'shc0a994ec, 32'shc0a92196, 32'shc0a8ae67, 32'shc0a83b5e, 32'shc0a7c87d, 32'shc0a755c3, 32'shc0a6e330, 
               32'shc0a670c4, 32'shc0a5fe7f, 32'shc0a58c62, 32'shc0a51a6b, 32'shc0a4a89b, 32'shc0a436f3, 32'shc0a3c571, 32'shc0a35417, 
               32'shc0a2e2e3, 32'shc0a271d7, 32'shc0a200f2, 32'shc0a19034, 32'shc0a11f9d, 32'shc0a0af2d, 32'shc0a03ee4, 32'shc09fcec3, 
               32'shc09f5ec8, 32'shc09eeef5, 32'shc09e7f48, 32'shc09e0fc3, 32'shc09da065, 32'shc09d312e, 32'shc09cc21e, 32'shc09c5335, 
               32'shc09be473, 32'shc09b75d8, 32'shc09b0765, 32'shc09a9918, 32'shc09a2af3, 32'shc099bcf5, 32'shc0994f1d, 32'shc098e16d, 
               32'shc09873e4, 32'shc0980683, 32'shc0979948, 32'shc0972c34, 32'shc096bf48, 32'shc0965282, 32'shc095e5e4, 32'shc095796d, 
               32'shc0950d1d, 32'shc094a0f4, 32'shc09434f2, 32'shc093c917, 32'shc0935d64, 32'shc092f1d7, 32'shc0928672, 32'shc0921b34, 
               32'shc091b01d, 32'shc091452d, 32'shc090da64, 32'shc0906fc3, 32'shc0900548, 32'shc08f9af5, 32'shc08f30c8, 32'shc08ec6c3, 
               32'shc08e5ce5, 32'shc08df32e, 32'shc08d899f, 32'shc08d2036, 32'shc08cb6f5, 32'shc08c4dda, 32'shc08be4e7, 32'shc08b7c1b, 
               32'shc08b1376, 32'shc08aaaf8, 32'shc08a42a2, 32'shc089da72, 32'shc089726a, 32'shc0890a89, 32'shc088a2cf, 32'shc0883b3c, 
               32'shc087d3d0, 32'shc0876c8c, 32'shc087056e, 32'shc0869e78, 32'shc08637a9, 32'shc085d101, 32'shc0856a80, 32'shc0850426, 
               32'shc0849df4, 32'shc08437e9, 32'shc083d204, 32'shc0836c47, 32'shc08306b2, 32'shc082a143, 32'shc0823bfb, 32'shc081d6db, 
               32'shc08171e2, 32'shc0810d10, 32'shc080a865, 32'shc08043e1, 32'shc07fdf85, 32'shc07f7b50, 32'shc07f1741, 32'shc07eb35a, 
               32'shc07e4f9b, 32'shc07dec02, 32'shc07d8890, 32'shc07d2546, 32'shc07cc223, 32'shc07c5f27, 32'shc07bfc52, 32'shc07b99a5, 
               32'shc07b371e, 32'shc07ad4bf, 32'shc07a7287, 32'shc07a1076, 32'shc079ae8c, 32'shc0794cca, 32'shc078eb2f, 32'shc07889bb, 
               32'shc078286e, 32'shc077c748, 32'shc0776649, 32'shc0770572, 32'shc076a4c2, 32'shc0764439, 32'shc075e3d7, 32'shc075839c, 
               32'shc0752389, 32'shc074c39d, 32'shc07463d8, 32'shc074043a, 32'shc073a4c3, 32'shc0734574, 32'shc072e64c, 32'shc072874b, 
               32'shc0722871, 32'shc071c9be, 32'shc0716b33, 32'shc0710ccf, 32'shc070ae92, 32'shc070507c, 32'shc06ff28e, 32'shc06f94c6, 
               32'shc06f3726, 32'shc06ed9ad, 32'shc06e7c5b, 32'shc06e1f31, 32'shc06dc22e, 32'shc06d6551, 32'shc06d089d, 32'shc06cac0f, 
               32'shc06c4fa8, 32'shc06bf369, 32'shc06b9751, 32'shc06b3b60, 32'shc06adf97, 32'shc06a83f5, 32'shc06a2879, 32'shc069cd26, 
               32'shc06971f9, 32'shc06916f3, 32'shc068bc15, 32'shc068615e, 32'shc06806ce, 32'shc067ac66, 32'shc0675225, 32'shc066f80a, 
               32'shc0669e18, 32'shc066444c, 32'shc065eaa8, 32'shc065912a, 32'shc06537d4, 32'shc064dea6, 32'shc064859e, 32'shc0642cbe, 
               32'shc063d405, 32'shc0637b73, 32'shc0632309, 32'shc062cac6, 32'shc06272aa, 32'shc0621ab5, 32'shc061c2e7, 32'shc0616b41, 
               32'shc06113c2, 32'shc060bc6a, 32'shc060653a, 32'shc0600e30, 32'shc05fb74e, 32'shc05f6093, 32'shc05f0a00, 32'shc05eb393, 
               32'shc05e5d4e, 32'shc05e0730, 32'shc05db13a, 32'shc05d5b6b, 32'shc05d05c3, 32'shc05cb042, 32'shc05c5ae8, 32'shc05c05b6, 
               32'shc05bb0ab, 32'shc05b5bc7, 32'shc05b070a, 32'shc05ab275, 32'shc05a5e07, 32'shc05a09c0, 32'shc059b5a1, 32'shc05961a9, 
               32'shc0590dd8, 32'shc058ba2e, 32'shc05866ac, 32'shc0581350, 32'shc057c01d, 32'shc0576d10, 32'shc0571a2b, 32'shc056c76c, 
               32'shc05674d6, 32'shc0562266, 32'shc055d01e, 32'shc0557dfd, 32'shc0552c03, 32'shc054da30, 32'shc0548885, 32'shc0543701, 
               32'shc053e5a5, 32'shc053946f, 32'shc0534361, 32'shc052f27a, 32'shc052a1bb, 32'shc0525123, 32'shc05200b2, 32'shc051b068, 
               32'shc0516045, 32'shc051104a, 32'shc050c077, 32'shc05070ca, 32'shc0502145, 32'shc04fd1e7, 32'shc04f82b0, 32'shc04f33a1, 
               32'shc04ee4b8, 32'shc04e95f8, 32'shc04e475e, 32'shc04df8ec, 32'shc04daaa1, 32'shc04d5c7d, 32'shc04d0e81, 32'shc04cc0ac, 
               32'shc04c72fe, 32'shc04c2577, 32'shc04bd818, 32'shc04b8ae0, 32'shc04b3dcf, 32'shc04af0e6, 32'shc04aa424, 32'shc04a5789, 
               32'shc04a0b16, 32'shc049beca, 32'shc04972a5, 32'shc04926a7, 32'shc048dad1, 32'shc0488f22, 32'shc048439b, 32'shc047f83a, 
               32'shc047ad01, 32'shc04761ef, 32'shc0471705, 32'shc046cc42, 32'shc04681a6, 32'shc0463732, 32'shc045ece5, 32'shc045a2bf, 
               32'shc04558c0, 32'shc0450ee9, 32'shc044c539, 32'shc0447bb0, 32'shc044324f, 32'shc043e915, 32'shc043a002, 32'shc0435717, 
               32'shc0430e53, 32'shc042c5b6, 32'shc0427d41, 32'shc04234f3, 32'shc041eccc, 32'shc041a4cd, 32'shc0415cf4, 32'shc0411544, 
               32'shc040cdba, 32'shc0408658, 32'shc0403f1d, 32'shc03ff80a, 32'shc03fb11d, 32'shc03f6a58, 32'shc03f23bb, 32'shc03edd45, 
               32'shc03e96f6, 32'shc03e50ce, 32'shc03e0ace, 32'shc03dc4f5, 32'shc03d7f44, 32'shc03d39b9, 32'shc03cf456, 32'shc03caf1b, 
               32'shc03c6a07, 32'shc03c251a, 32'shc03be054, 32'shc03b9bb6, 32'shc03b573f, 32'shc03b12ef, 32'shc03acec7, 32'shc03a8ac6, 
               32'shc03a46ed, 32'shc03a033a, 32'shc039bfaf, 32'shc0397c4c, 32'shc0393910, 32'shc038f5fb, 32'shc038b30d, 32'shc0387047, 
               32'shc0382da8, 32'shc037eb31, 32'shc037a8e1, 32'shc03766b8, 32'shc03724b6, 32'shc036e2dc, 32'shc036a129, 32'shc0365f9e, 
               32'shc0361e3a, 32'shc035dcfd, 32'shc0359be8, 32'shc0355afa, 32'shc0351a33, 32'shc034d994, 32'shc034991c, 32'shc03458cb, 
               32'shc03418a2, 32'shc033d8a0, 32'shc03398c5, 32'shc0335912, 32'shc0331986, 32'shc032da22, 32'shc0329ae4, 32'shc0325bcf, 
               32'shc0321ce0, 32'shc031de19, 32'shc0319f79, 32'shc0316101, 32'shc03122b0, 32'shc030e486, 32'shc030a684, 32'shc03068a9, 
               32'shc0302af5, 32'shc02fed69, 32'shc02fb004, 32'shc02f72c7, 32'shc02f35b1, 32'shc02ef8c2, 32'shc02ebbfb, 32'shc02e7f5b, 
               32'shc02e42e2, 32'shc02e0691, 32'shc02dca67, 32'shc02d8e64, 32'shc02d5289, 32'shc02d16d5, 32'shc02cdb49, 32'shc02c9fe4, 
               32'shc02c64a6, 32'shc02c2990, 32'shc02beea1, 32'shc02bb3d9, 32'shc02b7939, 32'shc02b3ec0, 32'shc02b046f, 32'shc02aca44, 
               32'shc02a9042, 32'shc02a5666, 32'shc02a1cb2, 32'shc029e326, 32'shc029a9c1, 32'shc0297083, 32'shc029376c, 32'shc028fe7d, 
               32'shc028c5b6, 32'shc0288d15, 32'shc028549c, 32'shc0281c4b, 32'shc027e421, 32'shc027ac1e, 32'shc0277442, 32'shc0273c8e, 
               32'shc0270502, 32'shc026cd9d, 32'shc026965f, 32'shc0265f48, 32'shc0262859, 32'shc025f191, 32'shc025baf1, 32'shc0258478, 
               32'shc0254e27, 32'shc02517fc, 32'shc024e1fa, 32'shc024ac1e, 32'shc024766a, 32'shc02440de, 32'shc0240b78, 32'shc023d63b, 
               32'shc023a124, 32'shc0236c35, 32'shc023376e, 32'shc02302cd, 32'shc022ce54, 32'shc0229a03, 32'shc02265d9, 32'shc02231d6, 
               32'shc021fdfb, 32'shc021ca47, 32'shc02196bb, 32'shc0216356, 32'shc0213018, 32'shc020fd02, 32'shc020ca13, 32'shc020974b, 
               32'shc02064ab, 32'shc0203232, 32'shc01fffe1, 32'shc01fcdb7, 32'shc01f9bb5, 32'shc01f69da, 32'shc01f3826, 32'shc01f069a, 
               32'shc01ed535, 32'shc01ea3f7, 32'shc01e72e1, 32'shc01e41f3, 32'shc01e112b, 32'shc01de08c, 32'shc01db013, 32'shc01d7fc2, 
               32'shc01d4f99, 32'shc01d1f96, 32'shc01cefbb, 32'shc01cc008, 32'shc01c907c, 32'shc01c6118, 32'shc01c31da, 32'shc01c02c5, 
               32'shc01bd3d6, 32'shc01ba50f, 32'shc01b7670, 32'shc01b47f8, 32'shc01b19a7, 32'shc01aeb7e, 32'shc01abd7c, 32'shc01a8fa1, 
               32'shc01a61ee, 32'shc01a3463, 32'shc01a06fe, 32'shc019d9c2, 32'shc019acac, 32'shc0197fbe, 32'shc01952f8, 32'shc0192659, 
               32'shc018f9e1, 32'shc018cd91, 32'shc018a168, 32'shc0187566, 32'shc018498c, 32'shc0181dda, 32'shc017f24e, 32'shc017c6eb, 
               32'shc0179bae, 32'shc0177099, 32'shc01745ac, 32'shc0171ae6, 32'shc016f047, 32'shc016c5d0, 32'shc0169b80, 32'shc0167158, 
               32'shc0164757, 32'shc0161d7d, 32'shc015f3cb, 32'shc015ca40, 32'shc015a0dd, 32'shc01577a1, 32'shc0154e8d, 32'shc01525a0, 
               32'shc014fcda, 32'shc014d43c, 32'shc014abc5, 32'shc0148376, 32'shc0145b4e, 32'shc014334e, 32'shc0140b75, 32'shc013e3c3, 
               32'shc013bc39, 32'shc01394d6, 32'shc0136d9b, 32'shc0134687, 32'shc0131f9b, 32'shc012f8d6, 32'shc012d238, 32'shc012abc2, 
               32'shc0128574, 32'shc0125f4c, 32'shc012394c, 32'shc0121374, 32'shc011edc3, 32'shc011c83a, 32'shc011a2d8, 32'shc0117d9d, 
               32'shc011588a, 32'shc011339e, 32'shc0110eda, 32'shc010ea3d, 32'shc010c5c7, 32'shc010a179, 32'shc0107d53, 32'shc0105954, 
               32'shc010357c, 32'shc01011cc, 32'shc00fee43, 32'shc00fcae2, 32'shc00fa7a8, 32'shc00f8495, 32'shc00f61aa, 32'shc00f3ee6, 
               32'shc00f1c4a, 32'shc00ef9d6, 32'shc00ed788, 32'shc00eb562, 32'shc00e9364, 32'shc00e718d, 32'shc00e4fde, 32'shc00e2e56, 
               32'shc00e0cf5, 32'shc00debbc, 32'shc00dcaaa, 32'shc00da9c0, 32'shc00d88fd, 32'shc00d6861, 32'shc00d47ed, 32'shc00d27a1, 
               32'shc00d077c, 32'shc00ce77e, 32'shc00cc7a8, 32'shc00ca7f9, 32'shc00c8872, 32'shc00c6912, 32'shc00c49da, 32'shc00c2ac9, 
               32'shc00c0be0, 32'shc00bed1e, 32'shc00bce83, 32'shc00bb010, 32'shc00b91c4, 32'shc00b73a0, 32'shc00b55a3, 32'shc00b37ce, 
               32'shc00b1a20, 32'shc00afc9a, 32'shc00adf3b, 32'shc00ac203, 32'shc00aa4f3, 32'shc00a880a, 32'shc00a6b49, 32'shc00a4eb0, 
               32'shc00a323d, 32'shc00a15f3, 32'shc009f9cf, 32'shc009ddd3, 32'shc009c1ff, 32'shc009a652, 32'shc0098acc, 32'shc0096f6e, 
               32'shc0095438, 32'shc0093929, 32'shc0091e41, 32'shc0090381, 32'shc008e8e8, 32'shc008ce76, 32'shc008b42d, 32'shc0089a0a, 
               32'shc008800f, 32'shc008663c, 32'shc0084c90, 32'shc008330b, 32'shc00819ae, 32'shc0080078, 32'shc007e76a, 32'shc007ce83, 
               32'shc007b5c4, 32'shc0079d2c, 32'shc00784bc, 32'shc0076c73, 32'shc0075452, 32'shc0073c58, 32'shc0072485, 32'shc0070cda, 
               32'shc006f556, 32'shc006ddfa, 32'shc006c6c6, 32'shc006afb8, 32'shc00698d3, 32'shc0068214, 32'shc0066b7d, 32'shc006550e, 
               32'shc0063ec6, 32'shc00628a6, 32'shc00612ad, 32'shc005fcdb, 32'shc005e731, 32'shc005d1af, 32'shc005bc54, 32'shc005a720, 
               32'shc0059214, 32'shc0057d2f, 32'shc0056872, 32'shc00553dc, 32'shc0053f6e, 32'shc0052b27, 32'shc0051707, 32'shc005030f, 
               32'shc004ef3f, 32'shc004db96, 32'shc004c814, 32'shc004b4ba, 32'shc004a188, 32'shc0048e7d, 32'shc0047b99, 32'shc00468dd, 
               32'shc0045648, 32'shc00443db, 32'shc0043195, 32'shc0041f77, 32'shc0040d80, 32'shc003fbb0, 32'shc003ea09, 32'shc003d888, 
               32'shc003c72f, 32'shc003b5fe, 32'shc003a4f4, 32'shc0039411, 32'shc0038356, 32'shc00372c2, 32'shc0036256, 32'shc0035211, 
               32'shc00341f4, 32'shc00331fe, 32'shc0032230, 32'shc0031289, 32'shc003030a, 32'shc002f3b2, 32'shc002e482, 32'shc002d579, 
               32'shc002c697, 32'shc002b7dd, 32'shc002a94b, 32'shc0029ae0, 32'shc0028c9c, 32'shc0027e80, 32'shc002708c, 32'shc00262be, 
               32'shc0025519, 32'shc002479b, 32'shc0023a44, 32'shc0022d15, 32'shc002200d, 32'shc002132d, 32'shc0020674, 32'shc001f9e2, 
               32'shc001ed78, 32'shc001e136, 32'shc001d51b, 32'shc001c928, 32'shc001bd5c, 32'shc001b1b7, 32'shc001a63a, 32'shc0019ae5, 
               32'shc0018fb6, 32'shc00184b0, 32'shc00179d1, 32'shc0016f19, 32'shc0016489, 32'shc0015a20, 32'shc0014fdf, 32'shc00145c5, 
               32'shc0013bd3, 32'shc0013208, 32'shc0012865, 32'shc0011ee9, 32'shc0011594, 32'shc0010c67, 32'shc0010362, 32'shc000fa84, 
               32'shc000f1ce, 32'shc000e93f, 32'shc000e0d7, 32'shc000d897, 32'shc000d07e, 32'shc000c88d, 32'shc000c0c4, 32'shc000b921, 
               32'shc000b1a7, 32'shc000aa54, 32'shc000a328, 32'shc0009c24, 32'shc0009547, 32'shc0008e92, 32'shc0008804, 32'shc000819d, 
               32'shc0007b5f, 32'shc0007547, 32'shc0006f57, 32'shc000698f, 32'shc00063ee, 32'shc0005e74, 32'shc0005922, 32'shc00053f8, 
               32'shc0004ef5, 32'shc0004a19, 32'shc0004565, 32'shc00040d9, 32'shc0003c74, 32'shc0003836, 32'shc0003420, 32'shc0003031, 
               32'shc0002c6a, 32'shc00028ca, 32'shc0002552, 32'shc0002201, 32'shc0001ed8, 32'shc0001bd6, 32'shc00018fb, 32'shc0001649, 
               32'shc00013bd, 32'shc0001159, 32'shc0000f1d, 32'shc0000d08, 32'shc0000b1a, 32'shc0000954, 32'shc00007b6, 32'shc000063f, 
               32'shc00004ef, 32'shc00003c7, 32'shc00002c7, 32'shc00001ed, 32'shc000013c, 32'shc00000b2, 32'shc000004f, 32'shc0000014
            };

            reg signed [31:0] W_Im_table[16384] = '{
               32'sh00000000, 32'shfffcdbc1, 32'shfff9b781, 32'shfff69342, 32'shfff36f02, 32'shfff04ac3, 32'shffed2684, 32'shffea0245, 
               32'shffe6de05, 32'shffe3b9c6, 32'shffe09587, 32'shffdd7148, 32'shffda4d09, 32'shffd728ca, 32'shffd4048c, 32'shffd0e04d, 
               32'shffcdbc0f, 32'shffca97d0, 32'shffc77392, 32'shffc44f54, 32'shffc12b16, 32'shffbe06d8, 32'shffbae29a, 32'shffb7be5d, 
               32'shffb49a1f, 32'shffb175e2, 32'shffae51a5, 32'shffab2d69, 32'shffa8092c, 32'shffa4e4f0, 32'shffa1c0b4, 32'shff9e9c78, 
               32'shff9b783c, 32'shff985401, 32'shff952fc5, 32'shff920b8b, 32'shff8ee750, 32'shff8bc316, 32'shff889edb, 32'shff857aa2, 
               32'shff825668, 32'shff7f322f, 32'shff7c0df6, 32'shff78e9bd, 32'shff75c585, 32'shff72a14d, 32'shff6f7d16, 32'shff6c58de, 
               32'shff6934a8, 32'shff661071, 32'shff62ec3b, 32'shff5fc805, 32'shff5ca3d0, 32'shff597f9b, 32'shff565b66, 32'shff533732, 
               32'shff5012fe, 32'shff4ceecb, 32'shff49ca98, 32'shff46a666, 32'shff438234, 32'shff405e02, 32'shff3d39d1, 32'shff3a15a0, 
               32'shff36f170, 32'shff33cd40, 32'shff30a911, 32'shff2d84e3, 32'shff2a60b4, 32'shff273c87, 32'shff24185a, 32'shff20f42d, 
               32'shff1dd001, 32'shff1aabd5, 32'shff1787aa, 32'shff146380, 32'shff113f56, 32'shff0e1b2d, 32'shff0af704, 32'shff07d2dc, 
               32'shff04aeb5, 32'shff018a8e, 32'shfefe6668, 32'shfefb4242, 32'shfef81e1d, 32'shfef4f9f8, 32'shfef1d5d5, 32'shfeeeb1b2, 
               32'shfeeb8d8f, 32'shfee8696d, 32'shfee5454c, 32'shfee2212c, 32'shfedefd0c, 32'shfedbd8ed, 32'shfed8b4cf, 32'shfed590b1, 
               32'shfed26c94, 32'shfecf4878, 32'shfecc245d, 32'shfec90042, 32'shfec5dc28, 32'shfec2b80f, 32'shfebf93f6, 32'shfebc6fdf, 
               32'shfeb94bc8, 32'shfeb627b2, 32'shfeb3039d, 32'shfeafdf88, 32'shfeacbb74, 32'shfea99761, 32'shfea6734f, 32'shfea34f3e, 
               32'shfea02b2e, 32'shfe9d071e, 32'shfe99e310, 32'shfe96bf02, 32'shfe939af5, 32'shfe9076e9, 32'shfe8d52de, 32'shfe8a2ed4, 
               32'shfe870aca, 32'shfe83e6c2, 32'shfe80c2ba, 32'shfe7d9eb4, 32'shfe7a7aae, 32'shfe7756a9, 32'shfe7432a5, 32'shfe710ea2, 
               32'shfe6deaa1, 32'shfe6ac6a0, 32'shfe67a2a0, 32'shfe647ea1, 32'shfe615aa3, 32'shfe5e36a6, 32'shfe5b12aa, 32'shfe57eeaf, 
               32'shfe54cab5, 32'shfe51a6bc, 32'shfe4e82c4, 32'shfe4b5ecd, 32'shfe483ad8, 32'shfe4516e3, 32'shfe41f2ef, 32'shfe3ecefd, 
               32'shfe3bab0b, 32'shfe38871b, 32'shfe35632c, 32'shfe323f3d, 32'shfe2f1b50, 32'shfe2bf764, 32'shfe28d379, 32'shfe25af90, 
               32'shfe228ba7, 32'shfe1f67c0, 32'shfe1c43da, 32'shfe191ff5, 32'shfe15fc11, 32'shfe12d82e, 32'shfe0fb44c, 32'shfe0c906c, 
               32'shfe096c8d, 32'shfe0648af, 32'shfe0324d2, 32'shfe0000f7, 32'shfdfcdd1d, 32'shfdf9b944, 32'shfdf6956c, 32'shfdf37195, 
               32'shfdf04dc0, 32'shfded29ec, 32'shfdea0619, 32'shfde6e248, 32'shfde3be78, 32'shfde09aa9, 32'shfddd76dc, 32'shfdda530f, 
               32'shfdd72f45, 32'shfdd40b7b, 32'shfdd0e7b3, 32'shfdcdc3ec, 32'shfdcaa027, 32'shfdc77c62, 32'shfdc458a0, 32'shfdc134de, 
               32'shfdbe111e, 32'shfdbaed60, 32'shfdb7c9a3, 32'shfdb4a5e7, 32'shfdb1822c, 32'shfdae5e74, 32'shfdab3abc, 32'shfda81706, 
               32'shfda4f351, 32'shfda1cf9e, 32'shfd9eabec, 32'shfd9b883c, 32'shfd98648d, 32'shfd9540e0, 32'shfd921d34, 32'shfd8ef98a, 
               32'shfd8bd5e1, 32'shfd88b23a, 32'shfd858e94, 32'shfd826af0, 32'shfd7f474d, 32'shfd7c23ac, 32'shfd79000d, 32'shfd75dc6e, 
               32'shfd72b8d2, 32'shfd6f9537, 32'shfd6c719e, 32'shfd694e06, 32'shfd662a70, 32'shfd6306db, 32'shfd5fe348, 32'shfd5cbfb7, 
               32'shfd599c28, 32'shfd56789a, 32'shfd53550d, 32'shfd503182, 32'shfd4d0df9, 32'shfd49ea72, 32'shfd46c6ec, 32'shfd43a368, 
               32'shfd407fe6, 32'shfd3d5c65, 32'shfd3a38e6, 32'shfd371569, 32'shfd33f1ed, 32'shfd30ce73, 32'shfd2daafb, 32'shfd2a8785, 
               32'shfd276410, 32'shfd24409d, 32'shfd211d2c, 32'shfd1df9bd, 32'shfd1ad650, 32'shfd17b2e4, 32'shfd148f7a, 32'shfd116c12, 
               32'shfd0e48ab, 32'shfd0b2547, 32'shfd0801e4, 32'shfd04de83, 32'shfd01bb24, 32'shfcfe97c7, 32'shfcfb746c, 32'shfcf85112, 
               32'shfcf52dbb, 32'shfcf20a65, 32'shfceee711, 32'shfcebc3bf, 32'shfce8a06f, 32'shfce57d21, 32'shfce259d5, 32'shfcdf368a, 
               32'shfcdc1342, 32'shfcd8effb, 32'shfcd5ccb7, 32'shfcd2a974, 32'shfccf8634, 32'shfccc62f5, 32'shfcc93fb9, 32'shfcc61c7e, 
               32'shfcc2f945, 32'shfcbfd60e, 32'shfcbcb2da, 32'shfcb98fa7, 32'shfcb66c77, 32'shfcb34948, 32'shfcb0261b, 32'shfcad02f1, 
               32'shfca9dfc8, 32'shfca6bca2, 32'shfca3997e, 32'shfca0765b, 32'shfc9d533b, 32'shfc9a301d, 32'shfc970d01, 32'shfc93e9e7, 
               32'shfc90c6cf, 32'shfc8da3ba, 32'shfc8a80a6, 32'shfc875d95, 32'shfc843a85, 32'shfc811778, 32'shfc7df46d, 32'shfc7ad164, 
               32'shfc77ae5e, 32'shfc748b59, 32'shfc716857, 32'shfc6e4557, 32'shfc6b2259, 32'shfc67ff5d, 32'shfc64dc64, 32'shfc61b96d, 
               32'shfc5e9678, 32'shfc5b7385, 32'shfc585094, 32'shfc552da6, 32'shfc520aba, 32'shfc4ee7d0, 32'shfc4bc4e9, 32'shfc48a204, 
               32'shfc457f21, 32'shfc425c40, 32'shfc3f3962, 32'shfc3c1686, 32'shfc38f3ac, 32'shfc35d0d5, 32'shfc32ae00, 32'shfc2f8b2e, 
               32'shfc2c685d, 32'shfc29458f, 32'shfc2622c4, 32'shfc22fffb, 32'shfc1fdd34, 32'shfc1cba6f, 32'shfc1997ae, 32'shfc1674ee, 
               32'shfc135231, 32'shfc102f76, 32'shfc0d0cbe, 32'shfc09ea08, 32'shfc06c754, 32'shfc03a4a3, 32'shfc0081f5, 32'shfbfd5f49, 
               32'shfbfa3c9f, 32'shfbf719f8, 32'shfbf3f753, 32'shfbf0d4b1, 32'shfbedb212, 32'shfbea8f75, 32'shfbe76cda, 32'shfbe44a42, 
               32'shfbe127ac, 32'shfbde0519, 32'shfbdae289, 32'shfbd7bffb, 32'shfbd49d70, 32'shfbd17ae7, 32'shfbce5861, 32'shfbcb35dd, 
               32'shfbc8135c, 32'shfbc4f0de, 32'shfbc1ce62, 32'shfbbeabe9, 32'shfbbb8973, 32'shfbb866ff, 32'shfbb5448d, 32'shfbb2221f, 
               32'shfbaeffb3, 32'shfbabdd49, 32'shfba8bae3, 32'shfba5987f, 32'shfba2761e, 32'shfb9f53bf, 32'shfb9c3163, 32'shfb990f0a, 
               32'shfb95ecb4, 32'shfb92ca60, 32'shfb8fa80f, 32'shfb8c85c1, 32'shfb896375, 32'shfb86412c, 32'shfb831ee6, 32'shfb7ffca3, 
               32'shfb7cda63, 32'shfb79b825, 32'shfb7695ea, 32'shfb7373b2, 32'shfb70517d, 32'shfb6d2f4a, 32'shfb6a0d1b, 32'shfb66eaee, 
               32'shfb63c8c4, 32'shfb60a69d, 32'shfb5d8479, 32'shfb5a6257, 32'shfb574039, 32'shfb541e1d, 32'shfb50fc04, 32'shfb4dd9ee, 
               32'shfb4ab7db, 32'shfb4795cb, 32'shfb4473be, 32'shfb4151b4, 32'shfb3e2fac, 32'shfb3b0da8, 32'shfb37eba7, 32'shfb34c9a8, 
               32'shfb31a7ac, 32'shfb2e85b4, 32'shfb2b63be, 32'shfb2841cc, 32'shfb251fdc, 32'shfb21fdef, 32'shfb1edc06, 32'shfb1bba1f, 
               32'shfb18983b, 32'shfb15765b, 32'shfb12547d, 32'shfb0f32a3, 32'shfb0c10cb, 32'shfb08eef7, 32'shfb05cd25, 32'shfb02ab57, 
               32'shfaff898c, 32'shfafc67c4, 32'shfaf945ff, 32'shfaf6243d, 32'shfaf3027e, 32'shfaefe0c2, 32'shfaecbf0a, 32'shfae99d54, 
               32'shfae67ba2, 32'shfae359f3, 32'shfae03847, 32'shfadd169e, 32'shfad9f4f8, 32'shfad6d355, 32'shfad3b1b6, 32'shfad0901a, 
               32'shfacd6e81, 32'shfaca4ceb, 32'shfac72b59, 32'shfac409c9, 32'shfac0e83d, 32'shfabdc6b4, 32'shfabaa52f, 32'shfab783ad, 
               32'shfab4622d, 32'shfab140b2, 32'shfaae1f39, 32'shfaaafdc4, 32'shfaa7dc52, 32'shfaa4bae3, 32'shfaa19978, 32'shfa9e7810, 
               32'shfa9b56ab, 32'shfa98354a, 32'shfa9513eb, 32'shfa91f291, 32'shfa8ed139, 32'shfa8bafe5, 32'shfa888e95, 32'shfa856d47, 
               32'shfa824bfd, 32'shfa7f2ab7, 32'shfa7c0974, 32'shfa78e834, 32'shfa75c6f8, 32'shfa72a5bf, 32'shfa6f8489, 32'shfa6c6357, 
               32'shfa694229, 32'shfa6620fd, 32'shfa62ffd6, 32'shfa5fdeb1, 32'shfa5cbd91, 32'shfa599c73, 32'shfa567b5a, 32'shfa535a43, 
               32'shfa503930, 32'shfa4d1821, 32'shfa49f715, 32'shfa46d60d, 32'shfa43b508, 32'shfa409407, 32'shfa3d7309, 32'shfa3a520f, 
               32'shfa373119, 32'shfa341026, 32'shfa30ef36, 32'shfa2dce4b, 32'shfa2aad62, 32'shfa278c7e, 32'shfa246b9d, 32'shfa214abf, 
               32'shfa1e29e5, 32'shfa1b090f, 32'shfa17e83d, 32'shfa14c76e, 32'shfa11a6a3, 32'shfa0e85db, 32'shfa0b6517, 32'shfa084457, 
               32'shfa05239a, 32'shfa0202e1, 32'shf9fee22c, 32'shf9fbc17b, 32'shf9f8a0cd, 32'shf9f58023, 32'shf9f25f7d, 32'shf9ef3eda, 
               32'shf9ec1e3b, 32'shf9e8fda0, 32'shf9e5dd09, 32'shf9e2bc75, 32'shf9df9be6, 32'shf9dc7b5a, 32'shf9d95ad1, 32'shf9d63a4d, 
               32'shf9d319cc, 32'shf9cff94f, 32'shf9ccd8d6, 32'shf9c9b861, 32'shf9c697f0, 32'shf9c37782, 32'shf9c05719, 32'shf9bd36b3, 
               32'shf9ba1651, 32'shf9b6f5f3, 32'shf9b3d599, 32'shf9b0b542, 32'shf9ad94f0, 32'shf9aa74a1, 32'shf9a75457, 32'shf9a43410, 
               32'shf9a113cd, 32'shf99df38e, 32'shf99ad354, 32'shf997b31d, 32'shf99492ea, 32'shf99172bb, 32'shf98e528f, 32'shf98b3268, 
               32'shf9881245, 32'shf984f226, 32'shf981d20b, 32'shf97eb1f4, 32'shf97b91e1, 32'shf97871d2, 32'shf97551c6, 32'shf97231bf, 
               32'shf96f11bc, 32'shf96bf1be, 32'shf968d1c3, 32'shf965b1cc, 32'shf96291d9, 32'shf95f71ea, 32'shf95c5200, 32'shf9593219, 
               32'shf9561237, 32'shf952f259, 32'shf94fd27f, 32'shf94cb2a8, 32'shf94992d7, 32'shf9467309, 32'shf943533f, 32'shf940337a, 
               32'shf93d13b8, 32'shf939f3fb, 32'shf936d442, 32'shf933b48e, 32'shf93094dd, 32'shf92d7531, 32'shf92a5589, 32'shf92735e5, 
               32'shf9241645, 32'shf920f6a9, 32'shf91dd712, 32'shf91ab77f, 32'shf91797f0, 32'shf9147866, 32'shf91158e0, 32'shf90e395e, 
               32'shf90b19e0, 32'shf907fa67, 32'shf904daf2, 32'shf901bb81, 32'shf8fe9c15, 32'shf8fb7cac, 32'shf8f85d49, 32'shf8f53de9, 
               32'shf8f21e8e, 32'shf8eeff37, 32'shf8ebdfe5, 32'shf8e8c097, 32'shf8e5a14d, 32'shf8e28208, 32'shf8df62c7, 32'shf8dc438b, 
               32'shf8d92452, 32'shf8d6051f, 32'shf8d2e5f0, 32'shf8cfc6c5, 32'shf8cca79e, 32'shf8c9887c, 32'shf8c6695f, 32'shf8c34a46, 
               32'shf8c02b31, 32'shf8bd0c21, 32'shf8b9ed15, 32'shf8b6ce0e, 32'shf8b3af0c, 32'shf8b0900d, 32'shf8ad7114, 32'shf8aa521f, 
               32'shf8a7332e, 32'shf8a41442, 32'shf8a0f55b, 32'shf89dd678, 32'shf89ab799, 32'shf89798bf, 32'shf89479ea, 32'shf8915b19, 
               32'shf88e3c4d, 32'shf88b1d86, 32'shf887fec3, 32'shf884e004, 32'shf881c14b, 32'shf87ea295, 32'shf87b83e5, 32'shf8786539, 
               32'shf8754692, 32'shf87227ef, 32'shf86f0952, 32'shf86beab8, 32'shf868cc24, 32'shf865ad94, 32'shf8628f09, 32'shf85f7082, 
               32'shf85c5201, 32'shf8593383, 32'shf856150b, 32'shf852f698, 32'shf84fd829, 32'shf84cb9bf, 32'shf8499b59, 32'shf8467cf9, 
               32'shf8435e9d, 32'shf8404046, 32'shf83d21f3, 32'shf83a03a6, 32'shf836e55d, 32'shf833c719, 32'shf830a8da, 32'shf82d8aa0, 
               32'shf82a6c6a, 32'shf8274e3a, 32'shf824300e, 32'shf82111e7, 32'shf81df3c5, 32'shf81ad5a8, 32'shf817b78f, 32'shf814997c, 
               32'shf8117b6d, 32'shf80e5d64, 32'shf80b3f5f, 32'shf808215f, 32'shf8050364, 32'shf801e56e, 32'shf7fec77d, 32'shf7fba991, 
               32'shf7f88ba9, 32'shf7f56dc7, 32'shf7f24fea, 32'shf7ef3211, 32'shf7ec143e, 32'shf7e8f670, 32'shf7e5d8a6, 32'shf7e2bae2, 
               32'shf7df9d22, 32'shf7dc7f68, 32'shf7d961b3, 32'shf7d64402, 32'shf7d32657, 32'shf7d008b1, 32'shf7cceb0f, 32'shf7c9cd73, 
               32'shf7c6afdc, 32'shf7c3924a, 32'shf7c074bd, 32'shf7bd5735, 32'shf7ba39b3, 32'shf7b71c35, 32'shf7b3febc, 32'shf7b0e149, 
               32'shf7adc3db, 32'shf7aaa671, 32'shf7a7890d, 32'shf7a46baf, 32'shf7a14e55, 32'shf79e3100, 32'shf79b13b1, 32'shf797f667, 
               32'shf794d922, 32'shf791bbe2, 32'shf78e9ea7, 32'shf78b8172, 32'shf7886442, 32'shf7854717, 32'shf78229f1, 32'shf77f0cd0, 
               32'shf77befb5, 32'shf778d29f, 32'shf775b58e, 32'shf7729883, 32'shf76f7b7d, 32'shf76c5e7c, 32'shf7694180, 32'shf766248a, 
               32'shf7630799, 32'shf75feaad, 32'shf75ccdc6, 32'shf759b0e5, 32'shf756940a, 32'shf7537733, 32'shf7505a62, 32'shf74d3d96, 
               32'shf74a20d0, 32'shf747040f, 32'shf743e754, 32'shf740ca9d, 32'shf73daded, 32'shf73a9141, 32'shf737749b, 32'shf73457fb, 
               32'shf7313b60, 32'shf72e1eca, 32'shf72b023a, 32'shf727e5af, 32'shf724c92a, 32'shf721acaa, 32'shf71e902f, 32'shf71b73ba, 
               32'shf718574b, 32'shf7153ae1, 32'shf7121e7c, 32'shf70f021d, 32'shf70be5c4, 32'shf708c970, 32'shf705ad22, 32'shf70290d9, 
               32'shf6ff7496, 32'shf6fc5858, 32'shf6f93c20, 32'shf6f61fed, 32'shf6f303c0, 32'shf6efe798, 32'shf6eccb77, 32'shf6e9af5a, 
               32'shf6e69344, 32'shf6e37733, 32'shf6e05b27, 32'shf6dd3f21, 32'shf6da2321, 32'shf6d70727, 32'shf6d3eb32, 32'shf6d0cf43, 
               32'shf6cdb359, 32'shf6ca9775, 32'shf6c77b97, 32'shf6c45fbe, 32'shf6c143ec, 32'shf6be281e, 32'shf6bb0c57, 32'shf6b7f095, 
               32'shf6b4d4d9, 32'shf6b1b923, 32'shf6ae9d73, 32'shf6ab81c8, 32'shf6a86623, 32'shf6a54a84, 32'shf6a22eea, 32'shf69f1357, 
               32'shf69bf7c9, 32'shf698dc41, 32'shf695c0be, 32'shf692a542, 32'shf68f89cb, 32'shf68c6e5a, 32'shf68952ef, 32'shf686378a, 
               32'shf6831c2b, 32'shf68000d1, 32'shf67ce57e, 32'shf679ca30, 32'shf676aee8, 32'shf67393a6, 32'shf670786a, 32'shf66d5d34, 
               32'shf66a4203, 32'shf66726d9, 32'shf6640bb4, 32'shf660f096, 32'shf65dd57d, 32'shf65aba6b, 32'shf6579f5e, 32'shf6548457, 
               32'shf6516956, 32'shf64e4e5c, 32'shf64b3367, 32'shf6481878, 32'shf644fd8f, 32'shf641e2ac, 32'shf63ec7cf, 32'shf63bacf8, 
               32'shf6389228, 32'shf635775d, 32'shf6325c98, 32'shf62f41d9, 32'shf62c2721, 32'shf6290c6e, 32'shf625f1c2, 32'shf622d71b, 
               32'shf61fbc7b, 32'shf61ca1e1, 32'shf619874c, 32'shf6166cbe, 32'shf6135237, 32'shf61037b5, 32'shf60d1d39, 32'shf60a02c3, 
               32'shf606e854, 32'shf603cdeb, 32'shf600b388, 32'shf5fd992b, 32'shf5fa7ed4, 32'shf5f76484, 32'shf5f44a39, 32'shf5f12ff5, 
               32'shf5ee15b7, 32'shf5eafb7f, 32'shf5e7e14e, 32'shf5e4c722, 32'shf5e1acfd, 32'shf5de92de, 32'shf5db78c6, 32'shf5d85eb3, 
               32'shf5d544a7, 32'shf5d22aa2, 32'shf5cf10a2, 32'shf5cbf6a9, 32'shf5c8dcb6, 32'shf5c5c2c9, 32'shf5c2a8e3, 32'shf5bf8f03, 
               32'shf5bc7529, 32'shf5b95b56, 32'shf5b64189, 32'shf5b327c2, 32'shf5b00e02, 32'shf5acf448, 32'shf5a9da94, 32'shf5a6c0e7, 
               32'shf5a3a740, 32'shf5a08da0, 32'shf59d7406, 32'shf59a5a72, 32'shf59740e5, 32'shf594275e, 32'shf5910dde, 32'shf58df464, 
               32'shf58adaf0, 32'shf587c183, 32'shf584a81d, 32'shf5818ebd, 32'shf57e7563, 32'shf57b5c10, 32'shf57842c3, 32'shf575297d, 
               32'shf572103d, 32'shf56ef704, 32'shf56bddd1, 32'shf568c4a5, 32'shf565ab80, 32'shf5629261, 32'shf55f7948, 32'shf55c6036, 
               32'shf559472b, 32'shf5562e26, 32'shf5531528, 32'shf54ffc30, 32'shf54ce33f, 32'shf549ca55, 32'shf546b171, 32'shf5439893, 
               32'shf5407fbd, 32'shf53d66ed, 32'shf53a4e24, 32'shf5373561, 32'shf5341ca5, 32'shf53103ef, 32'shf52deb41, 32'shf52ad299, 
               32'shf527b9f7, 32'shf524a15d, 32'shf52188c9, 32'shf51e703b, 32'shf51b57b5, 32'shf5183f35, 32'shf51526bc, 32'shf5120e49, 
               32'shf50ef5de, 32'shf50bdd79, 32'shf508c51b, 32'shf505acc3, 32'shf5029473, 32'shf4ff7c29, 32'shf4fc63e6, 32'shf4f94baa, 
               32'shf4f63374, 32'shf4f31b46, 32'shf4f0031e, 32'shf4eceafd, 32'shf4e9d2e3, 32'shf4e6bacf, 32'shf4e3a2c3, 32'shf4e08abd, 
               32'shf4dd72be, 32'shf4da5ac7, 32'shf4d742d6, 32'shf4d42aeb, 32'shf4d11308, 32'shf4cdfb2c, 32'shf4cae356, 32'shf4c7cb88, 
               32'shf4c4b3c0, 32'shf4c19c00, 32'shf4be8446, 32'shf4bb6c93, 32'shf4b854e7, 32'shf4b53d42, 32'shf4b225a4, 32'shf4af0e0d, 
               32'shf4abf67e, 32'shf4a8def5, 32'shf4a5c773, 32'shf4a2aff8, 32'shf49f9884, 32'shf49c8117, 32'shf49969b1, 32'shf4965252, 
               32'shf4933afa, 32'shf49023a9, 32'shf48d0c5f, 32'shf489f51d, 32'shf486dde1, 32'shf483c6ad, 32'shf480af7f, 32'shf47d9859, 
               32'shf47a8139, 32'shf4776a21, 32'shf4745310, 32'shf4713c06, 32'shf46e2504, 32'shf46b0e08, 32'shf467f713, 32'shf464e026, 
               32'shf461c940, 32'shf45eb261, 32'shf45b9b89, 32'shf45884b8, 32'shf4556def, 32'shf452572c, 32'shf44f4071, 32'shf44c29be, 
               32'shf4491311, 32'shf445fc6b, 32'shf442e5cd, 32'shf43fcf36, 32'shf43cb8a7, 32'shf439a21e, 32'shf4368b9d, 32'shf4337523, 
               32'shf4305eb0, 32'shf42d4845, 32'shf42a31e1, 32'shf4271b84, 32'shf424052f, 32'shf420eee1, 32'shf41dd89a, 32'shf41ac25a, 
               32'shf417ac22, 32'shf41495f1, 32'shf4117fc8, 32'shf40e69a6, 32'shf40b538b, 32'shf4083d78, 32'shf405276c, 32'shf4021167, 
               32'shf3fefb6a, 32'shf3fbe574, 32'shf3f8cf86, 32'shf3f5b99f, 32'shf3f2a3bf, 32'shf3ef8de7, 32'shf3ec7817, 32'shf3e9624d, 
               32'shf3e64c8c, 32'shf3e336d1, 32'shf3e0211f, 32'shf3dd0b73, 32'shf3d9f5cf, 32'shf3d6e033, 32'shf3d3ca9e, 32'shf3d0b511, 
               32'shf3cd9f8b, 32'shf3ca8a0d, 32'shf3c77496, 32'shf3c45f27, 32'shf3c149bf, 32'shf3be345f, 32'shf3bb1f07, 32'shf3b809b6, 
               32'shf3b4f46c, 32'shf3b1df2a, 32'shf3aec9f0, 32'shf3abb4bd, 32'shf3a89f92, 32'shf3a58a6f, 32'shf3a27553, 32'shf39f603f, 
               32'shf39c4b32, 32'shf399362d, 32'shf3962130, 32'shf3930c3b, 32'shf38ff74d, 32'shf38ce266, 32'shf389cd88, 32'shf386b8b1, 
               32'shf383a3e2, 32'shf3808f1a, 32'shf37d7a5b, 32'shf37a65a2, 32'shf37750f2, 32'shf3743c49, 32'shf37127a9, 32'shf36e130f, 
               32'shf36afe7e, 32'shf367e9f4, 32'shf364d573, 32'shf361c0f9, 32'shf35eac86, 32'shf35b981c, 32'shf35883b9, 32'shf3556f5e, 
               32'shf3525b0b, 32'shf34f46c0, 32'shf34c327c, 32'shf3491e41, 32'shf3460a0d, 32'shf342f5e1, 32'shf33fe1bd, 32'shf33ccda1, 
               32'shf339b98d, 32'shf336a580, 32'shf333917c, 32'shf3307d7f, 32'shf32d698a, 32'shf32a559e, 32'shf32741b9, 32'shf3242ddc, 
               32'shf3211a07, 32'shf31e0639, 32'shf31af274, 32'shf317deb7, 32'shf314cb02, 32'shf311b755, 32'shf30ea3af, 32'shf30b9012, 
               32'shf3087c7d, 32'shf30568ef, 32'shf302556a, 32'shf2ff41ed, 32'shf2fc2e77, 32'shf2f91b0a, 32'shf2f607a5, 32'shf2f2f448, 
               32'shf2efe0f2, 32'shf2eccda5, 32'shf2e9ba60, 32'shf2e6a723, 32'shf2e393ef, 32'shf2e080c2, 32'shf2dd6d9d, 32'shf2da5a81, 
               32'shf2d7476c, 32'shf2d43460, 32'shf2d1215b, 32'shf2ce0e5f, 32'shf2cafb6b, 32'shf2c7e880, 32'shf2c4d59c, 32'shf2c1c2c0, 
               32'shf2beafed, 32'shf2bb9d22, 32'shf2b88a5f, 32'shf2b577a4, 32'shf2b264f2, 32'shf2af5247, 32'shf2ac3fa5, 32'shf2a92d0b, 
               32'shf2a61a7a, 32'shf2a307f0, 32'shf29ff56f, 32'shf29ce2f6, 32'shf299d085, 32'shf296be1d, 32'shf293abbd, 32'shf2909965, 
               32'shf28d8715, 32'shf28a74ce, 32'shf287628f, 32'shf2845058, 32'shf2813e2a, 32'shf27e2c04, 32'shf27b19e6, 32'shf27807d0, 
               32'shf274f5c3, 32'shf271e3bf, 32'shf26ed1c2, 32'shf26bbfce, 32'shf268ade3, 32'shf2659c00, 32'shf2628a25, 32'shf25f7852, 
               32'shf25c6688, 32'shf25954c7, 32'shf256430e, 32'shf253315d, 32'shf2501fb5, 32'shf24d0e15, 32'shf249fc7d, 32'shf246eaee, 
               32'shf243d968, 32'shf240c7ea, 32'shf23db674, 32'shf23aa507, 32'shf23793a3, 32'shf2348247, 32'shf23170f3, 32'shf22e5fa8, 
               32'shf22b4e66, 32'shf2283d2c, 32'shf2252bfa, 32'shf2221ad1, 32'shf21f09b1, 32'shf21bf899, 32'shf218e78a, 32'shf215d683, 
               32'shf212c585, 32'shf20fb490, 32'shf20ca3a3, 32'shf20992bf, 32'shf20681e3, 32'shf2037110, 32'shf2006046, 32'shf1fd4f84, 
               32'shf1fa3ecb, 32'shf1f72e1a, 32'shf1f41d72, 32'shf1f10cd3, 32'shf1edfc3d, 32'shf1eaebaf, 32'shf1e7db2a, 32'shf1e4caae, 
               32'shf1e1ba3a, 32'shf1dea9cf, 32'shf1db996d, 32'shf1d88913, 32'shf1d578c2, 32'shf1d2687a, 32'shf1cf583b, 32'shf1cc4804, 
               32'shf1c937d6, 32'shf1c627b1, 32'shf1c31795, 32'shf1c00781, 32'shf1bcf777, 32'shf1b9e775, 32'shf1b6d77c, 32'shf1b3c78b, 
               32'shf1b0b7a4, 32'shf1ada7c5, 32'shf1aa97ef, 32'shf1a78822, 32'shf1a4785e, 32'shf1a168a3, 32'shf19e58f1, 32'shf19b4947, 
               32'shf19839a6, 32'shf1952a0f, 32'shf1921a80, 32'shf18f0afa, 32'shf18bfb7d, 32'shf188ec09, 32'shf185dc9d, 32'shf182cd3b, 
               32'shf17fbde2, 32'shf17cae91, 32'shf1799f4a, 32'shf176900b, 32'shf17380d6, 32'shf17071a9, 32'shf16d6286, 32'shf16a536b, 
               32'shf1674459, 32'shf1643551, 32'shf1612651, 32'shf15e175b, 32'shf15b086d, 32'shf157f989, 32'shf154eaad, 32'shf151dbdb, 
               32'shf14ecd11, 32'shf14bbe51, 32'shf148af9a, 32'shf145a0ec, 32'shf1429247, 32'shf13f83ab, 32'shf13c7518, 32'shf139668e, 
               32'shf136580d, 32'shf1334996, 32'shf1303b27, 32'shf12d2cc2, 32'shf12a1e66, 32'shf1271013, 32'shf12401c9, 32'shf120f389, 
               32'shf11de551, 32'shf11ad723, 32'shf117c8fe, 32'shf114bae2, 32'shf111accf, 32'shf10e9ec6, 32'shf10b90c5, 32'shf10882ce, 
               32'shf10574e0, 32'shf10266fc, 32'shf0ff5921, 32'shf0fc4b4f, 32'shf0f93d86, 32'shf0f62fc6, 32'shf0f32210, 32'shf0f01463, 
               32'shf0ed06bf, 32'shf0e9f925, 32'shf0e6eb94, 32'shf0e3de0c, 32'shf0e0d08d, 32'shf0ddc318, 32'shf0dab5ad, 32'shf0d7a84a, 
               32'shf0d49af1, 32'shf0d18da1, 32'shf0ce805b, 32'shf0cb731e, 32'shf0c865ea, 32'shf0c558c0, 32'shf0c24b9f, 32'shf0bf3e88, 
               32'shf0bc317a, 32'shf0b92475, 32'shf0b6177a, 32'shf0b30a88, 32'shf0affda0, 32'shf0acf0c1, 32'shf0a9e3eb, 32'shf0a6d71f, 
               32'shf0a3ca5d, 32'shf0a0bda4, 32'shf09db0f4, 32'shf09aa44e, 32'shf09797b2, 32'shf0948b1f, 32'shf0917e95, 32'shf08e7215, 
               32'shf08b659f, 32'shf0885932, 32'shf0854cce, 32'shf0824074, 32'shf07f3424, 32'shf07c27dd, 32'shf0791ba0, 32'shf0760f6c, 
               32'shf0730342, 32'shf06ff722, 32'shf06ceb0b, 32'shf069defe, 32'shf066d2fa, 32'shf063c700, 32'shf060bb10, 32'shf05daf29, 
               32'shf05aa34c, 32'shf0579779, 32'shf0548baf, 32'shf0517fef, 32'shf04e7438, 32'shf04b688c, 32'shf0485ce9, 32'shf045514f, 
               32'shf04245c0, 32'shf03f3a3a, 32'shf03c2ebd, 32'shf039234b, 32'shf03617e2, 32'shf0330c83, 32'shf030012e, 32'shf02cf5e2, 
               32'shf029eaa1, 32'shf026df68, 32'shf023d43a, 32'shf020c916, 32'shf01dbdfb, 32'shf01ab2ea, 32'shf017a7e3, 32'shf0149ce6, 
               32'shf01191f3, 32'shf00e8709, 32'shf00b7c29, 32'shf0087153, 32'shf0056687, 32'shf0025bc5, 32'shefff510d, 32'sheffc465e, 
               32'sheff93bba, 32'sheff6311f, 32'sheff3268e, 32'sheff01c07, 32'shefed118a, 32'shefea0717, 32'shefe6fcae, 32'shefe3f24f, 
               32'shefe0e7f9, 32'shefddddae, 32'shefdad36c, 32'shefd7c935, 32'shefd4bf08, 32'shefd1b4e4, 32'shefceaacb, 32'shefcba0bb, 
               32'shefc896b5, 32'shefc58cba, 32'shefc282c8, 32'shefbf78e1, 32'shefbc6f03, 32'shefb96530, 32'shefb65b66, 32'shefb351a7, 
               32'shefb047f2, 32'shefad3e47, 32'shefaa34a5, 32'shefa72b0e, 32'shefa42181, 32'shefa117fe, 32'shef9e0e85, 32'shef9b0517, 
               32'shef97fbb2, 32'shef94f258, 32'shef91e907, 32'shef8edfc1, 32'shef8bd685, 32'shef88cd53, 32'shef85c42b, 32'shef82bb0e, 
               32'shef7fb1fa, 32'shef7ca8f1, 32'shef799ff2, 32'shef7696fd, 32'shef738e12, 32'shef708532, 32'shef6d7c5b, 32'shef6a738f, 
               32'shef676ace, 32'shef646216, 32'shef615969, 32'shef5e50c6, 32'shef5b482d, 32'shef583f9e, 32'shef55371a, 32'shef522ea0, 
               32'shef4f2630, 32'shef4c1dcb, 32'shef491570, 32'shef460d1f, 32'shef4304d8, 32'shef3ffc9c, 32'shef3cf46a, 32'shef39ec43, 
               32'shef36e426, 32'shef33dc13, 32'shef30d40a, 32'shef2dcc0c, 32'shef2ac419, 32'shef27bc2f, 32'shef24b451, 32'shef21ac7c, 
               32'shef1ea4b2, 32'shef1b9cf2, 32'shef18953d, 32'shef158d92, 32'shef1285f2, 32'shef0f7e5c, 32'shef0c76d0, 32'shef096f4f, 
               32'shef0667d9, 32'shef03606c, 32'shef00590b, 32'sheefd51b4, 32'sheefa4a67, 32'sheef74325, 32'sheef43bed, 32'sheef134c0, 
               32'sheeee2d9d, 32'sheeeb2685, 32'sheee81f78, 32'sheee51875, 32'sheee2117c, 32'sheedf0a8e, 32'sheedc03ab, 32'sheed8fcd2, 
               32'sheed5f604, 32'sheed2ef40, 32'sheecfe887, 32'sheecce1d9, 32'sheec9db35, 32'sheec6d49c, 32'sheec3ce0d, 32'sheec0c78a, 
               32'sheebdc110, 32'sheebabaa2, 32'sheeb7b43e, 32'sheeb4ade4, 32'sheeb1a796, 32'sheeaea152, 32'sheeab9b18, 32'sheea894ea, 
               32'sheea58ec6, 32'sheea288ad, 32'shee9f829e, 32'shee9c7c9a, 32'shee9976a1, 32'shee9670b3, 32'shee936acf, 32'shee9064f7, 
               32'shee8d5f29, 32'shee8a5965, 32'shee8753ad, 32'shee844dff, 32'shee81485c, 32'shee7e42c4, 32'shee7b3d36, 32'shee7837b4, 
               32'shee75323c, 32'shee722ccf, 32'shee6f276d, 32'shee6c2216, 32'shee691cc9, 32'shee661788, 32'shee631251, 32'shee600d25, 
               32'shee5d0804, 32'shee5a02ee, 32'shee56fde3, 32'shee53f8e2, 32'shee50f3ed, 32'shee4def02, 32'shee4aea23, 32'shee47e54e, 
               32'shee44e084, 32'shee41dbc6, 32'shee3ed712, 32'shee3bd269, 32'shee38cdcb, 32'shee35c938, 32'shee32c4b0, 32'shee2fc033, 
               32'shee2cbbc1, 32'shee29b75a, 32'shee26b2fe, 32'shee23aead, 32'shee20aa67, 32'shee1da62c, 32'shee1aa1fc, 32'shee179dd7, 
               32'shee1499bd, 32'shee1195ae, 32'shee0e91aa, 32'shee0b8db1, 32'shee0889c4, 32'shee0585e1, 32'shee02820a, 32'shedff7e3d, 
               32'shedfc7a7c, 32'shedf976c6, 32'shedf6731b, 32'shedf36f7b, 32'shedf06be6, 32'sheded685d, 32'shedea64de, 32'shede7616b, 
               32'shede45e03, 32'shede15aa6, 32'shedde5754, 32'sheddb540d, 32'shedd850d2, 32'shedd54da2, 32'shedd24a7d, 32'shedcf4763, 
               32'shedcc4454, 32'shedc94151, 32'shedc63e59, 32'shedc33b6c, 32'shedc0388a, 32'shedbd35b4, 32'shedba32e9, 32'shedb73029, 
               32'shedb42d74, 32'shedb12acb, 32'shedae282d, 32'shedab259a, 32'sheda82313, 32'sheda52097, 32'sheda21e26, 32'shed9f1bc1, 
               32'shed9c1967, 32'shed991718, 32'shed9614d5, 32'shed93129d, 32'shed901070, 32'shed8d0e4f, 32'shed8a0c39, 32'shed870a2e, 
               32'shed84082f, 32'shed81063b, 32'shed7e0453, 32'shed7b0276, 32'shed7800a5, 32'shed74fedf, 32'shed71fd24, 32'shed6efb75, 
               32'shed6bf9d1, 32'shed68f839, 32'shed65f6ac, 32'shed62f52b, 32'shed5ff3b5, 32'shed5cf24b, 32'shed59f0ec, 32'shed56ef99, 
               32'shed53ee51, 32'shed50ed14, 32'shed4debe4, 32'shed4aeabe, 32'shed47e9a5, 32'shed44e897, 32'shed41e794, 32'shed3ee69d, 
               32'shed3be5b1, 32'shed38e4d2, 32'shed35e3fd, 32'shed32e334, 32'shed2fe277, 32'shed2ce1c6, 32'shed29e120, 32'shed26e086, 
               32'shed23dff7, 32'shed20df74, 32'shed1ddefd, 32'shed1ade91, 32'shed17de31, 32'shed14dddc, 32'shed11dd94, 32'shed0edd56, 
               32'shed0bdd25, 32'shed08dcff, 32'shed05dce5, 32'shed02dcd7, 32'shecffdcd4, 32'shecfcdcde, 32'shecf9dcf3, 32'shecf6dd13, 
               32'shecf3dd3f, 32'shecf0dd78, 32'shecedddbb, 32'sheceade0b, 32'shece7de66, 32'shece4dece, 32'shece1df40, 32'shecdedfbf, 
               32'shecdbe04a, 32'shecd8e0e0, 32'shecd5e182, 32'shecd2e230, 32'sheccfe2ea, 32'sheccce3b0, 32'shecc9e481, 32'shecc6e55f, 
               32'shecc3e648, 32'shecc0e73d, 32'shecbde83e, 32'shecbae94b, 32'shecb7ea63, 32'shecb4eb88, 32'shecb1ecb8, 32'shecaeedf5, 
               32'shecabef3d, 32'sheca8f091, 32'sheca5f1f2, 32'sheca2f35e, 32'shec9ff4d6, 32'shec9cf65a, 32'shec99f7ea, 32'shec96f986, 
               32'shec93fb2e, 32'shec90fce1, 32'shec8dfea1, 32'shec8b006d, 32'shec880245, 32'shec850429, 32'shec820619, 32'shec7f0815, 
               32'shec7c0a1d, 32'shec790c31, 32'shec760e51, 32'shec73107d, 32'shec7012b5, 32'shec6d14f9, 32'shec6a1749, 32'shec6719a6, 
               32'shec641c0e, 32'shec611e83, 32'shec5e2103, 32'shec5b2390, 32'shec582629, 32'shec5528ce, 32'shec522b7f, 32'shec4f2e3d, 
               32'shec4c3106, 32'shec4933dc, 32'shec4636bd, 32'shec4339ab, 32'shec403ca5, 32'shec3d3fac, 32'shec3a42be, 32'shec3745dd, 
               32'shec344908, 32'shec314c3f, 32'shec2e4f82, 32'shec2b52d1, 32'shec28562d, 32'shec255995, 32'shec225d09, 32'shec1f608a, 
               32'shec1c6417, 32'shec1967b0, 32'shec166b55, 32'shec136f06, 32'shec1072c4, 32'shec0d768e, 32'shec0a7a65, 32'shec077e48, 
               32'shec048237, 32'shec018632, 32'shebfe8a3a, 32'shebfb8e4e, 32'shebf8926f, 32'shebf5969b, 32'shebf29ad4, 32'shebef9f1a, 
               32'shebeca36c, 32'shebe9a7ca, 32'shebe6ac35, 32'shebe3b0ac, 32'shebe0b52f, 32'shebddb9bf, 32'shebdabe5c, 32'shebd7c304, 
               32'shebd4c7ba, 32'shebd1cc7b, 32'shebced149, 32'shebcbd624, 32'shebc8db0b, 32'shebc5dffe, 32'shebc2e4fe, 32'shebbfea0b, 
               32'shebbcef23, 32'shebb9f449, 32'shebb6f97b, 32'shebb3feb9, 32'shebb10404, 32'shebae095c, 32'shebab0ec0, 32'sheba81430, 
               32'sheba519ad, 32'sheba21f37, 32'sheb9f24cd, 32'sheb9c2a70, 32'sheb99301f, 32'sheb9635db, 32'sheb933ba4, 32'sheb904179, 
               32'sheb8d475b, 32'sheb8a4d49, 32'sheb875344, 32'sheb84594c, 32'sheb815f60, 32'sheb7e6581, 32'sheb7b6bae, 32'sheb7871e8, 
               32'sheb75782f, 32'sheb727e83, 32'sheb6f84e3, 32'sheb6c8b50, 32'sheb6991ca, 32'sheb669850, 32'sheb639ee3, 32'sheb60a582, 
               32'sheb5dac2f, 32'sheb5ab2e8, 32'sheb57b9ae, 32'sheb54c081, 32'sheb51c760, 32'sheb4ece4c, 32'sheb4bd545, 32'sheb48dc4b, 
               32'sheb45e35d, 32'sheb42ea7c, 32'sheb3ff1a8, 32'sheb3cf8e1, 32'sheb3a0027, 32'sheb370779, 32'sheb340ed9, 32'sheb311645, 
               32'sheb2e1dbe, 32'sheb2b2543, 32'sheb282cd6, 32'sheb253475, 32'sheb223c22, 32'sheb1f43db, 32'sheb1c4ba1, 32'sheb195374, 
               32'sheb165b54, 32'sheb136341, 32'sheb106b3a, 32'sheb0d7341, 32'sheb0a7b54, 32'sheb078375, 32'sheb048ba2, 32'sheb0193dd, 
               32'sheafe9c24, 32'sheafba478, 32'sheaf8acd9, 32'sheaf5b547, 32'sheaf2bdc3, 32'sheaefc64b, 32'sheaeccee0, 32'sheae9d782, 
               32'sheae6e031, 32'sheae3e8ed, 32'sheae0f1b6, 32'sheaddfa8d, 32'sheadb0370, 32'shead80c60, 32'shead5155d, 32'shead21e68, 
               32'sheacf277f, 32'sheacc30a4, 32'sheac939d5, 32'sheac64314, 32'sheac34c60, 32'sheac055b9, 32'sheabd5f1f, 32'sheaba6892, 
               32'sheab77212, 32'sheab47b9f, 32'sheab1853a, 32'sheaae8ee2, 32'sheaab9896, 32'sheaa8a258, 32'sheaa5ac27, 32'sheaa2b604, 
               32'shea9fbfed, 32'shea9cc9e4, 32'shea99d3e8, 32'shea96ddf9, 32'shea93e817, 32'shea90f242, 32'shea8dfc7b, 32'shea8b06c1, 
               32'shea881114, 32'shea851b74, 32'shea8225e2, 32'shea7f305d, 32'shea7c3ae5, 32'shea79457a, 32'shea76501d, 32'shea735acd, 
               32'shea70658a, 32'shea6d7055, 32'shea6a7b2d, 32'shea678612, 32'shea649105, 32'shea619c04, 32'shea5ea712, 32'shea5bb22c, 
               32'shea58bd54, 32'shea55c889, 32'shea52d3cc, 32'shea4fdf1c, 32'shea4cea79, 32'shea49f5e4, 32'shea47015c, 32'shea440ce1, 
               32'shea411874, 32'shea3e2415, 32'shea3b2fc2, 32'shea383b7e, 32'shea354746, 32'shea32531c, 32'shea2f5f00, 32'shea2c6af1, 
               32'shea2976ef, 32'shea2682fb, 32'shea238f15, 32'shea209b3b, 32'shea1da770, 32'shea1ab3b2, 32'shea17c001, 32'shea14cc5e, 
               32'shea11d8c8, 32'shea0ee540, 32'shea0bf1c6, 32'shea08fe59, 32'shea060af9, 32'shea0317a7, 32'shea002463, 32'she9fd312c, 
               32'she9fa3e03, 32'she9f74ae8, 32'she9f457da, 32'she9f164d9, 32'she9ee71e6, 32'she9eb7f01, 32'she9e88c2a, 32'she9e59960, 
               32'she9e2a6a3, 32'she9dfb3f5, 32'she9dcc154, 32'she9d9cec0, 32'she9d6dc3b, 32'she9d3e9c3, 32'she9d0f758, 32'she9ce04fc, 
               32'she9cb12ad, 32'she9c8206b, 32'she9c52e38, 32'she9c23c12, 32'she9bf49fa, 32'she9bc57f0, 32'she9b965f3, 32'she9b67404, 
               32'she9b38223, 32'she9b0904f, 32'she9ad9e8a, 32'she9aaacd2, 32'she9a7bb28, 32'she9a4c98b, 32'she9a1d7fd, 32'she99ee67c, 
               32'she99bf509, 32'she99903a4, 32'she996124d, 32'she9932103, 32'she9902fc7, 32'she98d3e9a, 32'she98a4d7a, 32'she9875c68, 
               32'she9846b63, 32'she9817a6d, 32'she97e8984, 32'she97b98aa, 32'she978a7dd, 32'she975b71e, 32'she972c66d, 32'she96fd5ca, 
               32'she96ce535, 32'she969f4ae, 32'she9670435, 32'she96413c9, 32'she961236c, 32'she95e331d, 32'she95b42db, 32'she95852a8, 
               32'she9556282, 32'she952726b, 32'she94f8261, 32'she94c9266, 32'she949a278, 32'she946b299, 32'she943c2c7, 32'she940d304, 
               32'she93de34e, 32'she93af3a7, 32'she938040d, 32'she9351482, 32'she9322505, 32'she92f3596, 32'she92c4634, 32'she92956e1, 
               32'she926679c, 32'she9237866, 32'she920893d, 32'she91d9a22, 32'she91aab16, 32'she917bc17, 32'she914cd27, 32'she911de45, 
               32'she90eef71, 32'she90c00ab, 32'she90911f3, 32'she906234a, 32'she90334af, 32'she9004621, 32'she8fd57a2, 32'she8fa6932, 
               32'she8f77acf, 32'she8f48c7b, 32'she8f19e34, 32'she8eeaffd, 32'she8ebc1d3, 32'she8e8d3b7, 32'she8e5e5aa, 32'she8e2f7ab, 
               32'she8e009ba, 32'she8dd1bd8, 32'she8da2e04, 32'she8d7403e, 32'she8d45286, 32'she8d164dd, 32'she8ce7742, 32'she8cb89b5, 
               32'she8c89c37, 32'she8c5aec7, 32'she8c2c165, 32'she8bfd412, 32'she8bce6cd, 32'she8b9f996, 32'she8b70c6d, 32'she8b41f53, 
               32'she8b13248, 32'she8ae454b, 32'she8ab585c, 32'she8a86b7b, 32'she8a57ea9, 32'she8a291e5, 32'she89fa530, 32'she89cb889, 
               32'she899cbf1, 32'she896df67, 32'she893f2eb, 32'she891067e, 32'she88e1a20, 32'she88b2dcf, 32'she888418e, 32'she885555a, 
               32'she8826936, 32'she87f7d1f, 32'she87c9118, 32'she879a51e, 32'she876b934, 32'she873cd57, 32'she870e18a, 32'she86df5cb, 
               32'she86b0a1a, 32'she8681e78, 32'she86532e4, 32'she862475f, 32'she85f5be9, 32'she85c7081, 32'she8598528, 32'she85699dd, 
               32'she853aea1, 32'she850c374, 32'she84dd855, 32'she84aed45, 32'she8480243, 32'she8451750, 32'she8422c6c, 32'she83f4196, 
               32'she83c56cf, 32'she8396c16, 32'she836816d, 32'she83396d2, 32'she830ac45, 32'she82dc1c8, 32'she82ad759, 32'she827ecf8, 
               32'she82502a7, 32'she8221864, 32'she81f2e30, 32'she81c440a, 32'she81959f4, 32'she8166fec, 32'she81385f3, 32'she8109c08, 
               32'she80db22d, 32'she80ac860, 32'she807dea2, 32'she804f4f2, 32'she8020b52, 32'she7ff21c0, 32'she7fc383d, 32'she7f94ec9, 
               32'she7f66564, 32'she7f37c0d, 32'she7f092c6, 32'she7eda98d, 32'she7eac063, 32'she7e7d748, 32'she7e4ee3c, 32'she7e2053e, 
               32'she7df1c50, 32'she7dc3370, 32'she7d94a9f, 32'she7d661de, 32'she7d3792b, 32'she7d09087, 32'she7cda7f2, 32'she7cabf6c, 
               32'she7c7d6f4, 32'she7c4ee8c, 32'she7c20633, 32'she7bf1de8, 32'she7bc35ad, 32'she7b94d80, 32'she7b66563, 32'she7b37d55, 
               32'she7b09555, 32'she7adad65, 32'she7aac583, 32'she7a7ddb1, 32'she7a4f5ed, 32'she7a20e39, 32'she79f2693, 32'she79c3efd, 
               32'she7995776, 32'she7966ffd, 32'she7938894, 32'she790a13a, 32'she78db9ef, 32'she78ad2b3, 32'she787eb86, 32'she7850468, 
               32'she7821d59, 32'she77f365a, 32'she77c4f69, 32'she7796888, 32'she77681b6, 32'she7739af2, 32'she770b43e, 32'she76dcd9a, 
               32'she76ae704, 32'she768007e, 32'she7651a06, 32'she762339e, 32'she75f4d45, 32'she75c66fb, 32'she75980c1, 32'she7569a95, 
               32'she753b479, 32'she750ce6c, 32'she74de86f, 32'she74b0280, 32'she7481ca1, 32'she74536d1, 32'she7425110, 32'she73f6b5f, 
               32'she73c85bc, 32'she739a029, 32'she736baa6, 32'she733d531, 32'she730efcc, 32'she72e0a77, 32'she72b2530, 32'she7283ff9, 
               32'she7255ad1, 32'she72275b9, 32'she71f90b0, 32'she71cabb6, 32'she719c6cb, 32'she716e1f0, 32'she713fd25, 32'she7111868, 
               32'she70e33bb, 32'she70b4f1e, 32'she7086a8f, 32'she7058611, 32'she702a1a1, 32'she6ffbd41, 32'she6fcd8f1, 32'she6f9f4b0, 
               32'she6f7107e, 32'she6f42c5c, 32'she6f14849, 32'she6ee6446, 32'she6eb8052, 32'she6e89c6d, 32'she6e5b899, 32'she6e2d4d3, 
               32'she6dff11d, 32'she6dd0d77, 32'she6da29e0, 32'she6d74658, 32'she6d462e1, 32'she6d17f78, 32'she6ce9c1f, 32'she6cbb8d6, 
               32'she6c8d59c, 32'she6c5f272, 32'she6c30f57, 32'she6c02c4c, 32'she6bd4951, 32'she6ba6665, 32'she6b78389, 32'she6b4a0bc, 
               32'she6b1bdff, 32'she6aedb51, 32'she6abf8b3, 32'she6a91625, 32'she6a633a6, 32'she6a35137, 32'she6a06ed8, 32'she69d8c88, 
               32'she69aaa48, 32'she697c818, 32'she694e5f7, 32'she69203e6, 32'she68f21e5, 32'she68c3ff3, 32'she6895e11, 32'she6867c3f, 
               32'she6839a7c, 32'she680b8ca, 32'she67dd727, 32'she67af593, 32'she6781410, 32'she675329c, 32'she6725138, 32'she66f6fe3, 
               32'she66c8e9f, 32'she669ad6a, 32'she666cc45, 32'she663eb30, 32'she6610a2a, 32'she65e2935, 32'she65b484f, 32'she6586779, 
               32'she65586b3, 32'she652a5fc, 32'she64fc556, 32'she64ce4bf, 32'she64a0438, 32'she64723c2, 32'she644435a, 32'she6416303, 
               32'she63e82bc, 32'she63ba285, 32'she638c25d, 32'she635e245, 32'she633023e, 32'she6302246, 32'she62d425e, 32'she62a6286, 
               32'she62782be, 32'she624a306, 32'she621c35e, 32'she61ee3c6, 32'she61c043d, 32'she61924c5, 32'she616455d, 32'she6136605, 
               32'she61086bc, 32'she60da784, 32'she60ac85c, 32'she607e944, 32'she6050a3b, 32'she6022b43, 32'she5ff4c5b, 32'she5fc6d83, 
               32'she5f98ebb, 32'she5f6b003, 32'she5f3d15b, 32'she5f0f2c3, 32'she5ee143b, 32'she5eb35c3, 32'she5e8575b, 32'she5e57904, 
               32'she5e29abc, 32'she5dfbc85, 32'she5dcde5e, 32'she5da0047, 32'she5d72240, 32'she5d44449, 32'she5d16662, 32'she5ce888b, 
               32'she5cbaac5, 32'she5c8cd0f, 32'she5c5ef69, 32'she5c311d3, 32'she5c0344d, 32'she5bd56d7, 32'she5ba7972, 32'she5b79c1d, 
               32'she5b4bed8, 32'she5b1e1a3, 32'she5af047f, 32'she5ac276b, 32'she5a94a67, 32'she5a66d73, 32'she5a39090, 32'she5a0b3bc, 
               32'she59dd6f9, 32'she59afa47, 32'she5981da4, 32'she5954112, 32'she5926490, 32'she58f881f, 32'she58cabbe, 32'she589cf6d, 
               32'she586f32c, 32'she58416fc, 32'she5813adc, 32'she57e5ecc, 32'she57b82cd, 32'she578a6de, 32'she575cb00, 32'she572ef32, 
               32'she5701374, 32'she56d37c7, 32'she56a5c2a, 32'she567809d, 32'she564a521, 32'she561c9b5, 32'she55eee5a, 32'she55c130f, 
               32'she55937d5, 32'she5565cab, 32'she5538191, 32'she550a688, 32'she54dcb8f, 32'she54af0a7, 32'she54815cf, 32'she5453b08, 
               32'she5426051, 32'she53f85ab, 32'she53cab15, 32'she539d090, 32'she536f61b, 32'she5341bb7, 32'she5314163, 32'she52e6720, 
               32'she52b8cee, 32'she528b2cc, 32'she525d8ba, 32'she522feb9, 32'she52024c9, 32'she51d4ae9, 32'she51a711a, 32'she517975b, 
               32'she514bdad, 32'she511e410, 32'she50f0a83, 32'she50c3107, 32'she509579b, 32'she5067e40, 32'she503a4f6, 32'she500cbbc, 
               32'she4fdf294, 32'she4fb197b, 32'she4f84074, 32'she4f5677d, 32'she4f28e96, 32'she4efb5c1, 32'she4ecdcfc, 32'she4ea0448, 
               32'she4e72ba4, 32'she4e45311, 32'she4e17a8f, 32'she4dea21e, 32'she4dbc9bd, 32'she4d8f16d, 32'she4d6192e, 32'she4d34100, 
               32'she4d068e2, 32'she4cd90d5, 32'she4cab8d9, 32'she4c7e0ee, 32'she4c50914, 32'she4c2314a, 32'she4bf5991, 32'she4bc81e9, 
               32'she4b9aa52, 32'she4b6d2cb, 32'she4b3fb56, 32'she4b123f1, 32'she4ae4c9d, 32'she4ab755a, 32'she4a89e28, 32'she4a5c707, 
               32'she4a2eff6, 32'she4a018f7, 32'she49d4208, 32'she49a6b2a, 32'she497945d, 32'she494bda1, 32'she491e6f6, 32'she48f105c, 
               32'she48c39d3, 32'she489635a, 32'she4868cf3, 32'she483b69d, 32'she480e057, 32'she47e0a23, 32'she47b33ff, 32'she4785ded, 
               32'she47587eb, 32'she472b1fa, 32'she46fdc1b, 32'she46d064c, 32'she46a308f, 32'she4675ae2, 32'she4648547, 32'she461afbc, 
               32'she45eda43, 32'she45c04da, 32'she4592f83, 32'she4565a3c, 32'she4538507, 32'she450afe3, 32'she44ddad0, 32'she44b05ce, 
               32'she44830dd, 32'she4455bfd, 32'she442872e, 32'she43fb271, 32'she43cddc4, 32'she43a0929, 32'she437349f, 32'she4346026, 
               32'she4318bbe, 32'she42eb767, 32'she42be321, 32'she4290eed, 32'she4263ac9, 32'she42366b7, 32'she42092b6, 32'she41dbec7, 
               32'she41aeae8, 32'she418171b, 32'she415435f, 32'she4126fb4, 32'she40f9c1a, 32'she40cc891, 32'she409f51a, 32'she40721b4, 
               32'she4044e60, 32'she4017b1c, 32'she3fea7ea, 32'she3fbd4c9, 32'she3f901ba, 32'she3f62ebb, 32'she3f35bce, 32'she3f088f2, 
               32'she3edb628, 32'she3eae36f, 32'she3e810c7, 32'she3e53e31, 32'she3e26bac, 32'she3df9938, 32'she3dcc6d5, 32'she3d9f484, 
               32'she3d72245, 32'she3d45016, 32'she3d17df9, 32'she3ceabee, 32'she3cbd9f4, 32'she3c9080b, 32'she3c63633, 32'she3c3646d, 
               32'she3c092b9, 32'she3bdc116, 32'she3baef84, 32'she3b81e04, 32'she3b54c95, 32'she3b27b38, 32'she3afa9ec, 32'she3acd8b1, 
               32'she3aa0788, 32'she3a73671, 32'she3a4656b, 32'she3a19476, 32'she39ec393, 32'she39bf2c2, 32'she3992202, 32'she3965153, 
               32'she39380b6, 32'she390b02b, 32'she38ddfb1, 32'she38b0f49, 32'she3883ef2, 32'she3856ead, 32'she3829e79, 32'she37fce57, 
               32'she37cfe47, 32'she37a2e48, 32'she3775e5a, 32'she3748e7f, 32'she371beb5, 32'she36eeefc, 32'she36c1f55, 32'she3694fc0, 
               32'she366803c, 32'she363b0cb, 32'she360e16a, 32'she35e121c, 32'she35b42df, 32'she35873b3, 32'she355a49a, 32'she352d592, 
               32'she350069b, 32'she34d37b7, 32'she34a68e4, 32'she3479a23, 32'she344cb73, 32'she341fcd6, 32'she33f2e4a, 32'she33c5fcf, 
               32'she3399167, 32'she336c310, 32'she333f4cb, 32'she3312698, 32'she32e5876, 32'she32b8a67, 32'she328bc69, 32'she325ee7d, 
               32'she32320a2, 32'she32052da, 32'she31d8523, 32'she31ab77e, 32'she317e9eb, 32'she3151c6a, 32'she3124efa, 32'she30f819d, 
               32'she30cb451, 32'she309e717, 32'she30719ef, 32'she3044cd9, 32'she3017fd5, 32'she2feb2e3, 32'she2fbe602, 32'she2f91934, 
               32'she2f64c77, 32'she2f37fcc, 32'she2f0b333, 32'she2ede6ac, 32'she2eb1a37, 32'she2e84dd4, 32'she2e58183, 32'she2e2b544, 
               32'she2dfe917, 32'she2dd1cfc, 32'she2da50f3, 32'she2d784fb, 32'she2d4b916, 32'she2d1ed43, 32'she2cf2182, 32'she2cc55d2, 
               32'she2c98a35, 32'she2c6beaa, 32'she2c3f331, 32'she2c127c9, 32'she2be5c74, 32'she2bb9131, 32'she2b8c600, 32'she2b5fae1, 
               32'she2b32fd4, 32'she2b064da, 32'she2ad99f1, 32'she2aacf1a, 32'she2a80456, 32'she2a539a3, 32'she2a26f03, 32'she29fa474, 
               32'she29cd9f8, 32'she29a0f8e, 32'she2974536, 32'she2947af1, 32'she291b0bd, 32'she28ee69c, 32'she28c1c8c, 32'she289528f, 
               32'she28688a4, 32'she283becc, 32'she280f505, 32'she27e2b51, 32'she27b61af, 32'she278981f, 32'she275cea1, 32'she2730536, 
               32'she2703bdc, 32'she26d7295, 32'she26aa960, 32'she267e03e, 32'she265172e, 32'she2624e2f, 32'she25f8544, 32'she25cbc6a, 
               32'she259f3a3, 32'she2572aee, 32'she254624b, 32'she25199bb, 32'she24ed13d, 32'she24c08d1, 32'she2494078, 32'she2467831, 
               32'she243affc, 32'she240e7da, 32'she23e1fca, 32'she23b57cc, 32'she2388fe1, 32'she235c808, 32'she2330041, 32'she230388d, 
               32'she22d70eb, 32'she22aa95c, 32'she227e1df, 32'she2251a75, 32'she222531c, 32'she21f8bd7, 32'she21cc4a3, 32'she219fd82, 
               32'she2173674, 32'she2146f78, 32'she211a88f, 32'she20ee1b7, 32'she20c1af3, 32'she2095441, 32'she2068da1, 32'she203c714, 
               32'she2010099, 32'she1fe3a31, 32'she1fb73dc, 32'she1f8ad98, 32'she1f5e768, 32'she1f3214a, 32'she1f05b3e, 32'she1ed9545, 
               32'she1eacf5f, 32'she1e8098b, 32'she1e543ca, 32'she1e27e1b, 32'she1dfb87f, 32'she1dcf2f5, 32'she1da2d7e, 32'she1d7681a, 
               32'she1d4a2c8, 32'she1d1dd89, 32'she1cf185c, 32'she1cc5342, 32'she1c98e3b, 32'she1c6c946, 32'she1c40464, 32'she1c13f95, 
               32'she1be7ad8, 32'she1bbb62e, 32'she1b8f197, 32'she1b62d12, 32'she1b368a0, 32'she1b0a441, 32'she1addff4, 32'she1ab1bba, 
               32'she1a85793, 32'she1a5937e, 32'she1a2cf7c, 32'she1a00b8d, 32'she19d47b1, 32'she19a83e7, 32'she197c031, 32'she194fc8d, 
               32'she19238fb, 32'she18f757d, 32'she18cb211, 32'she189eeb8, 32'she1872b72, 32'she184683e, 32'she181a51e, 32'she17ee210, 
               32'she17c1f15, 32'she1795c2d, 32'she1769958, 32'she173d695, 32'she17113e5, 32'she16e5149, 32'she16b8ebf, 32'she168cc48, 
               32'she16609e3, 32'she1634792, 32'she1608554, 32'she15dc328, 32'she15b0110, 32'she1583f0a, 32'she1557d17, 32'she152bb37, 
               32'she14ff96a, 32'she14d37b0, 32'she14a7609, 32'she147b475, 32'she144f2f3, 32'she1423185, 32'she13f702a, 32'she13caee1, 
               32'she139edac, 32'she1372c8a, 32'she1346b7a, 32'she131aa7e, 32'she12ee995, 32'she12c28be, 32'she12967fb, 32'she126a74a, 
               32'she123e6ad, 32'she1212623, 32'she11e65ac, 32'she11ba547, 32'she118e4f6, 32'she11624b8, 32'she113648d, 32'she110a475, 
               32'she10de470, 32'she10b247f, 32'she10864a0, 32'she105a4d4, 32'she102e51c, 32'she1002577, 32'she0fd65e4, 32'she0faa665, 
               32'she0f7e6f9, 32'she0f527a0, 32'she0f2685b, 32'she0efa928, 32'she0ecea09, 32'she0ea2afd, 32'she0e76c04, 32'she0e4ad1e, 
               32'she0e1ee4b, 32'she0df2f8c, 32'she0dc70e0, 32'she0d9b247, 32'she0d6f3c1, 32'she0d4354e, 32'she0d176ef, 32'she0ceb8a3, 
               32'she0cbfa6a, 32'she0c93c44, 32'she0c67e32, 32'she0c3c033, 32'she0c10247, 32'she0be446e, 32'she0bb86a9, 32'she0b8c8f7, 
               32'she0b60b58, 32'she0b34dcd, 32'she0b09055, 32'she0add2f0, 32'she0ab159e, 32'she0a85860, 32'she0a59b35, 32'she0a2de1e, 
               32'she0a0211a, 32'she09d6429, 32'she09aa74b, 32'she097ea81, 32'she0952dcb, 32'she0927127, 32'she08fb497, 32'she08cf81b, 
               32'she08a3bb2, 32'she0877f5c, 32'she084c31a, 32'she08206eb, 32'she07f4acf, 32'she07c8ec7, 32'she079d2d3, 32'she07716f2, 
               32'she0745b24, 32'she0719f6a, 32'she06ee3c3, 32'she06c2830, 32'she0696cb0, 32'she066b144, 32'she063f5eb, 32'she0613aa5, 
               32'she05e7f74, 32'she05bc455, 32'she059094a, 32'she0564e53, 32'she053936f, 32'she050d89f, 32'she04e1de3, 32'she04b6339, 
               32'she048a8a4, 32'she045ee22, 32'she04333b3, 32'she0407959, 32'she03dbf11, 32'she03b04de, 32'she0384abe, 32'she03590b1, 
               32'she032d6b8, 32'she0301cd3, 32'she02d6301, 32'she02aa943, 32'she027ef99, 32'she0253602, 32'she0227c7f, 32'she01fc310, 
               32'she01d09b4, 32'she01a506c, 32'she0179738, 32'she014de17, 32'she012250a, 32'she00f6c11, 32'she00cb32b, 32'she009fa59, 
               32'she007419b, 32'she00488f0, 32'she001d05a, 32'shdfff17d7, 32'shdffc5f67, 32'shdff9a70c, 32'shdff6eec4, 32'shdff43690, 
               32'shdff17e70, 32'shdfeec663, 32'shdfec0e6a, 32'shdfe95686, 32'shdfe69eb4, 32'shdfe3e6f7, 32'shdfe12f4e, 32'shdfde77b8, 
               32'shdfdbc036, 32'shdfd908c8, 32'shdfd6516e, 32'shdfd39a27, 32'shdfd0e2f5, 32'shdfce2bd6, 32'shdfcb74cb, 32'shdfc8bdd4, 
               32'shdfc606f1, 32'shdfc35022, 32'shdfc09967, 32'shdfbde2bf, 32'shdfbb2c2c, 32'shdfb875ac, 32'shdfb5bf41, 32'shdfb308e9, 
               32'shdfb052a5, 32'shdfad9c75, 32'shdfaae659, 32'shdfa83051, 32'shdfa57a5d, 32'shdfa2c47d, 32'shdfa00eb1, 32'shdf9d58f8, 
               32'shdf9aa354, 32'shdf97edc4, 32'shdf953848, 32'shdf9282df, 32'shdf8fcd8b, 32'shdf8d184b, 32'shdf8a631f, 32'shdf87ae06, 
               32'shdf84f902, 32'shdf824412, 32'shdf7f8f36, 32'shdf7cda6e, 32'shdf7a25ba, 32'shdf77711a, 32'shdf74bc8e, 32'shdf720816, 
               32'shdf6f53b3, 32'shdf6c9f63, 32'shdf69eb27, 32'shdf673700, 32'shdf6482ed, 32'shdf61ceee, 32'shdf5f1b02, 32'shdf5c672b, 
               32'shdf59b369, 32'shdf56ffba, 32'shdf544c1f, 32'shdf519899, 32'shdf4ee527, 32'shdf4c31c9, 32'shdf497e7f, 32'shdf46cb49, 
               32'shdf441828, 32'shdf41651a, 32'shdf3eb221, 32'shdf3bff3c, 32'shdf394c6b, 32'shdf3699af, 32'shdf33e707, 32'shdf313473, 
               32'shdf2e81f3, 32'shdf2bcf87, 32'shdf291d30, 32'shdf266aed, 32'shdf23b8be, 32'shdf2106a4, 32'shdf1e549d, 32'shdf1ba2ab, 
               32'shdf18f0ce, 32'shdf163f04, 32'shdf138d4f, 32'shdf10dbaf, 32'shdf0e2a22, 32'shdf0b78aa, 32'shdf08c746, 32'shdf0615f7, 
               32'shdf0364bc, 32'shdf00b395, 32'shdefe0282, 32'shdefb5184, 32'shdef8a09b, 32'shdef5efc5, 32'shdef33f04, 32'shdef08e58, 
               32'shdeedddc0, 32'shdeeb2d3c, 32'shdee87ccc, 32'shdee5cc72, 32'shdee31c2b, 32'shdee06bf9, 32'shdeddbbdb, 32'shdedb0bd2, 
               32'shded85bdd, 32'shded5abfd, 32'shded2fc31, 32'shded04c7a, 32'shdecd9cd7, 32'shdecaed48, 32'shdec83dce, 32'shdec58e69, 
               32'shdec2df18, 32'shdec02fdb, 32'shdebd80b3, 32'shdebad1a0, 32'shdeb822a1, 32'shdeb573b7, 32'shdeb2c4e1, 32'shdeb0161f, 
               32'shdead6773, 32'shdeaab8da, 32'shdea80a57, 32'shdea55be8, 32'shdea2ad8d, 32'shde9fff47, 32'shde9d5116, 32'shde9aa2f9, 
               32'shde97f4f1, 32'shde9546fd, 32'shde92991e, 32'shde8feb54, 32'shde8d3d9e, 32'shde8a8ffd, 32'shde87e271, 32'shde8534f9, 
               32'shde828796, 32'shde7fda48, 32'shde7d2d0e, 32'shde7a7fe9, 32'shde77d2d8, 32'shde7525dc, 32'shde7278f5, 32'shde6fcc23, 
               32'shde6d1f65, 32'shde6a72bc, 32'shde67c628, 32'shde6519a9, 32'shde626d3e, 32'shde5fc0e8, 32'shde5d14a6, 32'shde5a687a, 
               32'shde57bc62, 32'shde55105f, 32'shde526471, 32'shde4fb897, 32'shde4d0cd2, 32'shde4a6122, 32'shde47b587, 32'shde450a01, 
               32'shde425e8f, 32'shde3fb333, 32'shde3d07eb, 32'shde3a5cb8, 32'shde37b199, 32'shde350690, 32'shde325b9b, 32'shde2fb0bc, 
               32'shde2d05f1, 32'shde2a5b3b, 32'shde27b09a, 32'shde25060e, 32'shde225b96, 32'shde1fb134, 32'shde1d06e6, 32'shde1a5cad, 
               32'shde17b28a, 32'shde15087b, 32'shde125e81, 32'shde0fb49c, 32'shde0d0acc, 32'shde0a6111, 32'shde07b76b, 32'shde050dd9, 
               32'shde02645d, 32'shddffbaf6, 32'shddfd11a3, 32'shddfa6866, 32'shddf7bf3e, 32'shddf5162a, 32'shddf26d2c, 32'shddefc443, 
               32'shdded1b6e, 32'shddea72af, 32'shdde7ca05, 32'shdde5216f, 32'shdde278ef, 32'shdddfd084, 32'shdddd282e, 32'shddda7fed, 
               32'shddd7d7c1, 32'shddd52faa, 32'shddd287a8, 32'shddcfdfbb, 32'shddcd37e4, 32'shddca9021, 32'shddc7e873, 32'shddc540db, 
               32'shddc29958, 32'shddbff1ea, 32'shddbd4a91, 32'shddbaa34d, 32'shddb7fc1e, 32'shddb55504, 32'shddb2ae00, 32'shddb00711, 
               32'shddad6036, 32'shddaab972, 32'shdda812c2, 32'shdda56c27, 32'shdda2c5a2, 32'shdda01f32, 32'shdd9d78d7, 32'shdd9ad291, 
               32'shdd982c60, 32'shdd958645, 32'shdd92e03f, 32'shdd903a4e, 32'shdd8d9472, 32'shdd8aeeac, 32'shdd8848fb, 32'shdd85a35f, 
               32'shdd82fdd8, 32'shdd805867, 32'shdd7db30b, 32'shdd7b0dc4, 32'shdd786892, 32'shdd75c376, 32'shdd731e6f, 32'shdd70797e, 
               32'shdd6dd4a2, 32'shdd6b2fdb, 32'shdd688b29, 32'shdd65e68d, 32'shdd634206, 32'shdd609d94, 32'shdd5df938, 32'shdd5b54f1, 
               32'shdd58b0c0, 32'shdd560ca4, 32'shdd53689d, 32'shdd50c4ac, 32'shdd4e20d0, 32'shdd4b7d09, 32'shdd48d958, 32'shdd4635bd, 
               32'shdd439236, 32'shdd40eec5, 32'shdd3e4b6a, 32'shdd3ba824, 32'shdd3904f4, 32'shdd3661d8, 32'shdd33bed3, 32'shdd311be3, 
               32'shdd2e7908, 32'shdd2bd643, 32'shdd293393, 32'shdd2690f9, 32'shdd23ee74, 32'shdd214c05, 32'shdd1ea9ab, 32'shdd1c0767, 
               32'shdd196538, 32'shdd16c31f, 32'shdd14211b, 32'shdd117f2d, 32'shdd0edd55, 32'shdd0c3b92, 32'shdd0999e4, 32'shdd06f84d, 
               32'shdd0456ca, 32'shdd01b55e, 32'shdcff1407, 32'shdcfc72c5, 32'shdcf9d199, 32'shdcf73083, 32'shdcf48f82, 32'shdcf1ee97, 
               32'shdcef4dc2, 32'shdcecad02, 32'shdcea0c58, 32'shdce76bc3, 32'shdce4cb44, 32'shdce22adb, 32'shdcdf8a87, 32'shdcdcea49, 
               32'shdcda4a21, 32'shdcd7aa0e, 32'shdcd50a12, 32'shdcd26a2a, 32'shdccfca59, 32'shdccd2a9d, 32'shdcca8af7, 32'shdcc7eb67, 
               32'shdcc54bec, 32'shdcc2ac87, 32'shdcc00d38, 32'shdcbd6dff, 32'shdcbacedb, 32'shdcb82fcd, 32'shdcb590d5, 32'shdcb2f1f3, 
               32'shdcb05326, 32'shdcadb46f, 32'shdcab15ce, 32'shdca87743, 32'shdca5d8cd, 32'shdca33a6e, 32'shdca09c24, 32'shdc9dfdf0, 
               32'shdc9b5fd2, 32'shdc98c1ca, 32'shdc9623d7, 32'shdc9385fa, 32'shdc90e834, 32'shdc8e4a83, 32'shdc8bace8, 32'shdc890f62, 
               32'shdc8671f3, 32'shdc83d49a, 32'shdc813756, 32'shdc7e9a28, 32'shdc7bfd11, 32'shdc79600f, 32'shdc76c323, 32'shdc74264d, 
               32'shdc71898d, 32'shdc6eece2, 32'shdc6c504e, 32'shdc69b3d0, 32'shdc671768, 32'shdc647b15, 32'shdc61ded9, 32'shdc5f42b2, 
               32'shdc5ca6a2, 32'shdc5a0aa8, 32'shdc576ec3, 32'shdc54d2f5, 32'shdc52373c, 32'shdc4f9b9a, 32'shdc4d000d, 32'shdc4a6497, 
               32'shdc47c936, 32'shdc452dec, 32'shdc4292b8, 32'shdc3ff799, 32'shdc3d5c91, 32'shdc3ac19f, 32'shdc3826c3, 32'shdc358bfd, 
               32'shdc32f14d, 32'shdc3056b3, 32'shdc2dbc2f, 32'shdc2b21c1, 32'shdc28876a, 32'shdc25ed28, 32'shdc2352fd, 32'shdc20b8e8, 
               32'shdc1e1ee9, 32'shdc1b8500, 32'shdc18eb2d, 32'shdc165170, 32'shdc13b7c9, 32'shdc111e39, 32'shdc0e84bf, 32'shdc0beb5b, 
               32'shdc09520d, 32'shdc06b8d5, 32'shdc041fb4, 32'shdc0186a8, 32'shdbfeedb3, 32'shdbfc54d4, 32'shdbf9bc0c, 32'shdbf72359, 
               32'shdbf48abd, 32'shdbf1f237, 32'shdbef59c7, 32'shdbecc16e, 32'shdbea292b, 32'shdbe790fe, 32'shdbe4f8e7, 32'shdbe260e6, 
               32'shdbdfc8fc, 32'shdbdd3128, 32'shdbda996b, 32'shdbd801c3, 32'shdbd56a32, 32'shdbd2d2b8, 32'shdbd03b53, 32'shdbcda405, 
               32'shdbcb0cce, 32'shdbc875ac, 32'shdbc5dea1, 32'shdbc347ac, 32'shdbc0b0ce, 32'shdbbe1a06, 32'shdbbb8354, 32'shdbb8ecb9, 
               32'shdbb65634, 32'shdbb3bfc6, 32'shdbb1296e, 32'shdbae932c, 32'shdbabfd01, 32'shdba966ec, 32'shdba6d0ed, 32'shdba43b05, 
               32'shdba1a534, 32'shdb9f0f78, 32'shdb9c79d4, 32'shdb99e445, 32'shdb974ece, 32'shdb94b96c, 32'shdb922421, 32'shdb8f8eed, 
               32'shdb8cf9cf, 32'shdb8a64c7, 32'shdb87cfd6, 32'shdb853afc, 32'shdb82a638, 32'shdb80118a, 32'shdb7d7cf3, 32'shdb7ae873, 
               32'shdb785409, 32'shdb75bfb5, 32'shdb732b79, 32'shdb709752, 32'shdb6e0342, 32'shdb6b6f49, 32'shdb68db67, 32'shdb66479b, 
               32'shdb63b3e5, 32'shdb612046, 32'shdb5e8cbe, 32'shdb5bf94c, 32'shdb5965f1, 32'shdb56d2ac, 32'shdb543f7e, 32'shdb51ac67, 
               32'shdb4f1967, 32'shdb4c867d, 32'shdb49f3a9, 32'shdb4760ec, 32'shdb44ce46, 32'shdb423bb7, 32'shdb3fa93e, 32'shdb3d16dc, 
               32'shdb3a8491, 32'shdb37f25c, 32'shdb35603e, 32'shdb32ce36, 32'shdb303c46, 32'shdb2daa6c, 32'shdb2b18a9, 32'shdb2886fc, 
               32'shdb25f566, 32'shdb2363e7, 32'shdb20d27f, 32'shdb1e412d, 32'shdb1baff2, 32'shdb191ece, 32'shdb168dc1, 32'shdb13fccb, 
               32'shdb116beb, 32'shdb0edb22, 32'shdb0c4a70, 32'shdb09b9d4, 32'shdb072950, 32'shdb0498e2, 32'shdb02088b, 32'shdaff784b, 
               32'shdafce821, 32'shdafa580f, 32'shdaf7c813, 32'shdaf5382e, 32'shdaf2a860, 32'shdaf018a9, 32'shdaed8909, 32'shdaeaf980, 
               32'shdae86a0d, 32'shdae5dab2, 32'shdae34b6d, 32'shdae0bc3f, 32'shdade2d28, 32'shdadb9e28, 32'shdad90f3f, 32'shdad6806d, 
               32'shdad3f1b1, 32'shdad1630d, 32'shdaced47f, 32'shdacc4609, 32'shdac9b7a9, 32'shdac72961, 32'shdac49b2f, 32'shdac20d15, 
               32'shdabf7f11, 32'shdabcf124, 32'shdaba634e, 32'shdab7d590, 32'shdab547e8, 32'shdab2ba57, 32'shdab02cdd, 32'shdaad9f7b, 
               32'shdaab122f, 32'shdaa884fa, 32'shdaa5f7dd, 32'shdaa36ad6, 32'shdaa0dde7, 32'shda9e510e, 32'shda9bc44d, 32'shda9937a2, 
               32'shda96ab0f, 32'shda941e93, 32'shda91922e, 32'shda8f05e0, 32'shda8c79a9, 32'shda89ed89, 32'shda876180, 32'shda84d58f, 
               32'shda8249b4, 32'shda7fbdf1, 32'shda7d3244, 32'shda7aa6af, 32'shda781b31, 32'shda758fcb, 32'shda73047b, 32'shda707942, 
               32'shda6dee21, 32'shda6b6317, 32'shda68d824, 32'shda664d48, 32'shda63c284, 32'shda6137d6, 32'shda5ead40, 32'shda5c22c1, 
               32'shda599859, 32'shda570e09, 32'shda5483d0, 32'shda51f9ae, 32'shda4f6fa3, 32'shda4ce5af, 32'shda4a5bd3, 32'shda47d20e, 
               32'shda454860, 32'shda42beca, 32'shda40354a, 32'shda3dabe2, 32'shda3b2292, 32'shda389958, 32'shda361036, 32'shda33872c, 
               32'shda30fe38, 32'shda2e755c, 32'shda2bec97, 32'shda2963ea, 32'shda26db54, 32'shda2452d5, 32'shda21ca6e, 32'shda1f421e, 
               32'shda1cb9e5, 32'shda1a31c4, 32'shda17a9ba, 32'shda1521c7, 32'shda1299ec, 32'shda101228, 32'shda0d8a7c, 32'shda0b02e7, 
               32'shda087b69, 32'shda05f403, 32'shda036cb5, 32'shda00e57d, 32'shd9fe5e5e, 32'shd9fbd755, 32'shd9f95064, 32'shd9f6c98b, 
               32'shd9f442c9, 32'shd9f1bc1e, 32'shd9ef358b, 32'shd9ecaf10, 32'shd9ea28ac, 32'shd9e7a25f, 32'shd9e51c2a, 32'shd9e2960c, 
               32'shd9e01006, 32'shd9dd8a18, 32'shd9db0441, 32'shd9d87e81, 32'shd9d5f8d9, 32'shd9d37349, 32'shd9d0edd0, 32'shd9ce686e, 
               32'shd9cbe325, 32'shd9c95df3, 32'shd9c6d8d8, 32'shd9c453d5, 32'shd9c1cee9, 32'shd9bf4a15, 32'shd9bcc559, 32'shd9ba40b5, 
               32'shd9b7bc27, 32'shd9b537b2, 32'shd9b2b354, 32'shd9b02f0e, 32'shd9adaadf, 32'shd9ab26c8, 32'shd9a8a2c9, 32'shd9a61ee1, 
               32'shd9a39b11, 32'shd9a11759, 32'shd99e93b8, 32'shd99c102f, 32'shd9998cbe, 32'shd9970965, 32'shd9948623, 32'shd99202f8, 
               32'shd98f7fe6, 32'shd98cfceb, 32'shd98a7a08, 32'shd987f73d, 32'shd9857489, 32'shd982f1ed, 32'shd9806f69, 32'shd97decfd, 
               32'shd97b6aa8, 32'shd978e86b, 32'shd9766646, 32'shd973e438, 32'shd9716243, 32'shd96ee065, 32'shd96c5e9f, 32'shd969dcf1, 
               32'shd9675b5a, 32'shd964d9dc, 32'shd9625875, 32'shd95fd726, 32'shd95d55ef, 32'shd95ad4d0, 32'shd95853c8, 32'shd955d2d9, 
               32'shd9535201, 32'shd950d141, 32'shd94e5099, 32'shd94bd009, 32'shd9494f90, 32'shd946cf30, 32'shd9444ee7, 32'shd941ceb7, 
               32'shd93f4e9e, 32'shd93cce9d, 32'shd93a4eb4, 32'shd937cee3, 32'shd9354f2a, 32'shd932cf89, 32'shd9305000, 32'shd92dd08e, 
               32'shd92b5135, 32'shd928d1f4, 32'shd92652ca, 32'shd923d3b9, 32'shd92154bf, 32'shd91ed5de, 32'shd91c5714, 32'shd919d863, 
               32'shd91759c9, 32'shd914db47, 32'shd9125cde, 32'shd90fde8c, 32'shd90d6053, 32'shd90ae231, 32'shd9086428, 32'shd905e636, 
               32'shd903685d, 32'shd900ea9c, 32'shd8fe6cf2, 32'shd8fbef61, 32'shd8f971e8, 32'shd8f6f487, 32'shd8f4773e, 32'shd8f1fa0d, 
               32'shd8ef7cf4, 32'shd8ecfff4, 32'shd8ea830b, 32'shd8e8063a, 32'shd8e58982, 32'shd8e30ce2, 32'shd8e0905a, 32'shd8de13ea, 
               32'shd8db9792, 32'shd8d91b52, 32'shd8d69f2a, 32'shd8d4231b, 32'shd8d1a724, 32'shd8cf2b45, 32'shd8ccaf7e, 32'shd8ca33cf, 
               32'shd8c7b838, 32'shd8c53cba, 32'shd8c2c154, 32'shd8c04606, 32'shd8bdcad0, 32'shd8bb4fb3, 32'shd8b8d4ad, 32'shd8b659c0, 
               32'shd8b3deeb, 32'shd8b1642f, 32'shd8aee98a, 32'shd8ac6efe, 32'shd8a9f48a, 32'shd8a77a2f, 32'shd8a4ffec, 32'shd8a285c0, 
               32'shd8a00bae, 32'shd89d91b3, 32'shd89b17d1, 32'shd8989e07, 32'shd8962456, 32'shd893aabc, 32'shd891313b, 32'shd88eb7d3, 
               32'shd88c3e83, 32'shd889c54b, 32'shd8874c2b, 32'shd884d324, 32'shd8825a35, 32'shd87fe15e, 32'shd87d68a0, 32'shd87aeffa, 
               32'shd878776d, 32'shd875fef8, 32'shd873869b, 32'shd8710e57, 32'shd86e962b, 32'shd86c1e18, 32'shd869a61d, 32'shd8672e3a, 
               32'shd864b670, 32'shd8623ebe, 32'shd85fc725, 32'shd85d4fa4, 32'shd85ad83c, 32'shd85860ec, 32'shd855e9b4, 32'shd8537295, 
               32'shd850fb8e, 32'shd84e84a0, 32'shd84c0dcb, 32'shd849970e, 32'shd8472069, 32'shd844a9dd, 32'shd8423369, 32'shd83fbd0e, 
               32'shd83d46cc, 32'shd83ad0a2, 32'shd8385a90, 32'shd835e497, 32'shd8336eb7, 32'shd830f8ef, 32'shd82e833f, 32'shd82c0da9, 
               32'shd829982b, 32'shd82722c5, 32'shd824ad78, 32'shd8223843, 32'shd81fc328, 32'shd81d4e24, 32'shd81ad93a, 32'shd8186468, 
               32'shd815efae, 32'shd8137b0d, 32'shd8110685, 32'shd80e9216, 32'shd80c1dbf, 32'shd809a980, 32'shd807355b, 32'shd804c14e, 
               32'shd8024d59, 32'shd7ffd97e, 32'shd7fd65bb, 32'shd7faf211, 32'shd7f87e7f, 32'shd7f60b06, 32'shd7f397a6, 32'shd7f1245e, 
               32'shd7eeb130, 32'shd7ec3e1a, 32'shd7e9cb1c, 32'shd7e75838, 32'shd7e4e56c, 32'shd7e272b8, 32'shd7e0001e, 32'shd7dd8d9c, 
               32'shd7db1b34, 32'shd7d8a8e3, 32'shd7d636ac, 32'shd7d3c48d, 32'shd7d15288, 32'shd7cee09b, 32'shd7cc6ec6, 32'shd7c9fd0b, 
               32'shd7c78b68, 32'shd7c519de, 32'shd7c2a86d, 32'shd7c03715, 32'shd7bdc5d6, 32'shd7bb54af, 32'shd7b8e3a2, 32'shd7b672ad, 
               32'shd7b401d1, 32'shd7b1910e, 32'shd7af2063, 32'shd7acafd2, 32'shd7aa3f5a, 32'shd7a7cefa, 32'shd7a55eb3, 32'shd7a2ee85, 
               32'shd7a07e70, 32'shd79e0e74, 32'shd79b9e91, 32'shd7992ec7, 32'shd796bf16, 32'shd7944f7d, 32'shd791dffe, 32'shd78f7097, 
               32'shd78d014a, 32'shd78a9215, 32'shd78822f9, 32'shd785b3f7, 32'shd783450d, 32'shd780d63c, 32'shd77e6784, 32'shd77bf8e6, 
               32'shd7798a60, 32'shd7771bf3, 32'shd774ad9f, 32'shd7723f64, 32'shd76fd143, 32'shd76d633a, 32'shd76af54a, 32'shd7688774, 
               32'shd76619b6, 32'shd763ac11, 32'shd7613e86, 32'shd75ed113, 32'shd75c63ba, 32'shd759f679, 32'shd7578952, 32'shd7551c44, 
               32'shd752af4f, 32'shd7504273, 32'shd74dd5b0, 32'shd74b6906, 32'shd748fc75, 32'shd7468ffe, 32'shd744239f, 32'shd741b75a, 
               32'shd73f4b2e, 32'shd73cdf1b, 32'shd73a7321, 32'shd7380740, 32'shd7359b78, 32'shd7332fca, 32'shd730c434, 32'shd72e58b8, 
               32'shd72bed55, 32'shd729820c, 32'shd72716db, 32'shd724abc4, 32'shd72240c5, 32'shd71fd5e0, 32'shd71d6b15, 32'shd71b0062, 
               32'shd71895c9, 32'shd7162b49, 32'shd713c0e2, 32'shd7115694, 32'shd70eec60, 32'shd70c8245, 32'shd70a1843, 32'shd707ae5a, 
               32'shd705448b, 32'shd702dad5, 32'shd7007138, 32'shd6fe07b5, 32'shd6fb9e4b, 32'shd6f934fa, 32'shd6f6cbc2, 32'shd6f462a4, 
               32'shd6f1f99f, 32'shd6ef90b4, 32'shd6ed27e1, 32'shd6eabf28, 32'shd6e85689, 32'shd6e5ee03, 32'shd6e38596, 32'shd6e11d42, 
               32'shd6deb508, 32'shd6dc4ce7, 32'shd6d9e4e0, 32'shd6d77cf2, 32'shd6d5151d, 32'shd6d2ad62, 32'shd6d045c0, 32'shd6cdde38, 
               32'shd6cb76c9, 32'shd6c90f73, 32'shd6c6a837, 32'shd6c44114, 32'shd6c1da0b, 32'shd6bf731b, 32'shd6bd0c45, 32'shd6baa588, 
               32'shd6b83ee4, 32'shd6b5d85a, 32'shd6b371ea, 32'shd6b10b92, 32'shd6aea555, 32'shd6ac3f31, 32'shd6a9d926, 32'shd6a77335, 
               32'shd6a50d5d, 32'shd6a2a79f, 32'shd6a041fa, 32'shd69ddc6f, 32'shd69b76fe, 32'shd69911a6, 32'shd696ac67, 32'shd6944742, 
               32'shd691e237, 32'shd68f7d45, 32'shd68d186d, 32'shd68ab3ae, 32'shd6884f09, 32'shd685ea7d, 32'shd683860b, 32'shd68121b3, 
               32'shd67ebd74, 32'shd67c594f, 32'shd679f543, 32'shd6779151, 32'shd6752d79, 32'shd672c9ba, 32'shd6706615, 32'shd66e028a, 
               32'shd66b9f18, 32'shd6693bc0, 32'shd666d881, 32'shd664755c, 32'shd6621251, 32'shd65faf60, 32'shd65d4c88, 32'shd65ae9ca, 
               32'shd6588725, 32'shd656249b, 32'shd653c229, 32'shd6515fd2, 32'shd64efd94, 32'shd64c9b71, 32'shd64a3966, 32'shd647d776, 
               32'shd645759f, 32'shd64313e2, 32'shd640b23f, 32'shd63e50b5, 32'shd63bef46, 32'shd6398df0, 32'shd6372cb3, 32'shd634cb91, 
               32'shd6326a88, 32'shd6300999, 32'shd62da8c4, 32'shd62b4809, 32'shd628e767, 32'shd62686e0, 32'shd6242672, 32'shd621c61e, 
               32'shd61f65e4, 32'shd61d05c3, 32'shd61aa5bd, 32'shd61845d0, 32'shd615e5fd, 32'shd6138644, 32'shd61126a5, 32'shd60ec720, 
               32'shd60c67b4, 32'shd60a0863, 32'shd607a92b, 32'shd6054a0d, 32'shd602eb0a, 32'shd6008c20, 32'shd5fe2d50, 32'shd5fbce9a, 
               32'shd5f96ffd, 32'shd5f7117b, 32'shd5f4b313, 32'shd5f254c4, 32'shd5eff690, 32'shd5ed9875, 32'shd5eb3a75, 32'shd5e8dc8e, 
               32'shd5e67ec1, 32'shd5e4210f, 32'shd5e1c376, 32'shd5df65f7, 32'shd5dd0892, 32'shd5daab48, 32'shd5d84e17, 32'shd5d5f100, 
               32'shd5d39403, 32'shd5d13721, 32'shd5ceda58, 32'shd5cc7da9, 32'shd5ca2115, 32'shd5c7c49a, 32'shd5c56839, 32'shd5c30bf3, 
               32'shd5c0afc6, 32'shd5be53b4, 32'shd5bbf7bc, 32'shd5b99bdd, 32'shd5b74019, 32'shd5b4e46f, 32'shd5b288df, 32'shd5b02d69, 
               32'shd5add20d, 32'shd5ab76cb, 32'shd5a91ba4, 32'shd5a6c096, 32'shd5a465a3, 32'shd5a20aca, 32'shd59fb00b, 32'shd59d5566, 
               32'shd59afadb, 32'shd598a06a, 32'shd5964614, 32'shd593ebd7, 32'shd59191b5, 32'shd58f37ad, 32'shd58cddbf, 32'shd58a83eb, 
               32'shd5882a32, 32'shd585d093, 32'shd583770e, 32'shd5811da3, 32'shd57ec452, 32'shd57c6b1c, 32'shd57a1200, 32'shd577b8fe, 
               32'shd5756016, 32'shd5730748, 32'shd570ae95, 32'shd56e55fc, 32'shd56bfd7d, 32'shd569a519, 32'shd5674ccf, 32'shd564f49f, 
               32'shd5629c89, 32'shd560448e, 32'shd55decad, 32'shd55b94e6, 32'shd5593d3a, 32'shd556e5a7, 32'shd5548e30, 32'shd55236d2, 
               32'shd54fdf8f, 32'shd54d8866, 32'shd54b3157, 32'shd548da63, 32'shd5468389, 32'shd5442cca, 32'shd541d625, 32'shd53f7f9a, 
               32'shd53d292a, 32'shd53ad2d4, 32'shd5387c98, 32'shd5362677, 32'shd533d070, 32'shd5317a84, 32'shd52f24b2, 32'shd52ccefa, 
               32'shd52a795d, 32'shd52823da, 32'shd525ce72, 32'shd5237924, 32'shd52123f0, 32'shd51eced7, 32'shd51c79d9, 32'shd51a24f5, 
               32'shd517d02b, 32'shd5157b7c, 32'shd51326e7, 32'shd510d26d, 32'shd50e7e0d, 32'shd50c29c8, 32'shd509d59d, 32'shd507818d, 
               32'shd5052d97, 32'shd502d9bc, 32'shd50085fb, 32'shd4fe3255, 32'shd4fbdec9, 32'shd4f98b58, 32'shd4f73801, 32'shd4f4e4c5, 
               32'shd4f291a4, 32'shd4f03e9d, 32'shd4edebb0, 32'shd4eb98de, 32'shd4e94627, 32'shd4e6f38b, 32'shd4e4a108, 32'shd4e24ea1, 
               32'shd4dffc54, 32'shd4ddaa22, 32'shd4db580a, 32'shd4d9060d, 32'shd4d6b42b, 32'shd4d46263, 32'shd4d210b5, 32'shd4cfbf23, 
               32'shd4cd6dab, 32'shd4cb1c4e, 32'shd4c8cb0b, 32'shd4c679e3, 32'shd4c428d6, 32'shd4c1d7e3, 32'shd4bf870b, 32'shd4bd364e, 
               32'shd4bae5ab, 32'shd4b89523, 32'shd4b644b6, 32'shd4b3f464, 32'shd4b1a42c, 32'shd4af540f, 32'shd4ad040c, 32'shd4aab425, 
               32'shd4a86458, 32'shd4a614a6, 32'shd4a3c50e, 32'shd4a17591, 32'shd49f2630, 32'shd49cd6e8, 32'shd49a87bc, 32'shd49838aa, 
               32'shd495e9b3, 32'shd4939ad7, 32'shd4914c16, 32'shd48efd6f, 32'shd48caee4, 32'shd48a6073, 32'shd488121d, 32'shd485c3e1, 
               32'shd48375c1, 32'shd48127bb, 32'shd47ed9d0, 32'shd47c8c00, 32'shd47a3e4b, 32'shd477f0b1, 32'shd475a332, 32'shd47355cd, 
               32'shd4710883, 32'shd46ebb54, 32'shd46c6e40, 32'shd46a2147, 32'shd467d469, 32'shd46587a6, 32'shd4633afd, 32'shd460ee70, 
               32'shd45ea1fd, 32'shd45c55a5, 32'shd45a0969, 32'shd457bd47, 32'shd4557140, 32'shd4532554, 32'shd450d983, 32'shd44e8dcd, 
               32'shd44c4232, 32'shd449f6b1, 32'shd447ab4c, 32'shd4456002, 32'shd44314d3, 32'shd440c9be, 32'shd43e7ec5, 32'shd43c33e7, 
               32'shd439e923, 32'shd4379e7b, 32'shd43553ee, 32'shd433097b, 32'shd430bf24, 32'shd42e74e8, 32'shd42c2ac6, 32'shd429e0c0, 
               32'shd42796d5, 32'shd4254d05, 32'shd4230350, 32'shd420b9b6, 32'shd41e7037, 32'shd41c26d3, 32'shd419dd8a, 32'shd417945c, 
               32'shd4154b4a, 32'shd4130252, 32'shd410b976, 32'shd40e70b4, 32'shd40c280e, 32'shd409df83, 32'shd4079713, 32'shd4054ebe, 
               32'shd4030684, 32'shd400be66, 32'shd3fe7662, 32'shd3fc2e7a, 32'shd3f9e6ad, 32'shd3f79efa, 32'shd3f55764, 32'shd3f30fe8, 
               32'shd3f0c887, 32'shd3ee8142, 32'shd3ec3a18, 32'shd3e9f309, 32'shd3e7ac15, 32'shd3e5653c, 32'shd3e31e7f, 32'shd3e0d7dd, 
               32'shd3de9156, 32'shd3dc4aea, 32'shd3da049a, 32'shd3d7be64, 32'shd3d5784a, 32'shd3d3324b, 32'shd3d0ec68, 32'shd3cea69f, 
               32'shd3cc60f2, 32'shd3ca1b61, 32'shd3c7d5ea, 32'shd3c5908f, 32'shd3c34b4f, 32'shd3c1062a, 32'shd3bec121, 32'shd3bc7c33, 
               32'shd3ba3760, 32'shd3b7f2a9, 32'shd3b5ae0d, 32'shd3b3698c, 32'shd3b12526, 32'shd3aee0dc, 32'shd3ac9cad, 32'shd3aa589a, 
               32'shd3a814a2, 32'shd3a5d0c5, 32'shd3a38d03, 32'shd3a1495d, 32'shd39f05d3, 32'shd39cc263, 32'shd39a7f0f, 32'shd3983bd7, 
               32'shd395f8ba, 32'shd393b5b8, 32'shd39172d2, 32'shd38f3007, 32'shd38ced57, 32'shd38aaac3, 32'shd388684a, 32'shd38625ed, 
               32'shd383e3ab, 32'shd381a185, 32'shd37f5f7a, 32'shd37d1d8a, 32'shd37adbb6, 32'shd37899fe, 32'shd3765861, 32'shd37416df, 
               32'shd371d579, 32'shd36f942e, 32'shd36d52ff, 32'shd36b11eb, 32'shd368d0f3, 32'shd3669017, 32'shd3644f55, 32'shd3620eb0, 
               32'shd35fce26, 32'shd35d8db7, 32'shd35b4d64, 32'shd3590d2c, 32'shd356cd11, 32'shd3548d10, 32'shd3524d2b, 32'shd3500d62, 
               32'shd34dcdb4, 32'shd34b8e22, 32'shd3494eab, 32'shd3470f50, 32'shd344d011, 32'shd34290ed, 32'shd34051e5, 32'shd33e12f8, 
               32'shd33bd427, 32'shd3399572, 32'shd33756d8, 32'shd335185a, 32'shd332d9f7, 32'shd3309bb0, 32'shd32e5d85, 32'shd32c1f75, 
               32'shd329e181, 32'shd327a3a9, 32'shd32565ec, 32'shd323284b, 32'shd320eac6, 32'shd31ead5c, 32'shd31c700f, 32'shd31a32dc, 
               32'shd317f5c6, 32'shd315b8cb, 32'shd3137bec, 32'shd3113f28, 32'shd30f0280, 32'shd30cc5f4, 32'shd30a8984, 32'shd3084d30, 
               32'shd30610f7, 32'shd303d4da, 32'shd30198d8, 32'shd2ff5cf3, 32'shd2fd2129, 32'shd2fae57b, 32'shd2f8a9e9, 32'shd2f66e72, 
               32'shd2f43318, 32'shd2f1f7d9, 32'shd2efbcb6, 32'shd2ed81ae, 32'shd2eb46c3, 32'shd2e90bf3, 32'shd2e6d13f, 32'shd2e496a7, 
               32'shd2e25c2b, 32'shd2e021ca, 32'shd2dde786, 32'shd2dbad5d, 32'shd2d97350, 32'shd2d7395f, 32'shd2d4ff8a, 32'shd2d2c5d0, 
               32'shd2d08c33, 32'shd2ce52b1, 32'shd2cc194c, 32'shd2c9e002, 32'shd2c7a6d4, 32'shd2c56dc2, 32'shd2c334cc, 32'shd2c0fbf1, 
               32'shd2bec333, 32'shd2bc8a91, 32'shd2ba520a, 32'shd2b8199f, 32'shd2b5e151, 32'shd2b3a91e, 32'shd2b17107, 32'shd2af390d, 
               32'shd2ad012e, 32'shd2aac96b, 32'shd2a891c4, 32'shd2a65a39, 32'shd2a422ca, 32'shd2a1eb77, 32'shd29fb440, 32'shd29d7d25, 
               32'shd29b4626, 32'shd2990f43, 32'shd296d87c, 32'shd294a1d0, 32'shd2926b41, 32'shd29034ce, 32'shd28dfe77, 32'shd28bc83d, 
               32'shd289921e, 32'shd2875c1b, 32'shd2852634, 32'shd282f069, 32'shd280babb, 32'shd27e8528, 32'shd27c4fb1, 32'shd27a1a57, 
               32'shd277e518, 32'shd275aff6, 32'shd2737af0, 32'shd2714606, 32'shd26f1138, 32'shd26cdc86, 32'shd26aa7f0, 32'shd2687376, 
               32'shd2663f19, 32'shd2640ad7, 32'shd261d6b2, 32'shd25fa2a9, 32'shd25d6ebc, 32'shd25b3aeb, 32'shd2590736, 32'shd256d39e, 
               32'shd254a021, 32'shd2526cc1, 32'shd250397d, 32'shd24e0655, 32'shd24bd34a, 32'shd249a05a, 32'shd2476d87, 32'shd2453ad0, 
               32'shd2430835, 32'shd240d5b6, 32'shd23ea354, 32'shd23c710e, 32'shd23a3ee4, 32'shd2380cd6, 32'shd235dae4, 32'shd233a90f, 
               32'shd2317756, 32'shd22f45b9, 32'shd22d1439, 32'shd22ae2d5, 32'shd228b18d, 32'shd2268061, 32'shd2244f52, 32'shd2221e5f, 
               32'shd21fed88, 32'shd21dbccd, 32'shd21b8c2f, 32'shd2195bad, 32'shd2172b48, 32'shd214fafe, 32'shd212cad1, 32'shd2109ac1, 
               32'shd20e6acc, 32'shd20c3af4, 32'shd20a0b39, 32'shd207db9a, 32'shd205ac17, 32'shd2037cb0, 32'shd2014d66, 32'shd1ff1e38, 
               32'shd1fcef27, 32'shd1fac032, 32'shd1f89159, 32'shd1f6629d, 32'shd1f433fd, 32'shd1f2057a, 32'shd1efd713, 32'shd1eda8c8, 
               32'shd1eb7a9a, 32'shd1e94c88, 32'shd1e71e93, 32'shd1e4f0ba, 32'shd1e2c2fd, 32'shd1e0955d, 32'shd1de67da, 32'shd1dc3a73, 
               32'shd1da0d28, 32'shd1d7dffa, 32'shd1d5b2e8, 32'shd1d385f3, 32'shd1d1591a, 32'shd1cf2c5e, 32'shd1ccffbe, 32'shd1cad33b, 
               32'shd1c8a6d4, 32'shd1c67a8a, 32'shd1c44e5c, 32'shd1c2224b, 32'shd1bff656, 32'shd1bdca7e, 32'shd1bb9ec2, 32'shd1b97323, 
               32'shd1b747a0, 32'shd1b51c3a, 32'shd1b2f0f1, 32'shd1b0c5c4, 32'shd1ae9ab4, 32'shd1ac6fc0, 32'shd1aa44e9, 32'shd1a81a2e, 
               32'shd1a5ef90, 32'shd1a3c50f, 32'shd1a19aaa, 32'shd19f7062, 32'shd19d4636, 32'shd19b1c27, 32'shd198f235, 32'shd196c85f, 
               32'shd1949ea6, 32'shd1927509, 32'shd1904b89, 32'shd18e2226, 32'shd18bf8e0, 32'shd189cfb6, 32'shd187a6a8, 32'shd1857db8, 
               32'shd18354e4, 32'shd1812c2d, 32'shd17f0392, 32'shd17cdb14, 32'shd17ab2b3, 32'shd1788a6f, 32'shd1766247, 32'shd1743a3c, 
               32'shd172124d, 32'shd16fea7c, 32'shd16dc2c7, 32'shd16b9b2f, 32'shd16973b3, 32'shd1674c54, 32'shd1652512, 32'shd162fded, 
               32'shd160d6e5, 32'shd15eaff9, 32'shd15c892a, 32'shd15a6278, 32'shd1583be2, 32'shd156156a, 32'shd153ef0e, 32'shd151c8cf, 
               32'shd14fa2ad, 32'shd14d7ca7, 32'shd14b56be, 32'shd14930f3, 32'shd1470b44, 32'shd144e5b1, 32'shd142c03c, 32'shd1409ae3, 
               32'shd13e75a8, 32'shd13c5089, 32'shd13a2b87, 32'shd13806a2, 32'shd135e1d9, 32'shd133bd2e, 32'shd131989f, 32'shd12f742d, 
               32'shd12d4fd9, 32'shd12b2ba1, 32'shd1290786, 32'shd126e387, 32'shd124bfa6, 32'shd1229be2, 32'shd120783a, 32'shd11e54b0, 
               32'shd11c3142, 32'shd11a0df1, 32'shd117eabd, 32'shd115c7a7, 32'shd113a4ad, 32'shd11181d0, 32'shd10f5f10, 32'shd10d3c6d, 
               32'shd10b19e7, 32'shd108f77d, 32'shd106d531, 32'shd104b302, 32'shd10290f0, 32'shd1006efb, 32'shd0fe4d22, 32'shd0fc2b67, 
               32'shd0fa09c9, 32'shd0f7e848, 32'shd0f5c6e3, 32'shd0f3a59c, 32'shd0f18472, 32'shd0ef6365, 32'shd0ed4275, 32'shd0eb21a2, 
               32'shd0e900ec, 32'shd0e6e053, 32'shd0e4bfd7, 32'shd0e29f78, 32'shd0e07f36, 32'shd0de5f11, 32'shd0dc3f0a, 32'shd0da1f1f, 
               32'shd0d7ff51, 32'shd0d5dfa1, 32'shd0d3c00e, 32'shd0d1a097, 32'shd0cf813e, 32'shd0cd6202, 32'shd0cb42e3, 32'shd0c923e1, 
               32'shd0c704fd, 32'shd0c4e635, 32'shd0c2c78b, 32'shd0c0a8fe, 32'shd0be8a8d, 32'shd0bc6c3a, 32'shd0ba4e05, 32'shd0b82fec, 
               32'shd0b611f1, 32'shd0b3f412, 32'shd0b1d651, 32'shd0afb8ad, 32'shd0ad9b26, 32'shd0ab7dbd, 32'shd0a96070, 32'shd0a74341, 
               32'shd0a5262f, 32'shd0a3093a, 32'shd0a0ec63, 32'shd09ecfa8, 32'shd09cb30b, 32'shd09a968b, 32'shd0987a29, 32'shd0965de3, 
               32'shd09441bb, 32'shd09225b0, 32'shd09009c3, 32'shd08dedf2, 32'shd08bd23f, 32'shd089b6a9, 32'shd0879b31, 32'shd0857fd5, 
               32'shd0836497, 32'shd0814977, 32'shd07f2e73, 32'shd07d138d, 32'shd07af8c4, 32'shd078de19, 32'shd076c38b, 32'shd074a91a, 
               32'shd0728ec6, 32'shd0707490, 32'shd06e5a77, 32'shd06c407c, 32'shd06a269d, 32'shd0680cdd, 32'shd065f339, 32'shd063d9b3, 
               32'shd061c04a, 32'shd05fa6ff, 32'shd05d8dd1, 32'shd05b74c0, 32'shd0595bcd, 32'shd05742f7, 32'shd0552a3f, 32'shd05311a4, 
               32'shd050f926, 32'shd04ee0c6, 32'shd04cc884, 32'shd04ab05e, 32'shd0489856, 32'shd046806c, 32'shd044689f, 32'shd04250ef, 
               32'shd040395d, 32'shd03e21e8, 32'shd03c0a91, 32'shd039f357, 32'shd037dc3b, 32'shd035c53c, 32'shd033ae5b, 32'shd0319797, 
               32'shd02f80f1, 32'shd02d6a68, 32'shd02b53fc, 32'shd0293dae, 32'shd027277e, 32'shd025116b, 32'shd022fb76, 32'shd020e59e, 
               32'shd01ecfe4, 32'shd01cba47, 32'shd01aa4c8, 32'shd0188f66, 32'shd0167a22, 32'shd01464fc, 32'shd0124ff3, 32'shd0103b07, 
               32'shd00e2639, 32'shd00c1189, 32'shd009fcf6, 32'shd007e881, 32'shd005d42a, 32'shd003bff0, 32'shd001abd3, 32'shcfff97d5, 
               32'shcffd83f4, 32'shcffb7030, 32'shcff95c8a, 32'shcff74902, 32'shcff53597, 32'shcff3224a, 32'shcff10f1b, 32'shcfeefc09, 
               32'shcfece915, 32'shcfead63f, 32'shcfe8c386, 32'shcfe6b0eb, 32'shcfe49e6d, 32'shcfe28c0e, 32'shcfe079cc, 32'shcfde67a7, 
               32'shcfdc55a1, 32'shcfda43b8, 32'shcfd831ec, 32'shcfd6203f, 32'shcfd40eaf, 32'shcfd1fd3d, 32'shcfcfebe8, 32'shcfcddab2, 
               32'shcfcbc999, 32'shcfc9b89d, 32'shcfc7a7c0, 32'shcfc59700, 32'shcfc3865e, 32'shcfc175da, 32'shcfbf6573, 32'shcfbd552b, 
               32'shcfbb4500, 32'shcfb934f2, 32'shcfb72503, 32'shcfb51531, 32'shcfb3057d, 32'shcfb0f5e7, 32'shcfaee66f, 32'shcfacd715, 
               32'shcfaac7d8, 32'shcfa8b8b9, 32'shcfa6a9b8, 32'shcfa49ad5, 32'shcfa28c10, 32'shcfa07d68, 32'shcf9e6edf, 32'shcf9c6073, 
               32'shcf9a5225, 32'shcf9843f5, 32'shcf9635e2, 32'shcf9427ee, 32'shcf921a17, 32'shcf900c5f, 32'shcf8dfec4, 32'shcf8bf147, 
               32'shcf89e3e8, 32'shcf87d6a7, 32'shcf85c984, 32'shcf83bc7e, 32'shcf81af97, 32'shcf7fa2cd, 32'shcf7d9622, 32'shcf7b8994, 
               32'shcf797d24, 32'shcf7770d3, 32'shcf75649f, 32'shcf735889, 32'shcf714c91, 32'shcf6f40b7, 32'shcf6d34fb, 32'shcf6b295d, 
               32'shcf691ddd, 32'shcf67127a, 32'shcf650736, 32'shcf62fc10, 32'shcf60f108, 32'shcf5ee61e, 32'shcf5cdb51, 32'shcf5ad0a3, 
               32'shcf58c613, 32'shcf56bba1, 32'shcf54b14d, 32'shcf52a716, 32'shcf509cfe, 32'shcf4e9304, 32'shcf4c8928, 32'shcf4a7f6a, 
               32'shcf4875ca, 32'shcf466c48, 32'shcf4462e4, 32'shcf42599f, 32'shcf405077, 32'shcf3e476d, 32'shcf3c3e82, 32'shcf3a35b4, 
               32'shcf382d05, 32'shcf362473, 32'shcf341c00, 32'shcf3213ab, 32'shcf300b74, 32'shcf2e035b, 32'shcf2bfb60, 32'shcf29f383, 
               32'shcf27ebc5, 32'shcf25e424, 32'shcf23dca2, 32'shcf21d53e, 32'shcf1fcdf8, 32'shcf1dc6d0, 32'shcf1bbfc6, 32'shcf19b8db, 
               32'shcf17b20d, 32'shcf15ab5e, 32'shcf13a4cd, 32'shcf119e5a, 32'shcf0f9805, 32'shcf0d91cf, 32'shcf0b8bb7, 32'shcf0985bc, 
               32'shcf077fe1, 32'shcf057a23, 32'shcf037483, 32'shcf016f02, 32'shceff699f, 32'shcefd645a, 32'shcefb5f34, 32'shcef95a2b, 
               32'shcef75541, 32'shcef55075, 32'shcef34bc8, 32'shcef14738, 32'shceef42c7, 32'shceed3e74, 32'shceeb3a40, 32'shcee93629, 
               32'shcee73231, 32'shcee52e58, 32'shcee32a9c, 32'shcee126ff, 32'shcedf2380, 32'shcedd2020, 32'shcedb1cde, 32'shced919ba, 
               32'shced716b4, 32'shced513cd, 32'shced31104, 32'shced10e59, 32'shcecf0bcd, 32'shcecd095f, 32'shcecb070f, 32'shcec904de, 
               32'shcec702cb, 32'shcec500d7, 32'shcec2ff01, 32'shcec0fd49, 32'shcebefbb0, 32'shcebcfa35, 32'shcebaf8d8, 32'shceb8f79a, 
               32'shceb6f67a, 32'shceb4f579, 32'shceb2f496, 32'shceb0f3d1, 32'shceaef32b, 32'shceacf2a3, 32'shceaaf23a, 32'shcea8f1ef, 
               32'shcea6f1c2, 32'shcea4f1b4, 32'shcea2f1c5, 32'shcea0f1f4, 32'shce9ef241, 32'shce9cf2ad, 32'shce9af337, 32'shce98f3e0, 
               32'shce96f4a7, 32'shce94f58c, 32'shce92f691, 32'shce90f7b3, 32'shce8ef8f4, 32'shce8cfa54, 32'shce8afbd2, 32'shce88fd6f, 
               32'shce86ff2a, 32'shce850104, 32'shce8302fc, 32'shce810512, 32'shce7f0748, 32'shce7d099b, 32'shce7b0c0e, 32'shce790e9f, 
               32'shce77114e, 32'shce75141c, 32'shce731709, 32'shce711a14, 32'shce6f1d3d, 32'shce6d2086, 32'shce6b23ec, 32'shce692772, 
               32'shce672b16, 32'shce652ed8, 32'shce6332ba, 32'shce6136b9, 32'shce5f3ad8, 32'shce5d3f15, 32'shce5b4370, 32'shce5947eb, 
               32'shce574c84, 32'shce55513b, 32'shce535611, 32'shce515b06, 32'shce4f6019, 32'shce4d654c, 32'shce4b6a9c, 32'shce49700c, 
               32'shce47759a, 32'shce457b47, 32'shce438112, 32'shce4186fc, 32'shce3f8d05, 32'shce3d932c, 32'shce3b9973, 32'shce399fd7, 
               32'shce37a65b, 32'shce35acfd, 32'shce33b3be, 32'shce31ba9e, 32'shce2fc19c, 32'shce2dc8ba, 32'shce2bcff5, 32'shce29d750, 
               32'shce27dec9, 32'shce25e662, 32'shce23ee18, 32'shce21f5ee, 32'shce1ffde2, 32'shce1e05f6, 32'shce1c0e28, 32'shce1a1678, 
               32'shce181ee8, 32'shce162776, 32'shce143023, 32'shce1238ef, 32'shce1041d9, 32'shce0e4ae3, 32'shce0c540b, 32'shce0a5d52, 
               32'shce0866b8, 32'shce06703d, 32'shce0479e0, 32'shce0283a3, 32'shce008d84, 32'shcdfe9784, 32'shcdfca1a3, 32'shcdfaabe1, 
               32'shcdf8b63d, 32'shcdf6c0b9, 32'shcdf4cb53, 32'shcdf2d60c, 32'shcdf0e0e4, 32'shcdeeebdb, 32'shcdecf6f1, 32'shcdeb0226, 
               32'shcde90d79, 32'shcde718ec, 32'shcde5247d, 32'shcde3302e, 32'shcde13bfd, 32'shcddf47eb, 32'shcddd53f8, 32'shcddb6024, 
               32'shcdd96c6f, 32'shcdd778d9, 32'shcdd58562, 32'shcdd39209, 32'shcdd19ed0, 32'shcdcfabb6, 32'shcdcdb8ba, 32'shcdcbc5de, 
               32'shcdc9d320, 32'shcdc7e082, 32'shcdc5ee02, 32'shcdc3fba2, 32'shcdc20960, 32'shcdc0173e, 32'shcdbe253a, 32'shcdbc3356, 
               32'shcdba4190, 32'shcdb84fea, 32'shcdb65e62, 32'shcdb46cfa, 32'shcdb27bb0, 32'shcdb08a86, 32'shcdae997a, 32'shcdaca88e, 
               32'shcdaab7c0, 32'shcda8c712, 32'shcda6d683, 32'shcda4e613, 32'shcda2f5c2, 32'shcda10590, 32'shcd9f157d, 32'shcd9d2589, 
               32'shcd9b35b4, 32'shcd9945fe, 32'shcd975668, 32'shcd9566f0, 32'shcd937798, 32'shcd91885e, 32'shcd8f9944, 32'shcd8daa49, 
               32'shcd8bbb6d, 32'shcd89ccb0, 32'shcd87de12, 32'shcd85ef94, 32'shcd840134, 32'shcd8212f4, 32'shcd8024d3, 32'shcd7e36d1, 
               32'shcd7c48ee, 32'shcd7a5b2a, 32'shcd786d85, 32'shcd768000, 32'shcd74929a, 32'shcd72a553, 32'shcd70b82b, 32'shcd6ecb22, 
               32'shcd6cde39, 32'shcd6af16e, 32'shcd6904c3, 32'shcd671837, 32'shcd652bcb, 32'shcd633f7d, 32'shcd61534f, 32'shcd5f6740, 
               32'shcd5d7b50, 32'shcd5b8f80, 32'shcd59a3ce, 32'shcd57b83c, 32'shcd55ccca, 32'shcd53e176, 32'shcd51f642, 32'shcd500b2d, 
               32'shcd4e2037, 32'shcd4c3560, 32'shcd4a4aa9, 32'shcd486011, 32'shcd467599, 32'shcd448b3f, 32'shcd42a105, 32'shcd40b6ea, 
               32'shcd3eccef, 32'shcd3ce313, 32'shcd3af956, 32'shcd390fb8, 32'shcd37263a, 32'shcd353cdb, 32'shcd33539c, 32'shcd316a7b, 
               32'shcd2f817b, 32'shcd2d9899, 32'shcd2bafd7, 32'shcd29c734, 32'shcd27deb0, 32'shcd25f64c, 32'shcd240e08, 32'shcd2225e2, 
               32'shcd203ddc, 32'shcd1e55f6, 32'shcd1c6e2e, 32'shcd1a8687, 32'shcd189efe, 32'shcd16b795, 32'shcd14d04b, 32'shcd12e921, 
               32'shcd110216, 32'shcd0f1b2b, 32'shcd0d345f, 32'shcd0b4db3, 32'shcd096725, 32'shcd0780b8, 32'shcd059a6a, 32'shcd03b43b, 
               32'shcd01ce2b, 32'shccffe83c, 32'shccfe026b, 32'shccfc1cba, 32'shccfa3729, 32'shccf851b7, 32'shccf66c64, 32'shccf48731, 
               32'shccf2a21d, 32'shccf0bd29, 32'shcceed855, 32'shccecf3a0, 32'shcceb0f0a, 32'shcce92a94, 32'shcce7463e, 32'shcce56206, 
               32'shcce37def, 32'shcce199f7, 32'shccdfb61f, 32'shccddd266, 32'shccdbeecc, 32'shccda0b52, 32'shccd827f8, 32'shccd644bd, 
               32'shccd461a2, 32'shccd27ea7, 32'shccd09bcb, 32'shccceb90e, 32'shccccd671, 32'shcccaf3f4, 32'shccc91196, 32'shccc72f58, 
               32'shccc54d3a, 32'shccc36b3b, 32'shccc1895c, 32'shccbfa79c, 32'shccbdc5fc, 32'shccbbe47b, 32'shccba031a, 32'shccb821d9, 
               32'shccb640b8, 32'shccb45fb6, 32'shccb27ed3, 32'shccb09e11, 32'shccaebd6e, 32'shccacdcea, 32'shccaafc87, 32'shcca91c43, 
               32'shcca73c1e, 32'shcca55c1a, 32'shcca37c35, 32'shcca19c6f, 32'shcc9fbcca, 32'shcc9ddd44, 32'shcc9bfddd, 32'shcc9a1e97, 
               32'shcc983f70, 32'shcc966069, 32'shcc948182, 32'shcc92a2ba, 32'shcc90c412, 32'shcc8ee58a, 32'shcc8d0721, 32'shcc8b28d8, 
               32'shcc894aaf, 32'shcc876ca6, 32'shcc858ebc, 32'shcc83b0f3, 32'shcc81d349, 32'shcc7ff5be, 32'shcc7e1854, 32'shcc7c3b09, 
               32'shcc7a5dde, 32'shcc7880d3, 32'shcc76a3e8, 32'shcc74c71c, 32'shcc72ea70, 32'shcc710de4, 32'shcc6f3178, 32'shcc6d552c, 
               32'shcc6b78ff, 32'shcc699cf2, 32'shcc67c105, 32'shcc65e538, 32'shcc64098b, 32'shcc622dfd, 32'shcc605290, 32'shcc5e7742, 
               32'shcc5c9c14, 32'shcc5ac106, 32'shcc58e618, 32'shcc570b4a, 32'shcc55309b, 32'shcc53560c, 32'shcc517b9e, 32'shcc4fa14f, 
               32'shcc4dc720, 32'shcc4bed11, 32'shcc4a1322, 32'shcc483952, 32'shcc465fa3, 32'shcc448614, 32'shcc42aca4, 32'shcc40d354, 
               32'shcc3efa25, 32'shcc3d2115, 32'shcc3b4825, 32'shcc396f55, 32'shcc3796a5, 32'shcc35be15, 32'shcc33e5a5, 32'shcc320d55, 
               32'shcc303524, 32'shcc2e5d14, 32'shcc2c8524, 32'shcc2aad54, 32'shcc28d5a3, 32'shcc26fe13, 32'shcc2526a2, 32'shcc234f52, 
               32'shcc217822, 32'shcc1fa111, 32'shcc1dca21, 32'shcc1bf350, 32'shcc1a1ca0, 32'shcc184610, 32'shcc166f9f, 32'shcc14994f, 
               32'shcc12c31f, 32'shcc10ed0e, 32'shcc0f171e, 32'shcc0d414e, 32'shcc0b6b9e, 32'shcc09960e, 32'shcc07c09e, 32'shcc05eb4e, 
               32'shcc04161e, 32'shcc02410e, 32'shcc006c1e, 32'shcbfe974e, 32'shcbfcc29f, 32'shcbfaee0f, 32'shcbf919a0, 32'shcbf74550, 
               32'shcbf57121, 32'shcbf39d12, 32'shcbf1c923, 32'shcbeff554, 32'shcbee21a5, 32'shcbec4e16, 32'shcbea7aa7, 32'shcbe8a759, 
               32'shcbe6d42b, 32'shcbe5011c, 32'shcbe32e2e, 32'shcbe15b60, 32'shcbdf88b3, 32'shcbddb625, 32'shcbdbe3b7, 32'shcbda116a, 
               32'shcbd83f3d, 32'shcbd66d30, 32'shcbd49b43, 32'shcbd2c977, 32'shcbd0f7ca, 32'shcbcf263e, 32'shcbcd54d2, 32'shcbcb8386, 
               32'shcbc9b25a, 32'shcbc7e14f, 32'shcbc61064, 32'shcbc43f99, 32'shcbc26eee, 32'shcbc09e64, 32'shcbbecdf9, 32'shcbbcfdaf, 
               32'shcbbb2d85, 32'shcbb95d7c, 32'shcbb78d92, 32'shcbb5bdc9, 32'shcbb3ee20, 32'shcbb21e98, 32'shcbb04f2f, 32'shcbae7fe7, 
               32'shcbacb0bf, 32'shcbaae1b8, 32'shcba912d1, 32'shcba7440a, 32'shcba57563, 32'shcba3a6dd, 32'shcba1d877, 32'shcba00a31, 
               32'shcb9e3c0b, 32'shcb9c6e06, 32'shcb9aa021, 32'shcb98d25d, 32'shcb9704b9, 32'shcb953735, 32'shcb9369d1, 32'shcb919c8e, 
               32'shcb8fcf6b, 32'shcb8e0269, 32'shcb8c3587, 32'shcb8a68c5, 32'shcb889c23, 32'shcb86cfa2, 32'shcb850342, 32'shcb833701, 
               32'shcb816ae1, 32'shcb7f9ee2, 32'shcb7dd303, 32'shcb7c0744, 32'shcb7a3ba5, 32'shcb787027, 32'shcb76a4ca, 32'shcb74d98d, 
               32'shcb730e70, 32'shcb714373, 32'shcb6f7898, 32'shcb6daddc, 32'shcb6be341, 32'shcb6a18c6, 32'shcb684e6c, 32'shcb668432, 
               32'shcb64ba19, 32'shcb62f020, 32'shcb612648, 32'shcb5f5c90, 32'shcb5d92f8, 32'shcb5bc981, 32'shcb5a002b, 32'shcb5836f4, 
               32'shcb566ddf, 32'shcb54a4ea, 32'shcb52dc15, 32'shcb511361, 32'shcb4f4acd, 32'shcb4d825a, 32'shcb4bba08, 32'shcb49f1d5, 
               32'shcb4829c4, 32'shcb4661d3, 32'shcb449a02, 32'shcb42d252, 32'shcb410ac3, 32'shcb3f4354, 32'shcb3d7c05, 32'shcb3bb4d7, 
               32'shcb39edca, 32'shcb3826dd, 32'shcb366011, 32'shcb349965, 32'shcb32d2da, 32'shcb310c70, 32'shcb2f4626, 32'shcb2d7ffc, 
               32'shcb2bb9f4, 32'shcb29f40b, 32'shcb282e44, 32'shcb26689d, 32'shcb24a316, 32'shcb22ddb1, 32'shcb21186b, 32'shcb1f5347, 
               32'shcb1d8e43, 32'shcb1bc95f, 32'shcb1a049d, 32'shcb183ffb, 32'shcb167b79, 32'shcb14b718, 32'shcb12f2d8, 32'shcb112eb9, 
               32'shcb0f6aba, 32'shcb0da6dc, 32'shcb0be31e, 32'shcb0a1f81, 32'shcb085c05, 32'shcb0698a9, 32'shcb04d56e, 32'shcb031254, 
               32'shcb014f5b, 32'shcaff8c82, 32'shcafdc9ca, 32'shcafc0732, 32'shcafa44bc, 32'shcaf88266, 32'shcaf6c030, 32'shcaf4fe1c, 
               32'shcaf33c28, 32'shcaf17a55, 32'shcaefb8a2, 32'shcaedf711, 32'shcaec35a0, 32'shcaea744f, 32'shcae8b320, 32'shcae6f211, 
               32'shcae53123, 32'shcae37056, 32'shcae1afaa, 32'shcadfef1e, 32'shcade2eb3, 32'shcadc6e69, 32'shcadaae40, 32'shcad8ee37, 
               32'shcad72e4f, 32'shcad56e88, 32'shcad3aee2, 32'shcad1ef5d, 32'shcad02ff8, 32'shcace70b4, 32'shcaccb191, 32'shcacaf28f, 
               32'shcac933ae, 32'shcac774ed, 32'shcac5b64e, 32'shcac3f7cf, 32'shcac23971, 32'shcac07b34, 32'shcabebd17, 32'shcabcff1c, 
               32'shcabb4141, 32'shcab98388, 32'shcab7c5ef, 32'shcab60877, 32'shcab44b1f, 32'shcab28de9, 32'shcab0d0d4, 32'shcaaf13df, 
               32'shcaad570c, 32'shcaab9a59, 32'shcaa9ddc7, 32'shcaa82156, 32'shcaa66506, 32'shcaa4a8d7, 32'shcaa2ecc9, 32'shcaa130db, 
               32'shca9f750f, 32'shca9db964, 32'shca9bfdd9, 32'shca9a4270, 32'shca988727, 32'shca96cbff, 32'shca9510f8, 32'shca935613, 
               32'shca919b4e, 32'shca8fe0aa, 32'shca8e2627, 32'shca8c6bc5, 32'shca8ab184, 32'shca88f764, 32'shca873d65, 32'shca858387, 
               32'shca83c9ca, 32'shca82102e, 32'shca8056b3, 32'shca7e9d59, 32'shca7ce420, 32'shca7b2b08, 32'shca797211, 32'shca77b93b, 
               32'shca760086, 32'shca7447f2, 32'shca728f7f, 32'shca70d72d, 32'shca6f1efc, 32'shca6d66ec, 32'shca6baefd, 32'shca69f72f, 
               32'shca683f83, 32'shca6687f7, 32'shca64d08d, 32'shca631943, 32'shca61621b, 32'shca5fab13, 32'shca5df42d, 32'shca5c3d68, 
               32'shca5a86c4, 32'shca58d041, 32'shca5719df, 32'shca55639e, 32'shca53ad7e, 32'shca51f780, 32'shca5041a2, 32'shca4e8be6, 
               32'shca4cd64b, 32'shca4b20d0, 32'shca496b77, 32'shca47b640, 32'shca460129, 32'shca444c33, 32'shca42975f, 32'shca40e2ac, 
               32'shca3f2e19, 32'shca3d79a8, 32'shca3bc559, 32'shca3a112a, 32'shca385d1d, 32'shca36a930, 32'shca34f565, 32'shca3341bb, 
               32'shca318e32, 32'shca2fdacb, 32'shca2e2784, 32'shca2c745f, 32'shca2ac15b, 32'shca290e79, 32'shca275bb7, 32'shca25a917, 
               32'shca23f698, 32'shca22443a, 32'shca2091fd, 32'shca1edfe2, 32'shca1d2de7, 32'shca1b7c0e, 32'shca19ca57, 32'shca1818c0, 
               32'shca16674b, 32'shca14b5f7, 32'shca1304c4, 32'shca1153b3, 32'shca0fa2c3, 32'shca0df1f4, 32'shca0c4146, 32'shca0a90ba, 
               32'shca08e04f, 32'shca073005, 32'shca057fdd, 32'shca03cfd5, 32'shca021fef, 32'shca00702b, 32'shc9fec088, 32'shc9fd1106, 
               32'shc9fb61a5, 32'shc9f9b266, 32'shc9f80348, 32'shc9f6544b, 32'shc9f4a570, 32'shc9f2f6b6, 32'shc9f1481d, 32'shc9ef99a6, 
               32'shc9edeb50, 32'shc9ec3d1b, 32'shc9ea8f08, 32'shc9e8e116, 32'shc9e73346, 32'shc9e58596, 32'shc9e3d809, 32'shc9e22a9c, 
               32'shc9e07d51, 32'shc9ded028, 32'shc9dd231f, 32'shc9db7639, 32'shc9d9c973, 32'shc9d81ccf, 32'shc9d6704c, 32'shc9d4c3eb, 
               32'shc9d317ab, 32'shc9d16b8d, 32'shc9cfbf90, 32'shc9ce13b4, 32'shc9cc67fa, 32'shc9cabc62, 32'shc9c910ea, 32'shc9c76595, 
               32'shc9c5ba60, 32'shc9c40f4d, 32'shc9c2645c, 32'shc9c0b98c, 32'shc9bf0edd, 32'shc9bd6450, 32'shc9bbb9e5, 32'shc9ba0f9b, 
               32'shc9b86572, 32'shc9b6bb6b, 32'shc9b51185, 32'shc9b367c1, 32'shc9b1be1e, 32'shc9b0149d, 32'shc9ae6b3d, 32'shc9acc1ff, 
               32'shc9ab18e3, 32'shc9a96fe7, 32'shc9a7c70e, 32'shc9a61e56, 32'shc9a475bf, 32'shc9a2cd4a, 32'shc9a124f7, 32'shc99f7cc5, 
               32'shc99dd4b4, 32'shc99c2cc5, 32'shc99a84f8, 32'shc998dd4c, 32'shc99735c2, 32'shc9958e59, 32'shc993e712, 32'shc9923fed, 
               32'shc99098e9, 32'shc98ef206, 32'shc98d4b45, 32'shc98ba4a6, 32'shc989fe29, 32'shc98857cd, 32'shc986b192, 32'shc9850b79, 
               32'shc9836582, 32'shc981bfac, 32'shc98019f8, 32'shc97e7466, 32'shc97ccef5, 32'shc97b29a6, 32'shc9798479, 32'shc977df6d, 
               32'shc9763a83, 32'shc97495ba, 32'shc972f113, 32'shc9714c8e, 32'shc96fa82a, 32'shc96e03e8, 32'shc96c5fc8, 32'shc96abbc9, 
               32'shc96917ec, 32'shc9677431, 32'shc965d097, 32'shc9642d1f, 32'shc96289c9, 32'shc960e695, 32'shc95f4382, 32'shc95da090, 
               32'shc95bfdc1, 32'shc95a5b13, 32'shc958b887, 32'shc957161d, 32'shc95573d4, 32'shc953d1ad, 32'shc9522fa8, 32'shc9508dc5, 
               32'shc94eec03, 32'shc94d4a63, 32'shc94ba8e5, 32'shc94a0788, 32'shc948664d, 32'shc946c534, 32'shc945243d, 32'shc9438368, 
               32'shc941e2b4, 32'shc9404222, 32'shc93ea1b2, 32'shc93d0163, 32'shc93b6137, 32'shc939c12c, 32'shc9382143, 32'shc936817b, 
               32'shc934e1d6, 32'shc9334252, 32'shc931a2f0, 32'shc93003b0, 32'shc92e6492, 32'shc92cc596, 32'shc92b26bb, 32'shc9298802, 
               32'shc927e96b, 32'shc9264af6, 32'shc924aca3, 32'shc9230e71, 32'shc9217062, 32'shc91fd274, 32'shc91e34a8, 32'shc91c96fe, 
               32'shc91af976, 32'shc9195c0f, 32'shc917becb, 32'shc91621a8, 32'shc91484a8, 32'shc912e7c9, 32'shc9114b0c, 32'shc90fae71, 
               32'shc90e11f7, 32'shc90c75a0, 32'shc90ad96b, 32'shc9093d57, 32'shc907a166, 32'shc9060596, 32'shc90469e8, 32'shc902ce5c, 
               32'shc90132f2, 32'shc8ff97aa, 32'shc8fdfc84, 32'shc8fc6180, 32'shc8fac69e, 32'shc8f92bdd, 32'shc8f7913f, 32'shc8f5f6c3, 
               32'shc8f45c68, 32'shc8f2c230, 32'shc8f12819, 32'shc8ef8e24, 32'shc8edf452, 32'shc8ec5aa1, 32'shc8eac112, 32'shc8e927a6, 
               32'shc8e78e5b, 32'shc8e5f532, 32'shc8e45c2c, 32'shc8e2c347, 32'shc8e12a84, 32'shc8df91e3, 32'shc8ddf965, 32'shc8dc6108, 
               32'shc8dac8cd, 32'shc8d930b4, 32'shc8d798be, 32'shc8d600e9, 32'shc8d46936, 32'shc8d2d1a6, 32'shc8d13a37, 32'shc8cfa2eb, 
               32'shc8ce0bc0, 32'shc8cc74b8, 32'shc8caddd1, 32'shc8c9470d, 32'shc8c7b06b, 32'shc8c619eb, 32'shc8c4838d, 32'shc8c2ed50, 
               32'shc8c15736, 32'shc8bfc13f, 32'shc8be2b69, 32'shc8bc95b5, 32'shc8bb0023, 32'shc8b96ab4, 32'shc8b7d566, 32'shc8b6403b, 
               32'shc8b4ab32, 32'shc8b3164a, 32'shc8b18185, 32'shc8afece2, 32'shc8ae5862, 32'shc8acc403, 32'shc8ab2fc6, 32'shc8a99bac, 
               32'shc8a807b4, 32'shc8a673dd, 32'shc8a4e029, 32'shc8a34c98, 32'shc8a1b928, 32'shc8a025da, 32'shc89e92af, 32'shc89cffa6, 
               32'shc89b6cbf, 32'shc899d9fa, 32'shc8984757, 32'shc896b4d6, 32'shc8952278, 32'shc893903c, 32'shc891fe22, 32'shc8906c2a, 
               32'shc88eda54, 32'shc88d48a1, 32'shc88bb710, 32'shc88a25a1, 32'shc8889454, 32'shc8870329, 32'shc8857221, 32'shc883e13b, 
               32'shc8825077, 32'shc880bfd5, 32'shc87f2f56, 32'shc87d9ef8, 32'shc87c0ebd, 32'shc87a7ea5, 32'shc878eeae, 32'shc8775eda, 
               32'shc875cf28, 32'shc8743f98, 32'shc872b02b, 32'shc87120e0, 32'shc86f91b7, 32'shc86e02b0, 32'shc86c73cc, 32'shc86ae50a, 
               32'shc869566a, 32'shc867c7ec, 32'shc8663991, 32'shc864ab58, 32'shc8631d42, 32'shc8618f4d, 32'shc860017b, 32'shc85e73cc, 
               32'shc85ce63e, 32'shc85b58d3, 32'shc859cb8a, 32'shc8583e64, 32'shc856b160, 32'shc855247e, 32'shc85397bf, 32'shc8520b22, 
               32'shc8507ea7, 32'shc84ef24f, 32'shc84d6619, 32'shc84bda05, 32'shc84a4e14, 32'shc848c245, 32'shc8473698, 32'shc845ab0e, 
               32'shc8441fa6, 32'shc8429461, 32'shc841093e, 32'shc83f7e3d, 32'shc83df35f, 32'shc83c68a3, 32'shc83ade0a, 32'shc8395393, 
               32'shc837c93e, 32'shc8363f0c, 32'shc834b4fc, 32'shc8332b0e, 32'shc831a143, 32'shc830179b, 32'shc82e8e15, 32'shc82d04b1, 
               32'shc82b7b70, 32'shc829f251, 32'shc8286954, 32'shc826e07a, 32'shc82557c3, 32'shc823cf2e, 32'shc82246bb, 32'shc820be6b, 
               32'shc81f363d, 32'shc81dae32, 32'shc81c2649, 32'shc81a9e83, 32'shc81916df, 32'shc8178f5e, 32'shc81607ff, 32'shc81480c3, 
               32'shc812f9a9, 32'shc81172b2, 32'shc80febdd, 32'shc80e652b, 32'shc80cde9b, 32'shc80b582e, 32'shc809d1e3, 32'shc8084bba, 
               32'shc806c5b5, 32'shc8053fd2, 32'shc803ba11, 32'shc8023473, 32'shc800aef7, 32'shc7ff299e, 32'shc7fda468, 32'shc7fc1f54, 
               32'shc7fa9a62, 32'shc7f91593, 32'shc7f790e7, 32'shc7f60c5d, 32'shc7f487f6, 32'shc7f303b1, 32'shc7f17f8f, 32'shc7effb90, 
               32'shc7ee77b3, 32'shc7ecf3f9, 32'shc7eb7061, 32'shc7e9ecec, 32'shc7e8699a, 32'shc7e6e66a, 32'shc7e5635c, 32'shc7e3e072, 
               32'shc7e25daa, 32'shc7e0db04, 32'shc7df5881, 32'shc7ddd621, 32'shc7dc53e3, 32'shc7dad1c9, 32'shc7d94fd0, 32'shc7d7cdfb, 
               32'shc7d64c47, 32'shc7d4cab7, 32'shc7d34949, 32'shc7d1c7fe, 32'shc7d046d6, 32'shc7cec5d0, 32'shc7cd44ed, 32'shc7cbc42c, 
               32'shc7ca438f, 32'shc7c8c313, 32'shc7c742bb, 32'shc7c5c285, 32'shc7c44272, 32'shc7c2c282, 32'shc7c142b4, 32'shc7bfc309, 
               32'shc7be4381, 32'shc7bcc41b, 32'shc7bb44d8, 32'shc7b9c5b8, 32'shc7b846ba, 32'shc7b6c7e0, 32'shc7b54928, 32'shc7b3ca92, 
               32'shc7b24c20, 32'shc7b0cdd0, 32'shc7af4fa3, 32'shc7add198, 32'shc7ac53b1, 32'shc7aad5ec, 32'shc7a9584a, 32'shc7a7daca, 
               32'shc7a65d6e, 32'shc7a4e034, 32'shc7a3631d, 32'shc7a1e628, 32'shc7a06957, 32'shc79eeca8, 32'shc79d701c, 32'shc79bf3b3, 
               32'shc79a776c, 32'shc798fb48, 32'shc7977f48, 32'shc7960369, 32'shc79487ae, 32'shc7930c16, 32'shc79190a0, 32'shc790154d, 
               32'shc78e9a1d, 32'shc78d1f10, 32'shc78ba425, 32'shc78a295e, 32'shc788aeb9, 32'shc7873437, 32'shc785b9d8, 32'shc7843f9c, 
               32'shc782c582, 32'shc7814b8c, 32'shc77fd1b8, 32'shc77e5807, 32'shc77cde79, 32'shc77b650e, 32'shc779ebc5, 32'shc77872a0, 
               32'shc776f99d, 32'shc77580be, 32'shc7740801, 32'shc7728f67, 32'shc77116f0, 32'shc76f9e9c, 32'shc76e266b, 32'shc76cae5c, 
               32'shc76b3671, 32'shc769bea8, 32'shc7684702, 32'shc766cf80, 32'shc7655820, 32'shc763e0e3, 32'shc76269c9, 32'shc760f2d2, 
               32'shc75f7bfe, 32'shc75e054c, 32'shc75c8ebe, 32'shc75b1853, 32'shc759a20a, 32'shc7582be5, 32'shc756b5e2, 32'shc7554003, 
               32'shc753ca46, 32'shc75254ac, 32'shc750df36, 32'shc74f69e2, 32'shc74df4b1, 32'shc74c7fa4, 32'shc74b0ab9, 32'shc74995f1, 
               32'shc748214c, 32'shc746acca, 32'shc745386b, 32'shc743c42f, 32'shc7425016, 32'shc740dc21, 32'shc73f684e, 32'shc73df49e, 
               32'shc73c8111, 32'shc73b0da7, 32'shc7399a60, 32'shc738273d, 32'shc736b43c, 32'shc735415e, 32'shc733cea3, 32'shc7325c0c, 
               32'shc730e997, 32'shc72f7745, 32'shc72e0517, 32'shc72c930b, 32'shc72b2123, 32'shc729af5d, 32'shc7283dbb, 32'shc726cc3c, 
               32'shc7255ae0, 32'shc723e9a6, 32'shc7227890, 32'shc721079d, 32'shc71f96ce, 32'shc71e2621, 32'shc71cb597, 32'shc71b4530, 
               32'shc719d4ed, 32'shc71864cc, 32'shc716f4cf, 32'shc71584f5, 32'shc714153e, 32'shc712a5aa, 32'shc7113639, 32'shc70fc6eb, 
               32'shc70e57c0, 32'shc70ce8b9, 32'shc70b79d4, 32'shc70a0b13, 32'shc7089c75, 32'shc7072dfa, 32'shc705bfa2, 32'shc704516d, 
               32'shc702e35c, 32'shc701756d, 32'shc70007a2, 32'shc6fe99fa, 32'shc6fd2c75, 32'shc6fbbf13, 32'shc6fa51d5, 32'shc6f8e4b9, 
               32'shc6f777c1, 32'shc6f60aec, 32'shc6f49e3a, 32'shc6f331ab, 32'shc6f1c540, 32'shc6f058f8, 32'shc6eeecd3, 32'shc6ed80d1, 
               32'shc6ec14f2, 32'shc6eaa936, 32'shc6e93d9e, 32'shc6e7d229, 32'shc6e666d7, 32'shc6e4fba9, 32'shc6e3909d, 32'shc6e225b5, 
               32'shc6e0baf0, 32'shc6df504f, 32'shc6dde5d0, 32'shc6dc7b75, 32'shc6db113d, 32'shc6d9a728, 32'shc6d83d37, 32'shc6d6d369, 
               32'shc6d569be, 32'shc6d40036, 32'shc6d296d1, 32'shc6d12d90, 32'shc6cfc472, 32'shc6ce5b78, 32'shc6ccf2a1, 32'shc6cb89ed, 
               32'shc6ca215c, 32'shc6c8b8ee, 32'shc6c750a4, 32'shc6c5e87d, 32'shc6c4807a, 32'shc6c31899, 32'shc6c1b0dd, 32'shc6c04943, 
               32'shc6bee1cd, 32'shc6bd7a7a, 32'shc6bc134a, 32'shc6baac3d, 32'shc6b94554, 32'shc6b7de8f, 32'shc6b677ec, 32'shc6b5116d, 
               32'shc6b3ab12, 32'shc6b244d9, 32'shc6b0dec4, 32'shc6af78d3, 32'shc6ae1304, 32'shc6acad59, 32'shc6ab47d2, 32'shc6a9e26e, 
               32'shc6a87d2d, 32'shc6a7180f, 32'shc6a5b315, 32'shc6a44e3e, 32'shc6a2e98b, 32'shc6a184fb, 32'shc6a0208f, 32'shc69ebc45, 
               32'shc69d5820, 32'shc69bf41d, 32'shc69a903e, 32'shc6992c83, 32'shc697c8eb, 32'shc6966576, 32'shc6950224, 32'shc6939ef6, 
               32'shc6923bec, 32'shc690d905, 32'shc68f7641, 32'shc68e13a1, 32'shc68cb124, 32'shc68b4ecb, 32'shc689ec95, 32'shc6888a83, 
               32'shc6872894, 32'shc685c6c8, 32'shc6846520, 32'shc683039b, 32'shc681a23a, 32'shc68040fc, 32'shc67edfe2, 32'shc67d7eeb, 
               32'shc67c1e18, 32'shc67abd68, 32'shc6795cdc, 32'shc677fc73, 32'shc6769c2e, 32'shc6753c0c, 32'shc673dc0d, 32'shc6727c32, 
               32'shc6711c7b, 32'shc66fbce7, 32'shc66e5d77, 32'shc66cfe2a, 32'shc66b9f01, 32'shc66a3ffb, 32'shc668e119, 32'shc667825a, 
               32'shc66623be, 32'shc664c547, 32'shc66366f3, 32'shc66208c2, 32'shc660aab5, 32'shc65f4ccb, 32'shc65def05, 32'shc65c9163, 
               32'shc65b33e4, 32'shc659d688, 32'shc6587951, 32'shc6571c3c, 32'shc655bf4c, 32'shc654627f, 32'shc65305d5, 32'shc651a94f, 
               32'shc6504ced, 32'shc64ef0ae, 32'shc64d9493, 32'shc64c389b, 32'shc64adcc7, 32'shc6498117, 32'shc648258a, 32'shc646ca21, 
               32'shc6456edb, 32'shc64413b9, 32'shc642b8bb, 32'shc6415de0, 32'shc6400329, 32'shc63ea896, 32'shc63d4e26, 32'shc63bf3d9, 
               32'shc63a99b1, 32'shc6393fac, 32'shc637e5ca, 32'shc6368c0d, 32'shc6353273, 32'shc633d8fc, 32'shc6327faa, 32'shc631267a, 
               32'shc62fcd6f, 32'shc62e7487, 32'shc62d1bc3, 32'shc62bc323, 32'shc62a6aa6, 32'shc629124d, 32'shc627ba17, 32'shc6266206, 
               32'shc6250a18, 32'shc623b24d, 32'shc6225aa6, 32'shc6210323, 32'shc61fabc4, 32'shc61e5489, 32'shc61cfd71, 32'shc61ba67d, 
               32'shc61a4fac, 32'shc618f8ff, 32'shc617a276, 32'shc6164c11, 32'shc614f5cf, 32'shc6139fb2, 32'shc61249b7, 32'shc610f3e1, 
               32'shc60f9e2e, 32'shc60e489f, 32'shc60cf334, 32'shc60b9ded, 32'shc60a48c9, 32'shc608f3c9, 32'shc6079eed, 32'shc6064a35, 
               32'shc604f5a0, 32'shc603a12f, 32'shc6024ce2, 32'shc600f8b9, 32'shc5ffa4b3, 32'shc5fe50d1, 32'shc5fcfd13, 32'shc5fba979, 
               32'shc5fa5603, 32'shc5f902b0, 32'shc5f7af81, 32'shc5f65c76, 32'shc5f5098f, 32'shc5f3b6cb, 32'shc5f2642c, 32'shc5f111b0, 
               32'shc5efbf58, 32'shc5ee6d24, 32'shc5ed1b13, 32'shc5ebc927, 32'shc5ea775e, 32'shc5e925b9, 32'shc5e7d438, 32'shc5e682db, 
               32'shc5e531a1, 32'shc5e3e08c, 32'shc5e28f9a, 32'shc5e13ecc, 32'shc5dfee22, 32'shc5de9d9c, 32'shc5dd4d3a, 32'shc5dbfcfb, 
               32'shc5daace1, 32'shc5d95cea, 32'shc5d80d17, 32'shc5d6bd68, 32'shc5d56ddd, 32'shc5d41e76, 32'shc5d2cf33, 32'shc5d18013, 
               32'shc5d03118, 32'shc5cee240, 32'shc5cd938c, 32'shc5cc44fc, 32'shc5caf690, 32'shc5c9a848, 32'shc5c85a24, 32'shc5c70c24, 
               32'shc5c5be47, 32'shc5c4708f, 32'shc5c322fb, 32'shc5c1d58a, 32'shc5c0883d, 32'shc5bf3b15, 32'shc5bdee10, 32'shc5bca12f, 
               32'shc5bb5472, 32'shc5ba07d9, 32'shc5b8bb64, 32'shc5b76f13, 32'shc5b622e6, 32'shc5b4d6dd, 32'shc5b38af8, 32'shc5b23f37, 
               32'shc5b0f399, 32'shc5afa820, 32'shc5ae5ccb, 32'shc5ad1199, 32'shc5abc68c, 32'shc5aa7ba3, 32'shc5a930dd, 32'shc5a7e63c, 
               32'shc5a69bbe, 32'shc5a55165, 32'shc5a4072f, 32'shc5a2bd1e, 32'shc5a17330, 32'shc5a02967, 32'shc59edfc2, 32'shc59d9640, 
               32'shc59c4ce3, 32'shc59b03a9, 32'shc599ba94, 32'shc59871a3, 32'shc59728d5, 32'shc595e02c, 32'shc59497a7, 32'shc5934f46, 
               32'shc5920708, 32'shc590beef, 32'shc58f76fa, 32'shc58e2f29, 32'shc58ce77c, 32'shc58b9ff3, 32'shc58a588e, 32'shc589114e, 
               32'shc587ca31, 32'shc5868338, 32'shc5853c63, 32'shc583f5b3, 32'shc582af26, 32'shc58168be, 32'shc580227a, 32'shc57edc5a, 
               32'shc57d965d, 32'shc57c5085, 32'shc57b0ad1, 32'shc579c542, 32'shc5787fd6, 32'shc5773a8e, 32'shc575f56b, 32'shc574b06b, 
               32'shc5736b90, 32'shc57226d9, 32'shc570e246, 32'shc56f9dd7, 32'shc56e598c, 32'shc56d1565, 32'shc56bd163, 32'shc56a8d84, 
               32'shc56949ca, 32'shc5680634, 32'shc566c2c2, 32'shc5657f74, 32'shc5643c4a, 32'shc562f944, 32'shc561b663, 32'shc56073a6, 
               32'shc55f310d, 32'shc55dee98, 32'shc55cac47, 32'shc55b6a1a, 32'shc55a2812, 32'shc558e62e, 32'shc557a46e, 32'shc55662d2, 
               32'shc555215a, 32'shc553e007, 32'shc5529ed7, 32'shc5515dcc, 32'shc5501ce5, 32'shc54edc23, 32'shc54d9b84, 32'shc54c5b0a, 
               32'shc54b1ab4, 32'shc549da82, 32'shc5489a74, 32'shc5475a8b, 32'shc5461ac6, 32'shc544db25, 32'shc5439ba8, 32'shc5425c4f, 
               32'shc5411d1b, 32'shc53fde0b, 32'shc53e9f1f, 32'shc53d6057, 32'shc53c21b4, 32'shc53ae335, 32'shc539a4da, 32'shc53866a4, 
               32'shc5372891, 32'shc535eaa3, 32'shc534acd9, 32'shc5336f34, 32'shc53231b3, 32'shc530f456, 32'shc52fb71d, 32'shc52e7a09, 
               32'shc52d3d18, 32'shc52c004d, 32'shc52ac3a5, 32'shc5298722, 32'shc5284ac3, 32'shc5270e88, 32'shc525d272, 32'shc5249680, 
               32'shc5235ab2, 32'shc5221f08, 32'shc520e383, 32'shc51fa822, 32'shc51e6ce6, 32'shc51d31ce, 32'shc51bf6da, 32'shc51abc0a, 
               32'shc519815f, 32'shc51846d8, 32'shc5170c75, 32'shc515d237, 32'shc514981d, 32'shc5135e28, 32'shc5122457, 32'shc510eaaa, 
               32'shc50fb121, 32'shc50e77bd, 32'shc50d3e7d, 32'shc50c0562, 32'shc50acc6b, 32'shc5099398, 32'shc5085aea, 32'shc5072260, 
               32'shc505e9fb, 32'shc504b1b9, 32'shc503799d, 32'shc50241a4, 32'shc50109d0, 32'shc4ffd221, 32'shc4fe9a95, 32'shc4fd632f, 
               32'shc4fc2bec, 32'shc4faf4ce, 32'shc4f9bdd4, 32'shc4f886ff, 32'shc4f7504e, 32'shc4f619c2, 32'shc4f4e35a, 32'shc4f3ad17, 
               32'shc4f276f7, 32'shc4f140fd, 32'shc4f00b27, 32'shc4eed575, 32'shc4ed9fe7, 32'shc4ec6a7e, 32'shc4eb353a, 32'shc4ea001a, 
               32'shc4e8cb1e, 32'shc4e79647, 32'shc4e66194, 32'shc4e52d06, 32'shc4e3f89c, 32'shc4e2c457, 32'shc4e19036, 32'shc4e05c3a, 
               32'shc4df2862, 32'shc4ddf4ae, 32'shc4dcc11f, 32'shc4db8db5, 32'shc4da5a6f, 32'shc4d9274d, 32'shc4d7f450, 32'shc4d6c177, 
               32'shc4d58ec3, 32'shc4d45c34, 32'shc4d329c9, 32'shc4d1f782, 32'shc4d0c560, 32'shc4cf9363, 32'shc4ce6189, 32'shc4cd2fd5, 
               32'shc4cbfe45, 32'shc4caccd9, 32'shc4c99b92, 32'shc4c86a70, 32'shc4c73972, 32'shc4c60899, 32'shc4c4d7e4, 32'shc4c3a753, 
               32'shc4c276e8, 32'shc4c146a0, 32'shc4c0167e, 32'shc4bee680, 32'shc4bdb6a6, 32'shc4bc86f1, 32'shc4bb5760, 32'shc4ba27f5, 
               32'shc4b8f8ad, 32'shc4b7c98a, 32'shc4b69a8c, 32'shc4b56bb3, 32'shc4b43cfd, 32'shc4b30e6d, 32'shc4b1e001, 32'shc4b0b1ba, 
               32'shc4af8397, 32'shc4ae5599, 32'shc4ad27bf, 32'shc4abfa0a, 32'shc4aacc7a, 32'shc4a99f0e, 32'shc4a871c7, 32'shc4a744a4, 
               32'shc4a617a6, 32'shc4a4eacd, 32'shc4a3be18, 32'shc4a29188, 32'shc4a1651c, 32'shc4a038d6, 32'shc49f0cb3, 32'shc49de0b6, 
               32'shc49cb4dd, 32'shc49b8928, 32'shc49a5d98, 32'shc499322d, 32'shc49806e7, 32'shc496dbc5, 32'shc495b0c8, 32'shc49485ef, 
               32'shc4935b3c, 32'shc49230ac, 32'shc4910642, 32'shc48fdbfc, 32'shc48eb1db, 32'shc48d87de, 32'shc48c5e06, 32'shc48b3453, 
               32'shc48a0ac4, 32'shc488e15b, 32'shc487b815, 32'shc4868ef5, 32'shc48565f9, 32'shc4843d22, 32'shc4831470, 32'shc481ebe2, 
               32'shc480c379, 32'shc47f9b34, 32'shc47e7315, 32'shc47d4b1a, 32'shc47c2344, 32'shc47afb92, 32'shc479d405, 32'shc478ac9d, 
               32'shc477855a, 32'shc4765e3b, 32'shc4753741, 32'shc474106c, 32'shc472e9bc, 32'shc471c330, 32'shc4709cc9, 32'shc46f7687, 
               32'shc46e5069, 32'shc46d2a71, 32'shc46c049d, 32'shc46adeee, 32'shc469b963, 32'shc46893fd, 32'shc4676ebc, 32'shc46649a0, 
               32'shc46524a9, 32'shc463ffd6, 32'shc462db28, 32'shc461b69f, 32'shc460923b, 32'shc45f6dfb, 32'shc45e49e0, 32'shc45d25ea, 
               32'shc45c0219, 32'shc45ade6c, 32'shc459bae5, 32'shc4589782, 32'shc4577444, 32'shc456512b, 32'shc4552e36, 32'shc4540b67, 
               32'shc452e8bc, 32'shc451c636, 32'shc450a3d4, 32'shc44f8198, 32'shc44e5f80, 32'shc44d3d8e, 32'shc44c1bc0, 32'shc44afa17, 
               32'shc449d892, 32'shc448b733, 32'shc44795f8, 32'shc44674e3, 32'shc44553f2, 32'shc4443326, 32'shc443127e, 32'shc441f1fc, 
               32'shc440d19e, 32'shc43fb166, 32'shc43e9152, 32'shc43d7163, 32'shc43c5199, 32'shc43b31f4, 32'shc43a1273, 32'shc438f318, 
               32'shc437d3e1, 32'shc436b4cf, 32'shc43595e3, 32'shc434771b, 32'shc4335877, 32'shc43239f9, 32'shc4311ba0, 32'shc42ffd6b, 
               32'shc42edf5c, 32'shc42dc171, 32'shc42ca3ac, 32'shc42b860b, 32'shc42a688f, 32'shc4294b38, 32'shc4282e06, 32'shc42710f9, 
               32'shc425f410, 32'shc424d74d, 32'shc423baae, 32'shc4229e35, 32'shc42181e0, 32'shc42065b1, 32'shc41f49a6, 32'shc41e2dc0, 
               32'shc41d11ff, 32'shc41bf664, 32'shc41adaed, 32'shc419bf9b, 32'shc418a46d, 32'shc4178965, 32'shc4166e82, 32'shc41553c4, 
               32'shc414392b, 32'shc4131eb7, 32'shc4120467, 32'shc410ea3d, 32'shc40fd037, 32'shc40eb657, 32'shc40d9c9c, 32'shc40c8305, 
               32'shc40b6994, 32'shc40a5047, 32'shc4093720, 32'shc4081e1d, 32'shc4070540, 32'shc405ec87, 32'shc404d3f4, 32'shc403bb85, 
               32'shc402a33c, 32'shc4018b17, 32'shc4007318, 32'shc3ff5b3d, 32'shc3fe4388, 32'shc3fd2bf7, 32'shc3fc148c, 32'shc3fafd45, 
               32'shc3f9e624, 32'shc3f8cf27, 32'shc3f7b850, 32'shc3f6a19e, 32'shc3f58b10, 32'shc3f474a8, 32'shc3f35e65, 32'shc3f24847, 
               32'shc3f1324e, 32'shc3f01c7a, 32'shc3ef06cb, 32'shc3edf141, 32'shc3ecdbdc, 32'shc3ebc69c, 32'shc3eab181, 32'shc3e99c8b, 
               32'shc3e887bb, 32'shc3e7730f, 32'shc3e65e88, 32'shc3e54a27, 32'shc3e435ea, 32'shc3e321d3, 32'shc3e20de1, 32'shc3e0fa14, 
               32'shc3dfe66c, 32'shc3ded2e9, 32'shc3ddbf8b, 32'shc3dcac52, 32'shc3db993e, 32'shc3da8650, 32'shc3d97386, 32'shc3d860e2, 
               32'shc3d74e62, 32'shc3d63c08, 32'shc3d529d3, 32'shc3d417c3, 32'shc3d305d8, 32'shc3d1f413, 32'shc3d0e272, 32'shc3cfd0f7, 
               32'shc3cebfa0, 32'shc3cdae6f, 32'shc3cc9d63, 32'shc3cb8c7c, 32'shc3ca7bba, 32'shc3c96b1e, 32'shc3c85aa6, 32'shc3c74a54, 
               32'shc3c63a26, 32'shc3c52a1e, 32'shc3c41a3b, 32'shc3c30a7e, 32'shc3c1fae5, 32'shc3c0eb71, 32'shc3bfdc23, 32'shc3beccfa, 
               32'shc3bdbdf6, 32'shc3bcaf17, 32'shc3bba05e, 32'shc3ba91c9, 32'shc3b9835a, 32'shc3b87510, 32'shc3b766eb, 32'shc3b658eb, 
               32'shc3b54b11, 32'shc3b43d5b, 32'shc3b32fcb, 32'shc3b22260, 32'shc3b1151b, 32'shc3b007fa, 32'shc3aefaff, 32'shc3adee28, 
               32'shc3ace178, 32'shc3abd4ec, 32'shc3aac885, 32'shc3a9bc44, 32'shc3a8b028, 32'shc3a7a431, 32'shc3a6985f, 32'shc3a58cb3, 
               32'shc3a4812c, 32'shc3a375ca, 32'shc3a26a8d, 32'shc3a15f76, 32'shc3a05484, 32'shc39f49b7, 32'shc39e3f0f, 32'shc39d348c, 
               32'shc39c2a2f, 32'shc39b1ff7, 32'shc39a15e4, 32'shc3990bf7, 32'shc398022f, 32'shc396f88c, 32'shc395ef0e, 32'shc394e5b6, 
               32'shc393dc82, 32'shc392d375, 32'shc391ca8c, 32'shc390c1c9, 32'shc38fb92a, 32'shc38eb0b2, 32'shc38da85e, 32'shc38ca030, 
               32'shc38b9827, 32'shc38a9043, 32'shc3898885, 32'shc38880ec, 32'shc3877978, 32'shc386722a, 32'shc3856b01, 32'shc38463fd, 
               32'shc3835d1e, 32'shc3825665, 32'shc3814fd1, 32'shc3804963, 32'shc37f4319, 32'shc37e3cf6, 32'shc37d36f7, 32'shc37c311e, 
               32'shc37b2b6a, 32'shc37a25db, 32'shc3792072, 32'shc3781b2e, 32'shc377160f, 32'shc3761116, 32'shc3750c42, 32'shc3740793, 
               32'shc373030a, 32'shc371fea6, 32'shc370fa68, 32'shc36ff64e, 32'shc36ef25b, 32'shc36dee8c, 32'shc36ceae3, 32'shc36be75f, 
               32'shc36ae401, 32'shc369e0c8, 32'shc368ddb4, 32'shc367dac6, 32'shc366d7fd, 32'shc365d55a, 32'shc364d2dc, 32'shc363d083, 
               32'shc362ce50, 32'shc361cc42, 32'shc360ca59, 32'shc35fc896, 32'shc35ec6f8, 32'shc35dc580, 32'shc35cc42d, 32'shc35bc2ff, 
               32'shc35ac1f7, 32'shc359c114, 32'shc358c057, 32'shc357bfbf, 32'shc356bf4d, 32'shc355bf00, 32'shc354bed8, 32'shc353bed6, 
               32'shc352bef9, 32'shc351bf41, 32'shc350bfaf, 32'shc34fc043, 32'shc34ec0fc, 32'shc34dc1da, 32'shc34cc2de, 32'shc34bc407, 
               32'shc34ac556, 32'shc349c6ca, 32'shc348c864, 32'shc347ca23, 32'shc346cc07, 32'shc345ce11, 32'shc344d041, 32'shc343d295, 
               32'shc342d510, 32'shc341d7b0, 32'shc340da75, 32'shc33fdd60, 32'shc33ee070, 32'shc33de3a5, 32'shc33ce701, 32'shc33bea81, 
               32'shc33aee27, 32'shc339f1f3, 32'shc338f5e4, 32'shc337f9fb, 32'shc336fe37, 32'shc3360298, 32'shc3350720, 32'shc3340bcc, 
               32'shc333109e, 32'shc3321596, 32'shc3311ab3, 32'shc3301ff5, 32'shc32f255e, 32'shc32e2aeb, 32'shc32d309e, 32'shc32c3677, 
               32'shc32b3c75, 32'shc32a4299, 32'shc32948e2, 32'shc3284f51, 32'shc32755e5, 32'shc3265c9f, 32'shc325637f, 32'shc3246a83, 
               32'shc32371ae, 32'shc32278fe, 32'shc3218073, 32'shc320880e, 32'shc31f8fcf, 32'shc31e97b5, 32'shc31d9fc1, 32'shc31ca7f2, 
               32'shc31bb049, 32'shc31ab8c6, 32'shc319c168, 32'shc318ca2f, 32'shc317d31c, 32'shc316dc2f, 32'shc315e567, 32'shc314eec5, 
               32'shc313f848, 32'shc31301f1, 32'shc3120bc0, 32'shc31115b4, 32'shc3101fce, 32'shc30f2a0d, 32'shc30e3472, 32'shc30d3efd, 
               32'shc30c49ad, 32'shc30b5482, 32'shc30a5f7e, 32'shc3096a9f, 32'shc30875e5, 32'shc3078151, 32'shc3068ce3, 32'shc305989a, 
               32'shc304a477, 32'shc303b07a, 32'shc302bca2, 32'shc301c8f0, 32'shc300d563, 32'shc2ffe1fc, 32'shc2feeebb, 32'shc2fdfb9f, 
               32'shc2fd08a9, 32'shc2fc15d9, 32'shc2fb232e, 32'shc2fa30a9, 32'shc2f93e4a, 32'shc2f84c10, 32'shc2f759fc, 32'shc2f6680d, 
               32'shc2f57644, 32'shc2f484a1, 32'shc2f39323, 32'shc2f2a1cb, 32'shc2f1b099, 32'shc2f0bf8c, 32'shc2efcea6, 32'shc2eedde4, 
               32'shc2eded49, 32'shc2ecfcd3, 32'shc2ec0c82, 32'shc2eb1c58, 32'shc2ea2c53, 32'shc2e93c74, 32'shc2e84cba, 32'shc2e75d26, 
               32'shc2e66db8, 32'shc2e57e70, 32'shc2e48f4d, 32'shc2e3a050, 32'shc2e2b178, 32'shc2e1c2c7, 32'shc2e0d43b, 32'shc2dfe5d4, 
               32'shc2def794, 32'shc2de0979, 32'shc2dd1b84, 32'shc2dc2db4, 32'shc2db400a, 32'shc2da5286, 32'shc2d96528, 32'shc2d877f0, 
               32'shc2d78add, 32'shc2d69df0, 32'shc2d5b128, 32'shc2d4c486, 32'shc2d3d80a, 32'shc2d2ebb4, 32'shc2d1ff84, 32'shc2d11379, 
               32'shc2d02794, 32'shc2cf3bd5, 32'shc2ce503b, 32'shc2cd64c7, 32'shc2cc7979, 32'shc2cb8e51, 32'shc2caa34f, 32'shc2c9b872, 
               32'shc2c8cdbb, 32'shc2c7e32a, 32'shc2c6f8be, 32'shc2c60e78, 32'shc2c52459, 32'shc2c43a5e, 32'shc2c3508a, 32'shc2c266db, 
               32'shc2c17d52, 32'shc2c093ef, 32'shc2bfaab2, 32'shc2bec19b, 32'shc2bdd8a9, 32'shc2bcefdd, 32'shc2bc0737, 32'shc2bb1eb6, 
               32'shc2ba365c, 32'shc2b94e27, 32'shc2b86618, 32'shc2b77e2f, 32'shc2b6966c, 32'shc2b5aece, 32'shc2b4c756, 32'shc2b3e004, 
               32'shc2b2f8d8, 32'shc2b211d2, 32'shc2b12af1, 32'shc2b04437, 32'shc2af5da2, 32'shc2ae7733, 32'shc2ad90ea, 32'shc2acaac6, 
               32'shc2abc4c9, 32'shc2aadef1, 32'shc2a9f93f, 32'shc2a913b3, 32'shc2a82e4d, 32'shc2a7490c, 32'shc2a663f2, 32'shc2a57efd, 
               32'shc2a49a2e, 32'shc2a3b585, 32'shc2a2d102, 32'shc2a1eca5, 32'shc2a1086d, 32'shc2a0245c, 32'shc29f4070, 32'shc29e5caa, 
               32'shc29d790a, 32'shc29c9590, 32'shc29bb23c, 32'shc29acf0d, 32'shc299ec05, 32'shc2990922, 32'shc2982665, 32'shc29743ce, 
               32'shc296615d, 32'shc2957f12, 32'shc2949ced, 32'shc293baed, 32'shc292d914, 32'shc291f760, 32'shc29115d3, 32'shc290346b, 
               32'shc28f5329, 32'shc28e720d, 32'shc28d9117, 32'shc28cb047, 32'shc28bcf9c, 32'shc28aef18, 32'shc28a0eb9, 32'shc2892e81, 
               32'shc2884e6e, 32'shc2876e82, 32'shc2868ebb, 32'shc285af1a, 32'shc284cf9f, 32'shc283f04a, 32'shc283111b, 32'shc2823211, 
               32'shc281532e, 32'shc2807471, 32'shc27f95d9, 32'shc27eb768, 32'shc27dd91c, 32'shc27cfaf7, 32'shc27c1cf7, 32'shc27b3f1e, 
               32'shc27a616a, 32'shc27983dc, 32'shc278a674, 32'shc277c932, 32'shc276ec16, 32'shc2760f20, 32'shc2753250, 32'shc27455a6, 
               32'shc2737922, 32'shc2729cc4, 32'shc271c08c, 32'shc270e47a, 32'shc270088e, 32'shc26f2cc7, 32'shc26e5127, 32'shc26d75ad, 
               32'shc26c9a58, 32'shc26bbf2a, 32'shc26ae422, 32'shc26a093f, 32'shc2692e83, 32'shc26853ed, 32'shc267797c, 32'shc2669f32, 
               32'shc265c50e, 32'shc264eb0f, 32'shc2641137, 32'shc2633785, 32'shc2625df8, 32'shc2618492, 32'shc260ab51, 32'shc25fd237, 
               32'shc25ef943, 32'shc25e2074, 32'shc25d47cc, 32'shc25c6f4a, 32'shc25b96ee, 32'shc25abeb7, 32'shc259e6a7, 32'shc2590ebd, 
               32'shc25836f9, 32'shc2575f5b, 32'shc25687e3, 32'shc255b091, 32'shc254d965, 32'shc254025f, 32'shc2532b7f, 32'shc25254c5, 
               32'shc2517e31, 32'shc250a7c3, 32'shc24fd17c, 32'shc24efb5a, 32'shc24e255e, 32'shc24d4f89, 32'shc24c79d9, 32'shc24ba450, 
               32'shc24aceed, 32'shc249f9af, 32'shc2492498, 32'shc2484fa7, 32'shc2477adc, 32'shc246a637, 32'shc245d1b8, 32'shc244fd5f, 
               32'shc244292c, 32'shc243551f, 32'shc2428139, 32'shc241ad78, 32'shc240d9de, 32'shc2400669, 32'shc23f331b, 32'shc23e5ff3, 
               32'shc23d8cf1, 32'shc23cba15, 32'shc23be75f, 32'shc23b14cf, 32'shc23a4265, 32'shc2397021, 32'shc2389e04, 32'shc237cc0d, 
               32'shc236fa3b, 32'shc2362890, 32'shc235570b, 32'shc23485ac, 32'shc233b473, 32'shc232e361, 32'shc2321274, 32'shc23141ae, 
               32'shc230710d, 32'shc22fa093, 32'shc22ed03f, 32'shc22e0011, 32'shc22d3009, 32'shc22c6028, 32'shc22b906c, 32'shc22ac0d7, 
               32'shc229f167, 32'shc229221e, 32'shc22852fb, 32'shc22783fe, 32'shc226b528, 32'shc225e677, 32'shc22517ed, 32'shc2244989, 
               32'shc2237b4b, 32'shc222ad33, 32'shc221df41, 32'shc2211176, 32'shc22043d0, 32'shc21f7651, 32'shc21ea8f8, 32'shc21ddbc5, 
               32'shc21d0eb8, 32'shc21c41d2, 32'shc21b7511, 32'shc21aa877, 32'shc219dc03, 32'shc2190fb5, 32'shc218438e, 32'shc217778c, 
               32'shc216abb1, 32'shc215dffc, 32'shc215146d, 32'shc2144904, 32'shc2137dc2, 32'shc212b2a5, 32'shc211e7af, 32'shc2111cdf, 
               32'shc2105236, 32'shc20f87b2, 32'shc20ebd55, 32'shc20df31e, 32'shc20d290d, 32'shc20c5f22, 32'shc20b955e, 32'shc20acbc0, 
               32'shc20a0248, 32'shc20938f6, 32'shc2086fca, 32'shc207a6c5, 32'shc206dde6, 32'shc206152d, 32'shc2054c9b, 32'shc204842e, 
               32'shc203bbe8, 32'shc202f3c8, 32'shc2022bce, 32'shc20163fb, 32'shc2009c4e, 32'shc1ffd4c7, 32'shc1ff0d66, 32'shc1fe462b, 
               32'shc1fd7f17, 32'shc1fcb829, 32'shc1fbf161, 32'shc1fb2ac0, 32'shc1fa6445, 32'shc1f99df0, 32'shc1f8d7c1, 32'shc1f811b9, 
               32'shc1f74bd6, 32'shc1f6861a, 32'shc1f5c085, 32'shc1f4fb15, 32'shc1f435cc, 32'shc1f370a9, 32'shc1f2abad, 32'shc1f1e6d7, 
               32'shc1f12227, 32'shc1f05d9d, 32'shc1ef9939, 32'shc1eed4fc, 32'shc1ee10e5, 32'shc1ed4cf5, 32'shc1ec892b, 32'shc1ebc587, 
               32'shc1eb0209, 32'shc1ea3eb1, 32'shc1e97b80, 32'shc1e8b876, 32'shc1e7f591, 32'shc1e732d3, 32'shc1e6703b, 32'shc1e5adc9, 
               32'shc1e4eb7e, 32'shc1e42959, 32'shc1e3675a, 32'shc1e2a582, 32'shc1e1e3d0, 32'shc1e12244, 32'shc1e060df, 32'shc1df9fa0, 
               32'shc1dede87, 32'shc1de1d94, 32'shc1dd5cc8, 32'shc1dc9c23, 32'shc1dbdba3, 32'shc1db1b4a, 32'shc1da5b17, 32'shc1d99b0b, 
               32'shc1d8db25, 32'shc1d81b65, 32'shc1d75bcb, 32'shc1d69c58, 32'shc1d5dd0c, 32'shc1d51de5, 32'shc1d45ee5, 32'shc1d3a00b, 
               32'shc1d2e158, 32'shc1d222cb, 32'shc1d16464, 32'shc1d0a624, 32'shc1cfe80a, 32'shc1cf2a17, 32'shc1ce6c49, 32'shc1cdaea3, 
               32'shc1ccf122, 32'shc1cc33c8, 32'shc1cb7694, 32'shc1cab987, 32'shc1c9fca0, 32'shc1c93fdf, 32'shc1c88345, 32'shc1c7c6d1, 
               32'shc1c70a84, 32'shc1c64e5d, 32'shc1c5925c, 32'shc1c4d682, 32'shc1c41ace, 32'shc1c35f40, 32'shc1c2a3d9, 32'shc1c1e898, 
               32'shc1c12d7e, 32'shc1c0728a, 32'shc1bfb7bc, 32'shc1befd15, 32'shc1be4294, 32'shc1bd883a, 32'shc1bcce06, 32'shc1bc13f8, 
               32'shc1bb5a11, 32'shc1baa050, 32'shc1b9e6b6, 32'shc1b92d42, 32'shc1b873f5, 32'shc1b7bacd, 32'shc1b701cd, 32'shc1b648f3, 
               32'shc1b5903f, 32'shc1b4d7b1, 32'shc1b41f4a, 32'shc1b3670a, 32'shc1b2aef0, 32'shc1b1f6fc, 32'shc1b13f2f, 32'shc1b08788, 
               32'shc1afd007, 32'shc1af18ae, 32'shc1ae617a, 32'shc1adaa6d, 32'shc1acf386, 32'shc1ac3cc6, 32'shc1ab862c, 32'shc1aacfb9, 
               32'shc1aa196c, 32'shc1a96346, 32'shc1a8ad46, 32'shc1a7f76c, 32'shc1a741b9, 32'shc1a68c2d, 32'shc1a5d6c7, 32'shc1a52187, 
               32'shc1a46c6e, 32'shc1a3b77b, 32'shc1a302af, 32'shc1a24e09, 32'shc1a1998a, 32'shc1a0e531, 32'shc1a030ff, 32'shc19f7cf3, 
               32'shc19ec90d, 32'shc19e154e, 32'shc19d61b6, 32'shc19cae44, 32'shc19bfaf9, 32'shc19b47d4, 32'shc19a94d5, 32'shc199e1fd, 
               32'shc1992f4c, 32'shc1987cc1, 32'shc197ca5c, 32'shc197181e, 32'shc1966606, 32'shc195b415, 32'shc195024b, 32'shc19450a7, 
               32'shc1939f29, 32'shc192edd2, 32'shc1923ca2, 32'shc1918b98, 32'shc190dab4, 32'shc19029f7, 32'shc18f7961, 32'shc18ec8f1, 
               32'shc18e18a7, 32'shc18d6884, 32'shc18cb888, 32'shc18c08b2, 32'shc18b5903, 32'shc18aa97a, 32'shc189fa17, 32'shc1894adc, 
               32'shc1889bc6, 32'shc187ecd8, 32'shc1873e10, 32'shc1868f6e, 32'shc185e0f3, 32'shc185329e, 32'shc1848470, 32'shc183d669, 
               32'shc1832888, 32'shc1827acd, 32'shc181cd3a, 32'shc1811fcc, 32'shc1807285, 32'shc17fc565, 32'shc17f186c, 32'shc17e6b99, 
               32'shc17dbeec, 32'shc17d1266, 32'shc17c6607, 32'shc17bb9ce, 32'shc17b0dbb, 32'shc17a61d0, 32'shc179b60b, 32'shc1790a6c, 
               32'shc1785ef4, 32'shc177b3a3, 32'shc1770878, 32'shc1765d73, 32'shc175b296, 32'shc17507df, 32'shc1745d4e, 32'shc173b2e4, 
               32'shc17308a1, 32'shc1725e84, 32'shc171b48e, 32'shc1710abe, 32'shc1706115, 32'shc16fb792, 32'shc16f0e36, 32'shc16e6501, 
               32'shc16dbbf3, 32'shc16d130a, 32'shc16c6a49, 32'shc16bc1ae, 32'shc16b193a, 32'shc16a70ec, 32'shc169c8c5, 32'shc16920c5, 
               32'shc16878eb, 32'shc167d137, 32'shc16729ab, 32'shc1668245, 32'shc165db05, 32'shc16533ed, 32'shc1648cfa, 32'shc163e62f, 
               32'shc1633f8a, 32'shc162990c, 32'shc161f2b4, 32'shc1614c83, 32'shc160a678, 32'shc1600095, 32'shc15f5ad7, 32'shc15eb541, 
               32'shc15e0fd1, 32'shc15d6a88, 32'shc15cc565, 32'shc15c2069, 32'shc15b7b94, 32'shc15ad6e5, 32'shc15a325d, 32'shc1598dfb, 
               32'shc158e9c1, 32'shc15845ac, 32'shc157a1bf, 32'shc156fdf8, 32'shc1565a58, 32'shc155b6de, 32'shc155138c, 32'shc154705f, 
               32'shc153cd5a, 32'shc1532a7b, 32'shc15287c3, 32'shc151e531, 32'shc15142c6, 32'shc150a082, 32'shc14ffe64, 32'shc14f5c6d, 
               32'shc14eba9d, 32'shc14e18f3, 32'shc14d7771, 32'shc14cd614, 32'shc14c34df, 32'shc14b93d0, 32'shc14af2e8, 32'shc14a5226, 
               32'shc149b18b, 32'shc1491117, 32'shc14870ca, 32'shc147d0a3, 32'shc14730a3, 32'shc14690ca, 32'shc145f117, 32'shc145518b, 
               32'shc144b225, 32'shc14412e7, 32'shc14373cf, 32'shc142d4de, 32'shc1423613, 32'shc141976f, 32'shc140f8f2, 32'shc1405a9c, 
               32'shc13fbc6c, 32'shc13f1e63, 32'shc13e8081, 32'shc13de2c5, 32'shc13d4530, 32'shc13ca7c2, 32'shc13c0a7b, 32'shc13b6d5a, 
               32'shc13ad060, 32'shc13a338d, 32'shc13996e0, 32'shc138fa5a, 32'shc1385dfb, 32'shc137c1c3, 32'shc13725b1, 32'shc13689c6, 
               32'shc135ee02, 32'shc1355265, 32'shc134b6ee, 32'shc1341b9e, 32'shc1338075, 32'shc132e572, 32'shc1324a96, 32'shc131afe1, 
               32'shc1311553, 32'shc1307aeb, 32'shc12fe0ab, 32'shc12f4690, 32'shc12eac9d, 32'shc12e12d1, 32'shc12d792b, 32'shc12cdfac, 
               32'shc12c4653, 32'shc12bad22, 32'shc12b1417, 32'shc12a7b33, 32'shc129e276, 32'shc12949df, 32'shc128b16f, 32'shc1281926, 
               32'shc1278104, 32'shc126e909, 32'shc1265134, 32'shc125b986, 32'shc12521ff, 32'shc1248a9e, 32'shc123f365, 32'shc1235c52, 
               32'shc122c566, 32'shc1222ea1, 32'shc1219802, 32'shc121018a, 32'shc1206b39, 32'shc11fd50f, 32'shc11f3f0c, 32'shc11ea92f, 
               32'shc11e1379, 32'shc11d7dea, 32'shc11ce882, 32'shc11c5341, 32'shc11bbe26, 32'shc11b2932, 32'shc11a9465, 32'shc119ffbf, 
               32'shc1196b3f, 32'shc118d6e7, 32'shc11842b5, 32'shc117aeaa, 32'shc1171ac6, 32'shc1168708, 32'shc115f372, 32'shc1156002, 
               32'shc114ccb9, 32'shc1143997, 32'shc113a69b, 32'shc11313c7, 32'shc1128119, 32'shc111ee92, 32'shc1115c32, 32'shc110c9f8, 
               32'shc11037e6, 32'shc10fa5fa, 32'shc10f1435, 32'shc10e8297, 32'shc10df120, 32'shc10d5fd0, 32'shc10ccea6, 32'shc10c3da4, 
               32'shc10bacc8, 32'shc10b1c13, 32'shc10a8b85, 32'shc109fb1d, 32'shc1096add, 32'shc108dac3, 32'shc1084ad0, 32'shc107bb04, 
               32'shc1072b5f, 32'shc1069be1, 32'shc1060c89, 32'shc1057d59, 32'shc104ee4f, 32'shc1045f6c, 32'shc103d0b0, 32'shc103421b, 
               32'shc102b3ac, 32'shc1022565, 32'shc1019744, 32'shc101094a, 32'shc1007b77, 32'shc0ffedcb, 32'shc0ff6046, 32'shc0fed2e8, 
               32'shc0fe45b0, 32'shc0fdb8a0, 32'shc0fd2bb6, 32'shc0fc9ef3, 32'shc0fc1257, 32'shc0fb85e2, 32'shc0faf993, 32'shc0fa6d6c, 
               32'shc0f9e16b, 32'shc0f95592, 32'shc0f8c9df, 32'shc0f83e53, 32'shc0f7b2ee, 32'shc0f727b0, 32'shc0f69c99, 32'shc0f611a8, 
               32'shc0f586df, 32'shc0f4fc3c, 32'shc0f471c1, 32'shc0f3e76c, 32'shc0f35d3e, 32'shc0f2d337, 32'shc0f24957, 32'shc0f1bf9d, 
               32'shc0f1360b, 32'shc0f0aca0, 32'shc0f0235b, 32'shc0ef9a3d, 32'shc0ef1147, 32'shc0ee8877, 32'shc0edffce, 32'shc0ed774c, 
               32'shc0eceef1, 32'shc0ec66bc, 32'shc0ebdeaf, 32'shc0eb56c9, 32'shc0eacf09, 32'shc0ea4771, 32'shc0e9bfff, 32'shc0e938b4, 
               32'shc0e8b190, 32'shc0e82a93, 32'shc0e7a3bd, 32'shc0e71d0e, 32'shc0e69686, 32'shc0e61025, 32'shc0e589eb, 32'shc0e503d7, 
               32'shc0e47deb, 32'shc0e3f825, 32'shc0e37287, 32'shc0e2ed0f, 32'shc0e267be, 32'shc0e1e294, 32'shc0e15d92, 32'shc0e0d8b6, 
               32'shc0e05401, 32'shc0dfcf73, 32'shc0df4b0b, 32'shc0dec6cb, 32'shc0de42b2, 32'shc0ddbec0, 32'shc0dd3af4, 32'shc0dcb750, 
               32'shc0dc33d2, 32'shc0dbb07c, 32'shc0db2d4c, 32'shc0daaa44, 32'shc0da2762, 32'shc0d9a4a7, 32'shc0d92214, 32'shc0d89fa7, 
               32'shc0d81d61, 32'shc0d79b42, 32'shc0d7194a, 32'shc0d69779, 32'shc0d615cf, 32'shc0d5944c, 32'shc0d512f0, 32'shc0d491bb, 
               32'shc0d410ad, 32'shc0d38fc6, 32'shc0d30f05, 32'shc0d28e6c, 32'shc0d20dfa, 32'shc0d18dae, 32'shc0d10d8a, 32'shc0d08d8d, 
               32'shc0d00db6, 32'shc0cf8e07, 32'shc0cf0e7f, 32'shc0ce8f1d, 32'shc0ce0fe3, 32'shc0cd90cf, 32'shc0cd11e3, 32'shc0cc931d, 
               32'shc0cc147f, 32'shc0cb9607, 32'shc0cb17b7, 32'shc0ca998d, 32'shc0ca1b8a, 32'shc0c99daf, 32'shc0c91ffa, 32'shc0c8a26d, 
               32'shc0c82506, 32'shc0c7a7c6, 32'shc0c72aae, 32'shc0c6adbc, 32'shc0c630f2, 32'shc0c5b44e, 32'shc0c537d1, 32'shc0c4bb7c, 
               32'shc0c43f4d, 32'shc0c3c346, 32'shc0c34765, 32'shc0c2cbab, 32'shc0c25019, 32'shc0c1d4ad, 32'shc0c15969, 32'shc0c0de4b, 
               32'shc0c06355, 32'shc0bfe885, 32'shc0bf6ddd, 32'shc0bef35b, 32'shc0be7901, 32'shc0bdfecd, 32'shc0bd84c1, 32'shc0bd0adb, 
               32'shc0bc911d, 32'shc0bc1786, 32'shc0bb9e15, 32'shc0bb24cc, 32'shc0baabaa, 32'shc0ba32af, 32'shc0b9b9da, 32'shc0b9412d, 
               32'shc0b8c8a7, 32'shc0b85048, 32'shc0b7d810, 32'shc0b75fff, 32'shc0b6e815, 32'shc0b67052, 32'shc0b5f8b6, 32'shc0b58141, 
               32'shc0b509f3, 32'shc0b492cc, 32'shc0b41bcd, 32'shc0b3a4f4, 32'shc0b32e42, 32'shc0b2b7b8, 32'shc0b24154, 32'shc0b1cb17, 
               32'shc0b15502, 32'shc0b0df13, 32'shc0b0694c, 32'shc0aff3ac, 32'shc0af7e33, 32'shc0af08e0, 32'shc0ae93b5, 32'shc0ae1eb1, 
               32'shc0ada9d4, 32'shc0ad351e, 32'shc0acc08f, 32'shc0ac4c27, 32'shc0abd7e6, 32'shc0ab63cd, 32'shc0aaefda, 32'shc0aa7c0e, 
               32'shc0aa086a, 32'shc0a994ec, 32'shc0a92196, 32'shc0a8ae67, 32'shc0a83b5e, 32'shc0a7c87d, 32'shc0a755c3, 32'shc0a6e330, 
               32'shc0a670c4, 32'shc0a5fe7f, 32'shc0a58c62, 32'shc0a51a6b, 32'shc0a4a89b, 32'shc0a436f3, 32'shc0a3c571, 32'shc0a35417, 
               32'shc0a2e2e3, 32'shc0a271d7, 32'shc0a200f2, 32'shc0a19034, 32'shc0a11f9d, 32'shc0a0af2d, 32'shc0a03ee4, 32'shc09fcec3, 
               32'shc09f5ec8, 32'shc09eeef5, 32'shc09e7f48, 32'shc09e0fc3, 32'shc09da065, 32'shc09d312e, 32'shc09cc21e, 32'shc09c5335, 
               32'shc09be473, 32'shc09b75d8, 32'shc09b0765, 32'shc09a9918, 32'shc09a2af3, 32'shc099bcf5, 32'shc0994f1d, 32'shc098e16d, 
               32'shc09873e4, 32'shc0980683, 32'shc0979948, 32'shc0972c34, 32'shc096bf48, 32'shc0965282, 32'shc095e5e4, 32'shc095796d, 
               32'shc0950d1d, 32'shc094a0f4, 32'shc09434f2, 32'shc093c917, 32'shc0935d64, 32'shc092f1d7, 32'shc0928672, 32'shc0921b34, 
               32'shc091b01d, 32'shc091452d, 32'shc090da64, 32'shc0906fc3, 32'shc0900548, 32'shc08f9af5, 32'shc08f30c8, 32'shc08ec6c3, 
               32'shc08e5ce5, 32'shc08df32e, 32'shc08d899f, 32'shc08d2036, 32'shc08cb6f5, 32'shc08c4dda, 32'shc08be4e7, 32'shc08b7c1b, 
               32'shc08b1376, 32'shc08aaaf8, 32'shc08a42a2, 32'shc089da72, 32'shc089726a, 32'shc0890a89, 32'shc088a2cf, 32'shc0883b3c, 
               32'shc087d3d0, 32'shc0876c8c, 32'shc087056e, 32'shc0869e78, 32'shc08637a9, 32'shc085d101, 32'shc0856a80, 32'shc0850426, 
               32'shc0849df4, 32'shc08437e9, 32'shc083d204, 32'shc0836c47, 32'shc08306b2, 32'shc082a143, 32'shc0823bfb, 32'shc081d6db, 
               32'shc08171e2, 32'shc0810d10, 32'shc080a865, 32'shc08043e1, 32'shc07fdf85, 32'shc07f7b50, 32'shc07f1741, 32'shc07eb35a, 
               32'shc07e4f9b, 32'shc07dec02, 32'shc07d8890, 32'shc07d2546, 32'shc07cc223, 32'shc07c5f27, 32'shc07bfc52, 32'shc07b99a5, 
               32'shc07b371e, 32'shc07ad4bf, 32'shc07a7287, 32'shc07a1076, 32'shc079ae8c, 32'shc0794cca, 32'shc078eb2f, 32'shc07889bb, 
               32'shc078286e, 32'shc077c748, 32'shc0776649, 32'shc0770572, 32'shc076a4c2, 32'shc0764439, 32'shc075e3d7, 32'shc075839c, 
               32'shc0752389, 32'shc074c39d, 32'shc07463d8, 32'shc074043a, 32'shc073a4c3, 32'shc0734574, 32'shc072e64c, 32'shc072874b, 
               32'shc0722871, 32'shc071c9be, 32'shc0716b33, 32'shc0710ccf, 32'shc070ae92, 32'shc070507c, 32'shc06ff28e, 32'shc06f94c6, 
               32'shc06f3726, 32'shc06ed9ad, 32'shc06e7c5b, 32'shc06e1f31, 32'shc06dc22e, 32'shc06d6551, 32'shc06d089d, 32'shc06cac0f, 
               32'shc06c4fa8, 32'shc06bf369, 32'shc06b9751, 32'shc06b3b60, 32'shc06adf97, 32'shc06a83f5, 32'shc06a2879, 32'shc069cd26, 
               32'shc06971f9, 32'shc06916f3, 32'shc068bc15, 32'shc068615e, 32'shc06806ce, 32'shc067ac66, 32'shc0675225, 32'shc066f80a, 
               32'shc0669e18, 32'shc066444c, 32'shc065eaa8, 32'shc065912a, 32'shc06537d4, 32'shc064dea6, 32'shc064859e, 32'shc0642cbe, 
               32'shc063d405, 32'shc0637b73, 32'shc0632309, 32'shc062cac6, 32'shc06272aa, 32'shc0621ab5, 32'shc061c2e7, 32'shc0616b41, 
               32'shc06113c2, 32'shc060bc6a, 32'shc060653a, 32'shc0600e30, 32'shc05fb74e, 32'shc05f6093, 32'shc05f0a00, 32'shc05eb393, 
               32'shc05e5d4e, 32'shc05e0730, 32'shc05db13a, 32'shc05d5b6b, 32'shc05d05c3, 32'shc05cb042, 32'shc05c5ae8, 32'shc05c05b6, 
               32'shc05bb0ab, 32'shc05b5bc7, 32'shc05b070a, 32'shc05ab275, 32'shc05a5e07, 32'shc05a09c0, 32'shc059b5a1, 32'shc05961a9, 
               32'shc0590dd8, 32'shc058ba2e, 32'shc05866ac, 32'shc0581350, 32'shc057c01d, 32'shc0576d10, 32'shc0571a2b, 32'shc056c76c, 
               32'shc05674d6, 32'shc0562266, 32'shc055d01e, 32'shc0557dfd, 32'shc0552c03, 32'shc054da30, 32'shc0548885, 32'shc0543701, 
               32'shc053e5a5, 32'shc053946f, 32'shc0534361, 32'shc052f27a, 32'shc052a1bb, 32'shc0525123, 32'shc05200b2, 32'shc051b068, 
               32'shc0516045, 32'shc051104a, 32'shc050c077, 32'shc05070ca, 32'shc0502145, 32'shc04fd1e7, 32'shc04f82b0, 32'shc04f33a1, 
               32'shc04ee4b8, 32'shc04e95f8, 32'shc04e475e, 32'shc04df8ec, 32'shc04daaa1, 32'shc04d5c7d, 32'shc04d0e81, 32'shc04cc0ac, 
               32'shc04c72fe, 32'shc04c2577, 32'shc04bd818, 32'shc04b8ae0, 32'shc04b3dcf, 32'shc04af0e6, 32'shc04aa424, 32'shc04a5789, 
               32'shc04a0b16, 32'shc049beca, 32'shc04972a5, 32'shc04926a7, 32'shc048dad1, 32'shc0488f22, 32'shc048439b, 32'shc047f83a, 
               32'shc047ad01, 32'shc04761ef, 32'shc0471705, 32'shc046cc42, 32'shc04681a6, 32'shc0463732, 32'shc045ece5, 32'shc045a2bf, 
               32'shc04558c0, 32'shc0450ee9, 32'shc044c539, 32'shc0447bb0, 32'shc044324f, 32'shc043e915, 32'shc043a002, 32'shc0435717, 
               32'shc0430e53, 32'shc042c5b6, 32'shc0427d41, 32'shc04234f3, 32'shc041eccc, 32'shc041a4cd, 32'shc0415cf4, 32'shc0411544, 
               32'shc040cdba, 32'shc0408658, 32'shc0403f1d, 32'shc03ff80a, 32'shc03fb11d, 32'shc03f6a58, 32'shc03f23bb, 32'shc03edd45, 
               32'shc03e96f6, 32'shc03e50ce, 32'shc03e0ace, 32'shc03dc4f5, 32'shc03d7f44, 32'shc03d39b9, 32'shc03cf456, 32'shc03caf1b, 
               32'shc03c6a07, 32'shc03c251a, 32'shc03be054, 32'shc03b9bb6, 32'shc03b573f, 32'shc03b12ef, 32'shc03acec7, 32'shc03a8ac6, 
               32'shc03a46ed, 32'shc03a033a, 32'shc039bfaf, 32'shc0397c4c, 32'shc0393910, 32'shc038f5fb, 32'shc038b30d, 32'shc0387047, 
               32'shc0382da8, 32'shc037eb31, 32'shc037a8e1, 32'shc03766b8, 32'shc03724b6, 32'shc036e2dc, 32'shc036a129, 32'shc0365f9e, 
               32'shc0361e3a, 32'shc035dcfd, 32'shc0359be8, 32'shc0355afa, 32'shc0351a33, 32'shc034d994, 32'shc034991c, 32'shc03458cb, 
               32'shc03418a2, 32'shc033d8a0, 32'shc03398c5, 32'shc0335912, 32'shc0331986, 32'shc032da22, 32'shc0329ae4, 32'shc0325bcf, 
               32'shc0321ce0, 32'shc031de19, 32'shc0319f79, 32'shc0316101, 32'shc03122b0, 32'shc030e486, 32'shc030a684, 32'shc03068a9, 
               32'shc0302af5, 32'shc02fed69, 32'shc02fb004, 32'shc02f72c7, 32'shc02f35b1, 32'shc02ef8c2, 32'shc02ebbfb, 32'shc02e7f5b, 
               32'shc02e42e2, 32'shc02e0691, 32'shc02dca67, 32'shc02d8e64, 32'shc02d5289, 32'shc02d16d5, 32'shc02cdb49, 32'shc02c9fe4, 
               32'shc02c64a6, 32'shc02c2990, 32'shc02beea1, 32'shc02bb3d9, 32'shc02b7939, 32'shc02b3ec0, 32'shc02b046f, 32'shc02aca44, 
               32'shc02a9042, 32'shc02a5666, 32'shc02a1cb2, 32'shc029e326, 32'shc029a9c1, 32'shc0297083, 32'shc029376c, 32'shc028fe7d, 
               32'shc028c5b6, 32'shc0288d15, 32'shc028549c, 32'shc0281c4b, 32'shc027e421, 32'shc027ac1e, 32'shc0277442, 32'shc0273c8e, 
               32'shc0270502, 32'shc026cd9d, 32'shc026965f, 32'shc0265f48, 32'shc0262859, 32'shc025f191, 32'shc025baf1, 32'shc0258478, 
               32'shc0254e27, 32'shc02517fc, 32'shc024e1fa, 32'shc024ac1e, 32'shc024766a, 32'shc02440de, 32'shc0240b78, 32'shc023d63b, 
               32'shc023a124, 32'shc0236c35, 32'shc023376e, 32'shc02302cd, 32'shc022ce54, 32'shc0229a03, 32'shc02265d9, 32'shc02231d6, 
               32'shc021fdfb, 32'shc021ca47, 32'shc02196bb, 32'shc0216356, 32'shc0213018, 32'shc020fd02, 32'shc020ca13, 32'shc020974b, 
               32'shc02064ab, 32'shc0203232, 32'shc01fffe1, 32'shc01fcdb7, 32'shc01f9bb5, 32'shc01f69da, 32'shc01f3826, 32'shc01f069a, 
               32'shc01ed535, 32'shc01ea3f7, 32'shc01e72e1, 32'shc01e41f3, 32'shc01e112b, 32'shc01de08c, 32'shc01db013, 32'shc01d7fc2, 
               32'shc01d4f99, 32'shc01d1f96, 32'shc01cefbb, 32'shc01cc008, 32'shc01c907c, 32'shc01c6118, 32'shc01c31da, 32'shc01c02c5, 
               32'shc01bd3d6, 32'shc01ba50f, 32'shc01b7670, 32'shc01b47f8, 32'shc01b19a7, 32'shc01aeb7e, 32'shc01abd7c, 32'shc01a8fa1, 
               32'shc01a61ee, 32'shc01a3463, 32'shc01a06fe, 32'shc019d9c2, 32'shc019acac, 32'shc0197fbe, 32'shc01952f8, 32'shc0192659, 
               32'shc018f9e1, 32'shc018cd91, 32'shc018a168, 32'shc0187566, 32'shc018498c, 32'shc0181dda, 32'shc017f24e, 32'shc017c6eb, 
               32'shc0179bae, 32'shc0177099, 32'shc01745ac, 32'shc0171ae6, 32'shc016f047, 32'shc016c5d0, 32'shc0169b80, 32'shc0167158, 
               32'shc0164757, 32'shc0161d7d, 32'shc015f3cb, 32'shc015ca40, 32'shc015a0dd, 32'shc01577a1, 32'shc0154e8d, 32'shc01525a0, 
               32'shc014fcda, 32'shc014d43c, 32'shc014abc5, 32'shc0148376, 32'shc0145b4e, 32'shc014334e, 32'shc0140b75, 32'shc013e3c3, 
               32'shc013bc39, 32'shc01394d6, 32'shc0136d9b, 32'shc0134687, 32'shc0131f9b, 32'shc012f8d6, 32'shc012d238, 32'shc012abc2, 
               32'shc0128574, 32'shc0125f4c, 32'shc012394c, 32'shc0121374, 32'shc011edc3, 32'shc011c83a, 32'shc011a2d8, 32'shc0117d9d, 
               32'shc011588a, 32'shc011339e, 32'shc0110eda, 32'shc010ea3d, 32'shc010c5c7, 32'shc010a179, 32'shc0107d53, 32'shc0105954, 
               32'shc010357c, 32'shc01011cc, 32'shc00fee43, 32'shc00fcae2, 32'shc00fa7a8, 32'shc00f8495, 32'shc00f61aa, 32'shc00f3ee6, 
               32'shc00f1c4a, 32'shc00ef9d6, 32'shc00ed788, 32'shc00eb562, 32'shc00e9364, 32'shc00e718d, 32'shc00e4fde, 32'shc00e2e56, 
               32'shc00e0cf5, 32'shc00debbc, 32'shc00dcaaa, 32'shc00da9c0, 32'shc00d88fd, 32'shc00d6861, 32'shc00d47ed, 32'shc00d27a1, 
               32'shc00d077c, 32'shc00ce77e, 32'shc00cc7a8, 32'shc00ca7f9, 32'shc00c8872, 32'shc00c6912, 32'shc00c49da, 32'shc00c2ac9, 
               32'shc00c0be0, 32'shc00bed1e, 32'shc00bce83, 32'shc00bb010, 32'shc00b91c4, 32'shc00b73a0, 32'shc00b55a3, 32'shc00b37ce, 
               32'shc00b1a20, 32'shc00afc9a, 32'shc00adf3b, 32'shc00ac203, 32'shc00aa4f3, 32'shc00a880a, 32'shc00a6b49, 32'shc00a4eb0, 
               32'shc00a323d, 32'shc00a15f3, 32'shc009f9cf, 32'shc009ddd3, 32'shc009c1ff, 32'shc009a652, 32'shc0098acc, 32'shc0096f6e, 
               32'shc0095438, 32'shc0093929, 32'shc0091e41, 32'shc0090381, 32'shc008e8e8, 32'shc008ce76, 32'shc008b42d, 32'shc0089a0a, 
               32'shc008800f, 32'shc008663c, 32'shc0084c90, 32'shc008330b, 32'shc00819ae, 32'shc0080078, 32'shc007e76a, 32'shc007ce83, 
               32'shc007b5c4, 32'shc0079d2c, 32'shc00784bc, 32'shc0076c73, 32'shc0075452, 32'shc0073c58, 32'shc0072485, 32'shc0070cda, 
               32'shc006f556, 32'shc006ddfa, 32'shc006c6c6, 32'shc006afb8, 32'shc00698d3, 32'shc0068214, 32'shc0066b7d, 32'shc006550e, 
               32'shc0063ec6, 32'shc00628a6, 32'shc00612ad, 32'shc005fcdb, 32'shc005e731, 32'shc005d1af, 32'shc005bc54, 32'shc005a720, 
               32'shc0059214, 32'shc0057d2f, 32'shc0056872, 32'shc00553dc, 32'shc0053f6e, 32'shc0052b27, 32'shc0051707, 32'shc005030f, 
               32'shc004ef3f, 32'shc004db96, 32'shc004c814, 32'shc004b4ba, 32'shc004a188, 32'shc0048e7d, 32'shc0047b99, 32'shc00468dd, 
               32'shc0045648, 32'shc00443db, 32'shc0043195, 32'shc0041f77, 32'shc0040d80, 32'shc003fbb0, 32'shc003ea09, 32'shc003d888, 
               32'shc003c72f, 32'shc003b5fe, 32'shc003a4f4, 32'shc0039411, 32'shc0038356, 32'shc00372c2, 32'shc0036256, 32'shc0035211, 
               32'shc00341f4, 32'shc00331fe, 32'shc0032230, 32'shc0031289, 32'shc003030a, 32'shc002f3b2, 32'shc002e482, 32'shc002d579, 
               32'shc002c697, 32'shc002b7dd, 32'shc002a94b, 32'shc0029ae0, 32'shc0028c9c, 32'shc0027e80, 32'shc002708c, 32'shc00262be, 
               32'shc0025519, 32'shc002479b, 32'shc0023a44, 32'shc0022d15, 32'shc002200d, 32'shc002132d, 32'shc0020674, 32'shc001f9e2, 
               32'shc001ed78, 32'shc001e136, 32'shc001d51b, 32'shc001c928, 32'shc001bd5c, 32'shc001b1b7, 32'shc001a63a, 32'shc0019ae5, 
               32'shc0018fb6, 32'shc00184b0, 32'shc00179d1, 32'shc0016f19, 32'shc0016489, 32'shc0015a20, 32'shc0014fdf, 32'shc00145c5, 
               32'shc0013bd3, 32'shc0013208, 32'shc0012865, 32'shc0011ee9, 32'shc0011594, 32'shc0010c67, 32'shc0010362, 32'shc000fa84, 
               32'shc000f1ce, 32'shc000e93f, 32'shc000e0d7, 32'shc000d897, 32'shc000d07e, 32'shc000c88d, 32'shc000c0c4, 32'shc000b921, 
               32'shc000b1a7, 32'shc000aa54, 32'shc000a328, 32'shc0009c24, 32'shc0009547, 32'shc0008e92, 32'shc0008804, 32'shc000819d, 
               32'shc0007b5f, 32'shc0007547, 32'shc0006f57, 32'shc000698f, 32'shc00063ee, 32'shc0005e74, 32'shc0005922, 32'shc00053f8, 
               32'shc0004ef5, 32'shc0004a19, 32'shc0004565, 32'shc00040d9, 32'shc0003c74, 32'shc0003836, 32'shc0003420, 32'shc0003031, 
               32'shc0002c6a, 32'shc00028ca, 32'shc0002552, 32'shc0002201, 32'shc0001ed8, 32'shc0001bd6, 32'shc00018fb, 32'shc0001649, 
               32'shc00013bd, 32'shc0001159, 32'shc0000f1d, 32'shc0000d08, 32'shc0000b1a, 32'shc0000954, 32'shc00007b6, 32'shc000063f, 
               32'shc00004ef, 32'shc00003c7, 32'shc00002c7, 32'shc00001ed, 32'shc000013c, 32'shc00000b2, 32'shc000004f, 32'shc0000014, 
               32'shc0000000, 32'shc0000014, 32'shc000004f, 32'shc00000b2, 32'shc000013c, 32'shc00001ed, 32'shc00002c7, 32'shc00003c7, 
               32'shc00004ef, 32'shc000063f, 32'shc00007b6, 32'shc0000954, 32'shc0000b1a, 32'shc0000d08, 32'shc0000f1d, 32'shc0001159, 
               32'shc00013bd, 32'shc0001649, 32'shc00018fb, 32'shc0001bd6, 32'shc0001ed8, 32'shc0002201, 32'shc0002552, 32'shc00028ca, 
               32'shc0002c6a, 32'shc0003031, 32'shc0003420, 32'shc0003836, 32'shc0003c74, 32'shc00040d9, 32'shc0004565, 32'shc0004a19, 
               32'shc0004ef5, 32'shc00053f8, 32'shc0005922, 32'shc0005e74, 32'shc00063ee, 32'shc000698f, 32'shc0006f57, 32'shc0007547, 
               32'shc0007b5f, 32'shc000819d, 32'shc0008804, 32'shc0008e92, 32'shc0009547, 32'shc0009c24, 32'shc000a328, 32'shc000aa54, 
               32'shc000b1a7, 32'shc000b921, 32'shc000c0c4, 32'shc000c88d, 32'shc000d07e, 32'shc000d897, 32'shc000e0d7, 32'shc000e93f, 
               32'shc000f1ce, 32'shc000fa84, 32'shc0010362, 32'shc0010c67, 32'shc0011594, 32'shc0011ee9, 32'shc0012865, 32'shc0013208, 
               32'shc0013bd3, 32'shc00145c5, 32'shc0014fdf, 32'shc0015a20, 32'shc0016489, 32'shc0016f19, 32'shc00179d1, 32'shc00184b0, 
               32'shc0018fb6, 32'shc0019ae5, 32'shc001a63a, 32'shc001b1b7, 32'shc001bd5c, 32'shc001c928, 32'shc001d51b, 32'shc001e136, 
               32'shc001ed78, 32'shc001f9e2, 32'shc0020674, 32'shc002132d, 32'shc002200d, 32'shc0022d15, 32'shc0023a44, 32'shc002479b, 
               32'shc0025519, 32'shc00262be, 32'shc002708c, 32'shc0027e80, 32'shc0028c9c, 32'shc0029ae0, 32'shc002a94b, 32'shc002b7dd, 
               32'shc002c697, 32'shc002d579, 32'shc002e482, 32'shc002f3b2, 32'shc003030a, 32'shc0031289, 32'shc0032230, 32'shc00331fe, 
               32'shc00341f4, 32'shc0035211, 32'shc0036256, 32'shc00372c2, 32'shc0038356, 32'shc0039411, 32'shc003a4f4, 32'shc003b5fe, 
               32'shc003c72f, 32'shc003d888, 32'shc003ea09, 32'shc003fbb0, 32'shc0040d80, 32'shc0041f77, 32'shc0043195, 32'shc00443db, 
               32'shc0045648, 32'shc00468dd, 32'shc0047b99, 32'shc0048e7d, 32'shc004a188, 32'shc004b4ba, 32'shc004c814, 32'shc004db96, 
               32'shc004ef3f, 32'shc005030f, 32'shc0051707, 32'shc0052b27, 32'shc0053f6e, 32'shc00553dc, 32'shc0056872, 32'shc0057d2f, 
               32'shc0059214, 32'shc005a720, 32'shc005bc54, 32'shc005d1af, 32'shc005e731, 32'shc005fcdb, 32'shc00612ad, 32'shc00628a6, 
               32'shc0063ec6, 32'shc006550e, 32'shc0066b7d, 32'shc0068214, 32'shc00698d3, 32'shc006afb8, 32'shc006c6c6, 32'shc006ddfa, 
               32'shc006f556, 32'shc0070cda, 32'shc0072485, 32'shc0073c58, 32'shc0075452, 32'shc0076c73, 32'shc00784bc, 32'shc0079d2c, 
               32'shc007b5c4, 32'shc007ce83, 32'shc007e76a, 32'shc0080078, 32'shc00819ae, 32'shc008330b, 32'shc0084c90, 32'shc008663c, 
               32'shc008800f, 32'shc0089a0a, 32'shc008b42d, 32'shc008ce76, 32'shc008e8e8, 32'shc0090381, 32'shc0091e41, 32'shc0093929, 
               32'shc0095438, 32'shc0096f6e, 32'shc0098acc, 32'shc009a652, 32'shc009c1ff, 32'shc009ddd3, 32'shc009f9cf, 32'shc00a15f3, 
               32'shc00a323d, 32'shc00a4eb0, 32'shc00a6b49, 32'shc00a880a, 32'shc00aa4f3, 32'shc00ac203, 32'shc00adf3b, 32'shc00afc9a, 
               32'shc00b1a20, 32'shc00b37ce, 32'shc00b55a3, 32'shc00b73a0, 32'shc00b91c4, 32'shc00bb010, 32'shc00bce83, 32'shc00bed1e, 
               32'shc00c0be0, 32'shc00c2ac9, 32'shc00c49da, 32'shc00c6912, 32'shc00c8872, 32'shc00ca7f9, 32'shc00cc7a8, 32'shc00ce77e, 
               32'shc00d077c, 32'shc00d27a1, 32'shc00d47ed, 32'shc00d6861, 32'shc00d88fd, 32'shc00da9c0, 32'shc00dcaaa, 32'shc00debbc, 
               32'shc00e0cf5, 32'shc00e2e56, 32'shc00e4fde, 32'shc00e718d, 32'shc00e9364, 32'shc00eb562, 32'shc00ed788, 32'shc00ef9d6, 
               32'shc00f1c4a, 32'shc00f3ee6, 32'shc00f61aa, 32'shc00f8495, 32'shc00fa7a8, 32'shc00fcae2, 32'shc00fee43, 32'shc01011cc, 
               32'shc010357c, 32'shc0105954, 32'shc0107d53, 32'shc010a179, 32'shc010c5c7, 32'shc010ea3d, 32'shc0110eda, 32'shc011339e, 
               32'shc011588a, 32'shc0117d9d, 32'shc011a2d8, 32'shc011c83a, 32'shc011edc3, 32'shc0121374, 32'shc012394c, 32'shc0125f4c, 
               32'shc0128574, 32'shc012abc2, 32'shc012d238, 32'shc012f8d6, 32'shc0131f9b, 32'shc0134687, 32'shc0136d9b, 32'shc01394d6, 
               32'shc013bc39, 32'shc013e3c3, 32'shc0140b75, 32'shc014334e, 32'shc0145b4e, 32'shc0148376, 32'shc014abc5, 32'shc014d43c, 
               32'shc014fcda, 32'shc01525a0, 32'shc0154e8d, 32'shc01577a1, 32'shc015a0dd, 32'shc015ca40, 32'shc015f3cb, 32'shc0161d7d, 
               32'shc0164757, 32'shc0167158, 32'shc0169b80, 32'shc016c5d0, 32'shc016f047, 32'shc0171ae6, 32'shc01745ac, 32'shc0177099, 
               32'shc0179bae, 32'shc017c6eb, 32'shc017f24e, 32'shc0181dda, 32'shc018498c, 32'shc0187566, 32'shc018a168, 32'shc018cd91, 
               32'shc018f9e1, 32'shc0192659, 32'shc01952f8, 32'shc0197fbe, 32'shc019acac, 32'shc019d9c2, 32'shc01a06fe, 32'shc01a3463, 
               32'shc01a61ee, 32'shc01a8fa1, 32'shc01abd7c, 32'shc01aeb7e, 32'shc01b19a7, 32'shc01b47f8, 32'shc01b7670, 32'shc01ba50f, 
               32'shc01bd3d6, 32'shc01c02c5, 32'shc01c31da, 32'shc01c6118, 32'shc01c907c, 32'shc01cc008, 32'shc01cefbb, 32'shc01d1f96, 
               32'shc01d4f99, 32'shc01d7fc2, 32'shc01db013, 32'shc01de08c, 32'shc01e112b, 32'shc01e41f3, 32'shc01e72e1, 32'shc01ea3f7, 
               32'shc01ed535, 32'shc01f069a, 32'shc01f3826, 32'shc01f69da, 32'shc01f9bb5, 32'shc01fcdb7, 32'shc01fffe1, 32'shc0203232, 
               32'shc02064ab, 32'shc020974b, 32'shc020ca13, 32'shc020fd02, 32'shc0213018, 32'shc0216356, 32'shc02196bb, 32'shc021ca47, 
               32'shc021fdfb, 32'shc02231d6, 32'shc02265d9, 32'shc0229a03, 32'shc022ce54, 32'shc02302cd, 32'shc023376e, 32'shc0236c35, 
               32'shc023a124, 32'shc023d63b, 32'shc0240b78, 32'shc02440de, 32'shc024766a, 32'shc024ac1e, 32'shc024e1fa, 32'shc02517fc, 
               32'shc0254e27, 32'shc0258478, 32'shc025baf1, 32'shc025f191, 32'shc0262859, 32'shc0265f48, 32'shc026965f, 32'shc026cd9d, 
               32'shc0270502, 32'shc0273c8e, 32'shc0277442, 32'shc027ac1e, 32'shc027e421, 32'shc0281c4b, 32'shc028549c, 32'shc0288d15, 
               32'shc028c5b6, 32'shc028fe7d, 32'shc029376c, 32'shc0297083, 32'shc029a9c1, 32'shc029e326, 32'shc02a1cb2, 32'shc02a5666, 
               32'shc02a9042, 32'shc02aca44, 32'shc02b046f, 32'shc02b3ec0, 32'shc02b7939, 32'shc02bb3d9, 32'shc02beea1, 32'shc02c2990, 
               32'shc02c64a6, 32'shc02c9fe4, 32'shc02cdb49, 32'shc02d16d5, 32'shc02d5289, 32'shc02d8e64, 32'shc02dca67, 32'shc02e0691, 
               32'shc02e42e2, 32'shc02e7f5b, 32'shc02ebbfb, 32'shc02ef8c2, 32'shc02f35b1, 32'shc02f72c7, 32'shc02fb004, 32'shc02fed69, 
               32'shc0302af5, 32'shc03068a9, 32'shc030a684, 32'shc030e486, 32'shc03122b0, 32'shc0316101, 32'shc0319f79, 32'shc031de19, 
               32'shc0321ce0, 32'shc0325bcf, 32'shc0329ae4, 32'shc032da22, 32'shc0331986, 32'shc0335912, 32'shc03398c5, 32'shc033d8a0, 
               32'shc03418a2, 32'shc03458cb, 32'shc034991c, 32'shc034d994, 32'shc0351a33, 32'shc0355afa, 32'shc0359be8, 32'shc035dcfd, 
               32'shc0361e3a, 32'shc0365f9e, 32'shc036a129, 32'shc036e2dc, 32'shc03724b6, 32'shc03766b8, 32'shc037a8e1, 32'shc037eb31, 
               32'shc0382da8, 32'shc0387047, 32'shc038b30d, 32'shc038f5fb, 32'shc0393910, 32'shc0397c4c, 32'shc039bfaf, 32'shc03a033a, 
               32'shc03a46ed, 32'shc03a8ac6, 32'shc03acec7, 32'shc03b12ef, 32'shc03b573f, 32'shc03b9bb6, 32'shc03be054, 32'shc03c251a, 
               32'shc03c6a07, 32'shc03caf1b, 32'shc03cf456, 32'shc03d39b9, 32'shc03d7f44, 32'shc03dc4f5, 32'shc03e0ace, 32'shc03e50ce, 
               32'shc03e96f6, 32'shc03edd45, 32'shc03f23bb, 32'shc03f6a58, 32'shc03fb11d, 32'shc03ff80a, 32'shc0403f1d, 32'shc0408658, 
               32'shc040cdba, 32'shc0411544, 32'shc0415cf4, 32'shc041a4cd, 32'shc041eccc, 32'shc04234f3, 32'shc0427d41, 32'shc042c5b6, 
               32'shc0430e53, 32'shc0435717, 32'shc043a002, 32'shc043e915, 32'shc044324f, 32'shc0447bb0, 32'shc044c539, 32'shc0450ee9, 
               32'shc04558c0, 32'shc045a2bf, 32'shc045ece5, 32'shc0463732, 32'shc04681a6, 32'shc046cc42, 32'shc0471705, 32'shc04761ef, 
               32'shc047ad01, 32'shc047f83a, 32'shc048439b, 32'shc0488f22, 32'shc048dad1, 32'shc04926a7, 32'shc04972a5, 32'shc049beca, 
               32'shc04a0b16, 32'shc04a5789, 32'shc04aa424, 32'shc04af0e6, 32'shc04b3dcf, 32'shc04b8ae0, 32'shc04bd818, 32'shc04c2577, 
               32'shc04c72fe, 32'shc04cc0ac, 32'shc04d0e81, 32'shc04d5c7d, 32'shc04daaa1, 32'shc04df8ec, 32'shc04e475e, 32'shc04e95f8, 
               32'shc04ee4b8, 32'shc04f33a1, 32'shc04f82b0, 32'shc04fd1e7, 32'shc0502145, 32'shc05070ca, 32'shc050c077, 32'shc051104a, 
               32'shc0516045, 32'shc051b068, 32'shc05200b2, 32'shc0525123, 32'shc052a1bb, 32'shc052f27a, 32'shc0534361, 32'shc053946f, 
               32'shc053e5a5, 32'shc0543701, 32'shc0548885, 32'shc054da30, 32'shc0552c03, 32'shc0557dfd, 32'shc055d01e, 32'shc0562266, 
               32'shc05674d6, 32'shc056c76c, 32'shc0571a2b, 32'shc0576d10, 32'shc057c01d, 32'shc0581350, 32'shc05866ac, 32'shc058ba2e, 
               32'shc0590dd8, 32'shc05961a9, 32'shc059b5a1, 32'shc05a09c0, 32'shc05a5e07, 32'shc05ab275, 32'shc05b070a, 32'shc05b5bc7, 
               32'shc05bb0ab, 32'shc05c05b6, 32'shc05c5ae8, 32'shc05cb042, 32'shc05d05c3, 32'shc05d5b6b, 32'shc05db13a, 32'shc05e0730, 
               32'shc05e5d4e, 32'shc05eb393, 32'shc05f0a00, 32'shc05f6093, 32'shc05fb74e, 32'shc0600e30, 32'shc060653a, 32'shc060bc6a, 
               32'shc06113c2, 32'shc0616b41, 32'shc061c2e7, 32'shc0621ab5, 32'shc06272aa, 32'shc062cac6, 32'shc0632309, 32'shc0637b73, 
               32'shc063d405, 32'shc0642cbe, 32'shc064859e, 32'shc064dea6, 32'shc06537d4, 32'shc065912a, 32'shc065eaa8, 32'shc066444c, 
               32'shc0669e18, 32'shc066f80a, 32'shc0675225, 32'shc067ac66, 32'shc06806ce, 32'shc068615e, 32'shc068bc15, 32'shc06916f3, 
               32'shc06971f9, 32'shc069cd26, 32'shc06a2879, 32'shc06a83f5, 32'shc06adf97, 32'shc06b3b60, 32'shc06b9751, 32'shc06bf369, 
               32'shc06c4fa8, 32'shc06cac0f, 32'shc06d089d, 32'shc06d6551, 32'shc06dc22e, 32'shc06e1f31, 32'shc06e7c5b, 32'shc06ed9ad, 
               32'shc06f3726, 32'shc06f94c6, 32'shc06ff28e, 32'shc070507c, 32'shc070ae92, 32'shc0710ccf, 32'shc0716b33, 32'shc071c9be, 
               32'shc0722871, 32'shc072874b, 32'shc072e64c, 32'shc0734574, 32'shc073a4c3, 32'shc074043a, 32'shc07463d8, 32'shc074c39d, 
               32'shc0752389, 32'shc075839c, 32'shc075e3d7, 32'shc0764439, 32'shc076a4c2, 32'shc0770572, 32'shc0776649, 32'shc077c748, 
               32'shc078286e, 32'shc07889bb, 32'shc078eb2f, 32'shc0794cca, 32'shc079ae8c, 32'shc07a1076, 32'shc07a7287, 32'shc07ad4bf, 
               32'shc07b371e, 32'shc07b99a5, 32'shc07bfc52, 32'shc07c5f27, 32'shc07cc223, 32'shc07d2546, 32'shc07d8890, 32'shc07dec02, 
               32'shc07e4f9b, 32'shc07eb35a, 32'shc07f1741, 32'shc07f7b50, 32'shc07fdf85, 32'shc08043e1, 32'shc080a865, 32'shc0810d10, 
               32'shc08171e2, 32'shc081d6db, 32'shc0823bfb, 32'shc082a143, 32'shc08306b2, 32'shc0836c47, 32'shc083d204, 32'shc08437e9, 
               32'shc0849df4, 32'shc0850426, 32'shc0856a80, 32'shc085d101, 32'shc08637a9, 32'shc0869e78, 32'shc087056e, 32'shc0876c8c, 
               32'shc087d3d0, 32'shc0883b3c, 32'shc088a2cf, 32'shc0890a89, 32'shc089726a, 32'shc089da72, 32'shc08a42a2, 32'shc08aaaf8, 
               32'shc08b1376, 32'shc08b7c1b, 32'shc08be4e7, 32'shc08c4dda, 32'shc08cb6f5, 32'shc08d2036, 32'shc08d899f, 32'shc08df32e, 
               32'shc08e5ce5, 32'shc08ec6c3, 32'shc08f30c8, 32'shc08f9af5, 32'shc0900548, 32'shc0906fc3, 32'shc090da64, 32'shc091452d, 
               32'shc091b01d, 32'shc0921b34, 32'shc0928672, 32'shc092f1d7, 32'shc0935d64, 32'shc093c917, 32'shc09434f2, 32'shc094a0f4, 
               32'shc0950d1d, 32'shc095796d, 32'shc095e5e4, 32'shc0965282, 32'shc096bf48, 32'shc0972c34, 32'shc0979948, 32'shc0980683, 
               32'shc09873e4, 32'shc098e16d, 32'shc0994f1d, 32'shc099bcf5, 32'shc09a2af3, 32'shc09a9918, 32'shc09b0765, 32'shc09b75d8, 
               32'shc09be473, 32'shc09c5335, 32'shc09cc21e, 32'shc09d312e, 32'shc09da065, 32'shc09e0fc3, 32'shc09e7f48, 32'shc09eeef5, 
               32'shc09f5ec8, 32'shc09fcec3, 32'shc0a03ee4, 32'shc0a0af2d, 32'shc0a11f9d, 32'shc0a19034, 32'shc0a200f2, 32'shc0a271d7, 
               32'shc0a2e2e3, 32'shc0a35417, 32'shc0a3c571, 32'shc0a436f3, 32'shc0a4a89b, 32'shc0a51a6b, 32'shc0a58c62, 32'shc0a5fe7f, 
               32'shc0a670c4, 32'shc0a6e330, 32'shc0a755c3, 32'shc0a7c87d, 32'shc0a83b5e, 32'shc0a8ae67, 32'shc0a92196, 32'shc0a994ec, 
               32'shc0aa086a, 32'shc0aa7c0e, 32'shc0aaefda, 32'shc0ab63cd, 32'shc0abd7e6, 32'shc0ac4c27, 32'shc0acc08f, 32'shc0ad351e, 
               32'shc0ada9d4, 32'shc0ae1eb1, 32'shc0ae93b5, 32'shc0af08e0, 32'shc0af7e33, 32'shc0aff3ac, 32'shc0b0694c, 32'shc0b0df13, 
               32'shc0b15502, 32'shc0b1cb17, 32'shc0b24154, 32'shc0b2b7b8, 32'shc0b32e42, 32'shc0b3a4f4, 32'shc0b41bcd, 32'shc0b492cc, 
               32'shc0b509f3, 32'shc0b58141, 32'shc0b5f8b6, 32'shc0b67052, 32'shc0b6e815, 32'shc0b75fff, 32'shc0b7d810, 32'shc0b85048, 
               32'shc0b8c8a7, 32'shc0b9412d, 32'shc0b9b9da, 32'shc0ba32af, 32'shc0baabaa, 32'shc0bb24cc, 32'shc0bb9e15, 32'shc0bc1786, 
               32'shc0bc911d, 32'shc0bd0adb, 32'shc0bd84c1, 32'shc0bdfecd, 32'shc0be7901, 32'shc0bef35b, 32'shc0bf6ddd, 32'shc0bfe885, 
               32'shc0c06355, 32'shc0c0de4b, 32'shc0c15969, 32'shc0c1d4ad, 32'shc0c25019, 32'shc0c2cbab, 32'shc0c34765, 32'shc0c3c346, 
               32'shc0c43f4d, 32'shc0c4bb7c, 32'shc0c537d1, 32'shc0c5b44e, 32'shc0c630f2, 32'shc0c6adbc, 32'shc0c72aae, 32'shc0c7a7c6, 
               32'shc0c82506, 32'shc0c8a26d, 32'shc0c91ffa, 32'shc0c99daf, 32'shc0ca1b8a, 32'shc0ca998d, 32'shc0cb17b7, 32'shc0cb9607, 
               32'shc0cc147f, 32'shc0cc931d, 32'shc0cd11e3, 32'shc0cd90cf, 32'shc0ce0fe3, 32'shc0ce8f1d, 32'shc0cf0e7f, 32'shc0cf8e07, 
               32'shc0d00db6, 32'shc0d08d8d, 32'shc0d10d8a, 32'shc0d18dae, 32'shc0d20dfa, 32'shc0d28e6c, 32'shc0d30f05, 32'shc0d38fc6, 
               32'shc0d410ad, 32'shc0d491bb, 32'shc0d512f0, 32'shc0d5944c, 32'shc0d615cf, 32'shc0d69779, 32'shc0d7194a, 32'shc0d79b42, 
               32'shc0d81d61, 32'shc0d89fa7, 32'shc0d92214, 32'shc0d9a4a7, 32'shc0da2762, 32'shc0daaa44, 32'shc0db2d4c, 32'shc0dbb07c, 
               32'shc0dc33d2, 32'shc0dcb750, 32'shc0dd3af4, 32'shc0ddbec0, 32'shc0de42b2, 32'shc0dec6cb, 32'shc0df4b0b, 32'shc0dfcf73, 
               32'shc0e05401, 32'shc0e0d8b6, 32'shc0e15d92, 32'shc0e1e294, 32'shc0e267be, 32'shc0e2ed0f, 32'shc0e37287, 32'shc0e3f825, 
               32'shc0e47deb, 32'shc0e503d7, 32'shc0e589eb, 32'shc0e61025, 32'shc0e69686, 32'shc0e71d0e, 32'shc0e7a3bd, 32'shc0e82a93, 
               32'shc0e8b190, 32'shc0e938b4, 32'shc0e9bfff, 32'shc0ea4771, 32'shc0eacf09, 32'shc0eb56c9, 32'shc0ebdeaf, 32'shc0ec66bc, 
               32'shc0eceef1, 32'shc0ed774c, 32'shc0edffce, 32'shc0ee8877, 32'shc0ef1147, 32'shc0ef9a3d, 32'shc0f0235b, 32'shc0f0aca0, 
               32'shc0f1360b, 32'shc0f1bf9d, 32'shc0f24957, 32'shc0f2d337, 32'shc0f35d3e, 32'shc0f3e76c, 32'shc0f471c1, 32'shc0f4fc3c, 
               32'shc0f586df, 32'shc0f611a8, 32'shc0f69c99, 32'shc0f727b0, 32'shc0f7b2ee, 32'shc0f83e53, 32'shc0f8c9df, 32'shc0f95592, 
               32'shc0f9e16b, 32'shc0fa6d6c, 32'shc0faf993, 32'shc0fb85e2, 32'shc0fc1257, 32'shc0fc9ef3, 32'shc0fd2bb6, 32'shc0fdb8a0, 
               32'shc0fe45b0, 32'shc0fed2e8, 32'shc0ff6046, 32'shc0ffedcb, 32'shc1007b77, 32'shc101094a, 32'shc1019744, 32'shc1022565, 
               32'shc102b3ac, 32'shc103421b, 32'shc103d0b0, 32'shc1045f6c, 32'shc104ee4f, 32'shc1057d59, 32'shc1060c89, 32'shc1069be1, 
               32'shc1072b5f, 32'shc107bb04, 32'shc1084ad0, 32'shc108dac3, 32'shc1096add, 32'shc109fb1d, 32'shc10a8b85, 32'shc10b1c13, 
               32'shc10bacc8, 32'shc10c3da4, 32'shc10ccea6, 32'shc10d5fd0, 32'shc10df120, 32'shc10e8297, 32'shc10f1435, 32'shc10fa5fa, 
               32'shc11037e6, 32'shc110c9f8, 32'shc1115c32, 32'shc111ee92, 32'shc1128119, 32'shc11313c7, 32'shc113a69b, 32'shc1143997, 
               32'shc114ccb9, 32'shc1156002, 32'shc115f372, 32'shc1168708, 32'shc1171ac6, 32'shc117aeaa, 32'shc11842b5, 32'shc118d6e7, 
               32'shc1196b3f, 32'shc119ffbf, 32'shc11a9465, 32'shc11b2932, 32'shc11bbe26, 32'shc11c5341, 32'shc11ce882, 32'shc11d7dea, 
               32'shc11e1379, 32'shc11ea92f, 32'shc11f3f0c, 32'shc11fd50f, 32'shc1206b39, 32'shc121018a, 32'shc1219802, 32'shc1222ea1, 
               32'shc122c566, 32'shc1235c52, 32'shc123f365, 32'shc1248a9e, 32'shc12521ff, 32'shc125b986, 32'shc1265134, 32'shc126e909, 
               32'shc1278104, 32'shc1281926, 32'shc128b16f, 32'shc12949df, 32'shc129e276, 32'shc12a7b33, 32'shc12b1417, 32'shc12bad22, 
               32'shc12c4653, 32'shc12cdfac, 32'shc12d792b, 32'shc12e12d1, 32'shc12eac9d, 32'shc12f4690, 32'shc12fe0ab, 32'shc1307aeb, 
               32'shc1311553, 32'shc131afe1, 32'shc1324a96, 32'shc132e572, 32'shc1338075, 32'shc1341b9e, 32'shc134b6ee, 32'shc1355265, 
               32'shc135ee02, 32'shc13689c6, 32'shc13725b1, 32'shc137c1c3, 32'shc1385dfb, 32'shc138fa5a, 32'shc13996e0, 32'shc13a338d, 
               32'shc13ad060, 32'shc13b6d5a, 32'shc13c0a7b, 32'shc13ca7c2, 32'shc13d4530, 32'shc13de2c5, 32'shc13e8081, 32'shc13f1e63, 
               32'shc13fbc6c, 32'shc1405a9c, 32'shc140f8f2, 32'shc141976f, 32'shc1423613, 32'shc142d4de, 32'shc14373cf, 32'shc14412e7, 
               32'shc144b225, 32'shc145518b, 32'shc145f117, 32'shc14690ca, 32'shc14730a3, 32'shc147d0a3, 32'shc14870ca, 32'shc1491117, 
               32'shc149b18b, 32'shc14a5226, 32'shc14af2e8, 32'shc14b93d0, 32'shc14c34df, 32'shc14cd614, 32'shc14d7771, 32'shc14e18f3, 
               32'shc14eba9d, 32'shc14f5c6d, 32'shc14ffe64, 32'shc150a082, 32'shc15142c6, 32'shc151e531, 32'shc15287c3, 32'shc1532a7b, 
               32'shc153cd5a, 32'shc154705f, 32'shc155138c, 32'shc155b6de, 32'shc1565a58, 32'shc156fdf8, 32'shc157a1bf, 32'shc15845ac, 
               32'shc158e9c1, 32'shc1598dfb, 32'shc15a325d, 32'shc15ad6e5, 32'shc15b7b94, 32'shc15c2069, 32'shc15cc565, 32'shc15d6a88, 
               32'shc15e0fd1, 32'shc15eb541, 32'shc15f5ad7, 32'shc1600095, 32'shc160a678, 32'shc1614c83, 32'shc161f2b4, 32'shc162990c, 
               32'shc1633f8a, 32'shc163e62f, 32'shc1648cfa, 32'shc16533ed, 32'shc165db05, 32'shc1668245, 32'shc16729ab, 32'shc167d137, 
               32'shc16878eb, 32'shc16920c5, 32'shc169c8c5, 32'shc16a70ec, 32'shc16b193a, 32'shc16bc1ae, 32'shc16c6a49, 32'shc16d130a, 
               32'shc16dbbf3, 32'shc16e6501, 32'shc16f0e36, 32'shc16fb792, 32'shc1706115, 32'shc1710abe, 32'shc171b48e, 32'shc1725e84, 
               32'shc17308a1, 32'shc173b2e4, 32'shc1745d4e, 32'shc17507df, 32'shc175b296, 32'shc1765d73, 32'shc1770878, 32'shc177b3a3, 
               32'shc1785ef4, 32'shc1790a6c, 32'shc179b60b, 32'shc17a61d0, 32'shc17b0dbb, 32'shc17bb9ce, 32'shc17c6607, 32'shc17d1266, 
               32'shc17dbeec, 32'shc17e6b99, 32'shc17f186c, 32'shc17fc565, 32'shc1807285, 32'shc1811fcc, 32'shc181cd3a, 32'shc1827acd, 
               32'shc1832888, 32'shc183d669, 32'shc1848470, 32'shc185329e, 32'shc185e0f3, 32'shc1868f6e, 32'shc1873e10, 32'shc187ecd8, 
               32'shc1889bc6, 32'shc1894adc, 32'shc189fa17, 32'shc18aa97a, 32'shc18b5903, 32'shc18c08b2, 32'shc18cb888, 32'shc18d6884, 
               32'shc18e18a7, 32'shc18ec8f1, 32'shc18f7961, 32'shc19029f7, 32'shc190dab4, 32'shc1918b98, 32'shc1923ca2, 32'shc192edd2, 
               32'shc1939f29, 32'shc19450a7, 32'shc195024b, 32'shc195b415, 32'shc1966606, 32'shc197181e, 32'shc197ca5c, 32'shc1987cc1, 
               32'shc1992f4c, 32'shc199e1fd, 32'shc19a94d5, 32'shc19b47d4, 32'shc19bfaf9, 32'shc19cae44, 32'shc19d61b6, 32'shc19e154e, 
               32'shc19ec90d, 32'shc19f7cf3, 32'shc1a030ff, 32'shc1a0e531, 32'shc1a1998a, 32'shc1a24e09, 32'shc1a302af, 32'shc1a3b77b, 
               32'shc1a46c6e, 32'shc1a52187, 32'shc1a5d6c7, 32'shc1a68c2d, 32'shc1a741b9, 32'shc1a7f76c, 32'shc1a8ad46, 32'shc1a96346, 
               32'shc1aa196c, 32'shc1aacfb9, 32'shc1ab862c, 32'shc1ac3cc6, 32'shc1acf386, 32'shc1adaa6d, 32'shc1ae617a, 32'shc1af18ae, 
               32'shc1afd007, 32'shc1b08788, 32'shc1b13f2f, 32'shc1b1f6fc, 32'shc1b2aef0, 32'shc1b3670a, 32'shc1b41f4a, 32'shc1b4d7b1, 
               32'shc1b5903f, 32'shc1b648f3, 32'shc1b701cd, 32'shc1b7bacd, 32'shc1b873f5, 32'shc1b92d42, 32'shc1b9e6b6, 32'shc1baa050, 
               32'shc1bb5a11, 32'shc1bc13f8, 32'shc1bcce06, 32'shc1bd883a, 32'shc1be4294, 32'shc1befd15, 32'shc1bfb7bc, 32'shc1c0728a, 
               32'shc1c12d7e, 32'shc1c1e898, 32'shc1c2a3d9, 32'shc1c35f40, 32'shc1c41ace, 32'shc1c4d682, 32'shc1c5925c, 32'shc1c64e5d, 
               32'shc1c70a84, 32'shc1c7c6d1, 32'shc1c88345, 32'shc1c93fdf, 32'shc1c9fca0, 32'shc1cab987, 32'shc1cb7694, 32'shc1cc33c8, 
               32'shc1ccf122, 32'shc1cdaea3, 32'shc1ce6c49, 32'shc1cf2a17, 32'shc1cfe80a, 32'shc1d0a624, 32'shc1d16464, 32'shc1d222cb, 
               32'shc1d2e158, 32'shc1d3a00b, 32'shc1d45ee5, 32'shc1d51de5, 32'shc1d5dd0c, 32'shc1d69c58, 32'shc1d75bcb, 32'shc1d81b65, 
               32'shc1d8db25, 32'shc1d99b0b, 32'shc1da5b17, 32'shc1db1b4a, 32'shc1dbdba3, 32'shc1dc9c23, 32'shc1dd5cc8, 32'shc1de1d94, 
               32'shc1dede87, 32'shc1df9fa0, 32'shc1e060df, 32'shc1e12244, 32'shc1e1e3d0, 32'shc1e2a582, 32'shc1e3675a, 32'shc1e42959, 
               32'shc1e4eb7e, 32'shc1e5adc9, 32'shc1e6703b, 32'shc1e732d3, 32'shc1e7f591, 32'shc1e8b876, 32'shc1e97b80, 32'shc1ea3eb1, 
               32'shc1eb0209, 32'shc1ebc587, 32'shc1ec892b, 32'shc1ed4cf5, 32'shc1ee10e5, 32'shc1eed4fc, 32'shc1ef9939, 32'shc1f05d9d, 
               32'shc1f12227, 32'shc1f1e6d7, 32'shc1f2abad, 32'shc1f370a9, 32'shc1f435cc, 32'shc1f4fb15, 32'shc1f5c085, 32'shc1f6861a, 
               32'shc1f74bd6, 32'shc1f811b9, 32'shc1f8d7c1, 32'shc1f99df0, 32'shc1fa6445, 32'shc1fb2ac0, 32'shc1fbf161, 32'shc1fcb829, 
               32'shc1fd7f17, 32'shc1fe462b, 32'shc1ff0d66, 32'shc1ffd4c7, 32'shc2009c4e, 32'shc20163fb, 32'shc2022bce, 32'shc202f3c8, 
               32'shc203bbe8, 32'shc204842e, 32'shc2054c9b, 32'shc206152d, 32'shc206dde6, 32'shc207a6c5, 32'shc2086fca, 32'shc20938f6, 
               32'shc20a0248, 32'shc20acbc0, 32'shc20b955e, 32'shc20c5f22, 32'shc20d290d, 32'shc20df31e, 32'shc20ebd55, 32'shc20f87b2, 
               32'shc2105236, 32'shc2111cdf, 32'shc211e7af, 32'shc212b2a5, 32'shc2137dc2, 32'shc2144904, 32'shc215146d, 32'shc215dffc, 
               32'shc216abb1, 32'shc217778c, 32'shc218438e, 32'shc2190fb5, 32'shc219dc03, 32'shc21aa877, 32'shc21b7511, 32'shc21c41d2, 
               32'shc21d0eb8, 32'shc21ddbc5, 32'shc21ea8f8, 32'shc21f7651, 32'shc22043d0, 32'shc2211176, 32'shc221df41, 32'shc222ad33, 
               32'shc2237b4b, 32'shc2244989, 32'shc22517ed, 32'shc225e677, 32'shc226b528, 32'shc22783fe, 32'shc22852fb, 32'shc229221e, 
               32'shc229f167, 32'shc22ac0d7, 32'shc22b906c, 32'shc22c6028, 32'shc22d3009, 32'shc22e0011, 32'shc22ed03f, 32'shc22fa093, 
               32'shc230710d, 32'shc23141ae, 32'shc2321274, 32'shc232e361, 32'shc233b473, 32'shc23485ac, 32'shc235570b, 32'shc2362890, 
               32'shc236fa3b, 32'shc237cc0d, 32'shc2389e04, 32'shc2397021, 32'shc23a4265, 32'shc23b14cf, 32'shc23be75f, 32'shc23cba15, 
               32'shc23d8cf1, 32'shc23e5ff3, 32'shc23f331b, 32'shc2400669, 32'shc240d9de, 32'shc241ad78, 32'shc2428139, 32'shc243551f, 
               32'shc244292c, 32'shc244fd5f, 32'shc245d1b8, 32'shc246a637, 32'shc2477adc, 32'shc2484fa7, 32'shc2492498, 32'shc249f9af, 
               32'shc24aceed, 32'shc24ba450, 32'shc24c79d9, 32'shc24d4f89, 32'shc24e255e, 32'shc24efb5a, 32'shc24fd17c, 32'shc250a7c3, 
               32'shc2517e31, 32'shc25254c5, 32'shc2532b7f, 32'shc254025f, 32'shc254d965, 32'shc255b091, 32'shc25687e3, 32'shc2575f5b, 
               32'shc25836f9, 32'shc2590ebd, 32'shc259e6a7, 32'shc25abeb7, 32'shc25b96ee, 32'shc25c6f4a, 32'shc25d47cc, 32'shc25e2074, 
               32'shc25ef943, 32'shc25fd237, 32'shc260ab51, 32'shc2618492, 32'shc2625df8, 32'shc2633785, 32'shc2641137, 32'shc264eb0f, 
               32'shc265c50e, 32'shc2669f32, 32'shc267797c, 32'shc26853ed, 32'shc2692e83, 32'shc26a093f, 32'shc26ae422, 32'shc26bbf2a, 
               32'shc26c9a58, 32'shc26d75ad, 32'shc26e5127, 32'shc26f2cc7, 32'shc270088e, 32'shc270e47a, 32'shc271c08c, 32'shc2729cc4, 
               32'shc2737922, 32'shc27455a6, 32'shc2753250, 32'shc2760f20, 32'shc276ec16, 32'shc277c932, 32'shc278a674, 32'shc27983dc, 
               32'shc27a616a, 32'shc27b3f1e, 32'shc27c1cf7, 32'shc27cfaf7, 32'shc27dd91c, 32'shc27eb768, 32'shc27f95d9, 32'shc2807471, 
               32'shc281532e, 32'shc2823211, 32'shc283111b, 32'shc283f04a, 32'shc284cf9f, 32'shc285af1a, 32'shc2868ebb, 32'shc2876e82, 
               32'shc2884e6e, 32'shc2892e81, 32'shc28a0eb9, 32'shc28aef18, 32'shc28bcf9c, 32'shc28cb047, 32'shc28d9117, 32'shc28e720d, 
               32'shc28f5329, 32'shc290346b, 32'shc29115d3, 32'shc291f760, 32'shc292d914, 32'shc293baed, 32'shc2949ced, 32'shc2957f12, 
               32'shc296615d, 32'shc29743ce, 32'shc2982665, 32'shc2990922, 32'shc299ec05, 32'shc29acf0d, 32'shc29bb23c, 32'shc29c9590, 
               32'shc29d790a, 32'shc29e5caa, 32'shc29f4070, 32'shc2a0245c, 32'shc2a1086d, 32'shc2a1eca5, 32'shc2a2d102, 32'shc2a3b585, 
               32'shc2a49a2e, 32'shc2a57efd, 32'shc2a663f2, 32'shc2a7490c, 32'shc2a82e4d, 32'shc2a913b3, 32'shc2a9f93f, 32'shc2aadef1, 
               32'shc2abc4c9, 32'shc2acaac6, 32'shc2ad90ea, 32'shc2ae7733, 32'shc2af5da2, 32'shc2b04437, 32'shc2b12af1, 32'shc2b211d2, 
               32'shc2b2f8d8, 32'shc2b3e004, 32'shc2b4c756, 32'shc2b5aece, 32'shc2b6966c, 32'shc2b77e2f, 32'shc2b86618, 32'shc2b94e27, 
               32'shc2ba365c, 32'shc2bb1eb6, 32'shc2bc0737, 32'shc2bcefdd, 32'shc2bdd8a9, 32'shc2bec19b, 32'shc2bfaab2, 32'shc2c093ef, 
               32'shc2c17d52, 32'shc2c266db, 32'shc2c3508a, 32'shc2c43a5e, 32'shc2c52459, 32'shc2c60e78, 32'shc2c6f8be, 32'shc2c7e32a, 
               32'shc2c8cdbb, 32'shc2c9b872, 32'shc2caa34f, 32'shc2cb8e51, 32'shc2cc7979, 32'shc2cd64c7, 32'shc2ce503b, 32'shc2cf3bd5, 
               32'shc2d02794, 32'shc2d11379, 32'shc2d1ff84, 32'shc2d2ebb4, 32'shc2d3d80a, 32'shc2d4c486, 32'shc2d5b128, 32'shc2d69df0, 
               32'shc2d78add, 32'shc2d877f0, 32'shc2d96528, 32'shc2da5286, 32'shc2db400a, 32'shc2dc2db4, 32'shc2dd1b84, 32'shc2de0979, 
               32'shc2def794, 32'shc2dfe5d4, 32'shc2e0d43b, 32'shc2e1c2c7, 32'shc2e2b178, 32'shc2e3a050, 32'shc2e48f4d, 32'shc2e57e70, 
               32'shc2e66db8, 32'shc2e75d26, 32'shc2e84cba, 32'shc2e93c74, 32'shc2ea2c53, 32'shc2eb1c58, 32'shc2ec0c82, 32'shc2ecfcd3, 
               32'shc2eded49, 32'shc2eedde4, 32'shc2efcea6, 32'shc2f0bf8c, 32'shc2f1b099, 32'shc2f2a1cb, 32'shc2f39323, 32'shc2f484a1, 
               32'shc2f57644, 32'shc2f6680d, 32'shc2f759fc, 32'shc2f84c10, 32'shc2f93e4a, 32'shc2fa30a9, 32'shc2fb232e, 32'shc2fc15d9, 
               32'shc2fd08a9, 32'shc2fdfb9f, 32'shc2feeebb, 32'shc2ffe1fc, 32'shc300d563, 32'shc301c8f0, 32'shc302bca2, 32'shc303b07a, 
               32'shc304a477, 32'shc305989a, 32'shc3068ce3, 32'shc3078151, 32'shc30875e5, 32'shc3096a9f, 32'shc30a5f7e, 32'shc30b5482, 
               32'shc30c49ad, 32'shc30d3efd, 32'shc30e3472, 32'shc30f2a0d, 32'shc3101fce, 32'shc31115b4, 32'shc3120bc0, 32'shc31301f1, 
               32'shc313f848, 32'shc314eec5, 32'shc315e567, 32'shc316dc2f, 32'shc317d31c, 32'shc318ca2f, 32'shc319c168, 32'shc31ab8c6, 
               32'shc31bb049, 32'shc31ca7f2, 32'shc31d9fc1, 32'shc31e97b5, 32'shc31f8fcf, 32'shc320880e, 32'shc3218073, 32'shc32278fe, 
               32'shc32371ae, 32'shc3246a83, 32'shc325637f, 32'shc3265c9f, 32'shc32755e5, 32'shc3284f51, 32'shc32948e2, 32'shc32a4299, 
               32'shc32b3c75, 32'shc32c3677, 32'shc32d309e, 32'shc32e2aeb, 32'shc32f255e, 32'shc3301ff5, 32'shc3311ab3, 32'shc3321596, 
               32'shc333109e, 32'shc3340bcc, 32'shc3350720, 32'shc3360298, 32'shc336fe37, 32'shc337f9fb, 32'shc338f5e4, 32'shc339f1f3, 
               32'shc33aee27, 32'shc33bea81, 32'shc33ce701, 32'shc33de3a5, 32'shc33ee070, 32'shc33fdd60, 32'shc340da75, 32'shc341d7b0, 
               32'shc342d510, 32'shc343d295, 32'shc344d041, 32'shc345ce11, 32'shc346cc07, 32'shc347ca23, 32'shc348c864, 32'shc349c6ca, 
               32'shc34ac556, 32'shc34bc407, 32'shc34cc2de, 32'shc34dc1da, 32'shc34ec0fc, 32'shc34fc043, 32'shc350bfaf, 32'shc351bf41, 
               32'shc352bef9, 32'shc353bed6, 32'shc354bed8, 32'shc355bf00, 32'shc356bf4d, 32'shc357bfbf, 32'shc358c057, 32'shc359c114, 
               32'shc35ac1f7, 32'shc35bc2ff, 32'shc35cc42d, 32'shc35dc580, 32'shc35ec6f8, 32'shc35fc896, 32'shc360ca59, 32'shc361cc42, 
               32'shc362ce50, 32'shc363d083, 32'shc364d2dc, 32'shc365d55a, 32'shc366d7fd, 32'shc367dac6, 32'shc368ddb4, 32'shc369e0c8, 
               32'shc36ae401, 32'shc36be75f, 32'shc36ceae3, 32'shc36dee8c, 32'shc36ef25b, 32'shc36ff64e, 32'shc370fa68, 32'shc371fea6, 
               32'shc373030a, 32'shc3740793, 32'shc3750c42, 32'shc3761116, 32'shc377160f, 32'shc3781b2e, 32'shc3792072, 32'shc37a25db, 
               32'shc37b2b6a, 32'shc37c311e, 32'shc37d36f7, 32'shc37e3cf6, 32'shc37f4319, 32'shc3804963, 32'shc3814fd1, 32'shc3825665, 
               32'shc3835d1e, 32'shc38463fd, 32'shc3856b01, 32'shc386722a, 32'shc3877978, 32'shc38880ec, 32'shc3898885, 32'shc38a9043, 
               32'shc38b9827, 32'shc38ca030, 32'shc38da85e, 32'shc38eb0b2, 32'shc38fb92a, 32'shc390c1c9, 32'shc391ca8c, 32'shc392d375, 
               32'shc393dc82, 32'shc394e5b6, 32'shc395ef0e, 32'shc396f88c, 32'shc398022f, 32'shc3990bf7, 32'shc39a15e4, 32'shc39b1ff7, 
               32'shc39c2a2f, 32'shc39d348c, 32'shc39e3f0f, 32'shc39f49b7, 32'shc3a05484, 32'shc3a15f76, 32'shc3a26a8d, 32'shc3a375ca, 
               32'shc3a4812c, 32'shc3a58cb3, 32'shc3a6985f, 32'shc3a7a431, 32'shc3a8b028, 32'shc3a9bc44, 32'shc3aac885, 32'shc3abd4ec, 
               32'shc3ace178, 32'shc3adee28, 32'shc3aefaff, 32'shc3b007fa, 32'shc3b1151b, 32'shc3b22260, 32'shc3b32fcb, 32'shc3b43d5b, 
               32'shc3b54b11, 32'shc3b658eb, 32'shc3b766eb, 32'shc3b87510, 32'shc3b9835a, 32'shc3ba91c9, 32'shc3bba05e, 32'shc3bcaf17, 
               32'shc3bdbdf6, 32'shc3beccfa, 32'shc3bfdc23, 32'shc3c0eb71, 32'shc3c1fae5, 32'shc3c30a7e, 32'shc3c41a3b, 32'shc3c52a1e, 
               32'shc3c63a26, 32'shc3c74a54, 32'shc3c85aa6, 32'shc3c96b1e, 32'shc3ca7bba, 32'shc3cb8c7c, 32'shc3cc9d63, 32'shc3cdae6f, 
               32'shc3cebfa0, 32'shc3cfd0f7, 32'shc3d0e272, 32'shc3d1f413, 32'shc3d305d8, 32'shc3d417c3, 32'shc3d529d3, 32'shc3d63c08, 
               32'shc3d74e62, 32'shc3d860e2, 32'shc3d97386, 32'shc3da8650, 32'shc3db993e, 32'shc3dcac52, 32'shc3ddbf8b, 32'shc3ded2e9, 
               32'shc3dfe66c, 32'shc3e0fa14, 32'shc3e20de1, 32'shc3e321d3, 32'shc3e435ea, 32'shc3e54a27, 32'shc3e65e88, 32'shc3e7730f, 
               32'shc3e887bb, 32'shc3e99c8b, 32'shc3eab181, 32'shc3ebc69c, 32'shc3ecdbdc, 32'shc3edf141, 32'shc3ef06cb, 32'shc3f01c7a, 
               32'shc3f1324e, 32'shc3f24847, 32'shc3f35e65, 32'shc3f474a8, 32'shc3f58b10, 32'shc3f6a19e, 32'shc3f7b850, 32'shc3f8cf27, 
               32'shc3f9e624, 32'shc3fafd45, 32'shc3fc148c, 32'shc3fd2bf7, 32'shc3fe4388, 32'shc3ff5b3d, 32'shc4007318, 32'shc4018b17, 
               32'shc402a33c, 32'shc403bb85, 32'shc404d3f4, 32'shc405ec87, 32'shc4070540, 32'shc4081e1d, 32'shc4093720, 32'shc40a5047, 
               32'shc40b6994, 32'shc40c8305, 32'shc40d9c9c, 32'shc40eb657, 32'shc40fd037, 32'shc410ea3d, 32'shc4120467, 32'shc4131eb7, 
               32'shc414392b, 32'shc41553c4, 32'shc4166e82, 32'shc4178965, 32'shc418a46d, 32'shc419bf9b, 32'shc41adaed, 32'shc41bf664, 
               32'shc41d11ff, 32'shc41e2dc0, 32'shc41f49a6, 32'shc42065b1, 32'shc42181e0, 32'shc4229e35, 32'shc423baae, 32'shc424d74d, 
               32'shc425f410, 32'shc42710f9, 32'shc4282e06, 32'shc4294b38, 32'shc42a688f, 32'shc42b860b, 32'shc42ca3ac, 32'shc42dc171, 
               32'shc42edf5c, 32'shc42ffd6b, 32'shc4311ba0, 32'shc43239f9, 32'shc4335877, 32'shc434771b, 32'shc43595e3, 32'shc436b4cf, 
               32'shc437d3e1, 32'shc438f318, 32'shc43a1273, 32'shc43b31f4, 32'shc43c5199, 32'shc43d7163, 32'shc43e9152, 32'shc43fb166, 
               32'shc440d19e, 32'shc441f1fc, 32'shc443127e, 32'shc4443326, 32'shc44553f2, 32'shc44674e3, 32'shc44795f8, 32'shc448b733, 
               32'shc449d892, 32'shc44afa17, 32'shc44c1bc0, 32'shc44d3d8e, 32'shc44e5f80, 32'shc44f8198, 32'shc450a3d4, 32'shc451c636, 
               32'shc452e8bc, 32'shc4540b67, 32'shc4552e36, 32'shc456512b, 32'shc4577444, 32'shc4589782, 32'shc459bae5, 32'shc45ade6c, 
               32'shc45c0219, 32'shc45d25ea, 32'shc45e49e0, 32'shc45f6dfb, 32'shc460923b, 32'shc461b69f, 32'shc462db28, 32'shc463ffd6, 
               32'shc46524a9, 32'shc46649a0, 32'shc4676ebc, 32'shc46893fd, 32'shc469b963, 32'shc46adeee, 32'shc46c049d, 32'shc46d2a71, 
               32'shc46e5069, 32'shc46f7687, 32'shc4709cc9, 32'shc471c330, 32'shc472e9bc, 32'shc474106c, 32'shc4753741, 32'shc4765e3b, 
               32'shc477855a, 32'shc478ac9d, 32'shc479d405, 32'shc47afb92, 32'shc47c2344, 32'shc47d4b1a, 32'shc47e7315, 32'shc47f9b34, 
               32'shc480c379, 32'shc481ebe2, 32'shc4831470, 32'shc4843d22, 32'shc48565f9, 32'shc4868ef5, 32'shc487b815, 32'shc488e15b, 
               32'shc48a0ac4, 32'shc48b3453, 32'shc48c5e06, 32'shc48d87de, 32'shc48eb1db, 32'shc48fdbfc, 32'shc4910642, 32'shc49230ac, 
               32'shc4935b3c, 32'shc49485ef, 32'shc495b0c8, 32'shc496dbc5, 32'shc49806e7, 32'shc499322d, 32'shc49a5d98, 32'shc49b8928, 
               32'shc49cb4dd, 32'shc49de0b6, 32'shc49f0cb3, 32'shc4a038d6, 32'shc4a1651c, 32'shc4a29188, 32'shc4a3be18, 32'shc4a4eacd, 
               32'shc4a617a6, 32'shc4a744a4, 32'shc4a871c7, 32'shc4a99f0e, 32'shc4aacc7a, 32'shc4abfa0a, 32'shc4ad27bf, 32'shc4ae5599, 
               32'shc4af8397, 32'shc4b0b1ba, 32'shc4b1e001, 32'shc4b30e6d, 32'shc4b43cfd, 32'shc4b56bb3, 32'shc4b69a8c, 32'shc4b7c98a, 
               32'shc4b8f8ad, 32'shc4ba27f5, 32'shc4bb5760, 32'shc4bc86f1, 32'shc4bdb6a6, 32'shc4bee680, 32'shc4c0167e, 32'shc4c146a0, 
               32'shc4c276e8, 32'shc4c3a753, 32'shc4c4d7e4, 32'shc4c60899, 32'shc4c73972, 32'shc4c86a70, 32'shc4c99b92, 32'shc4caccd9, 
               32'shc4cbfe45, 32'shc4cd2fd5, 32'shc4ce6189, 32'shc4cf9363, 32'shc4d0c560, 32'shc4d1f782, 32'shc4d329c9, 32'shc4d45c34, 
               32'shc4d58ec3, 32'shc4d6c177, 32'shc4d7f450, 32'shc4d9274d, 32'shc4da5a6f, 32'shc4db8db5, 32'shc4dcc11f, 32'shc4ddf4ae, 
               32'shc4df2862, 32'shc4e05c3a, 32'shc4e19036, 32'shc4e2c457, 32'shc4e3f89c, 32'shc4e52d06, 32'shc4e66194, 32'shc4e79647, 
               32'shc4e8cb1e, 32'shc4ea001a, 32'shc4eb353a, 32'shc4ec6a7e, 32'shc4ed9fe7, 32'shc4eed575, 32'shc4f00b27, 32'shc4f140fd, 
               32'shc4f276f7, 32'shc4f3ad17, 32'shc4f4e35a, 32'shc4f619c2, 32'shc4f7504e, 32'shc4f886ff, 32'shc4f9bdd4, 32'shc4faf4ce, 
               32'shc4fc2bec, 32'shc4fd632f, 32'shc4fe9a95, 32'shc4ffd221, 32'shc50109d0, 32'shc50241a4, 32'shc503799d, 32'shc504b1b9, 
               32'shc505e9fb, 32'shc5072260, 32'shc5085aea, 32'shc5099398, 32'shc50acc6b, 32'shc50c0562, 32'shc50d3e7d, 32'shc50e77bd, 
               32'shc50fb121, 32'shc510eaaa, 32'shc5122457, 32'shc5135e28, 32'shc514981d, 32'shc515d237, 32'shc5170c75, 32'shc51846d8, 
               32'shc519815f, 32'shc51abc0a, 32'shc51bf6da, 32'shc51d31ce, 32'shc51e6ce6, 32'shc51fa822, 32'shc520e383, 32'shc5221f08, 
               32'shc5235ab2, 32'shc5249680, 32'shc525d272, 32'shc5270e88, 32'shc5284ac3, 32'shc5298722, 32'shc52ac3a5, 32'shc52c004d, 
               32'shc52d3d18, 32'shc52e7a09, 32'shc52fb71d, 32'shc530f456, 32'shc53231b3, 32'shc5336f34, 32'shc534acd9, 32'shc535eaa3, 
               32'shc5372891, 32'shc53866a4, 32'shc539a4da, 32'shc53ae335, 32'shc53c21b4, 32'shc53d6057, 32'shc53e9f1f, 32'shc53fde0b, 
               32'shc5411d1b, 32'shc5425c4f, 32'shc5439ba8, 32'shc544db25, 32'shc5461ac6, 32'shc5475a8b, 32'shc5489a74, 32'shc549da82, 
               32'shc54b1ab4, 32'shc54c5b0a, 32'shc54d9b84, 32'shc54edc23, 32'shc5501ce5, 32'shc5515dcc, 32'shc5529ed7, 32'shc553e007, 
               32'shc555215a, 32'shc55662d2, 32'shc557a46e, 32'shc558e62e, 32'shc55a2812, 32'shc55b6a1a, 32'shc55cac47, 32'shc55dee98, 
               32'shc55f310d, 32'shc56073a6, 32'shc561b663, 32'shc562f944, 32'shc5643c4a, 32'shc5657f74, 32'shc566c2c2, 32'shc5680634, 
               32'shc56949ca, 32'shc56a8d84, 32'shc56bd163, 32'shc56d1565, 32'shc56e598c, 32'shc56f9dd7, 32'shc570e246, 32'shc57226d9, 
               32'shc5736b90, 32'shc574b06b, 32'shc575f56b, 32'shc5773a8e, 32'shc5787fd6, 32'shc579c542, 32'shc57b0ad1, 32'shc57c5085, 
               32'shc57d965d, 32'shc57edc5a, 32'shc580227a, 32'shc58168be, 32'shc582af26, 32'shc583f5b3, 32'shc5853c63, 32'shc5868338, 
               32'shc587ca31, 32'shc589114e, 32'shc58a588e, 32'shc58b9ff3, 32'shc58ce77c, 32'shc58e2f29, 32'shc58f76fa, 32'shc590beef, 
               32'shc5920708, 32'shc5934f46, 32'shc59497a7, 32'shc595e02c, 32'shc59728d5, 32'shc59871a3, 32'shc599ba94, 32'shc59b03a9, 
               32'shc59c4ce3, 32'shc59d9640, 32'shc59edfc2, 32'shc5a02967, 32'shc5a17330, 32'shc5a2bd1e, 32'shc5a4072f, 32'shc5a55165, 
               32'shc5a69bbe, 32'shc5a7e63c, 32'shc5a930dd, 32'shc5aa7ba3, 32'shc5abc68c, 32'shc5ad1199, 32'shc5ae5ccb, 32'shc5afa820, 
               32'shc5b0f399, 32'shc5b23f37, 32'shc5b38af8, 32'shc5b4d6dd, 32'shc5b622e6, 32'shc5b76f13, 32'shc5b8bb64, 32'shc5ba07d9, 
               32'shc5bb5472, 32'shc5bca12f, 32'shc5bdee10, 32'shc5bf3b15, 32'shc5c0883d, 32'shc5c1d58a, 32'shc5c322fb, 32'shc5c4708f, 
               32'shc5c5be47, 32'shc5c70c24, 32'shc5c85a24, 32'shc5c9a848, 32'shc5caf690, 32'shc5cc44fc, 32'shc5cd938c, 32'shc5cee240, 
               32'shc5d03118, 32'shc5d18013, 32'shc5d2cf33, 32'shc5d41e76, 32'shc5d56ddd, 32'shc5d6bd68, 32'shc5d80d17, 32'shc5d95cea, 
               32'shc5daace1, 32'shc5dbfcfb, 32'shc5dd4d3a, 32'shc5de9d9c, 32'shc5dfee22, 32'shc5e13ecc, 32'shc5e28f9a, 32'shc5e3e08c, 
               32'shc5e531a1, 32'shc5e682db, 32'shc5e7d438, 32'shc5e925b9, 32'shc5ea775e, 32'shc5ebc927, 32'shc5ed1b13, 32'shc5ee6d24, 
               32'shc5efbf58, 32'shc5f111b0, 32'shc5f2642c, 32'shc5f3b6cb, 32'shc5f5098f, 32'shc5f65c76, 32'shc5f7af81, 32'shc5f902b0, 
               32'shc5fa5603, 32'shc5fba979, 32'shc5fcfd13, 32'shc5fe50d1, 32'shc5ffa4b3, 32'shc600f8b9, 32'shc6024ce2, 32'shc603a12f, 
               32'shc604f5a0, 32'shc6064a35, 32'shc6079eed, 32'shc608f3c9, 32'shc60a48c9, 32'shc60b9ded, 32'shc60cf334, 32'shc60e489f, 
               32'shc60f9e2e, 32'shc610f3e1, 32'shc61249b7, 32'shc6139fb2, 32'shc614f5cf, 32'shc6164c11, 32'shc617a276, 32'shc618f8ff, 
               32'shc61a4fac, 32'shc61ba67d, 32'shc61cfd71, 32'shc61e5489, 32'shc61fabc4, 32'shc6210323, 32'shc6225aa6, 32'shc623b24d, 
               32'shc6250a18, 32'shc6266206, 32'shc627ba17, 32'shc629124d, 32'shc62a6aa6, 32'shc62bc323, 32'shc62d1bc3, 32'shc62e7487, 
               32'shc62fcd6f, 32'shc631267a, 32'shc6327faa, 32'shc633d8fc, 32'shc6353273, 32'shc6368c0d, 32'shc637e5ca, 32'shc6393fac, 
               32'shc63a99b1, 32'shc63bf3d9, 32'shc63d4e26, 32'shc63ea896, 32'shc6400329, 32'shc6415de0, 32'shc642b8bb, 32'shc64413b9, 
               32'shc6456edb, 32'shc646ca21, 32'shc648258a, 32'shc6498117, 32'shc64adcc7, 32'shc64c389b, 32'shc64d9493, 32'shc64ef0ae, 
               32'shc6504ced, 32'shc651a94f, 32'shc65305d5, 32'shc654627f, 32'shc655bf4c, 32'shc6571c3c, 32'shc6587951, 32'shc659d688, 
               32'shc65b33e4, 32'shc65c9163, 32'shc65def05, 32'shc65f4ccb, 32'shc660aab5, 32'shc66208c2, 32'shc66366f3, 32'shc664c547, 
               32'shc66623be, 32'shc667825a, 32'shc668e119, 32'shc66a3ffb, 32'shc66b9f01, 32'shc66cfe2a, 32'shc66e5d77, 32'shc66fbce7, 
               32'shc6711c7b, 32'shc6727c32, 32'shc673dc0d, 32'shc6753c0c, 32'shc6769c2e, 32'shc677fc73, 32'shc6795cdc, 32'shc67abd68, 
               32'shc67c1e18, 32'shc67d7eeb, 32'shc67edfe2, 32'shc68040fc, 32'shc681a23a, 32'shc683039b, 32'shc6846520, 32'shc685c6c8, 
               32'shc6872894, 32'shc6888a83, 32'shc689ec95, 32'shc68b4ecb, 32'shc68cb124, 32'shc68e13a1, 32'shc68f7641, 32'shc690d905, 
               32'shc6923bec, 32'shc6939ef6, 32'shc6950224, 32'shc6966576, 32'shc697c8eb, 32'shc6992c83, 32'shc69a903e, 32'shc69bf41d, 
               32'shc69d5820, 32'shc69ebc45, 32'shc6a0208f, 32'shc6a184fb, 32'shc6a2e98b, 32'shc6a44e3e, 32'shc6a5b315, 32'shc6a7180f, 
               32'shc6a87d2d, 32'shc6a9e26e, 32'shc6ab47d2, 32'shc6acad59, 32'shc6ae1304, 32'shc6af78d3, 32'shc6b0dec4, 32'shc6b244d9, 
               32'shc6b3ab12, 32'shc6b5116d, 32'shc6b677ec, 32'shc6b7de8f, 32'shc6b94554, 32'shc6baac3d, 32'shc6bc134a, 32'shc6bd7a7a, 
               32'shc6bee1cd, 32'shc6c04943, 32'shc6c1b0dd, 32'shc6c31899, 32'shc6c4807a, 32'shc6c5e87d, 32'shc6c750a4, 32'shc6c8b8ee, 
               32'shc6ca215c, 32'shc6cb89ed, 32'shc6ccf2a1, 32'shc6ce5b78, 32'shc6cfc472, 32'shc6d12d90, 32'shc6d296d1, 32'shc6d40036, 
               32'shc6d569be, 32'shc6d6d369, 32'shc6d83d37, 32'shc6d9a728, 32'shc6db113d, 32'shc6dc7b75, 32'shc6dde5d0, 32'shc6df504f, 
               32'shc6e0baf0, 32'shc6e225b5, 32'shc6e3909d, 32'shc6e4fba9, 32'shc6e666d7, 32'shc6e7d229, 32'shc6e93d9e, 32'shc6eaa936, 
               32'shc6ec14f2, 32'shc6ed80d1, 32'shc6eeecd3, 32'shc6f058f8, 32'shc6f1c540, 32'shc6f331ab, 32'shc6f49e3a, 32'shc6f60aec, 
               32'shc6f777c1, 32'shc6f8e4b9, 32'shc6fa51d5, 32'shc6fbbf13, 32'shc6fd2c75, 32'shc6fe99fa, 32'shc70007a2, 32'shc701756d, 
               32'shc702e35c, 32'shc704516d, 32'shc705bfa2, 32'shc7072dfa, 32'shc7089c75, 32'shc70a0b13, 32'shc70b79d4, 32'shc70ce8b9, 
               32'shc70e57c0, 32'shc70fc6eb, 32'shc7113639, 32'shc712a5aa, 32'shc714153e, 32'shc71584f5, 32'shc716f4cf, 32'shc71864cc, 
               32'shc719d4ed, 32'shc71b4530, 32'shc71cb597, 32'shc71e2621, 32'shc71f96ce, 32'shc721079d, 32'shc7227890, 32'shc723e9a6, 
               32'shc7255ae0, 32'shc726cc3c, 32'shc7283dbb, 32'shc729af5d, 32'shc72b2123, 32'shc72c930b, 32'shc72e0517, 32'shc72f7745, 
               32'shc730e997, 32'shc7325c0c, 32'shc733cea3, 32'shc735415e, 32'shc736b43c, 32'shc738273d, 32'shc7399a60, 32'shc73b0da7, 
               32'shc73c8111, 32'shc73df49e, 32'shc73f684e, 32'shc740dc21, 32'shc7425016, 32'shc743c42f, 32'shc745386b, 32'shc746acca, 
               32'shc748214c, 32'shc74995f1, 32'shc74b0ab9, 32'shc74c7fa4, 32'shc74df4b1, 32'shc74f69e2, 32'shc750df36, 32'shc75254ac, 
               32'shc753ca46, 32'shc7554003, 32'shc756b5e2, 32'shc7582be5, 32'shc759a20a, 32'shc75b1853, 32'shc75c8ebe, 32'shc75e054c, 
               32'shc75f7bfe, 32'shc760f2d2, 32'shc76269c9, 32'shc763e0e3, 32'shc7655820, 32'shc766cf80, 32'shc7684702, 32'shc769bea8, 
               32'shc76b3671, 32'shc76cae5c, 32'shc76e266b, 32'shc76f9e9c, 32'shc77116f0, 32'shc7728f67, 32'shc7740801, 32'shc77580be, 
               32'shc776f99d, 32'shc77872a0, 32'shc779ebc5, 32'shc77b650e, 32'shc77cde79, 32'shc77e5807, 32'shc77fd1b8, 32'shc7814b8c, 
               32'shc782c582, 32'shc7843f9c, 32'shc785b9d8, 32'shc7873437, 32'shc788aeb9, 32'shc78a295e, 32'shc78ba425, 32'shc78d1f10, 
               32'shc78e9a1d, 32'shc790154d, 32'shc79190a0, 32'shc7930c16, 32'shc79487ae, 32'shc7960369, 32'shc7977f48, 32'shc798fb48, 
               32'shc79a776c, 32'shc79bf3b3, 32'shc79d701c, 32'shc79eeca8, 32'shc7a06957, 32'shc7a1e628, 32'shc7a3631d, 32'shc7a4e034, 
               32'shc7a65d6e, 32'shc7a7daca, 32'shc7a9584a, 32'shc7aad5ec, 32'shc7ac53b1, 32'shc7add198, 32'shc7af4fa3, 32'shc7b0cdd0, 
               32'shc7b24c20, 32'shc7b3ca92, 32'shc7b54928, 32'shc7b6c7e0, 32'shc7b846ba, 32'shc7b9c5b8, 32'shc7bb44d8, 32'shc7bcc41b, 
               32'shc7be4381, 32'shc7bfc309, 32'shc7c142b4, 32'shc7c2c282, 32'shc7c44272, 32'shc7c5c285, 32'shc7c742bb, 32'shc7c8c313, 
               32'shc7ca438f, 32'shc7cbc42c, 32'shc7cd44ed, 32'shc7cec5d0, 32'shc7d046d6, 32'shc7d1c7fe, 32'shc7d34949, 32'shc7d4cab7, 
               32'shc7d64c47, 32'shc7d7cdfb, 32'shc7d94fd0, 32'shc7dad1c9, 32'shc7dc53e3, 32'shc7ddd621, 32'shc7df5881, 32'shc7e0db04, 
               32'shc7e25daa, 32'shc7e3e072, 32'shc7e5635c, 32'shc7e6e66a, 32'shc7e8699a, 32'shc7e9ecec, 32'shc7eb7061, 32'shc7ecf3f9, 
               32'shc7ee77b3, 32'shc7effb90, 32'shc7f17f8f, 32'shc7f303b1, 32'shc7f487f6, 32'shc7f60c5d, 32'shc7f790e7, 32'shc7f91593, 
               32'shc7fa9a62, 32'shc7fc1f54, 32'shc7fda468, 32'shc7ff299e, 32'shc800aef7, 32'shc8023473, 32'shc803ba11, 32'shc8053fd2, 
               32'shc806c5b5, 32'shc8084bba, 32'shc809d1e3, 32'shc80b582e, 32'shc80cde9b, 32'shc80e652b, 32'shc80febdd, 32'shc81172b2, 
               32'shc812f9a9, 32'shc81480c3, 32'shc81607ff, 32'shc8178f5e, 32'shc81916df, 32'shc81a9e83, 32'shc81c2649, 32'shc81dae32, 
               32'shc81f363d, 32'shc820be6b, 32'shc82246bb, 32'shc823cf2e, 32'shc82557c3, 32'shc826e07a, 32'shc8286954, 32'shc829f251, 
               32'shc82b7b70, 32'shc82d04b1, 32'shc82e8e15, 32'shc830179b, 32'shc831a143, 32'shc8332b0e, 32'shc834b4fc, 32'shc8363f0c, 
               32'shc837c93e, 32'shc8395393, 32'shc83ade0a, 32'shc83c68a3, 32'shc83df35f, 32'shc83f7e3d, 32'shc841093e, 32'shc8429461, 
               32'shc8441fa6, 32'shc845ab0e, 32'shc8473698, 32'shc848c245, 32'shc84a4e14, 32'shc84bda05, 32'shc84d6619, 32'shc84ef24f, 
               32'shc8507ea7, 32'shc8520b22, 32'shc85397bf, 32'shc855247e, 32'shc856b160, 32'shc8583e64, 32'shc859cb8a, 32'shc85b58d3, 
               32'shc85ce63e, 32'shc85e73cc, 32'shc860017b, 32'shc8618f4d, 32'shc8631d42, 32'shc864ab58, 32'shc8663991, 32'shc867c7ec, 
               32'shc869566a, 32'shc86ae50a, 32'shc86c73cc, 32'shc86e02b0, 32'shc86f91b7, 32'shc87120e0, 32'shc872b02b, 32'shc8743f98, 
               32'shc875cf28, 32'shc8775eda, 32'shc878eeae, 32'shc87a7ea5, 32'shc87c0ebd, 32'shc87d9ef8, 32'shc87f2f56, 32'shc880bfd5, 
               32'shc8825077, 32'shc883e13b, 32'shc8857221, 32'shc8870329, 32'shc8889454, 32'shc88a25a1, 32'shc88bb710, 32'shc88d48a1, 
               32'shc88eda54, 32'shc8906c2a, 32'shc891fe22, 32'shc893903c, 32'shc8952278, 32'shc896b4d6, 32'shc8984757, 32'shc899d9fa, 
               32'shc89b6cbf, 32'shc89cffa6, 32'shc89e92af, 32'shc8a025da, 32'shc8a1b928, 32'shc8a34c98, 32'shc8a4e029, 32'shc8a673dd, 
               32'shc8a807b4, 32'shc8a99bac, 32'shc8ab2fc6, 32'shc8acc403, 32'shc8ae5862, 32'shc8afece2, 32'shc8b18185, 32'shc8b3164a, 
               32'shc8b4ab32, 32'shc8b6403b, 32'shc8b7d566, 32'shc8b96ab4, 32'shc8bb0023, 32'shc8bc95b5, 32'shc8be2b69, 32'shc8bfc13f, 
               32'shc8c15736, 32'shc8c2ed50, 32'shc8c4838d, 32'shc8c619eb, 32'shc8c7b06b, 32'shc8c9470d, 32'shc8caddd1, 32'shc8cc74b8, 
               32'shc8ce0bc0, 32'shc8cfa2eb, 32'shc8d13a37, 32'shc8d2d1a6, 32'shc8d46936, 32'shc8d600e9, 32'shc8d798be, 32'shc8d930b4, 
               32'shc8dac8cd, 32'shc8dc6108, 32'shc8ddf965, 32'shc8df91e3, 32'shc8e12a84, 32'shc8e2c347, 32'shc8e45c2c, 32'shc8e5f532, 
               32'shc8e78e5b, 32'shc8e927a6, 32'shc8eac112, 32'shc8ec5aa1, 32'shc8edf452, 32'shc8ef8e24, 32'shc8f12819, 32'shc8f2c230, 
               32'shc8f45c68, 32'shc8f5f6c3, 32'shc8f7913f, 32'shc8f92bdd, 32'shc8fac69e, 32'shc8fc6180, 32'shc8fdfc84, 32'shc8ff97aa, 
               32'shc90132f2, 32'shc902ce5c, 32'shc90469e8, 32'shc9060596, 32'shc907a166, 32'shc9093d57, 32'shc90ad96b, 32'shc90c75a0, 
               32'shc90e11f7, 32'shc90fae71, 32'shc9114b0c, 32'shc912e7c9, 32'shc91484a8, 32'shc91621a8, 32'shc917becb, 32'shc9195c0f, 
               32'shc91af976, 32'shc91c96fe, 32'shc91e34a8, 32'shc91fd274, 32'shc9217062, 32'shc9230e71, 32'shc924aca3, 32'shc9264af6, 
               32'shc927e96b, 32'shc9298802, 32'shc92b26bb, 32'shc92cc596, 32'shc92e6492, 32'shc93003b0, 32'shc931a2f0, 32'shc9334252, 
               32'shc934e1d6, 32'shc936817b, 32'shc9382143, 32'shc939c12c, 32'shc93b6137, 32'shc93d0163, 32'shc93ea1b2, 32'shc9404222, 
               32'shc941e2b4, 32'shc9438368, 32'shc945243d, 32'shc946c534, 32'shc948664d, 32'shc94a0788, 32'shc94ba8e5, 32'shc94d4a63, 
               32'shc94eec03, 32'shc9508dc5, 32'shc9522fa8, 32'shc953d1ad, 32'shc95573d4, 32'shc957161d, 32'shc958b887, 32'shc95a5b13, 
               32'shc95bfdc1, 32'shc95da090, 32'shc95f4382, 32'shc960e695, 32'shc96289c9, 32'shc9642d1f, 32'shc965d097, 32'shc9677431, 
               32'shc96917ec, 32'shc96abbc9, 32'shc96c5fc8, 32'shc96e03e8, 32'shc96fa82a, 32'shc9714c8e, 32'shc972f113, 32'shc97495ba, 
               32'shc9763a83, 32'shc977df6d, 32'shc9798479, 32'shc97b29a6, 32'shc97ccef5, 32'shc97e7466, 32'shc98019f8, 32'shc981bfac, 
               32'shc9836582, 32'shc9850b79, 32'shc986b192, 32'shc98857cd, 32'shc989fe29, 32'shc98ba4a6, 32'shc98d4b45, 32'shc98ef206, 
               32'shc99098e9, 32'shc9923fed, 32'shc993e712, 32'shc9958e59, 32'shc99735c2, 32'shc998dd4c, 32'shc99a84f8, 32'shc99c2cc5, 
               32'shc99dd4b4, 32'shc99f7cc5, 32'shc9a124f7, 32'shc9a2cd4a, 32'shc9a475bf, 32'shc9a61e56, 32'shc9a7c70e, 32'shc9a96fe7, 
               32'shc9ab18e3, 32'shc9acc1ff, 32'shc9ae6b3d, 32'shc9b0149d, 32'shc9b1be1e, 32'shc9b367c1, 32'shc9b51185, 32'shc9b6bb6b, 
               32'shc9b86572, 32'shc9ba0f9b, 32'shc9bbb9e5, 32'shc9bd6450, 32'shc9bf0edd, 32'shc9c0b98c, 32'shc9c2645c, 32'shc9c40f4d, 
               32'shc9c5ba60, 32'shc9c76595, 32'shc9c910ea, 32'shc9cabc62, 32'shc9cc67fa, 32'shc9ce13b4, 32'shc9cfbf90, 32'shc9d16b8d, 
               32'shc9d317ab, 32'shc9d4c3eb, 32'shc9d6704c, 32'shc9d81ccf, 32'shc9d9c973, 32'shc9db7639, 32'shc9dd231f, 32'shc9ded028, 
               32'shc9e07d51, 32'shc9e22a9c, 32'shc9e3d809, 32'shc9e58596, 32'shc9e73346, 32'shc9e8e116, 32'shc9ea8f08, 32'shc9ec3d1b, 
               32'shc9edeb50, 32'shc9ef99a6, 32'shc9f1481d, 32'shc9f2f6b6, 32'shc9f4a570, 32'shc9f6544b, 32'shc9f80348, 32'shc9f9b266, 
               32'shc9fb61a5, 32'shc9fd1106, 32'shc9fec088, 32'shca00702b, 32'shca021fef, 32'shca03cfd5, 32'shca057fdd, 32'shca073005, 
               32'shca08e04f, 32'shca0a90ba, 32'shca0c4146, 32'shca0df1f4, 32'shca0fa2c3, 32'shca1153b3, 32'shca1304c4, 32'shca14b5f7, 
               32'shca16674b, 32'shca1818c0, 32'shca19ca57, 32'shca1b7c0e, 32'shca1d2de7, 32'shca1edfe2, 32'shca2091fd, 32'shca22443a, 
               32'shca23f698, 32'shca25a917, 32'shca275bb7, 32'shca290e79, 32'shca2ac15b, 32'shca2c745f, 32'shca2e2784, 32'shca2fdacb, 
               32'shca318e32, 32'shca3341bb, 32'shca34f565, 32'shca36a930, 32'shca385d1d, 32'shca3a112a, 32'shca3bc559, 32'shca3d79a8, 
               32'shca3f2e19, 32'shca40e2ac, 32'shca42975f, 32'shca444c33, 32'shca460129, 32'shca47b640, 32'shca496b77, 32'shca4b20d0, 
               32'shca4cd64b, 32'shca4e8be6, 32'shca5041a2, 32'shca51f780, 32'shca53ad7e, 32'shca55639e, 32'shca5719df, 32'shca58d041, 
               32'shca5a86c4, 32'shca5c3d68, 32'shca5df42d, 32'shca5fab13, 32'shca61621b, 32'shca631943, 32'shca64d08d, 32'shca6687f7, 
               32'shca683f83, 32'shca69f72f, 32'shca6baefd, 32'shca6d66ec, 32'shca6f1efc, 32'shca70d72d, 32'shca728f7f, 32'shca7447f2, 
               32'shca760086, 32'shca77b93b, 32'shca797211, 32'shca7b2b08, 32'shca7ce420, 32'shca7e9d59, 32'shca8056b3, 32'shca82102e, 
               32'shca83c9ca, 32'shca858387, 32'shca873d65, 32'shca88f764, 32'shca8ab184, 32'shca8c6bc5, 32'shca8e2627, 32'shca8fe0aa, 
               32'shca919b4e, 32'shca935613, 32'shca9510f8, 32'shca96cbff, 32'shca988727, 32'shca9a4270, 32'shca9bfdd9, 32'shca9db964, 
               32'shca9f750f, 32'shcaa130db, 32'shcaa2ecc9, 32'shcaa4a8d7, 32'shcaa66506, 32'shcaa82156, 32'shcaa9ddc7, 32'shcaab9a59, 
               32'shcaad570c, 32'shcaaf13df, 32'shcab0d0d4, 32'shcab28de9, 32'shcab44b1f, 32'shcab60877, 32'shcab7c5ef, 32'shcab98388, 
               32'shcabb4141, 32'shcabcff1c, 32'shcabebd17, 32'shcac07b34, 32'shcac23971, 32'shcac3f7cf, 32'shcac5b64e, 32'shcac774ed, 
               32'shcac933ae, 32'shcacaf28f, 32'shcaccb191, 32'shcace70b4, 32'shcad02ff8, 32'shcad1ef5d, 32'shcad3aee2, 32'shcad56e88, 
               32'shcad72e4f, 32'shcad8ee37, 32'shcadaae40, 32'shcadc6e69, 32'shcade2eb3, 32'shcadfef1e, 32'shcae1afaa, 32'shcae37056, 
               32'shcae53123, 32'shcae6f211, 32'shcae8b320, 32'shcaea744f, 32'shcaec35a0, 32'shcaedf711, 32'shcaefb8a2, 32'shcaf17a55, 
               32'shcaf33c28, 32'shcaf4fe1c, 32'shcaf6c030, 32'shcaf88266, 32'shcafa44bc, 32'shcafc0732, 32'shcafdc9ca, 32'shcaff8c82, 
               32'shcb014f5b, 32'shcb031254, 32'shcb04d56e, 32'shcb0698a9, 32'shcb085c05, 32'shcb0a1f81, 32'shcb0be31e, 32'shcb0da6dc, 
               32'shcb0f6aba, 32'shcb112eb9, 32'shcb12f2d8, 32'shcb14b718, 32'shcb167b79, 32'shcb183ffb, 32'shcb1a049d, 32'shcb1bc95f, 
               32'shcb1d8e43, 32'shcb1f5347, 32'shcb21186b, 32'shcb22ddb1, 32'shcb24a316, 32'shcb26689d, 32'shcb282e44, 32'shcb29f40b, 
               32'shcb2bb9f4, 32'shcb2d7ffc, 32'shcb2f4626, 32'shcb310c70, 32'shcb32d2da, 32'shcb349965, 32'shcb366011, 32'shcb3826dd, 
               32'shcb39edca, 32'shcb3bb4d7, 32'shcb3d7c05, 32'shcb3f4354, 32'shcb410ac3, 32'shcb42d252, 32'shcb449a02, 32'shcb4661d3, 
               32'shcb4829c4, 32'shcb49f1d5, 32'shcb4bba08, 32'shcb4d825a, 32'shcb4f4acd, 32'shcb511361, 32'shcb52dc15, 32'shcb54a4ea, 
               32'shcb566ddf, 32'shcb5836f4, 32'shcb5a002b, 32'shcb5bc981, 32'shcb5d92f8, 32'shcb5f5c90, 32'shcb612648, 32'shcb62f020, 
               32'shcb64ba19, 32'shcb668432, 32'shcb684e6c, 32'shcb6a18c6, 32'shcb6be341, 32'shcb6daddc, 32'shcb6f7898, 32'shcb714373, 
               32'shcb730e70, 32'shcb74d98d, 32'shcb76a4ca, 32'shcb787027, 32'shcb7a3ba5, 32'shcb7c0744, 32'shcb7dd303, 32'shcb7f9ee2, 
               32'shcb816ae1, 32'shcb833701, 32'shcb850342, 32'shcb86cfa2, 32'shcb889c23, 32'shcb8a68c5, 32'shcb8c3587, 32'shcb8e0269, 
               32'shcb8fcf6b, 32'shcb919c8e, 32'shcb9369d1, 32'shcb953735, 32'shcb9704b9, 32'shcb98d25d, 32'shcb9aa021, 32'shcb9c6e06, 
               32'shcb9e3c0b, 32'shcba00a31, 32'shcba1d877, 32'shcba3a6dd, 32'shcba57563, 32'shcba7440a, 32'shcba912d1, 32'shcbaae1b8, 
               32'shcbacb0bf, 32'shcbae7fe7, 32'shcbb04f2f, 32'shcbb21e98, 32'shcbb3ee20, 32'shcbb5bdc9, 32'shcbb78d92, 32'shcbb95d7c, 
               32'shcbbb2d85, 32'shcbbcfdaf, 32'shcbbecdf9, 32'shcbc09e64, 32'shcbc26eee, 32'shcbc43f99, 32'shcbc61064, 32'shcbc7e14f, 
               32'shcbc9b25a, 32'shcbcb8386, 32'shcbcd54d2, 32'shcbcf263e, 32'shcbd0f7ca, 32'shcbd2c977, 32'shcbd49b43, 32'shcbd66d30, 
               32'shcbd83f3d, 32'shcbda116a, 32'shcbdbe3b7, 32'shcbddb625, 32'shcbdf88b3, 32'shcbe15b60, 32'shcbe32e2e, 32'shcbe5011c, 
               32'shcbe6d42b, 32'shcbe8a759, 32'shcbea7aa7, 32'shcbec4e16, 32'shcbee21a5, 32'shcbeff554, 32'shcbf1c923, 32'shcbf39d12, 
               32'shcbf57121, 32'shcbf74550, 32'shcbf919a0, 32'shcbfaee0f, 32'shcbfcc29f, 32'shcbfe974e, 32'shcc006c1e, 32'shcc02410e, 
               32'shcc04161e, 32'shcc05eb4e, 32'shcc07c09e, 32'shcc09960e, 32'shcc0b6b9e, 32'shcc0d414e, 32'shcc0f171e, 32'shcc10ed0e, 
               32'shcc12c31f, 32'shcc14994f, 32'shcc166f9f, 32'shcc184610, 32'shcc1a1ca0, 32'shcc1bf350, 32'shcc1dca21, 32'shcc1fa111, 
               32'shcc217822, 32'shcc234f52, 32'shcc2526a2, 32'shcc26fe13, 32'shcc28d5a3, 32'shcc2aad54, 32'shcc2c8524, 32'shcc2e5d14, 
               32'shcc303524, 32'shcc320d55, 32'shcc33e5a5, 32'shcc35be15, 32'shcc3796a5, 32'shcc396f55, 32'shcc3b4825, 32'shcc3d2115, 
               32'shcc3efa25, 32'shcc40d354, 32'shcc42aca4, 32'shcc448614, 32'shcc465fa3, 32'shcc483952, 32'shcc4a1322, 32'shcc4bed11, 
               32'shcc4dc720, 32'shcc4fa14f, 32'shcc517b9e, 32'shcc53560c, 32'shcc55309b, 32'shcc570b4a, 32'shcc58e618, 32'shcc5ac106, 
               32'shcc5c9c14, 32'shcc5e7742, 32'shcc605290, 32'shcc622dfd, 32'shcc64098b, 32'shcc65e538, 32'shcc67c105, 32'shcc699cf2, 
               32'shcc6b78ff, 32'shcc6d552c, 32'shcc6f3178, 32'shcc710de4, 32'shcc72ea70, 32'shcc74c71c, 32'shcc76a3e8, 32'shcc7880d3, 
               32'shcc7a5dde, 32'shcc7c3b09, 32'shcc7e1854, 32'shcc7ff5be, 32'shcc81d349, 32'shcc83b0f3, 32'shcc858ebc, 32'shcc876ca6, 
               32'shcc894aaf, 32'shcc8b28d8, 32'shcc8d0721, 32'shcc8ee58a, 32'shcc90c412, 32'shcc92a2ba, 32'shcc948182, 32'shcc966069, 
               32'shcc983f70, 32'shcc9a1e97, 32'shcc9bfddd, 32'shcc9ddd44, 32'shcc9fbcca, 32'shcca19c6f, 32'shcca37c35, 32'shcca55c1a, 
               32'shcca73c1e, 32'shcca91c43, 32'shccaafc87, 32'shccacdcea, 32'shccaebd6e, 32'shccb09e11, 32'shccb27ed3, 32'shccb45fb6, 
               32'shccb640b8, 32'shccb821d9, 32'shccba031a, 32'shccbbe47b, 32'shccbdc5fc, 32'shccbfa79c, 32'shccc1895c, 32'shccc36b3b, 
               32'shccc54d3a, 32'shccc72f58, 32'shccc91196, 32'shcccaf3f4, 32'shccccd671, 32'shccceb90e, 32'shccd09bcb, 32'shccd27ea7, 
               32'shccd461a2, 32'shccd644bd, 32'shccd827f8, 32'shccda0b52, 32'shccdbeecc, 32'shccddd266, 32'shccdfb61f, 32'shcce199f7, 
               32'shcce37def, 32'shcce56206, 32'shcce7463e, 32'shcce92a94, 32'shcceb0f0a, 32'shccecf3a0, 32'shcceed855, 32'shccf0bd29, 
               32'shccf2a21d, 32'shccf48731, 32'shccf66c64, 32'shccf851b7, 32'shccfa3729, 32'shccfc1cba, 32'shccfe026b, 32'shccffe83c, 
               32'shcd01ce2b, 32'shcd03b43b, 32'shcd059a6a, 32'shcd0780b8, 32'shcd096725, 32'shcd0b4db3, 32'shcd0d345f, 32'shcd0f1b2b, 
               32'shcd110216, 32'shcd12e921, 32'shcd14d04b, 32'shcd16b795, 32'shcd189efe, 32'shcd1a8687, 32'shcd1c6e2e, 32'shcd1e55f6, 
               32'shcd203ddc, 32'shcd2225e2, 32'shcd240e08, 32'shcd25f64c, 32'shcd27deb0, 32'shcd29c734, 32'shcd2bafd7, 32'shcd2d9899, 
               32'shcd2f817b, 32'shcd316a7b, 32'shcd33539c, 32'shcd353cdb, 32'shcd37263a, 32'shcd390fb8, 32'shcd3af956, 32'shcd3ce313, 
               32'shcd3eccef, 32'shcd40b6ea, 32'shcd42a105, 32'shcd448b3f, 32'shcd467599, 32'shcd486011, 32'shcd4a4aa9, 32'shcd4c3560, 
               32'shcd4e2037, 32'shcd500b2d, 32'shcd51f642, 32'shcd53e176, 32'shcd55ccca, 32'shcd57b83c, 32'shcd59a3ce, 32'shcd5b8f80, 
               32'shcd5d7b50, 32'shcd5f6740, 32'shcd61534f, 32'shcd633f7d, 32'shcd652bcb, 32'shcd671837, 32'shcd6904c3, 32'shcd6af16e, 
               32'shcd6cde39, 32'shcd6ecb22, 32'shcd70b82b, 32'shcd72a553, 32'shcd74929a, 32'shcd768000, 32'shcd786d85, 32'shcd7a5b2a, 
               32'shcd7c48ee, 32'shcd7e36d1, 32'shcd8024d3, 32'shcd8212f4, 32'shcd840134, 32'shcd85ef94, 32'shcd87de12, 32'shcd89ccb0, 
               32'shcd8bbb6d, 32'shcd8daa49, 32'shcd8f9944, 32'shcd91885e, 32'shcd937798, 32'shcd9566f0, 32'shcd975668, 32'shcd9945fe, 
               32'shcd9b35b4, 32'shcd9d2589, 32'shcd9f157d, 32'shcda10590, 32'shcda2f5c2, 32'shcda4e613, 32'shcda6d683, 32'shcda8c712, 
               32'shcdaab7c0, 32'shcdaca88e, 32'shcdae997a, 32'shcdb08a86, 32'shcdb27bb0, 32'shcdb46cfa, 32'shcdb65e62, 32'shcdb84fea, 
               32'shcdba4190, 32'shcdbc3356, 32'shcdbe253a, 32'shcdc0173e, 32'shcdc20960, 32'shcdc3fba2, 32'shcdc5ee02, 32'shcdc7e082, 
               32'shcdc9d320, 32'shcdcbc5de, 32'shcdcdb8ba, 32'shcdcfabb6, 32'shcdd19ed0, 32'shcdd39209, 32'shcdd58562, 32'shcdd778d9, 
               32'shcdd96c6f, 32'shcddb6024, 32'shcddd53f8, 32'shcddf47eb, 32'shcde13bfd, 32'shcde3302e, 32'shcde5247d, 32'shcde718ec, 
               32'shcde90d79, 32'shcdeb0226, 32'shcdecf6f1, 32'shcdeeebdb, 32'shcdf0e0e4, 32'shcdf2d60c, 32'shcdf4cb53, 32'shcdf6c0b9, 
               32'shcdf8b63d, 32'shcdfaabe1, 32'shcdfca1a3, 32'shcdfe9784, 32'shce008d84, 32'shce0283a3, 32'shce0479e0, 32'shce06703d, 
               32'shce0866b8, 32'shce0a5d52, 32'shce0c540b, 32'shce0e4ae3, 32'shce1041d9, 32'shce1238ef, 32'shce143023, 32'shce162776, 
               32'shce181ee8, 32'shce1a1678, 32'shce1c0e28, 32'shce1e05f6, 32'shce1ffde2, 32'shce21f5ee, 32'shce23ee18, 32'shce25e662, 
               32'shce27dec9, 32'shce29d750, 32'shce2bcff5, 32'shce2dc8ba, 32'shce2fc19c, 32'shce31ba9e, 32'shce33b3be, 32'shce35acfd, 
               32'shce37a65b, 32'shce399fd7, 32'shce3b9973, 32'shce3d932c, 32'shce3f8d05, 32'shce4186fc, 32'shce438112, 32'shce457b47, 
               32'shce47759a, 32'shce49700c, 32'shce4b6a9c, 32'shce4d654c, 32'shce4f6019, 32'shce515b06, 32'shce535611, 32'shce55513b, 
               32'shce574c84, 32'shce5947eb, 32'shce5b4370, 32'shce5d3f15, 32'shce5f3ad8, 32'shce6136b9, 32'shce6332ba, 32'shce652ed8, 
               32'shce672b16, 32'shce692772, 32'shce6b23ec, 32'shce6d2086, 32'shce6f1d3d, 32'shce711a14, 32'shce731709, 32'shce75141c, 
               32'shce77114e, 32'shce790e9f, 32'shce7b0c0e, 32'shce7d099b, 32'shce7f0748, 32'shce810512, 32'shce8302fc, 32'shce850104, 
               32'shce86ff2a, 32'shce88fd6f, 32'shce8afbd2, 32'shce8cfa54, 32'shce8ef8f4, 32'shce90f7b3, 32'shce92f691, 32'shce94f58c, 
               32'shce96f4a7, 32'shce98f3e0, 32'shce9af337, 32'shce9cf2ad, 32'shce9ef241, 32'shcea0f1f4, 32'shcea2f1c5, 32'shcea4f1b4, 
               32'shcea6f1c2, 32'shcea8f1ef, 32'shceaaf23a, 32'shceacf2a3, 32'shceaef32b, 32'shceb0f3d1, 32'shceb2f496, 32'shceb4f579, 
               32'shceb6f67a, 32'shceb8f79a, 32'shcebaf8d8, 32'shcebcfa35, 32'shcebefbb0, 32'shcec0fd49, 32'shcec2ff01, 32'shcec500d7, 
               32'shcec702cb, 32'shcec904de, 32'shcecb070f, 32'shcecd095f, 32'shcecf0bcd, 32'shced10e59, 32'shced31104, 32'shced513cd, 
               32'shced716b4, 32'shced919ba, 32'shcedb1cde, 32'shcedd2020, 32'shcedf2380, 32'shcee126ff, 32'shcee32a9c, 32'shcee52e58, 
               32'shcee73231, 32'shcee93629, 32'shceeb3a40, 32'shceed3e74, 32'shceef42c7, 32'shcef14738, 32'shcef34bc8, 32'shcef55075, 
               32'shcef75541, 32'shcef95a2b, 32'shcefb5f34, 32'shcefd645a, 32'shceff699f, 32'shcf016f02, 32'shcf037483, 32'shcf057a23, 
               32'shcf077fe1, 32'shcf0985bc, 32'shcf0b8bb7, 32'shcf0d91cf, 32'shcf0f9805, 32'shcf119e5a, 32'shcf13a4cd, 32'shcf15ab5e, 
               32'shcf17b20d, 32'shcf19b8db, 32'shcf1bbfc6, 32'shcf1dc6d0, 32'shcf1fcdf8, 32'shcf21d53e, 32'shcf23dca2, 32'shcf25e424, 
               32'shcf27ebc5, 32'shcf29f383, 32'shcf2bfb60, 32'shcf2e035b, 32'shcf300b74, 32'shcf3213ab, 32'shcf341c00, 32'shcf362473, 
               32'shcf382d05, 32'shcf3a35b4, 32'shcf3c3e82, 32'shcf3e476d, 32'shcf405077, 32'shcf42599f, 32'shcf4462e4, 32'shcf466c48, 
               32'shcf4875ca, 32'shcf4a7f6a, 32'shcf4c8928, 32'shcf4e9304, 32'shcf509cfe, 32'shcf52a716, 32'shcf54b14d, 32'shcf56bba1, 
               32'shcf58c613, 32'shcf5ad0a3, 32'shcf5cdb51, 32'shcf5ee61e, 32'shcf60f108, 32'shcf62fc10, 32'shcf650736, 32'shcf67127a, 
               32'shcf691ddd, 32'shcf6b295d, 32'shcf6d34fb, 32'shcf6f40b7, 32'shcf714c91, 32'shcf735889, 32'shcf75649f, 32'shcf7770d3, 
               32'shcf797d24, 32'shcf7b8994, 32'shcf7d9622, 32'shcf7fa2cd, 32'shcf81af97, 32'shcf83bc7e, 32'shcf85c984, 32'shcf87d6a7, 
               32'shcf89e3e8, 32'shcf8bf147, 32'shcf8dfec4, 32'shcf900c5f, 32'shcf921a17, 32'shcf9427ee, 32'shcf9635e2, 32'shcf9843f5, 
               32'shcf9a5225, 32'shcf9c6073, 32'shcf9e6edf, 32'shcfa07d68, 32'shcfa28c10, 32'shcfa49ad5, 32'shcfa6a9b8, 32'shcfa8b8b9, 
               32'shcfaac7d8, 32'shcfacd715, 32'shcfaee66f, 32'shcfb0f5e7, 32'shcfb3057d, 32'shcfb51531, 32'shcfb72503, 32'shcfb934f2, 
               32'shcfbb4500, 32'shcfbd552b, 32'shcfbf6573, 32'shcfc175da, 32'shcfc3865e, 32'shcfc59700, 32'shcfc7a7c0, 32'shcfc9b89d, 
               32'shcfcbc999, 32'shcfcddab2, 32'shcfcfebe8, 32'shcfd1fd3d, 32'shcfd40eaf, 32'shcfd6203f, 32'shcfd831ec, 32'shcfda43b8, 
               32'shcfdc55a1, 32'shcfde67a7, 32'shcfe079cc, 32'shcfe28c0e, 32'shcfe49e6d, 32'shcfe6b0eb, 32'shcfe8c386, 32'shcfead63f, 
               32'shcfece915, 32'shcfeefc09, 32'shcff10f1b, 32'shcff3224a, 32'shcff53597, 32'shcff74902, 32'shcff95c8a, 32'shcffb7030, 
               32'shcffd83f4, 32'shcfff97d5, 32'shd001abd3, 32'shd003bff0, 32'shd005d42a, 32'shd007e881, 32'shd009fcf6, 32'shd00c1189, 
               32'shd00e2639, 32'shd0103b07, 32'shd0124ff3, 32'shd01464fc, 32'shd0167a22, 32'shd0188f66, 32'shd01aa4c8, 32'shd01cba47, 
               32'shd01ecfe4, 32'shd020e59e, 32'shd022fb76, 32'shd025116b, 32'shd027277e, 32'shd0293dae, 32'shd02b53fc, 32'shd02d6a68, 
               32'shd02f80f1, 32'shd0319797, 32'shd033ae5b, 32'shd035c53c, 32'shd037dc3b, 32'shd039f357, 32'shd03c0a91, 32'shd03e21e8, 
               32'shd040395d, 32'shd04250ef, 32'shd044689f, 32'shd046806c, 32'shd0489856, 32'shd04ab05e, 32'shd04cc884, 32'shd04ee0c6, 
               32'shd050f926, 32'shd05311a4, 32'shd0552a3f, 32'shd05742f7, 32'shd0595bcd, 32'shd05b74c0, 32'shd05d8dd1, 32'shd05fa6ff, 
               32'shd061c04a, 32'shd063d9b3, 32'shd065f339, 32'shd0680cdd, 32'shd06a269d, 32'shd06c407c, 32'shd06e5a77, 32'shd0707490, 
               32'shd0728ec6, 32'shd074a91a, 32'shd076c38b, 32'shd078de19, 32'shd07af8c4, 32'shd07d138d, 32'shd07f2e73, 32'shd0814977, 
               32'shd0836497, 32'shd0857fd5, 32'shd0879b31, 32'shd089b6a9, 32'shd08bd23f, 32'shd08dedf2, 32'shd09009c3, 32'shd09225b0, 
               32'shd09441bb, 32'shd0965de3, 32'shd0987a29, 32'shd09a968b, 32'shd09cb30b, 32'shd09ecfa8, 32'shd0a0ec63, 32'shd0a3093a, 
               32'shd0a5262f, 32'shd0a74341, 32'shd0a96070, 32'shd0ab7dbd, 32'shd0ad9b26, 32'shd0afb8ad, 32'shd0b1d651, 32'shd0b3f412, 
               32'shd0b611f1, 32'shd0b82fec, 32'shd0ba4e05, 32'shd0bc6c3a, 32'shd0be8a8d, 32'shd0c0a8fe, 32'shd0c2c78b, 32'shd0c4e635, 
               32'shd0c704fd, 32'shd0c923e1, 32'shd0cb42e3, 32'shd0cd6202, 32'shd0cf813e, 32'shd0d1a097, 32'shd0d3c00e, 32'shd0d5dfa1, 
               32'shd0d7ff51, 32'shd0da1f1f, 32'shd0dc3f0a, 32'shd0de5f11, 32'shd0e07f36, 32'shd0e29f78, 32'shd0e4bfd7, 32'shd0e6e053, 
               32'shd0e900ec, 32'shd0eb21a2, 32'shd0ed4275, 32'shd0ef6365, 32'shd0f18472, 32'shd0f3a59c, 32'shd0f5c6e3, 32'shd0f7e848, 
               32'shd0fa09c9, 32'shd0fc2b67, 32'shd0fe4d22, 32'shd1006efb, 32'shd10290f0, 32'shd104b302, 32'shd106d531, 32'shd108f77d, 
               32'shd10b19e7, 32'shd10d3c6d, 32'shd10f5f10, 32'shd11181d0, 32'shd113a4ad, 32'shd115c7a7, 32'shd117eabd, 32'shd11a0df1, 
               32'shd11c3142, 32'shd11e54b0, 32'shd120783a, 32'shd1229be2, 32'shd124bfa6, 32'shd126e387, 32'shd1290786, 32'shd12b2ba1, 
               32'shd12d4fd9, 32'shd12f742d, 32'shd131989f, 32'shd133bd2e, 32'shd135e1d9, 32'shd13806a2, 32'shd13a2b87, 32'shd13c5089, 
               32'shd13e75a8, 32'shd1409ae3, 32'shd142c03c, 32'shd144e5b1, 32'shd1470b44, 32'shd14930f3, 32'shd14b56be, 32'shd14d7ca7, 
               32'shd14fa2ad, 32'shd151c8cf, 32'shd153ef0e, 32'shd156156a, 32'shd1583be2, 32'shd15a6278, 32'shd15c892a, 32'shd15eaff9, 
               32'shd160d6e5, 32'shd162fded, 32'shd1652512, 32'shd1674c54, 32'shd16973b3, 32'shd16b9b2f, 32'shd16dc2c7, 32'shd16fea7c, 
               32'shd172124d, 32'shd1743a3c, 32'shd1766247, 32'shd1788a6f, 32'shd17ab2b3, 32'shd17cdb14, 32'shd17f0392, 32'shd1812c2d, 
               32'shd18354e4, 32'shd1857db8, 32'shd187a6a8, 32'shd189cfb6, 32'shd18bf8e0, 32'shd18e2226, 32'shd1904b89, 32'shd1927509, 
               32'shd1949ea6, 32'shd196c85f, 32'shd198f235, 32'shd19b1c27, 32'shd19d4636, 32'shd19f7062, 32'shd1a19aaa, 32'shd1a3c50f, 
               32'shd1a5ef90, 32'shd1a81a2e, 32'shd1aa44e9, 32'shd1ac6fc0, 32'shd1ae9ab4, 32'shd1b0c5c4, 32'shd1b2f0f1, 32'shd1b51c3a, 
               32'shd1b747a0, 32'shd1b97323, 32'shd1bb9ec2, 32'shd1bdca7e, 32'shd1bff656, 32'shd1c2224b, 32'shd1c44e5c, 32'shd1c67a8a, 
               32'shd1c8a6d4, 32'shd1cad33b, 32'shd1ccffbe, 32'shd1cf2c5e, 32'shd1d1591a, 32'shd1d385f3, 32'shd1d5b2e8, 32'shd1d7dffa, 
               32'shd1da0d28, 32'shd1dc3a73, 32'shd1de67da, 32'shd1e0955d, 32'shd1e2c2fd, 32'shd1e4f0ba, 32'shd1e71e93, 32'shd1e94c88, 
               32'shd1eb7a9a, 32'shd1eda8c8, 32'shd1efd713, 32'shd1f2057a, 32'shd1f433fd, 32'shd1f6629d, 32'shd1f89159, 32'shd1fac032, 
               32'shd1fcef27, 32'shd1ff1e38, 32'shd2014d66, 32'shd2037cb0, 32'shd205ac17, 32'shd207db9a, 32'shd20a0b39, 32'shd20c3af4, 
               32'shd20e6acc, 32'shd2109ac1, 32'shd212cad1, 32'shd214fafe, 32'shd2172b48, 32'shd2195bad, 32'shd21b8c2f, 32'shd21dbccd, 
               32'shd21fed88, 32'shd2221e5f, 32'shd2244f52, 32'shd2268061, 32'shd228b18d, 32'shd22ae2d5, 32'shd22d1439, 32'shd22f45b9, 
               32'shd2317756, 32'shd233a90f, 32'shd235dae4, 32'shd2380cd6, 32'shd23a3ee4, 32'shd23c710e, 32'shd23ea354, 32'shd240d5b6, 
               32'shd2430835, 32'shd2453ad0, 32'shd2476d87, 32'shd249a05a, 32'shd24bd34a, 32'shd24e0655, 32'shd250397d, 32'shd2526cc1, 
               32'shd254a021, 32'shd256d39e, 32'shd2590736, 32'shd25b3aeb, 32'shd25d6ebc, 32'shd25fa2a9, 32'shd261d6b2, 32'shd2640ad7, 
               32'shd2663f19, 32'shd2687376, 32'shd26aa7f0, 32'shd26cdc86, 32'shd26f1138, 32'shd2714606, 32'shd2737af0, 32'shd275aff6, 
               32'shd277e518, 32'shd27a1a57, 32'shd27c4fb1, 32'shd27e8528, 32'shd280babb, 32'shd282f069, 32'shd2852634, 32'shd2875c1b, 
               32'shd289921e, 32'shd28bc83d, 32'shd28dfe77, 32'shd29034ce, 32'shd2926b41, 32'shd294a1d0, 32'shd296d87c, 32'shd2990f43, 
               32'shd29b4626, 32'shd29d7d25, 32'shd29fb440, 32'shd2a1eb77, 32'shd2a422ca, 32'shd2a65a39, 32'shd2a891c4, 32'shd2aac96b, 
               32'shd2ad012e, 32'shd2af390d, 32'shd2b17107, 32'shd2b3a91e, 32'shd2b5e151, 32'shd2b8199f, 32'shd2ba520a, 32'shd2bc8a91, 
               32'shd2bec333, 32'shd2c0fbf1, 32'shd2c334cc, 32'shd2c56dc2, 32'shd2c7a6d4, 32'shd2c9e002, 32'shd2cc194c, 32'shd2ce52b1, 
               32'shd2d08c33, 32'shd2d2c5d0, 32'shd2d4ff8a, 32'shd2d7395f, 32'shd2d97350, 32'shd2dbad5d, 32'shd2dde786, 32'shd2e021ca, 
               32'shd2e25c2b, 32'shd2e496a7, 32'shd2e6d13f, 32'shd2e90bf3, 32'shd2eb46c3, 32'shd2ed81ae, 32'shd2efbcb6, 32'shd2f1f7d9, 
               32'shd2f43318, 32'shd2f66e72, 32'shd2f8a9e9, 32'shd2fae57b, 32'shd2fd2129, 32'shd2ff5cf3, 32'shd30198d8, 32'shd303d4da, 
               32'shd30610f7, 32'shd3084d30, 32'shd30a8984, 32'shd30cc5f4, 32'shd30f0280, 32'shd3113f28, 32'shd3137bec, 32'shd315b8cb, 
               32'shd317f5c6, 32'shd31a32dc, 32'shd31c700f, 32'shd31ead5c, 32'shd320eac6, 32'shd323284b, 32'shd32565ec, 32'shd327a3a9, 
               32'shd329e181, 32'shd32c1f75, 32'shd32e5d85, 32'shd3309bb0, 32'shd332d9f7, 32'shd335185a, 32'shd33756d8, 32'shd3399572, 
               32'shd33bd427, 32'shd33e12f8, 32'shd34051e5, 32'shd34290ed, 32'shd344d011, 32'shd3470f50, 32'shd3494eab, 32'shd34b8e22, 
               32'shd34dcdb4, 32'shd3500d62, 32'shd3524d2b, 32'shd3548d10, 32'shd356cd11, 32'shd3590d2c, 32'shd35b4d64, 32'shd35d8db7, 
               32'shd35fce26, 32'shd3620eb0, 32'shd3644f55, 32'shd3669017, 32'shd368d0f3, 32'shd36b11eb, 32'shd36d52ff, 32'shd36f942e, 
               32'shd371d579, 32'shd37416df, 32'shd3765861, 32'shd37899fe, 32'shd37adbb6, 32'shd37d1d8a, 32'shd37f5f7a, 32'shd381a185, 
               32'shd383e3ab, 32'shd38625ed, 32'shd388684a, 32'shd38aaac3, 32'shd38ced57, 32'shd38f3007, 32'shd39172d2, 32'shd393b5b8, 
               32'shd395f8ba, 32'shd3983bd7, 32'shd39a7f0f, 32'shd39cc263, 32'shd39f05d3, 32'shd3a1495d, 32'shd3a38d03, 32'shd3a5d0c5, 
               32'shd3a814a2, 32'shd3aa589a, 32'shd3ac9cad, 32'shd3aee0dc, 32'shd3b12526, 32'shd3b3698c, 32'shd3b5ae0d, 32'shd3b7f2a9, 
               32'shd3ba3760, 32'shd3bc7c33, 32'shd3bec121, 32'shd3c1062a, 32'shd3c34b4f, 32'shd3c5908f, 32'shd3c7d5ea, 32'shd3ca1b61, 
               32'shd3cc60f2, 32'shd3cea69f, 32'shd3d0ec68, 32'shd3d3324b, 32'shd3d5784a, 32'shd3d7be64, 32'shd3da049a, 32'shd3dc4aea, 
               32'shd3de9156, 32'shd3e0d7dd, 32'shd3e31e7f, 32'shd3e5653c, 32'shd3e7ac15, 32'shd3e9f309, 32'shd3ec3a18, 32'shd3ee8142, 
               32'shd3f0c887, 32'shd3f30fe8, 32'shd3f55764, 32'shd3f79efa, 32'shd3f9e6ad, 32'shd3fc2e7a, 32'shd3fe7662, 32'shd400be66, 
               32'shd4030684, 32'shd4054ebe, 32'shd4079713, 32'shd409df83, 32'shd40c280e, 32'shd40e70b4, 32'shd410b976, 32'shd4130252, 
               32'shd4154b4a, 32'shd417945c, 32'shd419dd8a, 32'shd41c26d3, 32'shd41e7037, 32'shd420b9b6, 32'shd4230350, 32'shd4254d05, 
               32'shd42796d5, 32'shd429e0c0, 32'shd42c2ac6, 32'shd42e74e8, 32'shd430bf24, 32'shd433097b, 32'shd43553ee, 32'shd4379e7b, 
               32'shd439e923, 32'shd43c33e7, 32'shd43e7ec5, 32'shd440c9be, 32'shd44314d3, 32'shd4456002, 32'shd447ab4c, 32'shd449f6b1, 
               32'shd44c4232, 32'shd44e8dcd, 32'shd450d983, 32'shd4532554, 32'shd4557140, 32'shd457bd47, 32'shd45a0969, 32'shd45c55a5, 
               32'shd45ea1fd, 32'shd460ee70, 32'shd4633afd, 32'shd46587a6, 32'shd467d469, 32'shd46a2147, 32'shd46c6e40, 32'shd46ebb54, 
               32'shd4710883, 32'shd47355cd, 32'shd475a332, 32'shd477f0b1, 32'shd47a3e4b, 32'shd47c8c00, 32'shd47ed9d0, 32'shd48127bb, 
               32'shd48375c1, 32'shd485c3e1, 32'shd488121d, 32'shd48a6073, 32'shd48caee4, 32'shd48efd6f, 32'shd4914c16, 32'shd4939ad7, 
               32'shd495e9b3, 32'shd49838aa, 32'shd49a87bc, 32'shd49cd6e8, 32'shd49f2630, 32'shd4a17591, 32'shd4a3c50e, 32'shd4a614a6, 
               32'shd4a86458, 32'shd4aab425, 32'shd4ad040c, 32'shd4af540f, 32'shd4b1a42c, 32'shd4b3f464, 32'shd4b644b6, 32'shd4b89523, 
               32'shd4bae5ab, 32'shd4bd364e, 32'shd4bf870b, 32'shd4c1d7e3, 32'shd4c428d6, 32'shd4c679e3, 32'shd4c8cb0b, 32'shd4cb1c4e, 
               32'shd4cd6dab, 32'shd4cfbf23, 32'shd4d210b5, 32'shd4d46263, 32'shd4d6b42b, 32'shd4d9060d, 32'shd4db580a, 32'shd4ddaa22, 
               32'shd4dffc54, 32'shd4e24ea1, 32'shd4e4a108, 32'shd4e6f38b, 32'shd4e94627, 32'shd4eb98de, 32'shd4edebb0, 32'shd4f03e9d, 
               32'shd4f291a4, 32'shd4f4e4c5, 32'shd4f73801, 32'shd4f98b58, 32'shd4fbdec9, 32'shd4fe3255, 32'shd50085fb, 32'shd502d9bc, 
               32'shd5052d97, 32'shd507818d, 32'shd509d59d, 32'shd50c29c8, 32'shd50e7e0d, 32'shd510d26d, 32'shd51326e7, 32'shd5157b7c, 
               32'shd517d02b, 32'shd51a24f5, 32'shd51c79d9, 32'shd51eced7, 32'shd52123f0, 32'shd5237924, 32'shd525ce72, 32'shd52823da, 
               32'shd52a795d, 32'shd52ccefa, 32'shd52f24b2, 32'shd5317a84, 32'shd533d070, 32'shd5362677, 32'shd5387c98, 32'shd53ad2d4, 
               32'shd53d292a, 32'shd53f7f9a, 32'shd541d625, 32'shd5442cca, 32'shd5468389, 32'shd548da63, 32'shd54b3157, 32'shd54d8866, 
               32'shd54fdf8f, 32'shd55236d2, 32'shd5548e30, 32'shd556e5a7, 32'shd5593d3a, 32'shd55b94e6, 32'shd55decad, 32'shd560448e, 
               32'shd5629c89, 32'shd564f49f, 32'shd5674ccf, 32'shd569a519, 32'shd56bfd7d, 32'shd56e55fc, 32'shd570ae95, 32'shd5730748, 
               32'shd5756016, 32'shd577b8fe, 32'shd57a1200, 32'shd57c6b1c, 32'shd57ec452, 32'shd5811da3, 32'shd583770e, 32'shd585d093, 
               32'shd5882a32, 32'shd58a83eb, 32'shd58cddbf, 32'shd58f37ad, 32'shd59191b5, 32'shd593ebd7, 32'shd5964614, 32'shd598a06a, 
               32'shd59afadb, 32'shd59d5566, 32'shd59fb00b, 32'shd5a20aca, 32'shd5a465a3, 32'shd5a6c096, 32'shd5a91ba4, 32'shd5ab76cb, 
               32'shd5add20d, 32'shd5b02d69, 32'shd5b288df, 32'shd5b4e46f, 32'shd5b74019, 32'shd5b99bdd, 32'shd5bbf7bc, 32'shd5be53b4, 
               32'shd5c0afc6, 32'shd5c30bf3, 32'shd5c56839, 32'shd5c7c49a, 32'shd5ca2115, 32'shd5cc7da9, 32'shd5ceda58, 32'shd5d13721, 
               32'shd5d39403, 32'shd5d5f100, 32'shd5d84e17, 32'shd5daab48, 32'shd5dd0892, 32'shd5df65f7, 32'shd5e1c376, 32'shd5e4210f, 
               32'shd5e67ec1, 32'shd5e8dc8e, 32'shd5eb3a75, 32'shd5ed9875, 32'shd5eff690, 32'shd5f254c4, 32'shd5f4b313, 32'shd5f7117b, 
               32'shd5f96ffd, 32'shd5fbce9a, 32'shd5fe2d50, 32'shd6008c20, 32'shd602eb0a, 32'shd6054a0d, 32'shd607a92b, 32'shd60a0863, 
               32'shd60c67b4, 32'shd60ec720, 32'shd61126a5, 32'shd6138644, 32'shd615e5fd, 32'shd61845d0, 32'shd61aa5bd, 32'shd61d05c3, 
               32'shd61f65e4, 32'shd621c61e, 32'shd6242672, 32'shd62686e0, 32'shd628e767, 32'shd62b4809, 32'shd62da8c4, 32'shd6300999, 
               32'shd6326a88, 32'shd634cb91, 32'shd6372cb3, 32'shd6398df0, 32'shd63bef46, 32'shd63e50b5, 32'shd640b23f, 32'shd64313e2, 
               32'shd645759f, 32'shd647d776, 32'shd64a3966, 32'shd64c9b71, 32'shd64efd94, 32'shd6515fd2, 32'shd653c229, 32'shd656249b, 
               32'shd6588725, 32'shd65ae9ca, 32'shd65d4c88, 32'shd65faf60, 32'shd6621251, 32'shd664755c, 32'shd666d881, 32'shd6693bc0, 
               32'shd66b9f18, 32'shd66e028a, 32'shd6706615, 32'shd672c9ba, 32'shd6752d79, 32'shd6779151, 32'shd679f543, 32'shd67c594f, 
               32'shd67ebd74, 32'shd68121b3, 32'shd683860b, 32'shd685ea7d, 32'shd6884f09, 32'shd68ab3ae, 32'shd68d186d, 32'shd68f7d45, 
               32'shd691e237, 32'shd6944742, 32'shd696ac67, 32'shd69911a6, 32'shd69b76fe, 32'shd69ddc6f, 32'shd6a041fa, 32'shd6a2a79f, 
               32'shd6a50d5d, 32'shd6a77335, 32'shd6a9d926, 32'shd6ac3f31, 32'shd6aea555, 32'shd6b10b92, 32'shd6b371ea, 32'shd6b5d85a, 
               32'shd6b83ee4, 32'shd6baa588, 32'shd6bd0c45, 32'shd6bf731b, 32'shd6c1da0b, 32'shd6c44114, 32'shd6c6a837, 32'shd6c90f73, 
               32'shd6cb76c9, 32'shd6cdde38, 32'shd6d045c0, 32'shd6d2ad62, 32'shd6d5151d, 32'shd6d77cf2, 32'shd6d9e4e0, 32'shd6dc4ce7, 
               32'shd6deb508, 32'shd6e11d42, 32'shd6e38596, 32'shd6e5ee03, 32'shd6e85689, 32'shd6eabf28, 32'shd6ed27e1, 32'shd6ef90b4, 
               32'shd6f1f99f, 32'shd6f462a4, 32'shd6f6cbc2, 32'shd6f934fa, 32'shd6fb9e4b, 32'shd6fe07b5, 32'shd7007138, 32'shd702dad5, 
               32'shd705448b, 32'shd707ae5a, 32'shd70a1843, 32'shd70c8245, 32'shd70eec60, 32'shd7115694, 32'shd713c0e2, 32'shd7162b49, 
               32'shd71895c9, 32'shd71b0062, 32'shd71d6b15, 32'shd71fd5e0, 32'shd72240c5, 32'shd724abc4, 32'shd72716db, 32'shd729820c, 
               32'shd72bed55, 32'shd72e58b8, 32'shd730c434, 32'shd7332fca, 32'shd7359b78, 32'shd7380740, 32'shd73a7321, 32'shd73cdf1b, 
               32'shd73f4b2e, 32'shd741b75a, 32'shd744239f, 32'shd7468ffe, 32'shd748fc75, 32'shd74b6906, 32'shd74dd5b0, 32'shd7504273, 
               32'shd752af4f, 32'shd7551c44, 32'shd7578952, 32'shd759f679, 32'shd75c63ba, 32'shd75ed113, 32'shd7613e86, 32'shd763ac11, 
               32'shd76619b6, 32'shd7688774, 32'shd76af54a, 32'shd76d633a, 32'shd76fd143, 32'shd7723f64, 32'shd774ad9f, 32'shd7771bf3, 
               32'shd7798a60, 32'shd77bf8e6, 32'shd77e6784, 32'shd780d63c, 32'shd783450d, 32'shd785b3f7, 32'shd78822f9, 32'shd78a9215, 
               32'shd78d014a, 32'shd78f7097, 32'shd791dffe, 32'shd7944f7d, 32'shd796bf16, 32'shd7992ec7, 32'shd79b9e91, 32'shd79e0e74, 
               32'shd7a07e70, 32'shd7a2ee85, 32'shd7a55eb3, 32'shd7a7cefa, 32'shd7aa3f5a, 32'shd7acafd2, 32'shd7af2063, 32'shd7b1910e, 
               32'shd7b401d1, 32'shd7b672ad, 32'shd7b8e3a2, 32'shd7bb54af, 32'shd7bdc5d6, 32'shd7c03715, 32'shd7c2a86d, 32'shd7c519de, 
               32'shd7c78b68, 32'shd7c9fd0b, 32'shd7cc6ec6, 32'shd7cee09b, 32'shd7d15288, 32'shd7d3c48d, 32'shd7d636ac, 32'shd7d8a8e3, 
               32'shd7db1b34, 32'shd7dd8d9c, 32'shd7e0001e, 32'shd7e272b8, 32'shd7e4e56c, 32'shd7e75838, 32'shd7e9cb1c, 32'shd7ec3e1a, 
               32'shd7eeb130, 32'shd7f1245e, 32'shd7f397a6, 32'shd7f60b06, 32'shd7f87e7f, 32'shd7faf211, 32'shd7fd65bb, 32'shd7ffd97e, 
               32'shd8024d59, 32'shd804c14e, 32'shd807355b, 32'shd809a980, 32'shd80c1dbf, 32'shd80e9216, 32'shd8110685, 32'shd8137b0d, 
               32'shd815efae, 32'shd8186468, 32'shd81ad93a, 32'shd81d4e24, 32'shd81fc328, 32'shd8223843, 32'shd824ad78, 32'shd82722c5, 
               32'shd829982b, 32'shd82c0da9, 32'shd82e833f, 32'shd830f8ef, 32'shd8336eb7, 32'shd835e497, 32'shd8385a90, 32'shd83ad0a2, 
               32'shd83d46cc, 32'shd83fbd0e, 32'shd8423369, 32'shd844a9dd, 32'shd8472069, 32'shd849970e, 32'shd84c0dcb, 32'shd84e84a0, 
               32'shd850fb8e, 32'shd8537295, 32'shd855e9b4, 32'shd85860ec, 32'shd85ad83c, 32'shd85d4fa4, 32'shd85fc725, 32'shd8623ebe, 
               32'shd864b670, 32'shd8672e3a, 32'shd869a61d, 32'shd86c1e18, 32'shd86e962b, 32'shd8710e57, 32'shd873869b, 32'shd875fef8, 
               32'shd878776d, 32'shd87aeffa, 32'shd87d68a0, 32'shd87fe15e, 32'shd8825a35, 32'shd884d324, 32'shd8874c2b, 32'shd889c54b, 
               32'shd88c3e83, 32'shd88eb7d3, 32'shd891313b, 32'shd893aabc, 32'shd8962456, 32'shd8989e07, 32'shd89b17d1, 32'shd89d91b3, 
               32'shd8a00bae, 32'shd8a285c0, 32'shd8a4ffec, 32'shd8a77a2f, 32'shd8a9f48a, 32'shd8ac6efe, 32'shd8aee98a, 32'shd8b1642f, 
               32'shd8b3deeb, 32'shd8b659c0, 32'shd8b8d4ad, 32'shd8bb4fb3, 32'shd8bdcad0, 32'shd8c04606, 32'shd8c2c154, 32'shd8c53cba, 
               32'shd8c7b838, 32'shd8ca33cf, 32'shd8ccaf7e, 32'shd8cf2b45, 32'shd8d1a724, 32'shd8d4231b, 32'shd8d69f2a, 32'shd8d91b52, 
               32'shd8db9792, 32'shd8de13ea, 32'shd8e0905a, 32'shd8e30ce2, 32'shd8e58982, 32'shd8e8063a, 32'shd8ea830b, 32'shd8ecfff4, 
               32'shd8ef7cf4, 32'shd8f1fa0d, 32'shd8f4773e, 32'shd8f6f487, 32'shd8f971e8, 32'shd8fbef61, 32'shd8fe6cf2, 32'shd900ea9c, 
               32'shd903685d, 32'shd905e636, 32'shd9086428, 32'shd90ae231, 32'shd90d6053, 32'shd90fde8c, 32'shd9125cde, 32'shd914db47, 
               32'shd91759c9, 32'shd919d863, 32'shd91c5714, 32'shd91ed5de, 32'shd92154bf, 32'shd923d3b9, 32'shd92652ca, 32'shd928d1f4, 
               32'shd92b5135, 32'shd92dd08e, 32'shd9305000, 32'shd932cf89, 32'shd9354f2a, 32'shd937cee3, 32'shd93a4eb4, 32'shd93cce9d, 
               32'shd93f4e9e, 32'shd941ceb7, 32'shd9444ee7, 32'shd946cf30, 32'shd9494f90, 32'shd94bd009, 32'shd94e5099, 32'shd950d141, 
               32'shd9535201, 32'shd955d2d9, 32'shd95853c8, 32'shd95ad4d0, 32'shd95d55ef, 32'shd95fd726, 32'shd9625875, 32'shd964d9dc, 
               32'shd9675b5a, 32'shd969dcf1, 32'shd96c5e9f, 32'shd96ee065, 32'shd9716243, 32'shd973e438, 32'shd9766646, 32'shd978e86b, 
               32'shd97b6aa8, 32'shd97decfd, 32'shd9806f69, 32'shd982f1ed, 32'shd9857489, 32'shd987f73d, 32'shd98a7a08, 32'shd98cfceb, 
               32'shd98f7fe6, 32'shd99202f8, 32'shd9948623, 32'shd9970965, 32'shd9998cbe, 32'shd99c102f, 32'shd99e93b8, 32'shd9a11759, 
               32'shd9a39b11, 32'shd9a61ee1, 32'shd9a8a2c9, 32'shd9ab26c8, 32'shd9adaadf, 32'shd9b02f0e, 32'shd9b2b354, 32'shd9b537b2, 
               32'shd9b7bc27, 32'shd9ba40b5, 32'shd9bcc559, 32'shd9bf4a15, 32'shd9c1cee9, 32'shd9c453d5, 32'shd9c6d8d8, 32'shd9c95df3, 
               32'shd9cbe325, 32'shd9ce686e, 32'shd9d0edd0, 32'shd9d37349, 32'shd9d5f8d9, 32'shd9d87e81, 32'shd9db0441, 32'shd9dd8a18, 
               32'shd9e01006, 32'shd9e2960c, 32'shd9e51c2a, 32'shd9e7a25f, 32'shd9ea28ac, 32'shd9ecaf10, 32'shd9ef358b, 32'shd9f1bc1e, 
               32'shd9f442c9, 32'shd9f6c98b, 32'shd9f95064, 32'shd9fbd755, 32'shd9fe5e5e, 32'shda00e57d, 32'shda036cb5, 32'shda05f403, 
               32'shda087b69, 32'shda0b02e7, 32'shda0d8a7c, 32'shda101228, 32'shda1299ec, 32'shda1521c7, 32'shda17a9ba, 32'shda1a31c4, 
               32'shda1cb9e5, 32'shda1f421e, 32'shda21ca6e, 32'shda2452d5, 32'shda26db54, 32'shda2963ea, 32'shda2bec97, 32'shda2e755c, 
               32'shda30fe38, 32'shda33872c, 32'shda361036, 32'shda389958, 32'shda3b2292, 32'shda3dabe2, 32'shda40354a, 32'shda42beca, 
               32'shda454860, 32'shda47d20e, 32'shda4a5bd3, 32'shda4ce5af, 32'shda4f6fa3, 32'shda51f9ae, 32'shda5483d0, 32'shda570e09, 
               32'shda599859, 32'shda5c22c1, 32'shda5ead40, 32'shda6137d6, 32'shda63c284, 32'shda664d48, 32'shda68d824, 32'shda6b6317, 
               32'shda6dee21, 32'shda707942, 32'shda73047b, 32'shda758fcb, 32'shda781b31, 32'shda7aa6af, 32'shda7d3244, 32'shda7fbdf1, 
               32'shda8249b4, 32'shda84d58f, 32'shda876180, 32'shda89ed89, 32'shda8c79a9, 32'shda8f05e0, 32'shda91922e, 32'shda941e93, 
               32'shda96ab0f, 32'shda9937a2, 32'shda9bc44d, 32'shda9e510e, 32'shdaa0dde7, 32'shdaa36ad6, 32'shdaa5f7dd, 32'shdaa884fa, 
               32'shdaab122f, 32'shdaad9f7b, 32'shdab02cdd, 32'shdab2ba57, 32'shdab547e8, 32'shdab7d590, 32'shdaba634e, 32'shdabcf124, 
               32'shdabf7f11, 32'shdac20d15, 32'shdac49b2f, 32'shdac72961, 32'shdac9b7a9, 32'shdacc4609, 32'shdaced47f, 32'shdad1630d, 
               32'shdad3f1b1, 32'shdad6806d, 32'shdad90f3f, 32'shdadb9e28, 32'shdade2d28, 32'shdae0bc3f, 32'shdae34b6d, 32'shdae5dab2, 
               32'shdae86a0d, 32'shdaeaf980, 32'shdaed8909, 32'shdaf018a9, 32'shdaf2a860, 32'shdaf5382e, 32'shdaf7c813, 32'shdafa580f, 
               32'shdafce821, 32'shdaff784b, 32'shdb02088b, 32'shdb0498e2, 32'shdb072950, 32'shdb09b9d4, 32'shdb0c4a70, 32'shdb0edb22, 
               32'shdb116beb, 32'shdb13fccb, 32'shdb168dc1, 32'shdb191ece, 32'shdb1baff2, 32'shdb1e412d, 32'shdb20d27f, 32'shdb2363e7, 
               32'shdb25f566, 32'shdb2886fc, 32'shdb2b18a9, 32'shdb2daa6c, 32'shdb303c46, 32'shdb32ce36, 32'shdb35603e, 32'shdb37f25c, 
               32'shdb3a8491, 32'shdb3d16dc, 32'shdb3fa93e, 32'shdb423bb7, 32'shdb44ce46, 32'shdb4760ec, 32'shdb49f3a9, 32'shdb4c867d, 
               32'shdb4f1967, 32'shdb51ac67, 32'shdb543f7e, 32'shdb56d2ac, 32'shdb5965f1, 32'shdb5bf94c, 32'shdb5e8cbe, 32'shdb612046, 
               32'shdb63b3e5, 32'shdb66479b, 32'shdb68db67, 32'shdb6b6f49, 32'shdb6e0342, 32'shdb709752, 32'shdb732b79, 32'shdb75bfb5, 
               32'shdb785409, 32'shdb7ae873, 32'shdb7d7cf3, 32'shdb80118a, 32'shdb82a638, 32'shdb853afc, 32'shdb87cfd6, 32'shdb8a64c7, 
               32'shdb8cf9cf, 32'shdb8f8eed, 32'shdb922421, 32'shdb94b96c, 32'shdb974ece, 32'shdb99e445, 32'shdb9c79d4, 32'shdb9f0f78, 
               32'shdba1a534, 32'shdba43b05, 32'shdba6d0ed, 32'shdba966ec, 32'shdbabfd01, 32'shdbae932c, 32'shdbb1296e, 32'shdbb3bfc6, 
               32'shdbb65634, 32'shdbb8ecb9, 32'shdbbb8354, 32'shdbbe1a06, 32'shdbc0b0ce, 32'shdbc347ac, 32'shdbc5dea1, 32'shdbc875ac, 
               32'shdbcb0cce, 32'shdbcda405, 32'shdbd03b53, 32'shdbd2d2b8, 32'shdbd56a32, 32'shdbd801c3, 32'shdbda996b, 32'shdbdd3128, 
               32'shdbdfc8fc, 32'shdbe260e6, 32'shdbe4f8e7, 32'shdbe790fe, 32'shdbea292b, 32'shdbecc16e, 32'shdbef59c7, 32'shdbf1f237, 
               32'shdbf48abd, 32'shdbf72359, 32'shdbf9bc0c, 32'shdbfc54d4, 32'shdbfeedb3, 32'shdc0186a8, 32'shdc041fb4, 32'shdc06b8d5, 
               32'shdc09520d, 32'shdc0beb5b, 32'shdc0e84bf, 32'shdc111e39, 32'shdc13b7c9, 32'shdc165170, 32'shdc18eb2d, 32'shdc1b8500, 
               32'shdc1e1ee9, 32'shdc20b8e8, 32'shdc2352fd, 32'shdc25ed28, 32'shdc28876a, 32'shdc2b21c1, 32'shdc2dbc2f, 32'shdc3056b3, 
               32'shdc32f14d, 32'shdc358bfd, 32'shdc3826c3, 32'shdc3ac19f, 32'shdc3d5c91, 32'shdc3ff799, 32'shdc4292b8, 32'shdc452dec, 
               32'shdc47c936, 32'shdc4a6497, 32'shdc4d000d, 32'shdc4f9b9a, 32'shdc52373c, 32'shdc54d2f5, 32'shdc576ec3, 32'shdc5a0aa8, 
               32'shdc5ca6a2, 32'shdc5f42b2, 32'shdc61ded9, 32'shdc647b15, 32'shdc671768, 32'shdc69b3d0, 32'shdc6c504e, 32'shdc6eece2, 
               32'shdc71898d, 32'shdc74264d, 32'shdc76c323, 32'shdc79600f, 32'shdc7bfd11, 32'shdc7e9a28, 32'shdc813756, 32'shdc83d49a, 
               32'shdc8671f3, 32'shdc890f62, 32'shdc8bace8, 32'shdc8e4a83, 32'shdc90e834, 32'shdc9385fa, 32'shdc9623d7, 32'shdc98c1ca, 
               32'shdc9b5fd2, 32'shdc9dfdf0, 32'shdca09c24, 32'shdca33a6e, 32'shdca5d8cd, 32'shdca87743, 32'shdcab15ce, 32'shdcadb46f, 
               32'shdcb05326, 32'shdcb2f1f3, 32'shdcb590d5, 32'shdcb82fcd, 32'shdcbacedb, 32'shdcbd6dff, 32'shdcc00d38, 32'shdcc2ac87, 
               32'shdcc54bec, 32'shdcc7eb67, 32'shdcca8af7, 32'shdccd2a9d, 32'shdccfca59, 32'shdcd26a2a, 32'shdcd50a12, 32'shdcd7aa0e, 
               32'shdcda4a21, 32'shdcdcea49, 32'shdcdf8a87, 32'shdce22adb, 32'shdce4cb44, 32'shdce76bc3, 32'shdcea0c58, 32'shdcecad02, 
               32'shdcef4dc2, 32'shdcf1ee97, 32'shdcf48f82, 32'shdcf73083, 32'shdcf9d199, 32'shdcfc72c5, 32'shdcff1407, 32'shdd01b55e, 
               32'shdd0456ca, 32'shdd06f84d, 32'shdd0999e4, 32'shdd0c3b92, 32'shdd0edd55, 32'shdd117f2d, 32'shdd14211b, 32'shdd16c31f, 
               32'shdd196538, 32'shdd1c0767, 32'shdd1ea9ab, 32'shdd214c05, 32'shdd23ee74, 32'shdd2690f9, 32'shdd293393, 32'shdd2bd643, 
               32'shdd2e7908, 32'shdd311be3, 32'shdd33bed3, 32'shdd3661d8, 32'shdd3904f4, 32'shdd3ba824, 32'shdd3e4b6a, 32'shdd40eec5, 
               32'shdd439236, 32'shdd4635bd, 32'shdd48d958, 32'shdd4b7d09, 32'shdd4e20d0, 32'shdd50c4ac, 32'shdd53689d, 32'shdd560ca4, 
               32'shdd58b0c0, 32'shdd5b54f1, 32'shdd5df938, 32'shdd609d94, 32'shdd634206, 32'shdd65e68d, 32'shdd688b29, 32'shdd6b2fdb, 
               32'shdd6dd4a2, 32'shdd70797e, 32'shdd731e6f, 32'shdd75c376, 32'shdd786892, 32'shdd7b0dc4, 32'shdd7db30b, 32'shdd805867, 
               32'shdd82fdd8, 32'shdd85a35f, 32'shdd8848fb, 32'shdd8aeeac, 32'shdd8d9472, 32'shdd903a4e, 32'shdd92e03f, 32'shdd958645, 
               32'shdd982c60, 32'shdd9ad291, 32'shdd9d78d7, 32'shdda01f32, 32'shdda2c5a2, 32'shdda56c27, 32'shdda812c2, 32'shddaab972, 
               32'shddad6036, 32'shddb00711, 32'shddb2ae00, 32'shddb55504, 32'shddb7fc1e, 32'shddbaa34d, 32'shddbd4a91, 32'shddbff1ea, 
               32'shddc29958, 32'shddc540db, 32'shddc7e873, 32'shddca9021, 32'shddcd37e4, 32'shddcfdfbb, 32'shddd287a8, 32'shddd52faa, 
               32'shddd7d7c1, 32'shddda7fed, 32'shdddd282e, 32'shdddfd084, 32'shdde278ef, 32'shdde5216f, 32'shdde7ca05, 32'shddea72af, 
               32'shdded1b6e, 32'shddefc443, 32'shddf26d2c, 32'shddf5162a, 32'shddf7bf3e, 32'shddfa6866, 32'shddfd11a3, 32'shddffbaf6, 
               32'shde02645d, 32'shde050dd9, 32'shde07b76b, 32'shde0a6111, 32'shde0d0acc, 32'shde0fb49c, 32'shde125e81, 32'shde15087b, 
               32'shde17b28a, 32'shde1a5cad, 32'shde1d06e6, 32'shde1fb134, 32'shde225b96, 32'shde25060e, 32'shde27b09a, 32'shde2a5b3b, 
               32'shde2d05f1, 32'shde2fb0bc, 32'shde325b9b, 32'shde350690, 32'shde37b199, 32'shde3a5cb8, 32'shde3d07eb, 32'shde3fb333, 
               32'shde425e8f, 32'shde450a01, 32'shde47b587, 32'shde4a6122, 32'shde4d0cd2, 32'shde4fb897, 32'shde526471, 32'shde55105f, 
               32'shde57bc62, 32'shde5a687a, 32'shde5d14a6, 32'shde5fc0e8, 32'shde626d3e, 32'shde6519a9, 32'shde67c628, 32'shde6a72bc, 
               32'shde6d1f65, 32'shde6fcc23, 32'shde7278f5, 32'shde7525dc, 32'shde77d2d8, 32'shde7a7fe9, 32'shde7d2d0e, 32'shde7fda48, 
               32'shde828796, 32'shde8534f9, 32'shde87e271, 32'shde8a8ffd, 32'shde8d3d9e, 32'shde8feb54, 32'shde92991e, 32'shde9546fd, 
               32'shde97f4f1, 32'shde9aa2f9, 32'shde9d5116, 32'shde9fff47, 32'shdea2ad8d, 32'shdea55be8, 32'shdea80a57, 32'shdeaab8da, 
               32'shdead6773, 32'shdeb0161f, 32'shdeb2c4e1, 32'shdeb573b7, 32'shdeb822a1, 32'shdebad1a0, 32'shdebd80b3, 32'shdec02fdb, 
               32'shdec2df18, 32'shdec58e69, 32'shdec83dce, 32'shdecaed48, 32'shdecd9cd7, 32'shded04c7a, 32'shded2fc31, 32'shded5abfd, 
               32'shded85bdd, 32'shdedb0bd2, 32'shdeddbbdb, 32'shdee06bf9, 32'shdee31c2b, 32'shdee5cc72, 32'shdee87ccc, 32'shdeeb2d3c, 
               32'shdeedddc0, 32'shdef08e58, 32'shdef33f04, 32'shdef5efc5, 32'shdef8a09b, 32'shdefb5184, 32'shdefe0282, 32'shdf00b395, 
               32'shdf0364bc, 32'shdf0615f7, 32'shdf08c746, 32'shdf0b78aa, 32'shdf0e2a22, 32'shdf10dbaf, 32'shdf138d4f, 32'shdf163f04, 
               32'shdf18f0ce, 32'shdf1ba2ab, 32'shdf1e549d, 32'shdf2106a4, 32'shdf23b8be, 32'shdf266aed, 32'shdf291d30, 32'shdf2bcf87, 
               32'shdf2e81f3, 32'shdf313473, 32'shdf33e707, 32'shdf3699af, 32'shdf394c6b, 32'shdf3bff3c, 32'shdf3eb221, 32'shdf41651a, 
               32'shdf441828, 32'shdf46cb49, 32'shdf497e7f, 32'shdf4c31c9, 32'shdf4ee527, 32'shdf519899, 32'shdf544c1f, 32'shdf56ffba, 
               32'shdf59b369, 32'shdf5c672b, 32'shdf5f1b02, 32'shdf61ceee, 32'shdf6482ed, 32'shdf673700, 32'shdf69eb27, 32'shdf6c9f63, 
               32'shdf6f53b3, 32'shdf720816, 32'shdf74bc8e, 32'shdf77711a, 32'shdf7a25ba, 32'shdf7cda6e, 32'shdf7f8f36, 32'shdf824412, 
               32'shdf84f902, 32'shdf87ae06, 32'shdf8a631f, 32'shdf8d184b, 32'shdf8fcd8b, 32'shdf9282df, 32'shdf953848, 32'shdf97edc4, 
               32'shdf9aa354, 32'shdf9d58f8, 32'shdfa00eb1, 32'shdfa2c47d, 32'shdfa57a5d, 32'shdfa83051, 32'shdfaae659, 32'shdfad9c75, 
               32'shdfb052a5, 32'shdfb308e9, 32'shdfb5bf41, 32'shdfb875ac, 32'shdfbb2c2c, 32'shdfbde2bf, 32'shdfc09967, 32'shdfc35022, 
               32'shdfc606f1, 32'shdfc8bdd4, 32'shdfcb74cb, 32'shdfce2bd6, 32'shdfd0e2f5, 32'shdfd39a27, 32'shdfd6516e, 32'shdfd908c8, 
               32'shdfdbc036, 32'shdfde77b8, 32'shdfe12f4e, 32'shdfe3e6f7, 32'shdfe69eb4, 32'shdfe95686, 32'shdfec0e6a, 32'shdfeec663, 
               32'shdff17e70, 32'shdff43690, 32'shdff6eec4, 32'shdff9a70c, 32'shdffc5f67, 32'shdfff17d7, 32'she001d05a, 32'she00488f0, 
               32'she007419b, 32'she009fa59, 32'she00cb32b, 32'she00f6c11, 32'she012250a, 32'she014de17, 32'she0179738, 32'she01a506c, 
               32'she01d09b4, 32'she01fc310, 32'she0227c7f, 32'she0253602, 32'she027ef99, 32'she02aa943, 32'she02d6301, 32'she0301cd3, 
               32'she032d6b8, 32'she03590b1, 32'she0384abe, 32'she03b04de, 32'she03dbf11, 32'she0407959, 32'she04333b3, 32'she045ee22, 
               32'she048a8a4, 32'she04b6339, 32'she04e1de3, 32'she050d89f, 32'she053936f, 32'she0564e53, 32'she059094a, 32'she05bc455, 
               32'she05e7f74, 32'she0613aa5, 32'she063f5eb, 32'she066b144, 32'she0696cb0, 32'she06c2830, 32'she06ee3c3, 32'she0719f6a, 
               32'she0745b24, 32'she07716f2, 32'she079d2d3, 32'she07c8ec7, 32'she07f4acf, 32'she08206eb, 32'she084c31a, 32'she0877f5c, 
               32'she08a3bb2, 32'she08cf81b, 32'she08fb497, 32'she0927127, 32'she0952dcb, 32'she097ea81, 32'she09aa74b, 32'she09d6429, 
               32'she0a0211a, 32'she0a2de1e, 32'she0a59b35, 32'she0a85860, 32'she0ab159e, 32'she0add2f0, 32'she0b09055, 32'she0b34dcd, 
               32'she0b60b58, 32'she0b8c8f7, 32'she0bb86a9, 32'she0be446e, 32'she0c10247, 32'she0c3c033, 32'she0c67e32, 32'she0c93c44, 
               32'she0cbfa6a, 32'she0ceb8a3, 32'she0d176ef, 32'she0d4354e, 32'she0d6f3c1, 32'she0d9b247, 32'she0dc70e0, 32'she0df2f8c, 
               32'she0e1ee4b, 32'she0e4ad1e, 32'she0e76c04, 32'she0ea2afd, 32'she0ecea09, 32'she0efa928, 32'she0f2685b, 32'she0f527a0, 
               32'she0f7e6f9, 32'she0faa665, 32'she0fd65e4, 32'she1002577, 32'she102e51c, 32'she105a4d4, 32'she10864a0, 32'she10b247f, 
               32'she10de470, 32'she110a475, 32'she113648d, 32'she11624b8, 32'she118e4f6, 32'she11ba547, 32'she11e65ac, 32'she1212623, 
               32'she123e6ad, 32'she126a74a, 32'she12967fb, 32'she12c28be, 32'she12ee995, 32'she131aa7e, 32'she1346b7a, 32'she1372c8a, 
               32'she139edac, 32'she13caee1, 32'she13f702a, 32'she1423185, 32'she144f2f3, 32'she147b475, 32'she14a7609, 32'she14d37b0, 
               32'she14ff96a, 32'she152bb37, 32'she1557d17, 32'she1583f0a, 32'she15b0110, 32'she15dc328, 32'she1608554, 32'she1634792, 
               32'she16609e3, 32'she168cc48, 32'she16b8ebf, 32'she16e5149, 32'she17113e5, 32'she173d695, 32'she1769958, 32'she1795c2d, 
               32'she17c1f15, 32'she17ee210, 32'she181a51e, 32'she184683e, 32'she1872b72, 32'she189eeb8, 32'she18cb211, 32'she18f757d, 
               32'she19238fb, 32'she194fc8d, 32'she197c031, 32'she19a83e7, 32'she19d47b1, 32'she1a00b8d, 32'she1a2cf7c, 32'she1a5937e, 
               32'she1a85793, 32'she1ab1bba, 32'she1addff4, 32'she1b0a441, 32'she1b368a0, 32'she1b62d12, 32'she1b8f197, 32'she1bbb62e, 
               32'she1be7ad8, 32'she1c13f95, 32'she1c40464, 32'she1c6c946, 32'she1c98e3b, 32'she1cc5342, 32'she1cf185c, 32'she1d1dd89, 
               32'she1d4a2c8, 32'she1d7681a, 32'she1da2d7e, 32'she1dcf2f5, 32'she1dfb87f, 32'she1e27e1b, 32'she1e543ca, 32'she1e8098b, 
               32'she1eacf5f, 32'she1ed9545, 32'she1f05b3e, 32'she1f3214a, 32'she1f5e768, 32'she1f8ad98, 32'she1fb73dc, 32'she1fe3a31, 
               32'she2010099, 32'she203c714, 32'she2068da1, 32'she2095441, 32'she20c1af3, 32'she20ee1b7, 32'she211a88f, 32'she2146f78, 
               32'she2173674, 32'she219fd82, 32'she21cc4a3, 32'she21f8bd7, 32'she222531c, 32'she2251a75, 32'she227e1df, 32'she22aa95c, 
               32'she22d70eb, 32'she230388d, 32'she2330041, 32'she235c808, 32'she2388fe1, 32'she23b57cc, 32'she23e1fca, 32'she240e7da, 
               32'she243affc, 32'she2467831, 32'she2494078, 32'she24c08d1, 32'she24ed13d, 32'she25199bb, 32'she254624b, 32'she2572aee, 
               32'she259f3a3, 32'she25cbc6a, 32'she25f8544, 32'she2624e2f, 32'she265172e, 32'she267e03e, 32'she26aa960, 32'she26d7295, 
               32'she2703bdc, 32'she2730536, 32'she275cea1, 32'she278981f, 32'she27b61af, 32'she27e2b51, 32'she280f505, 32'she283becc, 
               32'she28688a4, 32'she289528f, 32'she28c1c8c, 32'she28ee69c, 32'she291b0bd, 32'she2947af1, 32'she2974536, 32'she29a0f8e, 
               32'she29cd9f8, 32'she29fa474, 32'she2a26f03, 32'she2a539a3, 32'she2a80456, 32'she2aacf1a, 32'she2ad99f1, 32'she2b064da, 
               32'she2b32fd4, 32'she2b5fae1, 32'she2b8c600, 32'she2bb9131, 32'she2be5c74, 32'she2c127c9, 32'she2c3f331, 32'she2c6beaa, 
               32'she2c98a35, 32'she2cc55d2, 32'she2cf2182, 32'she2d1ed43, 32'she2d4b916, 32'she2d784fb, 32'she2da50f3, 32'she2dd1cfc, 
               32'she2dfe917, 32'she2e2b544, 32'she2e58183, 32'she2e84dd4, 32'she2eb1a37, 32'she2ede6ac, 32'she2f0b333, 32'she2f37fcc, 
               32'she2f64c77, 32'she2f91934, 32'she2fbe602, 32'she2feb2e3, 32'she3017fd5, 32'she3044cd9, 32'she30719ef, 32'she309e717, 
               32'she30cb451, 32'she30f819d, 32'she3124efa, 32'she3151c6a, 32'she317e9eb, 32'she31ab77e, 32'she31d8523, 32'she32052da, 
               32'she32320a2, 32'she325ee7d, 32'she328bc69, 32'she32b8a67, 32'she32e5876, 32'she3312698, 32'she333f4cb, 32'she336c310, 
               32'she3399167, 32'she33c5fcf, 32'she33f2e4a, 32'she341fcd6, 32'she344cb73, 32'she3479a23, 32'she34a68e4, 32'she34d37b7, 
               32'she350069b, 32'she352d592, 32'she355a49a, 32'she35873b3, 32'she35b42df, 32'she35e121c, 32'she360e16a, 32'she363b0cb, 
               32'she366803c, 32'she3694fc0, 32'she36c1f55, 32'she36eeefc, 32'she371beb5, 32'she3748e7f, 32'she3775e5a, 32'she37a2e48, 
               32'she37cfe47, 32'she37fce57, 32'she3829e79, 32'she3856ead, 32'she3883ef2, 32'she38b0f49, 32'she38ddfb1, 32'she390b02b, 
               32'she39380b6, 32'she3965153, 32'she3992202, 32'she39bf2c2, 32'she39ec393, 32'she3a19476, 32'she3a4656b, 32'she3a73671, 
               32'she3aa0788, 32'she3acd8b1, 32'she3afa9ec, 32'she3b27b38, 32'she3b54c95, 32'she3b81e04, 32'she3baef84, 32'she3bdc116, 
               32'she3c092b9, 32'she3c3646d, 32'she3c63633, 32'she3c9080b, 32'she3cbd9f4, 32'she3ceabee, 32'she3d17df9, 32'she3d45016, 
               32'she3d72245, 32'she3d9f484, 32'she3dcc6d5, 32'she3df9938, 32'she3e26bac, 32'she3e53e31, 32'she3e810c7, 32'she3eae36f, 
               32'she3edb628, 32'she3f088f2, 32'she3f35bce, 32'she3f62ebb, 32'she3f901ba, 32'she3fbd4c9, 32'she3fea7ea, 32'she4017b1c, 
               32'she4044e60, 32'she40721b4, 32'she409f51a, 32'she40cc891, 32'she40f9c1a, 32'she4126fb4, 32'she415435f, 32'she418171b, 
               32'she41aeae8, 32'she41dbec7, 32'she42092b6, 32'she42366b7, 32'she4263ac9, 32'she4290eed, 32'she42be321, 32'she42eb767, 
               32'she4318bbe, 32'she4346026, 32'she437349f, 32'she43a0929, 32'she43cddc4, 32'she43fb271, 32'she442872e, 32'she4455bfd, 
               32'she44830dd, 32'she44b05ce, 32'she44ddad0, 32'she450afe3, 32'she4538507, 32'she4565a3c, 32'she4592f83, 32'she45c04da, 
               32'she45eda43, 32'she461afbc, 32'she4648547, 32'she4675ae2, 32'she46a308f, 32'she46d064c, 32'she46fdc1b, 32'she472b1fa, 
               32'she47587eb, 32'she4785ded, 32'she47b33ff, 32'she47e0a23, 32'she480e057, 32'she483b69d, 32'she4868cf3, 32'she489635a, 
               32'she48c39d3, 32'she48f105c, 32'she491e6f6, 32'she494bda1, 32'she497945d, 32'she49a6b2a, 32'she49d4208, 32'she4a018f7, 
               32'she4a2eff6, 32'she4a5c707, 32'she4a89e28, 32'she4ab755a, 32'she4ae4c9d, 32'she4b123f1, 32'she4b3fb56, 32'she4b6d2cb, 
               32'she4b9aa52, 32'she4bc81e9, 32'she4bf5991, 32'she4c2314a, 32'she4c50914, 32'she4c7e0ee, 32'she4cab8d9, 32'she4cd90d5, 
               32'she4d068e2, 32'she4d34100, 32'she4d6192e, 32'she4d8f16d, 32'she4dbc9bd, 32'she4dea21e, 32'she4e17a8f, 32'she4e45311, 
               32'she4e72ba4, 32'she4ea0448, 32'she4ecdcfc, 32'she4efb5c1, 32'she4f28e96, 32'she4f5677d, 32'she4f84074, 32'she4fb197b, 
               32'she4fdf294, 32'she500cbbc, 32'she503a4f6, 32'she5067e40, 32'she509579b, 32'she50c3107, 32'she50f0a83, 32'she511e410, 
               32'she514bdad, 32'she517975b, 32'she51a711a, 32'she51d4ae9, 32'she52024c9, 32'she522feb9, 32'she525d8ba, 32'she528b2cc, 
               32'she52b8cee, 32'she52e6720, 32'she5314163, 32'she5341bb7, 32'she536f61b, 32'she539d090, 32'she53cab15, 32'she53f85ab, 
               32'she5426051, 32'she5453b08, 32'she54815cf, 32'she54af0a7, 32'she54dcb8f, 32'she550a688, 32'she5538191, 32'she5565cab, 
               32'she55937d5, 32'she55c130f, 32'she55eee5a, 32'she561c9b5, 32'she564a521, 32'she567809d, 32'she56a5c2a, 32'she56d37c7, 
               32'she5701374, 32'she572ef32, 32'she575cb00, 32'she578a6de, 32'she57b82cd, 32'she57e5ecc, 32'she5813adc, 32'she58416fc, 
               32'she586f32c, 32'she589cf6d, 32'she58cabbe, 32'she58f881f, 32'she5926490, 32'she5954112, 32'she5981da4, 32'she59afa47, 
               32'she59dd6f9, 32'she5a0b3bc, 32'she5a39090, 32'she5a66d73, 32'she5a94a67, 32'she5ac276b, 32'she5af047f, 32'she5b1e1a3, 
               32'she5b4bed8, 32'she5b79c1d, 32'she5ba7972, 32'she5bd56d7, 32'she5c0344d, 32'she5c311d3, 32'she5c5ef69, 32'she5c8cd0f, 
               32'she5cbaac5, 32'she5ce888b, 32'she5d16662, 32'she5d44449, 32'she5d72240, 32'she5da0047, 32'she5dcde5e, 32'she5dfbc85, 
               32'she5e29abc, 32'she5e57904, 32'she5e8575b, 32'she5eb35c3, 32'she5ee143b, 32'she5f0f2c3, 32'she5f3d15b, 32'she5f6b003, 
               32'she5f98ebb, 32'she5fc6d83, 32'she5ff4c5b, 32'she6022b43, 32'she6050a3b, 32'she607e944, 32'she60ac85c, 32'she60da784, 
               32'she61086bc, 32'she6136605, 32'she616455d, 32'she61924c5, 32'she61c043d, 32'she61ee3c6, 32'she621c35e, 32'she624a306, 
               32'she62782be, 32'she62a6286, 32'she62d425e, 32'she6302246, 32'she633023e, 32'she635e245, 32'she638c25d, 32'she63ba285, 
               32'she63e82bc, 32'she6416303, 32'she644435a, 32'she64723c2, 32'she64a0438, 32'she64ce4bf, 32'she64fc556, 32'she652a5fc, 
               32'she65586b3, 32'she6586779, 32'she65b484f, 32'she65e2935, 32'she6610a2a, 32'she663eb30, 32'she666cc45, 32'she669ad6a, 
               32'she66c8e9f, 32'she66f6fe3, 32'she6725138, 32'she675329c, 32'she6781410, 32'she67af593, 32'she67dd727, 32'she680b8ca, 
               32'she6839a7c, 32'she6867c3f, 32'she6895e11, 32'she68c3ff3, 32'she68f21e5, 32'she69203e6, 32'she694e5f7, 32'she697c818, 
               32'she69aaa48, 32'she69d8c88, 32'she6a06ed8, 32'she6a35137, 32'she6a633a6, 32'she6a91625, 32'she6abf8b3, 32'she6aedb51, 
               32'she6b1bdff, 32'she6b4a0bc, 32'she6b78389, 32'she6ba6665, 32'she6bd4951, 32'she6c02c4c, 32'she6c30f57, 32'she6c5f272, 
               32'she6c8d59c, 32'she6cbb8d6, 32'she6ce9c1f, 32'she6d17f78, 32'she6d462e1, 32'she6d74658, 32'she6da29e0, 32'she6dd0d77, 
               32'she6dff11d, 32'she6e2d4d3, 32'she6e5b899, 32'she6e89c6d, 32'she6eb8052, 32'she6ee6446, 32'she6f14849, 32'she6f42c5c, 
               32'she6f7107e, 32'she6f9f4b0, 32'she6fcd8f1, 32'she6ffbd41, 32'she702a1a1, 32'she7058611, 32'she7086a8f, 32'she70b4f1e, 
               32'she70e33bb, 32'she7111868, 32'she713fd25, 32'she716e1f0, 32'she719c6cb, 32'she71cabb6, 32'she71f90b0, 32'she72275b9, 
               32'she7255ad1, 32'she7283ff9, 32'she72b2530, 32'she72e0a77, 32'she730efcc, 32'she733d531, 32'she736baa6, 32'she739a029, 
               32'she73c85bc, 32'she73f6b5f, 32'she7425110, 32'she74536d1, 32'she7481ca1, 32'she74b0280, 32'she74de86f, 32'she750ce6c, 
               32'she753b479, 32'she7569a95, 32'she75980c1, 32'she75c66fb, 32'she75f4d45, 32'she762339e, 32'she7651a06, 32'she768007e, 
               32'she76ae704, 32'she76dcd9a, 32'she770b43e, 32'she7739af2, 32'she77681b6, 32'she7796888, 32'she77c4f69, 32'she77f365a, 
               32'she7821d59, 32'she7850468, 32'she787eb86, 32'she78ad2b3, 32'she78db9ef, 32'she790a13a, 32'she7938894, 32'she7966ffd, 
               32'she7995776, 32'she79c3efd, 32'she79f2693, 32'she7a20e39, 32'she7a4f5ed, 32'she7a7ddb1, 32'she7aac583, 32'she7adad65, 
               32'she7b09555, 32'she7b37d55, 32'she7b66563, 32'she7b94d80, 32'she7bc35ad, 32'she7bf1de8, 32'she7c20633, 32'she7c4ee8c, 
               32'she7c7d6f4, 32'she7cabf6c, 32'she7cda7f2, 32'she7d09087, 32'she7d3792b, 32'she7d661de, 32'she7d94a9f, 32'she7dc3370, 
               32'she7df1c50, 32'she7e2053e, 32'she7e4ee3c, 32'she7e7d748, 32'she7eac063, 32'she7eda98d, 32'she7f092c6, 32'she7f37c0d, 
               32'she7f66564, 32'she7f94ec9, 32'she7fc383d, 32'she7ff21c0, 32'she8020b52, 32'she804f4f2, 32'she807dea2, 32'she80ac860, 
               32'she80db22d, 32'she8109c08, 32'she81385f3, 32'she8166fec, 32'she81959f4, 32'she81c440a, 32'she81f2e30, 32'she8221864, 
               32'she82502a7, 32'she827ecf8, 32'she82ad759, 32'she82dc1c8, 32'she830ac45, 32'she83396d2, 32'she836816d, 32'she8396c16, 
               32'she83c56cf, 32'she83f4196, 32'she8422c6c, 32'she8451750, 32'she8480243, 32'she84aed45, 32'she84dd855, 32'she850c374, 
               32'she853aea1, 32'she85699dd, 32'she8598528, 32'she85c7081, 32'she85f5be9, 32'she862475f, 32'she86532e4, 32'she8681e78, 
               32'she86b0a1a, 32'she86df5cb, 32'she870e18a, 32'she873cd57, 32'she876b934, 32'she879a51e, 32'she87c9118, 32'she87f7d1f, 
               32'she8826936, 32'she885555a, 32'she888418e, 32'she88b2dcf, 32'she88e1a20, 32'she891067e, 32'she893f2eb, 32'she896df67, 
               32'she899cbf1, 32'she89cb889, 32'she89fa530, 32'she8a291e5, 32'she8a57ea9, 32'she8a86b7b, 32'she8ab585c, 32'she8ae454b, 
               32'she8b13248, 32'she8b41f53, 32'she8b70c6d, 32'she8b9f996, 32'she8bce6cd, 32'she8bfd412, 32'she8c2c165, 32'she8c5aec7, 
               32'she8c89c37, 32'she8cb89b5, 32'she8ce7742, 32'she8d164dd, 32'she8d45286, 32'she8d7403e, 32'she8da2e04, 32'she8dd1bd8, 
               32'she8e009ba, 32'she8e2f7ab, 32'she8e5e5aa, 32'she8e8d3b7, 32'she8ebc1d3, 32'she8eeaffd, 32'she8f19e34, 32'she8f48c7b, 
               32'she8f77acf, 32'she8fa6932, 32'she8fd57a2, 32'she9004621, 32'she90334af, 32'she906234a, 32'she90911f3, 32'she90c00ab, 
               32'she90eef71, 32'she911de45, 32'she914cd27, 32'she917bc17, 32'she91aab16, 32'she91d9a22, 32'she920893d, 32'she9237866, 
               32'she926679c, 32'she92956e1, 32'she92c4634, 32'she92f3596, 32'she9322505, 32'she9351482, 32'she938040d, 32'she93af3a7, 
               32'she93de34e, 32'she940d304, 32'she943c2c7, 32'she946b299, 32'she949a278, 32'she94c9266, 32'she94f8261, 32'she952726b, 
               32'she9556282, 32'she95852a8, 32'she95b42db, 32'she95e331d, 32'she961236c, 32'she96413c9, 32'she9670435, 32'she969f4ae, 
               32'she96ce535, 32'she96fd5ca, 32'she972c66d, 32'she975b71e, 32'she978a7dd, 32'she97b98aa, 32'she97e8984, 32'she9817a6d, 
               32'she9846b63, 32'she9875c68, 32'she98a4d7a, 32'she98d3e9a, 32'she9902fc7, 32'she9932103, 32'she996124d, 32'she99903a4, 
               32'she99bf509, 32'she99ee67c, 32'she9a1d7fd, 32'she9a4c98b, 32'she9a7bb28, 32'she9aaacd2, 32'she9ad9e8a, 32'she9b0904f, 
               32'she9b38223, 32'she9b67404, 32'she9b965f3, 32'she9bc57f0, 32'she9bf49fa, 32'she9c23c12, 32'she9c52e38, 32'she9c8206b, 
               32'she9cb12ad, 32'she9ce04fc, 32'she9d0f758, 32'she9d3e9c3, 32'she9d6dc3b, 32'she9d9cec0, 32'she9dcc154, 32'she9dfb3f5, 
               32'she9e2a6a3, 32'she9e59960, 32'she9e88c2a, 32'she9eb7f01, 32'she9ee71e6, 32'she9f164d9, 32'she9f457da, 32'she9f74ae8, 
               32'she9fa3e03, 32'she9fd312c, 32'shea002463, 32'shea0317a7, 32'shea060af9, 32'shea08fe59, 32'shea0bf1c6, 32'shea0ee540, 
               32'shea11d8c8, 32'shea14cc5e, 32'shea17c001, 32'shea1ab3b2, 32'shea1da770, 32'shea209b3b, 32'shea238f15, 32'shea2682fb, 
               32'shea2976ef, 32'shea2c6af1, 32'shea2f5f00, 32'shea32531c, 32'shea354746, 32'shea383b7e, 32'shea3b2fc2, 32'shea3e2415, 
               32'shea411874, 32'shea440ce1, 32'shea47015c, 32'shea49f5e4, 32'shea4cea79, 32'shea4fdf1c, 32'shea52d3cc, 32'shea55c889, 
               32'shea58bd54, 32'shea5bb22c, 32'shea5ea712, 32'shea619c04, 32'shea649105, 32'shea678612, 32'shea6a7b2d, 32'shea6d7055, 
               32'shea70658a, 32'shea735acd, 32'shea76501d, 32'shea79457a, 32'shea7c3ae5, 32'shea7f305d, 32'shea8225e2, 32'shea851b74, 
               32'shea881114, 32'shea8b06c1, 32'shea8dfc7b, 32'shea90f242, 32'shea93e817, 32'shea96ddf9, 32'shea99d3e8, 32'shea9cc9e4, 
               32'shea9fbfed, 32'sheaa2b604, 32'sheaa5ac27, 32'sheaa8a258, 32'sheaab9896, 32'sheaae8ee2, 32'sheab1853a, 32'sheab47b9f, 
               32'sheab77212, 32'sheaba6892, 32'sheabd5f1f, 32'sheac055b9, 32'sheac34c60, 32'sheac64314, 32'sheac939d5, 32'sheacc30a4, 
               32'sheacf277f, 32'shead21e68, 32'shead5155d, 32'shead80c60, 32'sheadb0370, 32'sheaddfa8d, 32'sheae0f1b6, 32'sheae3e8ed, 
               32'sheae6e031, 32'sheae9d782, 32'sheaeccee0, 32'sheaefc64b, 32'sheaf2bdc3, 32'sheaf5b547, 32'sheaf8acd9, 32'sheafba478, 
               32'sheafe9c24, 32'sheb0193dd, 32'sheb048ba2, 32'sheb078375, 32'sheb0a7b54, 32'sheb0d7341, 32'sheb106b3a, 32'sheb136341, 
               32'sheb165b54, 32'sheb195374, 32'sheb1c4ba1, 32'sheb1f43db, 32'sheb223c22, 32'sheb253475, 32'sheb282cd6, 32'sheb2b2543, 
               32'sheb2e1dbe, 32'sheb311645, 32'sheb340ed9, 32'sheb370779, 32'sheb3a0027, 32'sheb3cf8e1, 32'sheb3ff1a8, 32'sheb42ea7c, 
               32'sheb45e35d, 32'sheb48dc4b, 32'sheb4bd545, 32'sheb4ece4c, 32'sheb51c760, 32'sheb54c081, 32'sheb57b9ae, 32'sheb5ab2e8, 
               32'sheb5dac2f, 32'sheb60a582, 32'sheb639ee3, 32'sheb669850, 32'sheb6991ca, 32'sheb6c8b50, 32'sheb6f84e3, 32'sheb727e83, 
               32'sheb75782f, 32'sheb7871e8, 32'sheb7b6bae, 32'sheb7e6581, 32'sheb815f60, 32'sheb84594c, 32'sheb875344, 32'sheb8a4d49, 
               32'sheb8d475b, 32'sheb904179, 32'sheb933ba4, 32'sheb9635db, 32'sheb99301f, 32'sheb9c2a70, 32'sheb9f24cd, 32'sheba21f37, 
               32'sheba519ad, 32'sheba81430, 32'shebab0ec0, 32'shebae095c, 32'shebb10404, 32'shebb3feb9, 32'shebb6f97b, 32'shebb9f449, 
               32'shebbcef23, 32'shebbfea0b, 32'shebc2e4fe, 32'shebc5dffe, 32'shebc8db0b, 32'shebcbd624, 32'shebced149, 32'shebd1cc7b, 
               32'shebd4c7ba, 32'shebd7c304, 32'shebdabe5c, 32'shebddb9bf, 32'shebe0b52f, 32'shebe3b0ac, 32'shebe6ac35, 32'shebe9a7ca, 
               32'shebeca36c, 32'shebef9f1a, 32'shebf29ad4, 32'shebf5969b, 32'shebf8926f, 32'shebfb8e4e, 32'shebfe8a3a, 32'shec018632, 
               32'shec048237, 32'shec077e48, 32'shec0a7a65, 32'shec0d768e, 32'shec1072c4, 32'shec136f06, 32'shec166b55, 32'shec1967b0, 
               32'shec1c6417, 32'shec1f608a, 32'shec225d09, 32'shec255995, 32'shec28562d, 32'shec2b52d1, 32'shec2e4f82, 32'shec314c3f, 
               32'shec344908, 32'shec3745dd, 32'shec3a42be, 32'shec3d3fac, 32'shec403ca5, 32'shec4339ab, 32'shec4636bd, 32'shec4933dc, 
               32'shec4c3106, 32'shec4f2e3d, 32'shec522b7f, 32'shec5528ce, 32'shec582629, 32'shec5b2390, 32'shec5e2103, 32'shec611e83, 
               32'shec641c0e, 32'shec6719a6, 32'shec6a1749, 32'shec6d14f9, 32'shec7012b5, 32'shec73107d, 32'shec760e51, 32'shec790c31, 
               32'shec7c0a1d, 32'shec7f0815, 32'shec820619, 32'shec850429, 32'shec880245, 32'shec8b006d, 32'shec8dfea1, 32'shec90fce1, 
               32'shec93fb2e, 32'shec96f986, 32'shec99f7ea, 32'shec9cf65a, 32'shec9ff4d6, 32'sheca2f35e, 32'sheca5f1f2, 32'sheca8f091, 
               32'shecabef3d, 32'shecaeedf5, 32'shecb1ecb8, 32'shecb4eb88, 32'shecb7ea63, 32'shecbae94b, 32'shecbde83e, 32'shecc0e73d, 
               32'shecc3e648, 32'shecc6e55f, 32'shecc9e481, 32'sheccce3b0, 32'sheccfe2ea, 32'shecd2e230, 32'shecd5e182, 32'shecd8e0e0, 
               32'shecdbe04a, 32'shecdedfbf, 32'shece1df40, 32'shece4dece, 32'shece7de66, 32'sheceade0b, 32'shecedddbb, 32'shecf0dd78, 
               32'shecf3dd3f, 32'shecf6dd13, 32'shecf9dcf3, 32'shecfcdcde, 32'shecffdcd4, 32'shed02dcd7, 32'shed05dce5, 32'shed08dcff, 
               32'shed0bdd25, 32'shed0edd56, 32'shed11dd94, 32'shed14dddc, 32'shed17de31, 32'shed1ade91, 32'shed1ddefd, 32'shed20df74, 
               32'shed23dff7, 32'shed26e086, 32'shed29e120, 32'shed2ce1c6, 32'shed2fe277, 32'shed32e334, 32'shed35e3fd, 32'shed38e4d2, 
               32'shed3be5b1, 32'shed3ee69d, 32'shed41e794, 32'shed44e897, 32'shed47e9a5, 32'shed4aeabe, 32'shed4debe4, 32'shed50ed14, 
               32'shed53ee51, 32'shed56ef99, 32'shed59f0ec, 32'shed5cf24b, 32'shed5ff3b5, 32'shed62f52b, 32'shed65f6ac, 32'shed68f839, 
               32'shed6bf9d1, 32'shed6efb75, 32'shed71fd24, 32'shed74fedf, 32'shed7800a5, 32'shed7b0276, 32'shed7e0453, 32'shed81063b, 
               32'shed84082f, 32'shed870a2e, 32'shed8a0c39, 32'shed8d0e4f, 32'shed901070, 32'shed93129d, 32'shed9614d5, 32'shed991718, 
               32'shed9c1967, 32'shed9f1bc1, 32'sheda21e26, 32'sheda52097, 32'sheda82313, 32'shedab259a, 32'shedae282d, 32'shedb12acb, 
               32'shedb42d74, 32'shedb73029, 32'shedba32e9, 32'shedbd35b4, 32'shedc0388a, 32'shedc33b6c, 32'shedc63e59, 32'shedc94151, 
               32'shedcc4454, 32'shedcf4763, 32'shedd24a7d, 32'shedd54da2, 32'shedd850d2, 32'sheddb540d, 32'shedde5754, 32'shede15aa6, 
               32'shede45e03, 32'shede7616b, 32'shedea64de, 32'sheded685d, 32'shedf06be6, 32'shedf36f7b, 32'shedf6731b, 32'shedf976c6, 
               32'shedfc7a7c, 32'shedff7e3d, 32'shee02820a, 32'shee0585e1, 32'shee0889c4, 32'shee0b8db1, 32'shee0e91aa, 32'shee1195ae, 
               32'shee1499bd, 32'shee179dd7, 32'shee1aa1fc, 32'shee1da62c, 32'shee20aa67, 32'shee23aead, 32'shee26b2fe, 32'shee29b75a, 
               32'shee2cbbc1, 32'shee2fc033, 32'shee32c4b0, 32'shee35c938, 32'shee38cdcb, 32'shee3bd269, 32'shee3ed712, 32'shee41dbc6, 
               32'shee44e084, 32'shee47e54e, 32'shee4aea23, 32'shee4def02, 32'shee50f3ed, 32'shee53f8e2, 32'shee56fde3, 32'shee5a02ee, 
               32'shee5d0804, 32'shee600d25, 32'shee631251, 32'shee661788, 32'shee691cc9, 32'shee6c2216, 32'shee6f276d, 32'shee722ccf, 
               32'shee75323c, 32'shee7837b4, 32'shee7b3d36, 32'shee7e42c4, 32'shee81485c, 32'shee844dff, 32'shee8753ad, 32'shee8a5965, 
               32'shee8d5f29, 32'shee9064f7, 32'shee936acf, 32'shee9670b3, 32'shee9976a1, 32'shee9c7c9a, 32'shee9f829e, 32'sheea288ad, 
               32'sheea58ec6, 32'sheea894ea, 32'sheeab9b18, 32'sheeaea152, 32'sheeb1a796, 32'sheeb4ade4, 32'sheeb7b43e, 32'sheebabaa2, 
               32'sheebdc110, 32'sheec0c78a, 32'sheec3ce0d, 32'sheec6d49c, 32'sheec9db35, 32'sheecce1d9, 32'sheecfe887, 32'sheed2ef40, 
               32'sheed5f604, 32'sheed8fcd2, 32'sheedc03ab, 32'sheedf0a8e, 32'sheee2117c, 32'sheee51875, 32'sheee81f78, 32'sheeeb2685, 
               32'sheeee2d9d, 32'sheef134c0, 32'sheef43bed, 32'sheef74325, 32'sheefa4a67, 32'sheefd51b4, 32'shef00590b, 32'shef03606c, 
               32'shef0667d9, 32'shef096f4f, 32'shef0c76d0, 32'shef0f7e5c, 32'shef1285f2, 32'shef158d92, 32'shef18953d, 32'shef1b9cf2, 
               32'shef1ea4b2, 32'shef21ac7c, 32'shef24b451, 32'shef27bc2f, 32'shef2ac419, 32'shef2dcc0c, 32'shef30d40a, 32'shef33dc13, 
               32'shef36e426, 32'shef39ec43, 32'shef3cf46a, 32'shef3ffc9c, 32'shef4304d8, 32'shef460d1f, 32'shef491570, 32'shef4c1dcb, 
               32'shef4f2630, 32'shef522ea0, 32'shef55371a, 32'shef583f9e, 32'shef5b482d, 32'shef5e50c6, 32'shef615969, 32'shef646216, 
               32'shef676ace, 32'shef6a738f, 32'shef6d7c5b, 32'shef708532, 32'shef738e12, 32'shef7696fd, 32'shef799ff2, 32'shef7ca8f1, 
               32'shef7fb1fa, 32'shef82bb0e, 32'shef85c42b, 32'shef88cd53, 32'shef8bd685, 32'shef8edfc1, 32'shef91e907, 32'shef94f258, 
               32'shef97fbb2, 32'shef9b0517, 32'shef9e0e85, 32'shefa117fe, 32'shefa42181, 32'shefa72b0e, 32'shefaa34a5, 32'shefad3e47, 
               32'shefb047f2, 32'shefb351a7, 32'shefb65b66, 32'shefb96530, 32'shefbc6f03, 32'shefbf78e1, 32'shefc282c8, 32'shefc58cba, 
               32'shefc896b5, 32'shefcba0bb, 32'shefceaacb, 32'shefd1b4e4, 32'shefd4bf08, 32'shefd7c935, 32'shefdad36c, 32'shefddddae, 
               32'shefe0e7f9, 32'shefe3f24f, 32'shefe6fcae, 32'shefea0717, 32'shefed118a, 32'sheff01c07, 32'sheff3268e, 32'sheff6311f, 
               32'sheff93bba, 32'sheffc465e, 32'shefff510d, 32'shf0025bc5, 32'shf0056687, 32'shf0087153, 32'shf00b7c29, 32'shf00e8709, 
               32'shf01191f3, 32'shf0149ce6, 32'shf017a7e3, 32'shf01ab2ea, 32'shf01dbdfb, 32'shf020c916, 32'shf023d43a, 32'shf026df68, 
               32'shf029eaa1, 32'shf02cf5e2, 32'shf030012e, 32'shf0330c83, 32'shf03617e2, 32'shf039234b, 32'shf03c2ebd, 32'shf03f3a3a, 
               32'shf04245c0, 32'shf045514f, 32'shf0485ce9, 32'shf04b688c, 32'shf04e7438, 32'shf0517fef, 32'shf0548baf, 32'shf0579779, 
               32'shf05aa34c, 32'shf05daf29, 32'shf060bb10, 32'shf063c700, 32'shf066d2fa, 32'shf069defe, 32'shf06ceb0b, 32'shf06ff722, 
               32'shf0730342, 32'shf0760f6c, 32'shf0791ba0, 32'shf07c27dd, 32'shf07f3424, 32'shf0824074, 32'shf0854cce, 32'shf0885932, 
               32'shf08b659f, 32'shf08e7215, 32'shf0917e95, 32'shf0948b1f, 32'shf09797b2, 32'shf09aa44e, 32'shf09db0f4, 32'shf0a0bda4, 
               32'shf0a3ca5d, 32'shf0a6d71f, 32'shf0a9e3eb, 32'shf0acf0c1, 32'shf0affda0, 32'shf0b30a88, 32'shf0b6177a, 32'shf0b92475, 
               32'shf0bc317a, 32'shf0bf3e88, 32'shf0c24b9f, 32'shf0c558c0, 32'shf0c865ea, 32'shf0cb731e, 32'shf0ce805b, 32'shf0d18da1, 
               32'shf0d49af1, 32'shf0d7a84a, 32'shf0dab5ad, 32'shf0ddc318, 32'shf0e0d08d, 32'shf0e3de0c, 32'shf0e6eb94, 32'shf0e9f925, 
               32'shf0ed06bf, 32'shf0f01463, 32'shf0f32210, 32'shf0f62fc6, 32'shf0f93d86, 32'shf0fc4b4f, 32'shf0ff5921, 32'shf10266fc, 
               32'shf10574e0, 32'shf10882ce, 32'shf10b90c5, 32'shf10e9ec6, 32'shf111accf, 32'shf114bae2, 32'shf117c8fe, 32'shf11ad723, 
               32'shf11de551, 32'shf120f389, 32'shf12401c9, 32'shf1271013, 32'shf12a1e66, 32'shf12d2cc2, 32'shf1303b27, 32'shf1334996, 
               32'shf136580d, 32'shf139668e, 32'shf13c7518, 32'shf13f83ab, 32'shf1429247, 32'shf145a0ec, 32'shf148af9a, 32'shf14bbe51, 
               32'shf14ecd11, 32'shf151dbdb, 32'shf154eaad, 32'shf157f989, 32'shf15b086d, 32'shf15e175b, 32'shf1612651, 32'shf1643551, 
               32'shf1674459, 32'shf16a536b, 32'shf16d6286, 32'shf17071a9, 32'shf17380d6, 32'shf176900b, 32'shf1799f4a, 32'shf17cae91, 
               32'shf17fbde2, 32'shf182cd3b, 32'shf185dc9d, 32'shf188ec09, 32'shf18bfb7d, 32'shf18f0afa, 32'shf1921a80, 32'shf1952a0f, 
               32'shf19839a6, 32'shf19b4947, 32'shf19e58f1, 32'shf1a168a3, 32'shf1a4785e, 32'shf1a78822, 32'shf1aa97ef, 32'shf1ada7c5, 
               32'shf1b0b7a4, 32'shf1b3c78b, 32'shf1b6d77c, 32'shf1b9e775, 32'shf1bcf777, 32'shf1c00781, 32'shf1c31795, 32'shf1c627b1, 
               32'shf1c937d6, 32'shf1cc4804, 32'shf1cf583b, 32'shf1d2687a, 32'shf1d578c2, 32'shf1d88913, 32'shf1db996d, 32'shf1dea9cf, 
               32'shf1e1ba3a, 32'shf1e4caae, 32'shf1e7db2a, 32'shf1eaebaf, 32'shf1edfc3d, 32'shf1f10cd3, 32'shf1f41d72, 32'shf1f72e1a, 
               32'shf1fa3ecb, 32'shf1fd4f84, 32'shf2006046, 32'shf2037110, 32'shf20681e3, 32'shf20992bf, 32'shf20ca3a3, 32'shf20fb490, 
               32'shf212c585, 32'shf215d683, 32'shf218e78a, 32'shf21bf899, 32'shf21f09b1, 32'shf2221ad1, 32'shf2252bfa, 32'shf2283d2c, 
               32'shf22b4e66, 32'shf22e5fa8, 32'shf23170f3, 32'shf2348247, 32'shf23793a3, 32'shf23aa507, 32'shf23db674, 32'shf240c7ea, 
               32'shf243d968, 32'shf246eaee, 32'shf249fc7d, 32'shf24d0e15, 32'shf2501fb5, 32'shf253315d, 32'shf256430e, 32'shf25954c7, 
               32'shf25c6688, 32'shf25f7852, 32'shf2628a25, 32'shf2659c00, 32'shf268ade3, 32'shf26bbfce, 32'shf26ed1c2, 32'shf271e3bf, 
               32'shf274f5c3, 32'shf27807d0, 32'shf27b19e6, 32'shf27e2c04, 32'shf2813e2a, 32'shf2845058, 32'shf287628f, 32'shf28a74ce, 
               32'shf28d8715, 32'shf2909965, 32'shf293abbd, 32'shf296be1d, 32'shf299d085, 32'shf29ce2f6, 32'shf29ff56f, 32'shf2a307f0, 
               32'shf2a61a7a, 32'shf2a92d0b, 32'shf2ac3fa5, 32'shf2af5247, 32'shf2b264f2, 32'shf2b577a4, 32'shf2b88a5f, 32'shf2bb9d22, 
               32'shf2beafed, 32'shf2c1c2c0, 32'shf2c4d59c, 32'shf2c7e880, 32'shf2cafb6b, 32'shf2ce0e5f, 32'shf2d1215b, 32'shf2d43460, 
               32'shf2d7476c, 32'shf2da5a81, 32'shf2dd6d9d, 32'shf2e080c2, 32'shf2e393ef, 32'shf2e6a723, 32'shf2e9ba60, 32'shf2eccda5, 
               32'shf2efe0f2, 32'shf2f2f448, 32'shf2f607a5, 32'shf2f91b0a, 32'shf2fc2e77, 32'shf2ff41ed, 32'shf302556a, 32'shf30568ef, 
               32'shf3087c7d, 32'shf30b9012, 32'shf30ea3af, 32'shf311b755, 32'shf314cb02, 32'shf317deb7, 32'shf31af274, 32'shf31e0639, 
               32'shf3211a07, 32'shf3242ddc, 32'shf32741b9, 32'shf32a559e, 32'shf32d698a, 32'shf3307d7f, 32'shf333917c, 32'shf336a580, 
               32'shf339b98d, 32'shf33ccda1, 32'shf33fe1bd, 32'shf342f5e1, 32'shf3460a0d, 32'shf3491e41, 32'shf34c327c, 32'shf34f46c0, 
               32'shf3525b0b, 32'shf3556f5e, 32'shf35883b9, 32'shf35b981c, 32'shf35eac86, 32'shf361c0f9, 32'shf364d573, 32'shf367e9f4, 
               32'shf36afe7e, 32'shf36e130f, 32'shf37127a9, 32'shf3743c49, 32'shf37750f2, 32'shf37a65a2, 32'shf37d7a5b, 32'shf3808f1a, 
               32'shf383a3e2, 32'shf386b8b1, 32'shf389cd88, 32'shf38ce266, 32'shf38ff74d, 32'shf3930c3b, 32'shf3962130, 32'shf399362d, 
               32'shf39c4b32, 32'shf39f603f, 32'shf3a27553, 32'shf3a58a6f, 32'shf3a89f92, 32'shf3abb4bd, 32'shf3aec9f0, 32'shf3b1df2a, 
               32'shf3b4f46c, 32'shf3b809b6, 32'shf3bb1f07, 32'shf3be345f, 32'shf3c149bf, 32'shf3c45f27, 32'shf3c77496, 32'shf3ca8a0d, 
               32'shf3cd9f8b, 32'shf3d0b511, 32'shf3d3ca9e, 32'shf3d6e033, 32'shf3d9f5cf, 32'shf3dd0b73, 32'shf3e0211f, 32'shf3e336d1, 
               32'shf3e64c8c, 32'shf3e9624d, 32'shf3ec7817, 32'shf3ef8de7, 32'shf3f2a3bf, 32'shf3f5b99f, 32'shf3f8cf86, 32'shf3fbe574, 
               32'shf3fefb6a, 32'shf4021167, 32'shf405276c, 32'shf4083d78, 32'shf40b538b, 32'shf40e69a6, 32'shf4117fc8, 32'shf41495f1, 
               32'shf417ac22, 32'shf41ac25a, 32'shf41dd89a, 32'shf420eee1, 32'shf424052f, 32'shf4271b84, 32'shf42a31e1, 32'shf42d4845, 
               32'shf4305eb0, 32'shf4337523, 32'shf4368b9d, 32'shf439a21e, 32'shf43cb8a7, 32'shf43fcf36, 32'shf442e5cd, 32'shf445fc6b, 
               32'shf4491311, 32'shf44c29be, 32'shf44f4071, 32'shf452572c, 32'shf4556def, 32'shf45884b8, 32'shf45b9b89, 32'shf45eb261, 
               32'shf461c940, 32'shf464e026, 32'shf467f713, 32'shf46b0e08, 32'shf46e2504, 32'shf4713c06, 32'shf4745310, 32'shf4776a21, 
               32'shf47a8139, 32'shf47d9859, 32'shf480af7f, 32'shf483c6ad, 32'shf486dde1, 32'shf489f51d, 32'shf48d0c5f, 32'shf49023a9, 
               32'shf4933afa, 32'shf4965252, 32'shf49969b1, 32'shf49c8117, 32'shf49f9884, 32'shf4a2aff8, 32'shf4a5c773, 32'shf4a8def5, 
               32'shf4abf67e, 32'shf4af0e0d, 32'shf4b225a4, 32'shf4b53d42, 32'shf4b854e7, 32'shf4bb6c93, 32'shf4be8446, 32'shf4c19c00, 
               32'shf4c4b3c0, 32'shf4c7cb88, 32'shf4cae356, 32'shf4cdfb2c, 32'shf4d11308, 32'shf4d42aeb, 32'shf4d742d6, 32'shf4da5ac7, 
               32'shf4dd72be, 32'shf4e08abd, 32'shf4e3a2c3, 32'shf4e6bacf, 32'shf4e9d2e3, 32'shf4eceafd, 32'shf4f0031e, 32'shf4f31b46, 
               32'shf4f63374, 32'shf4f94baa, 32'shf4fc63e6, 32'shf4ff7c29, 32'shf5029473, 32'shf505acc3, 32'shf508c51b, 32'shf50bdd79, 
               32'shf50ef5de, 32'shf5120e49, 32'shf51526bc, 32'shf5183f35, 32'shf51b57b5, 32'shf51e703b, 32'shf52188c9, 32'shf524a15d, 
               32'shf527b9f7, 32'shf52ad299, 32'shf52deb41, 32'shf53103ef, 32'shf5341ca5, 32'shf5373561, 32'shf53a4e24, 32'shf53d66ed, 
               32'shf5407fbd, 32'shf5439893, 32'shf546b171, 32'shf549ca55, 32'shf54ce33f, 32'shf54ffc30, 32'shf5531528, 32'shf5562e26, 
               32'shf559472b, 32'shf55c6036, 32'shf55f7948, 32'shf5629261, 32'shf565ab80, 32'shf568c4a5, 32'shf56bddd1, 32'shf56ef704, 
               32'shf572103d, 32'shf575297d, 32'shf57842c3, 32'shf57b5c10, 32'shf57e7563, 32'shf5818ebd, 32'shf584a81d, 32'shf587c183, 
               32'shf58adaf0, 32'shf58df464, 32'shf5910dde, 32'shf594275e, 32'shf59740e5, 32'shf59a5a72, 32'shf59d7406, 32'shf5a08da0, 
               32'shf5a3a740, 32'shf5a6c0e7, 32'shf5a9da94, 32'shf5acf448, 32'shf5b00e02, 32'shf5b327c2, 32'shf5b64189, 32'shf5b95b56, 
               32'shf5bc7529, 32'shf5bf8f03, 32'shf5c2a8e3, 32'shf5c5c2c9, 32'shf5c8dcb6, 32'shf5cbf6a9, 32'shf5cf10a2, 32'shf5d22aa2, 
               32'shf5d544a7, 32'shf5d85eb3, 32'shf5db78c6, 32'shf5de92de, 32'shf5e1acfd, 32'shf5e4c722, 32'shf5e7e14e, 32'shf5eafb7f, 
               32'shf5ee15b7, 32'shf5f12ff5, 32'shf5f44a39, 32'shf5f76484, 32'shf5fa7ed4, 32'shf5fd992b, 32'shf600b388, 32'shf603cdeb, 
               32'shf606e854, 32'shf60a02c3, 32'shf60d1d39, 32'shf61037b5, 32'shf6135237, 32'shf6166cbe, 32'shf619874c, 32'shf61ca1e1, 
               32'shf61fbc7b, 32'shf622d71b, 32'shf625f1c2, 32'shf6290c6e, 32'shf62c2721, 32'shf62f41d9, 32'shf6325c98, 32'shf635775d, 
               32'shf6389228, 32'shf63bacf8, 32'shf63ec7cf, 32'shf641e2ac, 32'shf644fd8f, 32'shf6481878, 32'shf64b3367, 32'shf64e4e5c, 
               32'shf6516956, 32'shf6548457, 32'shf6579f5e, 32'shf65aba6b, 32'shf65dd57d, 32'shf660f096, 32'shf6640bb4, 32'shf66726d9, 
               32'shf66a4203, 32'shf66d5d34, 32'shf670786a, 32'shf67393a6, 32'shf676aee8, 32'shf679ca30, 32'shf67ce57e, 32'shf68000d1, 
               32'shf6831c2b, 32'shf686378a, 32'shf68952ef, 32'shf68c6e5a, 32'shf68f89cb, 32'shf692a542, 32'shf695c0be, 32'shf698dc41, 
               32'shf69bf7c9, 32'shf69f1357, 32'shf6a22eea, 32'shf6a54a84, 32'shf6a86623, 32'shf6ab81c8, 32'shf6ae9d73, 32'shf6b1b923, 
               32'shf6b4d4d9, 32'shf6b7f095, 32'shf6bb0c57, 32'shf6be281e, 32'shf6c143ec, 32'shf6c45fbe, 32'shf6c77b97, 32'shf6ca9775, 
               32'shf6cdb359, 32'shf6d0cf43, 32'shf6d3eb32, 32'shf6d70727, 32'shf6da2321, 32'shf6dd3f21, 32'shf6e05b27, 32'shf6e37733, 
               32'shf6e69344, 32'shf6e9af5a, 32'shf6eccb77, 32'shf6efe798, 32'shf6f303c0, 32'shf6f61fed, 32'shf6f93c20, 32'shf6fc5858, 
               32'shf6ff7496, 32'shf70290d9, 32'shf705ad22, 32'shf708c970, 32'shf70be5c4, 32'shf70f021d, 32'shf7121e7c, 32'shf7153ae1, 
               32'shf718574b, 32'shf71b73ba, 32'shf71e902f, 32'shf721acaa, 32'shf724c92a, 32'shf727e5af, 32'shf72b023a, 32'shf72e1eca, 
               32'shf7313b60, 32'shf73457fb, 32'shf737749b, 32'shf73a9141, 32'shf73daded, 32'shf740ca9d, 32'shf743e754, 32'shf747040f, 
               32'shf74a20d0, 32'shf74d3d96, 32'shf7505a62, 32'shf7537733, 32'shf756940a, 32'shf759b0e5, 32'shf75ccdc6, 32'shf75feaad, 
               32'shf7630799, 32'shf766248a, 32'shf7694180, 32'shf76c5e7c, 32'shf76f7b7d, 32'shf7729883, 32'shf775b58e, 32'shf778d29f, 
               32'shf77befb5, 32'shf77f0cd0, 32'shf78229f1, 32'shf7854717, 32'shf7886442, 32'shf78b8172, 32'shf78e9ea7, 32'shf791bbe2, 
               32'shf794d922, 32'shf797f667, 32'shf79b13b1, 32'shf79e3100, 32'shf7a14e55, 32'shf7a46baf, 32'shf7a7890d, 32'shf7aaa671, 
               32'shf7adc3db, 32'shf7b0e149, 32'shf7b3febc, 32'shf7b71c35, 32'shf7ba39b3, 32'shf7bd5735, 32'shf7c074bd, 32'shf7c3924a, 
               32'shf7c6afdc, 32'shf7c9cd73, 32'shf7cceb0f, 32'shf7d008b1, 32'shf7d32657, 32'shf7d64402, 32'shf7d961b3, 32'shf7dc7f68, 
               32'shf7df9d22, 32'shf7e2bae2, 32'shf7e5d8a6, 32'shf7e8f670, 32'shf7ec143e, 32'shf7ef3211, 32'shf7f24fea, 32'shf7f56dc7, 
               32'shf7f88ba9, 32'shf7fba991, 32'shf7fec77d, 32'shf801e56e, 32'shf8050364, 32'shf808215f, 32'shf80b3f5f, 32'shf80e5d64, 
               32'shf8117b6d, 32'shf814997c, 32'shf817b78f, 32'shf81ad5a8, 32'shf81df3c5, 32'shf82111e7, 32'shf824300e, 32'shf8274e3a, 
               32'shf82a6c6a, 32'shf82d8aa0, 32'shf830a8da, 32'shf833c719, 32'shf836e55d, 32'shf83a03a6, 32'shf83d21f3, 32'shf8404046, 
               32'shf8435e9d, 32'shf8467cf9, 32'shf8499b59, 32'shf84cb9bf, 32'shf84fd829, 32'shf852f698, 32'shf856150b, 32'shf8593383, 
               32'shf85c5201, 32'shf85f7082, 32'shf8628f09, 32'shf865ad94, 32'shf868cc24, 32'shf86beab8, 32'shf86f0952, 32'shf87227ef, 
               32'shf8754692, 32'shf8786539, 32'shf87b83e5, 32'shf87ea295, 32'shf881c14b, 32'shf884e004, 32'shf887fec3, 32'shf88b1d86, 
               32'shf88e3c4d, 32'shf8915b19, 32'shf89479ea, 32'shf89798bf, 32'shf89ab799, 32'shf89dd678, 32'shf8a0f55b, 32'shf8a41442, 
               32'shf8a7332e, 32'shf8aa521f, 32'shf8ad7114, 32'shf8b0900d, 32'shf8b3af0c, 32'shf8b6ce0e, 32'shf8b9ed15, 32'shf8bd0c21, 
               32'shf8c02b31, 32'shf8c34a46, 32'shf8c6695f, 32'shf8c9887c, 32'shf8cca79e, 32'shf8cfc6c5, 32'shf8d2e5f0, 32'shf8d6051f, 
               32'shf8d92452, 32'shf8dc438b, 32'shf8df62c7, 32'shf8e28208, 32'shf8e5a14d, 32'shf8e8c097, 32'shf8ebdfe5, 32'shf8eeff37, 
               32'shf8f21e8e, 32'shf8f53de9, 32'shf8f85d49, 32'shf8fb7cac, 32'shf8fe9c15, 32'shf901bb81, 32'shf904daf2, 32'shf907fa67, 
               32'shf90b19e0, 32'shf90e395e, 32'shf91158e0, 32'shf9147866, 32'shf91797f0, 32'shf91ab77f, 32'shf91dd712, 32'shf920f6a9, 
               32'shf9241645, 32'shf92735e5, 32'shf92a5589, 32'shf92d7531, 32'shf93094dd, 32'shf933b48e, 32'shf936d442, 32'shf939f3fb, 
               32'shf93d13b8, 32'shf940337a, 32'shf943533f, 32'shf9467309, 32'shf94992d7, 32'shf94cb2a8, 32'shf94fd27f, 32'shf952f259, 
               32'shf9561237, 32'shf9593219, 32'shf95c5200, 32'shf95f71ea, 32'shf96291d9, 32'shf965b1cc, 32'shf968d1c3, 32'shf96bf1be, 
               32'shf96f11bc, 32'shf97231bf, 32'shf97551c6, 32'shf97871d2, 32'shf97b91e1, 32'shf97eb1f4, 32'shf981d20b, 32'shf984f226, 
               32'shf9881245, 32'shf98b3268, 32'shf98e528f, 32'shf99172bb, 32'shf99492ea, 32'shf997b31d, 32'shf99ad354, 32'shf99df38e, 
               32'shf9a113cd, 32'shf9a43410, 32'shf9a75457, 32'shf9aa74a1, 32'shf9ad94f0, 32'shf9b0b542, 32'shf9b3d599, 32'shf9b6f5f3, 
               32'shf9ba1651, 32'shf9bd36b3, 32'shf9c05719, 32'shf9c37782, 32'shf9c697f0, 32'shf9c9b861, 32'shf9ccd8d6, 32'shf9cff94f, 
               32'shf9d319cc, 32'shf9d63a4d, 32'shf9d95ad1, 32'shf9dc7b5a, 32'shf9df9be6, 32'shf9e2bc75, 32'shf9e5dd09, 32'shf9e8fda0, 
               32'shf9ec1e3b, 32'shf9ef3eda, 32'shf9f25f7d, 32'shf9f58023, 32'shf9f8a0cd, 32'shf9fbc17b, 32'shf9fee22c, 32'shfa0202e1, 
               32'shfa05239a, 32'shfa084457, 32'shfa0b6517, 32'shfa0e85db, 32'shfa11a6a3, 32'shfa14c76e, 32'shfa17e83d, 32'shfa1b090f, 
               32'shfa1e29e5, 32'shfa214abf, 32'shfa246b9d, 32'shfa278c7e, 32'shfa2aad62, 32'shfa2dce4b, 32'shfa30ef36, 32'shfa341026, 
               32'shfa373119, 32'shfa3a520f, 32'shfa3d7309, 32'shfa409407, 32'shfa43b508, 32'shfa46d60d, 32'shfa49f715, 32'shfa4d1821, 
               32'shfa503930, 32'shfa535a43, 32'shfa567b5a, 32'shfa599c73, 32'shfa5cbd91, 32'shfa5fdeb1, 32'shfa62ffd6, 32'shfa6620fd, 
               32'shfa694229, 32'shfa6c6357, 32'shfa6f8489, 32'shfa72a5bf, 32'shfa75c6f8, 32'shfa78e834, 32'shfa7c0974, 32'shfa7f2ab7, 
               32'shfa824bfd, 32'shfa856d47, 32'shfa888e95, 32'shfa8bafe5, 32'shfa8ed139, 32'shfa91f291, 32'shfa9513eb, 32'shfa98354a, 
               32'shfa9b56ab, 32'shfa9e7810, 32'shfaa19978, 32'shfaa4bae3, 32'shfaa7dc52, 32'shfaaafdc4, 32'shfaae1f39, 32'shfab140b2, 
               32'shfab4622d, 32'shfab783ad, 32'shfabaa52f, 32'shfabdc6b4, 32'shfac0e83d, 32'shfac409c9, 32'shfac72b59, 32'shfaca4ceb, 
               32'shfacd6e81, 32'shfad0901a, 32'shfad3b1b6, 32'shfad6d355, 32'shfad9f4f8, 32'shfadd169e, 32'shfae03847, 32'shfae359f3, 
               32'shfae67ba2, 32'shfae99d54, 32'shfaecbf0a, 32'shfaefe0c2, 32'shfaf3027e, 32'shfaf6243d, 32'shfaf945ff, 32'shfafc67c4, 
               32'shfaff898c, 32'shfb02ab57, 32'shfb05cd25, 32'shfb08eef7, 32'shfb0c10cb, 32'shfb0f32a3, 32'shfb12547d, 32'shfb15765b, 
               32'shfb18983b, 32'shfb1bba1f, 32'shfb1edc06, 32'shfb21fdef, 32'shfb251fdc, 32'shfb2841cc, 32'shfb2b63be, 32'shfb2e85b4, 
               32'shfb31a7ac, 32'shfb34c9a8, 32'shfb37eba7, 32'shfb3b0da8, 32'shfb3e2fac, 32'shfb4151b4, 32'shfb4473be, 32'shfb4795cb, 
               32'shfb4ab7db, 32'shfb4dd9ee, 32'shfb50fc04, 32'shfb541e1d, 32'shfb574039, 32'shfb5a6257, 32'shfb5d8479, 32'shfb60a69d, 
               32'shfb63c8c4, 32'shfb66eaee, 32'shfb6a0d1b, 32'shfb6d2f4a, 32'shfb70517d, 32'shfb7373b2, 32'shfb7695ea, 32'shfb79b825, 
               32'shfb7cda63, 32'shfb7ffca3, 32'shfb831ee6, 32'shfb86412c, 32'shfb896375, 32'shfb8c85c1, 32'shfb8fa80f, 32'shfb92ca60, 
               32'shfb95ecb4, 32'shfb990f0a, 32'shfb9c3163, 32'shfb9f53bf, 32'shfba2761e, 32'shfba5987f, 32'shfba8bae3, 32'shfbabdd49, 
               32'shfbaeffb3, 32'shfbb2221f, 32'shfbb5448d, 32'shfbb866ff, 32'shfbbb8973, 32'shfbbeabe9, 32'shfbc1ce62, 32'shfbc4f0de, 
               32'shfbc8135c, 32'shfbcb35dd, 32'shfbce5861, 32'shfbd17ae7, 32'shfbd49d70, 32'shfbd7bffb, 32'shfbdae289, 32'shfbde0519, 
               32'shfbe127ac, 32'shfbe44a42, 32'shfbe76cda, 32'shfbea8f75, 32'shfbedb212, 32'shfbf0d4b1, 32'shfbf3f753, 32'shfbf719f8, 
               32'shfbfa3c9f, 32'shfbfd5f49, 32'shfc0081f5, 32'shfc03a4a3, 32'shfc06c754, 32'shfc09ea08, 32'shfc0d0cbe, 32'shfc102f76, 
               32'shfc135231, 32'shfc1674ee, 32'shfc1997ae, 32'shfc1cba6f, 32'shfc1fdd34, 32'shfc22fffb, 32'shfc2622c4, 32'shfc29458f, 
               32'shfc2c685d, 32'shfc2f8b2e, 32'shfc32ae00, 32'shfc35d0d5, 32'shfc38f3ac, 32'shfc3c1686, 32'shfc3f3962, 32'shfc425c40, 
               32'shfc457f21, 32'shfc48a204, 32'shfc4bc4e9, 32'shfc4ee7d0, 32'shfc520aba, 32'shfc552da6, 32'shfc585094, 32'shfc5b7385, 
               32'shfc5e9678, 32'shfc61b96d, 32'shfc64dc64, 32'shfc67ff5d, 32'shfc6b2259, 32'shfc6e4557, 32'shfc716857, 32'shfc748b59, 
               32'shfc77ae5e, 32'shfc7ad164, 32'shfc7df46d, 32'shfc811778, 32'shfc843a85, 32'shfc875d95, 32'shfc8a80a6, 32'shfc8da3ba, 
               32'shfc90c6cf, 32'shfc93e9e7, 32'shfc970d01, 32'shfc9a301d, 32'shfc9d533b, 32'shfca0765b, 32'shfca3997e, 32'shfca6bca2, 
               32'shfca9dfc8, 32'shfcad02f1, 32'shfcb0261b, 32'shfcb34948, 32'shfcb66c77, 32'shfcb98fa7, 32'shfcbcb2da, 32'shfcbfd60e, 
               32'shfcc2f945, 32'shfcc61c7e, 32'shfcc93fb9, 32'shfccc62f5, 32'shfccf8634, 32'shfcd2a974, 32'shfcd5ccb7, 32'shfcd8effb, 
               32'shfcdc1342, 32'shfcdf368a, 32'shfce259d5, 32'shfce57d21, 32'shfce8a06f, 32'shfcebc3bf, 32'shfceee711, 32'shfcf20a65, 
               32'shfcf52dbb, 32'shfcf85112, 32'shfcfb746c, 32'shfcfe97c7, 32'shfd01bb24, 32'shfd04de83, 32'shfd0801e4, 32'shfd0b2547, 
               32'shfd0e48ab, 32'shfd116c12, 32'shfd148f7a, 32'shfd17b2e4, 32'shfd1ad650, 32'shfd1df9bd, 32'shfd211d2c, 32'shfd24409d, 
               32'shfd276410, 32'shfd2a8785, 32'shfd2daafb, 32'shfd30ce73, 32'shfd33f1ed, 32'shfd371569, 32'shfd3a38e6, 32'shfd3d5c65, 
               32'shfd407fe6, 32'shfd43a368, 32'shfd46c6ec, 32'shfd49ea72, 32'shfd4d0df9, 32'shfd503182, 32'shfd53550d, 32'shfd56789a, 
               32'shfd599c28, 32'shfd5cbfb7, 32'shfd5fe348, 32'shfd6306db, 32'shfd662a70, 32'shfd694e06, 32'shfd6c719e, 32'shfd6f9537, 
               32'shfd72b8d2, 32'shfd75dc6e, 32'shfd79000d, 32'shfd7c23ac, 32'shfd7f474d, 32'shfd826af0, 32'shfd858e94, 32'shfd88b23a, 
               32'shfd8bd5e1, 32'shfd8ef98a, 32'shfd921d34, 32'shfd9540e0, 32'shfd98648d, 32'shfd9b883c, 32'shfd9eabec, 32'shfda1cf9e, 
               32'shfda4f351, 32'shfda81706, 32'shfdab3abc, 32'shfdae5e74, 32'shfdb1822c, 32'shfdb4a5e7, 32'shfdb7c9a3, 32'shfdbaed60, 
               32'shfdbe111e, 32'shfdc134de, 32'shfdc458a0, 32'shfdc77c62, 32'shfdcaa027, 32'shfdcdc3ec, 32'shfdd0e7b3, 32'shfdd40b7b, 
               32'shfdd72f45, 32'shfdda530f, 32'shfddd76dc, 32'shfde09aa9, 32'shfde3be78, 32'shfde6e248, 32'shfdea0619, 32'shfded29ec, 
               32'shfdf04dc0, 32'shfdf37195, 32'shfdf6956c, 32'shfdf9b944, 32'shfdfcdd1d, 32'shfe0000f7, 32'shfe0324d2, 32'shfe0648af, 
               32'shfe096c8d, 32'shfe0c906c, 32'shfe0fb44c, 32'shfe12d82e, 32'shfe15fc11, 32'shfe191ff5, 32'shfe1c43da, 32'shfe1f67c0, 
               32'shfe228ba7, 32'shfe25af90, 32'shfe28d379, 32'shfe2bf764, 32'shfe2f1b50, 32'shfe323f3d, 32'shfe35632c, 32'shfe38871b, 
               32'shfe3bab0b, 32'shfe3ecefd, 32'shfe41f2ef, 32'shfe4516e3, 32'shfe483ad8, 32'shfe4b5ecd, 32'shfe4e82c4, 32'shfe51a6bc, 
               32'shfe54cab5, 32'shfe57eeaf, 32'shfe5b12aa, 32'shfe5e36a6, 32'shfe615aa3, 32'shfe647ea1, 32'shfe67a2a0, 32'shfe6ac6a0, 
               32'shfe6deaa1, 32'shfe710ea2, 32'shfe7432a5, 32'shfe7756a9, 32'shfe7a7aae, 32'shfe7d9eb4, 32'shfe80c2ba, 32'shfe83e6c2, 
               32'shfe870aca, 32'shfe8a2ed4, 32'shfe8d52de, 32'shfe9076e9, 32'shfe939af5, 32'shfe96bf02, 32'shfe99e310, 32'shfe9d071e, 
               32'shfea02b2e, 32'shfea34f3e, 32'shfea6734f, 32'shfea99761, 32'shfeacbb74, 32'shfeafdf88, 32'shfeb3039d, 32'shfeb627b2, 
               32'shfeb94bc8, 32'shfebc6fdf, 32'shfebf93f6, 32'shfec2b80f, 32'shfec5dc28, 32'shfec90042, 32'shfecc245d, 32'shfecf4878, 
               32'shfed26c94, 32'shfed590b1, 32'shfed8b4cf, 32'shfedbd8ed, 32'shfedefd0c, 32'shfee2212c, 32'shfee5454c, 32'shfee8696d, 
               32'shfeeb8d8f, 32'shfeeeb1b2, 32'shfef1d5d5, 32'shfef4f9f8, 32'shfef81e1d, 32'shfefb4242, 32'shfefe6668, 32'shff018a8e, 
               32'shff04aeb5, 32'shff07d2dc, 32'shff0af704, 32'shff0e1b2d, 32'shff113f56, 32'shff146380, 32'shff1787aa, 32'shff1aabd5, 
               32'shff1dd001, 32'shff20f42d, 32'shff24185a, 32'shff273c87, 32'shff2a60b4, 32'shff2d84e3, 32'shff30a911, 32'shff33cd40, 
               32'shff36f170, 32'shff3a15a0, 32'shff3d39d1, 32'shff405e02, 32'shff438234, 32'shff46a666, 32'shff49ca98, 32'shff4ceecb, 
               32'shff5012fe, 32'shff533732, 32'shff565b66, 32'shff597f9b, 32'shff5ca3d0, 32'shff5fc805, 32'shff62ec3b, 32'shff661071, 
               32'shff6934a8, 32'shff6c58de, 32'shff6f7d16, 32'shff72a14d, 32'shff75c585, 32'shff78e9bd, 32'shff7c0df6, 32'shff7f322f, 
               32'shff825668, 32'shff857aa2, 32'shff889edb, 32'shff8bc316, 32'shff8ee750, 32'shff920b8b, 32'shff952fc5, 32'shff985401, 
               32'shff9b783c, 32'shff9e9c78, 32'shffa1c0b4, 32'shffa4e4f0, 32'shffa8092c, 32'shffab2d69, 32'shffae51a5, 32'shffb175e2, 
               32'shffb49a1f, 32'shffb7be5d, 32'shffbae29a, 32'shffbe06d8, 32'shffc12b16, 32'shffc44f54, 32'shffc77392, 32'shffca97d0, 
               32'shffcdbc0f, 32'shffd0e04d, 32'shffd4048c, 32'shffd728ca, 32'shffda4d09, 32'shffdd7148, 32'shffe09587, 32'shffe3b9c6, 
               32'shffe6de05, 32'shffea0245, 32'shffed2684, 32'shfff04ac3, 32'shfff36f02, 32'shfff69342, 32'shfff9b781, 32'shfffcdbc1
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
      else if (POW == 16)
         begin
            reg signed [31:0] W_Re_table[32768] = '{
               32'sh40000000, 32'sh3ffffffb, 32'sh3fffffec, 32'sh3fffffd4, 32'sh3fffffb1, 32'sh3fffff85, 32'sh3fffff4e, 32'sh3fffff0e, 
               32'sh3ffffec4, 32'sh3ffffe70, 32'sh3ffffe13, 32'sh3ffffdab, 32'sh3ffffd39, 32'sh3ffffcbe, 32'sh3ffffc39, 32'sh3ffffbaa, 
               32'sh3ffffb11, 32'sh3ffffa6e, 32'sh3ffff9c1, 32'sh3ffff90b, 32'sh3ffff84a, 32'sh3ffff780, 32'sh3ffff6ac, 32'sh3ffff5cd, 
               32'sh3ffff4e6, 32'sh3ffff3f4, 32'sh3ffff2f8, 32'sh3ffff1f3, 32'sh3ffff0e3, 32'sh3fffefca, 32'sh3fffeea7, 32'sh3fffed7a, 
               32'sh3fffec43, 32'sh3fffeb02, 32'sh3fffe9b7, 32'sh3fffe863, 32'sh3fffe705, 32'sh3fffe59c, 32'sh3fffe42a, 32'sh3fffe2ae, 
               32'sh3fffe128, 32'sh3fffdf99, 32'sh3fffddff, 32'sh3fffdc5c, 32'sh3fffdaae, 32'sh3fffd8f7, 32'sh3fffd736, 32'sh3fffd56b, 
               32'sh3fffd396, 32'sh3fffd1b8, 32'sh3fffcfcf, 32'sh3fffcddd, 32'sh3fffcbe0, 32'sh3fffc9da, 32'sh3fffc7ca, 32'sh3fffc5b0, 
               32'sh3fffc38c, 32'sh3fffc15f, 32'sh3fffbf27, 32'sh3fffbce6, 32'sh3fffba9b, 32'sh3fffb846, 32'sh3fffb5e7, 32'sh3fffb37e, 
               32'sh3fffb10b, 32'sh3fffae8f, 32'sh3fffac08, 32'sh3fffa978, 32'sh3fffa6de, 32'sh3fffa439, 32'sh3fffa18c, 32'sh3fff9ed4, 
               32'sh3fff9c12, 32'sh3fff9947, 32'sh3fff9671, 32'sh3fff9392, 32'sh3fff90a9, 32'sh3fff8db6, 32'sh3fff8ab9, 32'sh3fff87b2, 
               32'sh3fff84a1, 32'sh3fff8187, 32'sh3fff7e63, 32'sh3fff7b34, 32'sh3fff77fc, 32'sh3fff74ba, 32'sh3fff716e, 32'sh3fff6e19, 
               32'sh3fff6ab9, 32'sh3fff6750, 32'sh3fff63dc, 32'sh3fff605f, 32'sh3fff5cd8, 32'sh3fff5947, 32'sh3fff55ac, 32'sh3fff5208, 
               32'sh3fff4e59, 32'sh3fff4aa1, 32'sh3fff46df, 32'sh3fff4312, 32'sh3fff3f3c, 32'sh3fff3b5c, 32'sh3fff3773, 32'sh3fff337f, 
               32'sh3fff2f82, 32'sh3fff2b7a, 32'sh3fff2769, 32'sh3fff234e, 32'sh3fff1f29, 32'sh3fff1afa, 32'sh3fff16c1, 32'sh3fff127f, 
               32'sh3fff0e32, 32'sh3fff09dc, 32'sh3fff057c, 32'sh3fff0112, 32'sh3ffefc9e, 32'sh3ffef820, 32'sh3ffef399, 32'sh3ffeef07, 
               32'sh3ffeea6c, 32'sh3ffee5c6, 32'sh3ffee117, 32'sh3ffedc5e, 32'sh3ffed79b, 32'sh3ffed2cf, 32'sh3ffecdf8, 32'sh3ffec918, 
               32'sh3ffec42d, 32'sh3ffebf39, 32'sh3ffeba3b, 32'sh3ffeb533, 32'sh3ffeb021, 32'sh3ffeab05, 32'sh3ffea5e0, 32'sh3ffea0b0, 
               32'sh3ffe9b77, 32'sh3ffe9634, 32'sh3ffe90e7, 32'sh3ffe8b90, 32'sh3ffe862f, 32'sh3ffe80c5, 32'sh3ffe7b50, 32'sh3ffe75d2, 
               32'sh3ffe704a, 32'sh3ffe6ab7, 32'sh3ffe651b, 32'sh3ffe5f76, 32'sh3ffe59c6, 32'sh3ffe540c, 32'sh3ffe4e49, 32'sh3ffe487c, 
               32'sh3ffe42a4, 32'sh3ffe3cc3, 32'sh3ffe36d8, 32'sh3ffe30e4, 32'sh3ffe2ae5, 32'sh3ffe24dc, 32'sh3ffe1eca, 32'sh3ffe18ae, 
               32'sh3ffe1288, 32'sh3ffe0c58, 32'sh3ffe061e, 32'sh3ffdffda, 32'sh3ffdf98c, 32'sh3ffdf335, 32'sh3ffdecd3, 32'sh3ffde668, 
               32'sh3ffddff3, 32'sh3ffdd974, 32'sh3ffdd2eb, 32'sh3ffdcc59, 32'sh3ffdc5bc, 32'sh3ffdbf16, 32'sh3ffdb865, 32'sh3ffdb1ab, 
               32'sh3ffdaae7, 32'sh3ffda419, 32'sh3ffd9d42, 32'sh3ffd9660, 32'sh3ffd8f74, 32'sh3ffd887f, 32'sh3ffd8180, 32'sh3ffd7a77, 
               32'sh3ffd7364, 32'sh3ffd6c47, 32'sh3ffd6520, 32'sh3ffd5df0, 32'sh3ffd56b5, 32'sh3ffd4f71, 32'sh3ffd4823, 32'sh3ffd40cb, 
               32'sh3ffd3969, 32'sh3ffd31fd, 32'sh3ffd2a87, 32'sh3ffd2308, 32'sh3ffd1b7e, 32'sh3ffd13eb, 32'sh3ffd0c4e, 32'sh3ffd04a7, 
               32'sh3ffcfcf6, 32'sh3ffcf53b, 32'sh3ffced77, 32'sh3ffce5a8, 32'sh3ffcddd0, 32'sh3ffcd5ee, 32'sh3ffcce02, 32'sh3ffcc60c, 
               32'sh3ffcbe0c, 32'sh3ffcb602, 32'sh3ffcadef, 32'sh3ffca5d1, 32'sh3ffc9daa, 32'sh3ffc9579, 32'sh3ffc8d3e, 32'sh3ffc84f9, 
               32'sh3ffc7caa, 32'sh3ffc7451, 32'sh3ffc6bef, 32'sh3ffc6383, 32'sh3ffc5b0c, 32'sh3ffc528c, 32'sh3ffc4a02, 32'sh3ffc416f, 
               32'sh3ffc38d1, 32'sh3ffc3029, 32'sh3ffc2778, 32'sh3ffc1ebd, 32'sh3ffc15f7, 32'sh3ffc0d28, 32'sh3ffc0450, 32'sh3ffbfb6d, 
               32'sh3ffbf280, 32'sh3ffbe98a, 32'sh3ffbe089, 32'sh3ffbd77f, 32'sh3ffbce6b, 32'sh3ffbc54d, 32'sh3ffbbc25, 32'sh3ffbb2f3, 
               32'sh3ffba9b8, 32'sh3ffba073, 32'sh3ffb9723, 32'sh3ffb8dca, 32'sh3ffb8467, 32'sh3ffb7afa, 32'sh3ffb7183, 32'sh3ffb6803, 
               32'sh3ffb5e78, 32'sh3ffb54e4, 32'sh3ffb4b46, 32'sh3ffb419e, 32'sh3ffb37ec, 32'sh3ffb2e30, 32'sh3ffb246a, 32'sh3ffb1a9a, 
               32'sh3ffb10c1, 32'sh3ffb06de, 32'sh3ffafcf1, 32'sh3ffaf2fa, 32'sh3ffae8f9, 32'sh3ffadeee, 32'sh3ffad4d9, 32'sh3ffacabb, 
               32'sh3ffac092, 32'sh3ffab660, 32'sh3ffaac24, 32'sh3ffaa1de, 32'sh3ffa978e, 32'sh3ffa8d35, 32'sh3ffa82d1, 32'sh3ffa7864, 
               32'sh3ffa6dec, 32'sh3ffa636b, 32'sh3ffa58e0, 32'sh3ffa4e4b, 32'sh3ffa43ac, 32'sh3ffa3904, 32'sh3ffa2e51, 32'sh3ffa2395, 
               32'sh3ffa18cf, 32'sh3ffa0dff, 32'sh3ffa0325, 32'sh3ff9f841, 32'sh3ff9ed53, 32'sh3ff9e25c, 32'sh3ff9d75a, 32'sh3ff9cc4f, 
               32'sh3ff9c13a, 32'sh3ff9b61b, 32'sh3ff9aaf2, 32'sh3ff99fbf, 32'sh3ff99483, 32'sh3ff9893c, 32'sh3ff97dec, 32'sh3ff97291, 
               32'sh3ff9672d, 32'sh3ff95bbf, 32'sh3ff95048, 32'sh3ff944c6, 32'sh3ff9393a, 32'sh3ff92da5, 32'sh3ff92206, 32'sh3ff9165d, 
               32'sh3ff90aaa, 32'sh3ff8feed, 32'sh3ff8f326, 32'sh3ff8e755, 32'sh3ff8db7b, 32'sh3ff8cf97, 32'sh3ff8c3a8, 32'sh3ff8b7b0, 
               32'sh3ff8abae, 32'sh3ff89fa3, 32'sh3ff8938d, 32'sh3ff8876d, 32'sh3ff87b44, 32'sh3ff86f11, 32'sh3ff862d4, 32'sh3ff8568d, 
               32'sh3ff84a3c, 32'sh3ff83de1, 32'sh3ff8317d, 32'sh3ff8250e, 32'sh3ff81896, 32'sh3ff80c14, 32'sh3ff7ff88, 32'sh3ff7f2f2, 
               32'sh3ff7e652, 32'sh3ff7d9a8, 32'sh3ff7ccf5, 32'sh3ff7c038, 32'sh3ff7b370, 32'sh3ff7a69f, 32'sh3ff799c4, 32'sh3ff78cdf, 
               32'sh3ff77ff1, 32'sh3ff772f8, 32'sh3ff765f6, 32'sh3ff758ea, 32'sh3ff74bd3, 32'sh3ff73eb3, 32'sh3ff7318a, 32'sh3ff72456, 
               32'sh3ff71718, 32'sh3ff709d1, 32'sh3ff6fc7f, 32'sh3ff6ef24, 32'sh3ff6e1bf, 32'sh3ff6d450, 32'sh3ff6c6d7, 32'sh3ff6b955, 
               32'sh3ff6abc8, 32'sh3ff69e32, 32'sh3ff69092, 32'sh3ff682e8, 32'sh3ff67534, 32'sh3ff66776, 32'sh3ff659ae, 32'sh3ff64bdd, 
               32'sh3ff63e01, 32'sh3ff6301c, 32'sh3ff6222d, 32'sh3ff61434, 32'sh3ff60631, 32'sh3ff5f824, 32'sh3ff5ea0d, 32'sh3ff5dbed, 
               32'sh3ff5cdc3, 32'sh3ff5bf8e, 32'sh3ff5b150, 32'sh3ff5a308, 32'sh3ff594b7, 32'sh3ff5865b, 32'sh3ff577f6, 32'sh3ff56986, 
               32'sh3ff55b0d, 32'sh3ff54c8a, 32'sh3ff53dfd, 32'sh3ff52f66, 32'sh3ff520c5, 32'sh3ff5121b, 32'sh3ff50366, 32'sh3ff4f4a8, 
               32'sh3ff4e5e0, 32'sh3ff4d70e, 32'sh3ff4c832, 32'sh3ff4b94c, 32'sh3ff4aa5d, 32'sh3ff49b63, 32'sh3ff48c60, 32'sh3ff47d53, 
               32'sh3ff46e3c, 32'sh3ff45f1b, 32'sh3ff44ff0, 32'sh3ff440bc, 32'sh3ff4317d, 32'sh3ff42235, 32'sh3ff412e2, 32'sh3ff40386, 
               32'sh3ff3f420, 32'sh3ff3e4b1, 32'sh3ff3d537, 32'sh3ff3c5b3, 32'sh3ff3b626, 32'sh3ff3a68f, 32'sh3ff396ee, 32'sh3ff38743, 
               32'sh3ff3778e, 32'sh3ff367cf, 32'sh3ff35807, 32'sh3ff34834, 32'sh3ff33858, 32'sh3ff32872, 32'sh3ff31882, 32'sh3ff30888, 
               32'sh3ff2f884, 32'sh3ff2e876, 32'sh3ff2d85f, 32'sh3ff2c83e, 32'sh3ff2b813, 32'sh3ff2a7dd, 32'sh3ff2979f, 32'sh3ff28756, 
               32'sh3ff27703, 32'sh3ff266a7, 32'sh3ff25640, 32'sh3ff245d0, 32'sh3ff23556, 32'sh3ff224d2, 32'sh3ff21444, 32'sh3ff203ad, 
               32'sh3ff1f30b, 32'sh3ff1e260, 32'sh3ff1d1aa, 32'sh3ff1c0eb, 32'sh3ff1b022, 32'sh3ff19f50, 32'sh3ff18e73, 32'sh3ff17d8c, 
               32'sh3ff16c9c, 32'sh3ff15ba2, 32'sh3ff14a9e, 32'sh3ff13990, 32'sh3ff12878, 32'sh3ff11756, 32'sh3ff1062a, 32'sh3ff0f4f5, 
               32'sh3ff0e3b6, 32'sh3ff0d26d, 32'sh3ff0c11a, 32'sh3ff0afbd, 32'sh3ff09e56, 32'sh3ff08ce5, 32'sh3ff07b6b, 32'sh3ff069e7, 
               32'sh3ff05858, 32'sh3ff046c0, 32'sh3ff0351e, 32'sh3ff02373, 32'sh3ff011bd, 32'sh3feffffe, 32'sh3fefee34, 32'sh3fefdc61, 
               32'sh3fefca84, 32'sh3fefb89d, 32'sh3fefa6ac, 32'sh3fef94b2, 32'sh3fef82ad, 32'sh3fef709f, 32'sh3fef5e87, 32'sh3fef4c65, 
               32'sh3fef3a39, 32'sh3fef2803, 32'sh3fef15c3, 32'sh3fef037a, 32'sh3feef126, 32'sh3feedec9, 32'sh3feecc62, 32'sh3feeb9f1, 
               32'sh3feea776, 32'sh3fee94f2, 32'sh3fee8263, 32'sh3fee6fcb, 32'sh3fee5d28, 32'sh3fee4a7c, 32'sh3fee37c6, 32'sh3fee2507, 
               32'sh3fee123d, 32'sh3fedff69, 32'sh3fedec8c, 32'sh3fedd9a5, 32'sh3fedc6b4, 32'sh3fedb3b9, 32'sh3feda0b4, 32'sh3fed8da5, 
               32'sh3fed7a8c, 32'sh3fed676a, 32'sh3fed543e, 32'sh3fed4108, 32'sh3fed2dc8, 32'sh3fed1a7e, 32'sh3fed072a, 32'sh3fecf3cd, 
               32'sh3fece065, 32'sh3fecccf4, 32'sh3fecb979, 32'sh3feca5f4, 32'sh3fec9265, 32'sh3fec7ecc, 32'sh3fec6b2a, 32'sh3fec577d, 
               32'sh3fec43c7, 32'sh3fec3007, 32'sh3fec1c3d, 32'sh3fec0869, 32'sh3febf48b, 32'sh3febe0a4, 32'sh3febccb2, 32'sh3febb8b7, 
               32'sh3feba4b2, 32'sh3feb90a3, 32'sh3feb7c8a, 32'sh3feb6867, 32'sh3feb543b, 32'sh3feb4004, 32'sh3feb2bc4, 32'sh3feb177a, 
               32'sh3feb0326, 32'sh3feaeec8, 32'sh3feada60, 32'sh3feac5ef, 32'sh3feab173, 32'sh3fea9cee, 32'sh3fea885f, 32'sh3fea73c6, 
               32'sh3fea5f23, 32'sh3fea4a76, 32'sh3fea35c0, 32'sh3fea20ff, 32'sh3fea0c35, 32'sh3fe9f761, 32'sh3fe9e283, 32'sh3fe9cd9b, 
               32'sh3fe9b8a9, 32'sh3fe9a3ae, 32'sh3fe98ea8, 32'sh3fe97999, 32'sh3fe96480, 32'sh3fe94f5d, 32'sh3fe93a30, 32'sh3fe924f9, 
               32'sh3fe90fb9, 32'sh3fe8fa6f, 32'sh3fe8e51a, 32'sh3fe8cfbc, 32'sh3fe8ba54, 32'sh3fe8a4e2, 32'sh3fe88f67, 32'sh3fe879e1, 
               32'sh3fe86452, 32'sh3fe84eb8, 32'sh3fe83915, 32'sh3fe82368, 32'sh3fe80db2, 32'sh3fe7f7f1, 32'sh3fe7e226, 32'sh3fe7cc52, 
               32'sh3fe7b674, 32'sh3fe7a08c, 32'sh3fe78a9a, 32'sh3fe7749e, 32'sh3fe75e98, 32'sh3fe74889, 32'sh3fe7326f, 32'sh3fe71c4c, 
               32'sh3fe7061f, 32'sh3fe6efe8, 32'sh3fe6d9a7, 32'sh3fe6c35d, 32'sh3fe6ad08, 32'sh3fe696aa, 32'sh3fe68042, 32'sh3fe669d0, 
               32'sh3fe65354, 32'sh3fe63cce, 32'sh3fe6263e, 32'sh3fe60fa5, 32'sh3fe5f902, 32'sh3fe5e254, 32'sh3fe5cb9d, 32'sh3fe5b4dc, 
               32'sh3fe59e12, 32'sh3fe5873d, 32'sh3fe5705f, 32'sh3fe55976, 32'sh3fe54284, 32'sh3fe52b88, 32'sh3fe51482, 32'sh3fe4fd73, 
               32'sh3fe4e659, 32'sh3fe4cf36, 32'sh3fe4b808, 32'sh3fe4a0d1, 32'sh3fe48990, 32'sh3fe47245, 32'sh3fe45af1, 32'sh3fe44392, 
               32'sh3fe42c2a, 32'sh3fe414b8, 32'sh3fe3fd3b, 32'sh3fe3e5b5, 32'sh3fe3ce26, 32'sh3fe3b68c, 32'sh3fe39ee8, 32'sh3fe3873b, 
               32'sh3fe36f84, 32'sh3fe357c3, 32'sh3fe33ff8, 32'sh3fe32823, 32'sh3fe31045, 32'sh3fe2f85c, 32'sh3fe2e06a, 32'sh3fe2c86e, 
               32'sh3fe2b067, 32'sh3fe29858, 32'sh3fe2803e, 32'sh3fe2681a, 32'sh3fe24fed, 32'sh3fe237b6, 32'sh3fe21f74, 32'sh3fe20729, 
               32'sh3fe1eed5, 32'sh3fe1d676, 32'sh3fe1be0d, 32'sh3fe1a59b, 32'sh3fe18d1f, 32'sh3fe17499, 32'sh3fe15c09, 32'sh3fe1436f, 
               32'sh3fe12acb, 32'sh3fe1121e, 32'sh3fe0f966, 32'sh3fe0e0a5, 32'sh3fe0c7da, 32'sh3fe0af05, 32'sh3fe09626, 32'sh3fe07d3e, 
               32'sh3fe0644b, 32'sh3fe04b4f, 32'sh3fe03249, 32'sh3fe01939, 32'sh3fe0001f, 32'sh3fdfe6fb, 32'sh3fdfcdce, 32'sh3fdfb496, 
               32'sh3fdf9b55, 32'sh3fdf820a, 32'sh3fdf68b5, 32'sh3fdf4f56, 32'sh3fdf35ed, 32'sh3fdf1c7b, 32'sh3fdf02fe, 32'sh3fdee978, 
               32'sh3fdecfe8, 32'sh3fdeb64e, 32'sh3fde9caa, 32'sh3fde82fd, 32'sh3fde6945, 32'sh3fde4f84, 32'sh3fde35b9, 32'sh3fde1be4, 
               32'sh3fde0205, 32'sh3fdde81c, 32'sh3fddce2a, 32'sh3fddb42d, 32'sh3fdd9a27, 32'sh3fdd8017, 32'sh3fdd65fd, 32'sh3fdd4bd9, 
               32'sh3fdd31ac, 32'sh3fdd1774, 32'sh3fdcfd33, 32'sh3fdce2e8, 32'sh3fdcc892, 32'sh3fdcae34, 32'sh3fdc93cb, 32'sh3fdc7958, 
               32'sh3fdc5edc, 32'sh3fdc4455, 32'sh3fdc29c5, 32'sh3fdc0f2b, 32'sh3fdbf488, 32'sh3fdbd9da, 32'sh3fdbbf22, 32'sh3fdba461, 
               32'sh3fdb8996, 32'sh3fdb6ec1, 32'sh3fdb53e2, 32'sh3fdb38f9, 32'sh3fdb1e06, 32'sh3fdb030a, 32'sh3fdae804, 32'sh3fdaccf3, 
               32'sh3fdab1d9, 32'sh3fda96b6, 32'sh3fda7b88, 32'sh3fda6050, 32'sh3fda450f, 32'sh3fda29c4, 32'sh3fda0e6f, 32'sh3fd9f310, 
               32'sh3fd9d7a7, 32'sh3fd9bc34, 32'sh3fd9a0b8, 32'sh3fd98531, 32'sh3fd969a1, 32'sh3fd94e07, 32'sh3fd93263, 32'sh3fd916b6, 
               32'sh3fd8fafe, 32'sh3fd8df3d, 32'sh3fd8c372, 32'sh3fd8a79c, 32'sh3fd88bbe, 32'sh3fd86fd5, 32'sh3fd853e2, 32'sh3fd837e6, 
               32'sh3fd81bdf, 32'sh3fd7ffcf, 32'sh3fd7e3b5, 32'sh3fd7c791, 32'sh3fd7ab64, 32'sh3fd78f2c, 32'sh3fd772eb, 32'sh3fd7569f, 
               32'sh3fd73a4a, 32'sh3fd71deb, 32'sh3fd70183, 32'sh3fd6e510, 32'sh3fd6c894, 32'sh3fd6ac0d, 32'sh3fd68f7d, 32'sh3fd672e3, 
               32'sh3fd6563f, 32'sh3fd63992, 32'sh3fd61cda, 32'sh3fd60019, 32'sh3fd5e34e, 32'sh3fd5c678, 32'sh3fd5a99a, 32'sh3fd58cb1, 
               32'sh3fd56fbe, 32'sh3fd552c2, 32'sh3fd535bc, 32'sh3fd518ab, 32'sh3fd4fb91, 32'sh3fd4de6e, 32'sh3fd4c140, 32'sh3fd4a408, 
               32'sh3fd486c7, 32'sh3fd4697c, 32'sh3fd44c27, 32'sh3fd42ec8, 32'sh3fd4115f, 32'sh3fd3f3ed, 32'sh3fd3d670, 32'sh3fd3b8ea, 
               32'sh3fd39b5a, 32'sh3fd37dc0, 32'sh3fd3601c, 32'sh3fd3426f, 32'sh3fd324b7, 32'sh3fd306f6, 32'sh3fd2e92b, 32'sh3fd2cb56, 
               32'sh3fd2ad77, 32'sh3fd28f8e, 32'sh3fd2719c, 32'sh3fd2539f, 32'sh3fd23599, 32'sh3fd21789, 32'sh3fd1f96f, 32'sh3fd1db4c, 
               32'sh3fd1bd1e, 32'sh3fd19ee7, 32'sh3fd180a5, 32'sh3fd1625a, 32'sh3fd14405, 32'sh3fd125a7, 32'sh3fd1073e, 32'sh3fd0e8cc, 
               32'sh3fd0ca4f, 32'sh3fd0abc9, 32'sh3fd08d39, 32'sh3fd06e9f, 32'sh3fd04ffc, 32'sh3fd0314e, 32'sh3fd01297, 32'sh3fcff3d6, 
               32'sh3fcfd50b, 32'sh3fcfb636, 32'sh3fcf9757, 32'sh3fcf786e, 32'sh3fcf597c, 32'sh3fcf3a80, 32'sh3fcf1b7a, 32'sh3fcefc6a, 
               32'sh3fcedd50, 32'sh3fcebe2d, 32'sh3fce9eff, 32'sh3fce7fc8, 32'sh3fce6087, 32'sh3fce413c, 32'sh3fce21e7, 32'sh3fce0288, 
               32'sh3fcde320, 32'sh3fcdc3ae, 32'sh3fcda431, 32'sh3fcd84ab, 32'sh3fcd651c, 32'sh3fcd4582, 32'sh3fcd25de, 32'sh3fcd0631, 
               32'sh3fcce67a, 32'sh3fccc6b9, 32'sh3fcca6ee, 32'sh3fcc8719, 32'sh3fcc673b, 32'sh3fcc4753, 32'sh3fcc2760, 32'sh3fcc0764, 
               32'sh3fcbe75e, 32'sh3fcbc74f, 32'sh3fcba735, 32'sh3fcb8712, 32'sh3fcb66e4, 32'sh3fcb46ad, 32'sh3fcb266c, 32'sh3fcb0622, 
               32'sh3fcae5cd, 32'sh3fcac56f, 32'sh3fcaa506, 32'sh3fca8494, 32'sh3fca6418, 32'sh3fca4393, 32'sh3fca2303, 32'sh3fca026a, 
               32'sh3fc9e1c6, 32'sh3fc9c119, 32'sh3fc9a062, 32'sh3fc97fa1, 32'sh3fc95ed7, 32'sh3fc93e02, 32'sh3fc91d24, 32'sh3fc8fc3c, 
               32'sh3fc8db4a, 32'sh3fc8ba4e, 32'sh3fc89948, 32'sh3fc87839, 32'sh3fc8571f, 32'sh3fc835fc, 32'sh3fc814cf, 32'sh3fc7f398, 
               32'sh3fc7d258, 32'sh3fc7b10d, 32'sh3fc78fb9, 32'sh3fc76e5b, 32'sh3fc74cf3, 32'sh3fc72b81, 32'sh3fc70a05, 32'sh3fc6e880, 
               32'sh3fc6c6f0, 32'sh3fc6a557, 32'sh3fc683b4, 32'sh3fc66207, 32'sh3fc64051, 32'sh3fc61e90, 32'sh3fc5fcc6, 32'sh3fc5daf2, 
               32'sh3fc5b913, 32'sh3fc5972c, 32'sh3fc5753a, 32'sh3fc5533e, 32'sh3fc53139, 32'sh3fc50f2a, 32'sh3fc4ed11, 32'sh3fc4caee, 
               32'sh3fc4a8c1, 32'sh3fc4868b, 32'sh3fc4644a, 32'sh3fc44200, 32'sh3fc41fac, 32'sh3fc3fd4e, 32'sh3fc3dae6, 32'sh3fc3b875, 
               32'sh3fc395f9, 32'sh3fc37374, 32'sh3fc350e5, 32'sh3fc32e4c, 32'sh3fc30baa, 32'sh3fc2e8fd, 32'sh3fc2c647, 32'sh3fc2a387, 
               32'sh3fc280bc, 32'sh3fc25de9, 32'sh3fc23b0b, 32'sh3fc21823, 32'sh3fc1f532, 32'sh3fc1d237, 32'sh3fc1af32, 32'sh3fc18c23, 
               32'sh3fc1690a, 32'sh3fc145e8, 32'sh3fc122bb, 32'sh3fc0ff85, 32'sh3fc0dc45, 32'sh3fc0b8fb, 32'sh3fc095a8, 32'sh3fc0724a, 
               32'sh3fc04ee3, 32'sh3fc02b71, 32'sh3fc007f6, 32'sh3fbfe472, 32'sh3fbfc0e3, 32'sh3fbf9d4a, 32'sh3fbf79a8, 32'sh3fbf55fc, 
               32'sh3fbf3246, 32'sh3fbf0e86, 32'sh3fbeeabc, 32'sh3fbec6e9, 32'sh3fbea30c, 32'sh3fbe7f24, 32'sh3fbe5b33, 32'sh3fbe3739, 
               32'sh3fbe1334, 32'sh3fbdef26, 32'sh3fbdcb0d, 32'sh3fbda6eb, 32'sh3fbd82bf, 32'sh3fbd5e89, 32'sh3fbd3a4a, 32'sh3fbd1600, 
               32'sh3fbcf1ad, 32'sh3fbccd50, 32'sh3fbca8e9, 32'sh3fbc8478, 32'sh3fbc5ffe, 32'sh3fbc3b79, 32'sh3fbc16eb, 32'sh3fbbf253, 
               32'sh3fbbcdb1, 32'sh3fbba905, 32'sh3fbb8450, 32'sh3fbb5f90, 32'sh3fbb3ac7, 32'sh3fbb15f4, 32'sh3fbaf117, 32'sh3fbacc30, 
               32'sh3fbaa740, 32'sh3fba8246, 32'sh3fba5d41, 32'sh3fba3833, 32'sh3fba131b, 32'sh3fb9edfa, 32'sh3fb9c8ce, 32'sh3fb9a399, 
               32'sh3fb97e5a, 32'sh3fb95911, 32'sh3fb933be, 32'sh3fb90e61, 32'sh3fb8e8fb, 32'sh3fb8c38b, 32'sh3fb89e11, 32'sh3fb8788d, 
               32'sh3fb852ff, 32'sh3fb82d67, 32'sh3fb807c6, 32'sh3fb7e21b, 32'sh3fb7bc65, 32'sh3fb796a7, 32'sh3fb770de, 32'sh3fb74b0b, 
               32'sh3fb7252f, 32'sh3fb6ff49, 32'sh3fb6d959, 32'sh3fb6b35f, 32'sh3fb68d5b, 32'sh3fb6674e, 32'sh3fb64136, 32'sh3fb61b15, 
               32'sh3fb5f4ea, 32'sh3fb5ceb5, 32'sh3fb5a877, 32'sh3fb5822e, 32'sh3fb55bdc, 32'sh3fb53580, 32'sh3fb50f1a, 32'sh3fb4e8aa, 
               32'sh3fb4c231, 32'sh3fb49bad, 32'sh3fb47520, 32'sh3fb44e89, 32'sh3fb427e8, 32'sh3fb4013d, 32'sh3fb3da89, 32'sh3fb3b3ca, 
               32'sh3fb38d02, 32'sh3fb36630, 32'sh3fb33f54, 32'sh3fb3186f, 32'sh3fb2f17f, 32'sh3fb2ca86, 32'sh3fb2a383, 32'sh3fb27c76, 
               32'sh3fb2555f, 32'sh3fb22e3f, 32'sh3fb20714, 32'sh3fb1dfe0, 32'sh3fb1b8a2, 32'sh3fb1915a, 32'sh3fb16a08, 32'sh3fb142ad, 
               32'sh3fb11b48, 32'sh3fb0f3d8, 32'sh3fb0cc5f, 32'sh3fb0a4dd, 32'sh3fb07d50, 32'sh3fb055ba, 32'sh3fb02e19, 32'sh3fb0066f, 
               32'sh3fafdebb, 32'sh3fafb6fe, 32'sh3faf8f36, 32'sh3faf6765, 32'sh3faf3f89, 32'sh3faf17a4, 32'sh3faeefb6, 32'sh3faec7bd, 
               32'sh3fae9fbb, 32'sh3fae77ae, 32'sh3fae4f98, 32'sh3fae2778, 32'sh3fadff4e, 32'sh3fadd71b, 32'sh3fadaedd, 32'sh3fad8696, 
               32'sh3fad5e45, 32'sh3fad35ea, 32'sh3fad0d86, 32'sh3face517, 32'sh3facbc9f, 32'sh3fac941d, 32'sh3fac6b91, 32'sh3fac42fb, 
               32'sh3fac1a5b, 32'sh3fabf1b2, 32'sh3fabc8ff, 32'sh3faba042, 32'sh3fab777b, 32'sh3fab4eaa, 32'sh3fab25d0, 32'sh3faafceb, 
               32'sh3faad3fd, 32'sh3faaab05, 32'sh3faa8203, 32'sh3faa58f8, 32'sh3faa2fe2, 32'sh3faa06c3, 32'sh3fa9dd9a, 32'sh3fa9b467, 
               32'sh3fa98b2a, 32'sh3fa961e4, 32'sh3fa93894, 32'sh3fa90f39, 32'sh3fa8e5d5, 32'sh3fa8bc68, 32'sh3fa892f0, 32'sh3fa8696f, 
               32'sh3fa83fe3, 32'sh3fa8164e, 32'sh3fa7ecb0, 32'sh3fa7c307, 32'sh3fa79954, 32'sh3fa76f98, 32'sh3fa745d2, 32'sh3fa71c02, 
               32'sh3fa6f228, 32'sh3fa6c845, 32'sh3fa69e57, 32'sh3fa67460, 32'sh3fa64a5f, 32'sh3fa62054, 32'sh3fa5f640, 32'sh3fa5cc21, 
               32'sh3fa5a1f9, 32'sh3fa577c7, 32'sh3fa54d8b, 32'sh3fa52345, 32'sh3fa4f8f6, 32'sh3fa4ce9c, 32'sh3fa4a439, 32'sh3fa479cc, 
               32'sh3fa44f55, 32'sh3fa424d5, 32'sh3fa3fa4a, 32'sh3fa3cfb6, 32'sh3fa3a518, 32'sh3fa37a70, 32'sh3fa34fbe, 32'sh3fa32503, 
               32'sh3fa2fa3d, 32'sh3fa2cf6e, 32'sh3fa2a495, 32'sh3fa279b3, 32'sh3fa24ec6, 32'sh3fa223d0, 32'sh3fa1f8d0, 32'sh3fa1cdc6, 
               32'sh3fa1a2b2, 32'sh3fa17794, 32'sh3fa14c6d, 32'sh3fa1213b, 32'sh3fa0f600, 32'sh3fa0cabb, 32'sh3fa09f6d, 32'sh3fa07414, 
               32'sh3fa048b2, 32'sh3fa01d46, 32'sh3f9ff1d0, 32'sh3f9fc650, 32'sh3f9f9ac6, 32'sh3f9f6f33, 32'sh3f9f4396, 32'sh3f9f17ef, 
               32'sh3f9eec3e, 32'sh3f9ec083, 32'sh3f9e94bf, 32'sh3f9e68f1, 32'sh3f9e3d19, 32'sh3f9e1137, 32'sh3f9de54b, 32'sh3f9db956, 
               32'sh3f9d8d56, 32'sh3f9d614d, 32'sh3f9d353a, 32'sh3f9d091e, 32'sh3f9cdcf7, 32'sh3f9cb0c7, 32'sh3f9c848d, 32'sh3f9c5849, 
               32'sh3f9c2bfb, 32'sh3f9bffa3, 32'sh3f9bd342, 32'sh3f9ba6d7, 32'sh3f9b7a62, 32'sh3f9b4de3, 32'sh3f9b215a, 32'sh3f9af4c8, 
               32'sh3f9ac82c, 32'sh3f9a9b85, 32'sh3f9a6ed6, 32'sh3f9a421c, 32'sh3f9a1558, 32'sh3f99e88b, 32'sh3f99bbb4, 32'sh3f998ed3, 
               32'sh3f9961e8, 32'sh3f9934f4, 32'sh3f9907f6, 32'sh3f98daed, 32'sh3f98addb, 32'sh3f9880c0, 32'sh3f98539a, 32'sh3f98266b, 
               32'sh3f97f932, 32'sh3f97cbef, 32'sh3f979ea2, 32'sh3f97714b, 32'sh3f9743eb, 32'sh3f971681, 32'sh3f96e90d, 32'sh3f96bb8f, 
               32'sh3f968e07, 32'sh3f966076, 32'sh3f9632da, 32'sh3f960535, 32'sh3f95d787, 32'sh3f95a9ce, 32'sh3f957c0b, 32'sh3f954e3f, 
               32'sh3f952069, 32'sh3f94f289, 32'sh3f94c4a0, 32'sh3f9496ac, 32'sh3f9468af, 32'sh3f943aa8, 32'sh3f940c97, 32'sh3f93de7c, 
               32'sh3f93b058, 32'sh3f938229, 32'sh3f9353f1, 32'sh3f9325af, 32'sh3f92f763, 32'sh3f92c90e, 32'sh3f929aaf, 32'sh3f926c45, 
               32'sh3f923dd2, 32'sh3f920f56, 32'sh3f91e0cf, 32'sh3f91b23f, 32'sh3f9183a5, 32'sh3f915501, 32'sh3f912653, 32'sh3f90f79b, 
               32'sh3f90c8da, 32'sh3f909a0f, 32'sh3f906b3a, 32'sh3f903c5b, 32'sh3f900d72, 32'sh3f8fde80, 32'sh3f8faf84, 32'sh3f8f807e, 
               32'sh3f8f516e, 32'sh3f8f2255, 32'sh3f8ef331, 32'sh3f8ec404, 32'sh3f8e94cd, 32'sh3f8e658c, 32'sh3f8e3642, 32'sh3f8e06ed, 
               32'sh3f8dd78f, 32'sh3f8da827, 32'sh3f8d78b5, 32'sh3f8d493a, 32'sh3f8d19b4, 32'sh3f8cea25, 32'sh3f8cba8c, 32'sh3f8c8ae9, 
               32'sh3f8c5b3d, 32'sh3f8c2b86, 32'sh3f8bfbc6, 32'sh3f8bcbfc, 32'sh3f8b9c28, 32'sh3f8b6c4b, 32'sh3f8b3c63, 32'sh3f8b0c72, 
               32'sh3f8adc77, 32'sh3f8aac72, 32'sh3f8a7c64, 32'sh3f8a4c4b, 32'sh3f8a1c29, 32'sh3f89ebfd, 32'sh3f89bbc7, 32'sh3f898b88, 
               32'sh3f895b3e, 32'sh3f892aeb, 32'sh3f88fa8e, 32'sh3f88ca27, 32'sh3f8899b7, 32'sh3f88693c, 32'sh3f8838b8, 32'sh3f88082a, 
               32'sh3f87d792, 32'sh3f87a6f1, 32'sh3f877645, 32'sh3f874590, 32'sh3f8714d1, 32'sh3f86e409, 32'sh3f86b336, 32'sh3f86825a, 
               32'sh3f865174, 32'sh3f862084, 32'sh3f85ef8a, 32'sh3f85be86, 32'sh3f858d79, 32'sh3f855c62, 32'sh3f852b41, 32'sh3f84fa16, 
               32'sh3f84c8e2, 32'sh3f8497a3, 32'sh3f84665b, 32'sh3f843509, 32'sh3f8403ae, 32'sh3f83d248, 32'sh3f83a0d9, 32'sh3f836f60, 
               32'sh3f833ddd, 32'sh3f830c50, 32'sh3f82daba, 32'sh3f82a91a, 32'sh3f827770, 32'sh3f8245bc, 32'sh3f8213fe, 32'sh3f81e237, 
               32'sh3f81b065, 32'sh3f817e8a, 32'sh3f814ca6, 32'sh3f811ab7, 32'sh3f80e8bf, 32'sh3f80b6bc, 32'sh3f8084b0, 32'sh3f80529b, 
               32'sh3f80207b, 32'sh3f7fee52, 32'sh3f7fbc1f, 32'sh3f7f89e2, 32'sh3f7f579b, 32'sh3f7f254a, 32'sh3f7ef2f0, 32'sh3f7ec08c, 
               32'sh3f7e8e1e, 32'sh3f7e5ba6, 32'sh3f7e2925, 32'sh3f7df69a, 32'sh3f7dc405, 32'sh3f7d9166, 32'sh3f7d5ebd, 32'sh3f7d2c0b, 
               32'sh3f7cf94e, 32'sh3f7cc688, 32'sh3f7c93b9, 32'sh3f7c60df, 32'sh3f7c2dfc, 32'sh3f7bfb0e, 32'sh3f7bc817, 32'sh3f7b9517, 
               32'sh3f7b620c, 32'sh3f7b2ef8, 32'sh3f7afbda, 32'sh3f7ac8b2, 32'sh3f7a9580, 32'sh3f7a6244, 32'sh3f7a2eff, 32'sh3f79fbb0, 
               32'sh3f79c857, 32'sh3f7994f4, 32'sh3f796188, 32'sh3f792e12, 32'sh3f78fa92, 32'sh3f78c708, 32'sh3f789374, 32'sh3f785fd7, 
               32'sh3f782c30, 32'sh3f77f87f, 32'sh3f77c4c4, 32'sh3f779100, 32'sh3f775d31, 32'sh3f772959, 32'sh3f76f577, 32'sh3f76c18b, 
               32'sh3f768d96, 32'sh3f765997, 32'sh3f76258e, 32'sh3f75f17b, 32'sh3f75bd5e, 32'sh3f758938, 32'sh3f755508, 32'sh3f7520ce, 
               32'sh3f74ec8a, 32'sh3f74b83c, 32'sh3f7483e5, 32'sh3f744f84, 32'sh3f741b19, 32'sh3f73e6a4, 32'sh3f73b226, 32'sh3f737d9e, 
               32'sh3f73490b, 32'sh3f731470, 32'sh3f72dfca, 32'sh3f72ab1b, 32'sh3f727661, 32'sh3f72419e, 32'sh3f720cd2, 32'sh3f71d7fb, 
               32'sh3f71a31b, 32'sh3f716e31, 32'sh3f71393d, 32'sh3f71043f, 32'sh3f70cf38, 32'sh3f709a26, 32'sh3f70650b, 32'sh3f702fe7, 
               32'sh3f6ffab8, 32'sh3f6fc580, 32'sh3f6f903d, 32'sh3f6f5af2, 32'sh3f6f259c, 32'sh3f6ef03c, 32'sh3f6ebad3, 32'sh3f6e8560, 
               32'sh3f6e4fe3, 32'sh3f6e1a5c, 32'sh3f6de4cc, 32'sh3f6daf32, 32'sh3f6d798e, 32'sh3f6d43e0, 32'sh3f6d0e29, 32'sh3f6cd867, 
               32'sh3f6ca29c, 32'sh3f6c6cc7, 32'sh3f6c36e9, 32'sh3f6c0100, 32'sh3f6bcb0e, 32'sh3f6b9512, 32'sh3f6b5f0c, 32'sh3f6b28fd, 
               32'sh3f6af2e3, 32'sh3f6abcc0, 32'sh3f6a8693, 32'sh3f6a505c, 32'sh3f6a1a1c, 32'sh3f69e3d2, 32'sh3f69ad7e, 32'sh3f697720, 
               32'sh3f6940b8, 32'sh3f690a47, 32'sh3f68d3cc, 32'sh3f689d47, 32'sh3f6866b8, 32'sh3f683020, 32'sh3f67f97d, 32'sh3f67c2d1, 
               32'sh3f678c1c, 32'sh3f67555c, 32'sh3f671e93, 32'sh3f66e7c0, 32'sh3f66b0e3, 32'sh3f6679fc, 32'sh3f66430b, 32'sh3f660c11, 
               32'sh3f65d50d, 32'sh3f659dff, 32'sh3f6566e8, 32'sh3f652fc6, 32'sh3f64f89b, 32'sh3f64c166, 32'sh3f648a28, 32'sh3f6452df, 
               32'sh3f641b8d, 32'sh3f63e431, 32'sh3f63accb, 32'sh3f63755c, 32'sh3f633de2, 32'sh3f63065f, 32'sh3f62ced2, 32'sh3f62973c, 
               32'sh3f625f9b, 32'sh3f6227f1, 32'sh3f61f03d, 32'sh3f61b87f, 32'sh3f6180b8, 32'sh3f6148e6, 32'sh3f61110b, 32'sh3f60d926, 
               32'sh3f60a138, 32'sh3f60693f, 32'sh3f60313d, 32'sh3f5ff931, 32'sh3f5fc11c, 32'sh3f5f88fc, 32'sh3f5f50d3, 32'sh3f5f18a0, 
               32'sh3f5ee063, 32'sh3f5ea81c, 32'sh3f5e6fcc, 32'sh3f5e3772, 32'sh3f5dff0e, 32'sh3f5dc6a0, 32'sh3f5d8e29, 32'sh3f5d55a8, 
               32'sh3f5d1d1d, 32'sh3f5ce488, 32'sh3f5cabe9, 32'sh3f5c7341, 32'sh3f5c3a8f, 32'sh3f5c01d3, 32'sh3f5bc90d, 32'sh3f5b903e, 
               32'sh3f5b5765, 32'sh3f5b1e82, 32'sh3f5ae595, 32'sh3f5aac9f, 32'sh3f5a739e, 32'sh3f5a3a94, 32'sh3f5a0181, 32'sh3f59c863, 
               32'sh3f598f3c, 32'sh3f59560b, 32'sh3f591cd0, 32'sh3f58e38b, 32'sh3f58aa3d, 32'sh3f5870e5, 32'sh3f583783, 32'sh3f57fe17, 
               32'sh3f57c4a2, 32'sh3f578b22, 32'sh3f575199, 32'sh3f571807, 32'sh3f56de6a, 32'sh3f56a4c4, 32'sh3f566b14, 32'sh3f56315a, 
               32'sh3f55f796, 32'sh3f55bdc9, 32'sh3f5583f2, 32'sh3f554a11, 32'sh3f551026, 32'sh3f54d632, 32'sh3f549c33, 32'sh3f54622b, 
               32'sh3f54281a, 32'sh3f53edfe, 32'sh3f53b3d9, 32'sh3f5379aa, 32'sh3f533f71, 32'sh3f53052e, 32'sh3f52cae2, 32'sh3f52908c, 
               32'sh3f52562c, 32'sh3f521bc2, 32'sh3f51e14f, 32'sh3f51a6d2, 32'sh3f516c4b, 32'sh3f5131ba, 32'sh3f50f720, 32'sh3f50bc7b, 
               32'sh3f5081cd, 32'sh3f504716, 32'sh3f500c54, 32'sh3f4fd189, 32'sh3f4f96b4, 32'sh3f4f5bd5, 32'sh3f4f20ed, 32'sh3f4ee5fa, 
               32'sh3f4eaafe, 32'sh3f4e6ff8, 32'sh3f4e34e9, 32'sh3f4df9cf, 32'sh3f4dbeac, 32'sh3f4d837f, 32'sh3f4d4848, 32'sh3f4d0d08, 
               32'sh3f4cd1be, 32'sh3f4c966a, 32'sh3f4c5b0c, 32'sh3f4c1fa5, 32'sh3f4be433, 32'sh3f4ba8b8, 32'sh3f4b6d34, 32'sh3f4b31a5, 
               32'sh3f4af60d, 32'sh3f4aba6b, 32'sh3f4a7ebf, 32'sh3f4a4309, 32'sh3f4a074a, 32'sh3f49cb81, 32'sh3f498fae, 32'sh3f4953d2, 
               32'sh3f4917eb, 32'sh3f48dbfb, 32'sh3f48a001, 32'sh3f4863fe, 32'sh3f4827f0, 32'sh3f47ebd9, 32'sh3f47afb8, 32'sh3f47738d, 
               32'sh3f473759, 32'sh3f46fb1b, 32'sh3f46bed3, 32'sh3f468281, 32'sh3f464626, 32'sh3f4609c0, 32'sh3f45cd51, 32'sh3f4590d9, 
               32'sh3f455456, 32'sh3f4517ca, 32'sh3f44db34, 32'sh3f449e94, 32'sh3f4461eb, 32'sh3f442537, 32'sh3f43e87a, 32'sh3f43abb3, 
               32'sh3f436ee3, 32'sh3f433209, 32'sh3f42f525, 32'sh3f42b837, 32'sh3f427b3f, 32'sh3f423e3e, 32'sh3f420133, 32'sh3f41c41e, 
               32'sh3f4186ff, 32'sh3f4149d7, 32'sh3f410ca5, 32'sh3f40cf69, 32'sh3f409223, 32'sh3f4054d4, 32'sh3f40177b, 32'sh3f3fda18, 
               32'sh3f3f9cab, 32'sh3f3f5f35, 32'sh3f3f21b5, 32'sh3f3ee42b, 32'sh3f3ea697, 32'sh3f3e68fa, 32'sh3f3e2b53, 32'sh3f3deda2, 
               32'sh3f3dafe7, 32'sh3f3d7223, 32'sh3f3d3455, 32'sh3f3cf67d, 32'sh3f3cb89b, 32'sh3f3c7ab0, 32'sh3f3c3cba, 32'sh3f3bfebc, 
               32'sh3f3bc0b3, 32'sh3f3b82a0, 32'sh3f3b4484, 32'sh3f3b065e, 32'sh3f3ac82f, 32'sh3f3a89f5, 32'sh3f3a4bb2, 32'sh3f3a0d65, 
               32'sh3f39cf0e, 32'sh3f3990ae, 32'sh3f395244, 32'sh3f3913d0, 32'sh3f38d552, 32'sh3f3896cb, 32'sh3f38583a, 32'sh3f38199f, 
               32'sh3f37dafa, 32'sh3f379c4c, 32'sh3f375d93, 32'sh3f371ed1, 32'sh3f36e006, 32'sh3f36a130, 32'sh3f366251, 32'sh3f362368, 
               32'sh3f35e476, 32'sh3f35a579, 32'sh3f356673, 32'sh3f352763, 32'sh3f34e849, 32'sh3f34a926, 32'sh3f3469f9, 32'sh3f342ac2, 
               32'sh3f33eb81, 32'sh3f33ac37, 32'sh3f336ce3, 32'sh3f332d85, 32'sh3f32ee1d, 32'sh3f32aeac, 32'sh3f326f31, 32'sh3f322fac, 
               32'sh3f31f01d, 32'sh3f31b085, 32'sh3f3170e3, 32'sh3f313137, 32'sh3f30f181, 32'sh3f30b1c2, 32'sh3f3071f9, 32'sh3f303226, 
               32'sh3f2ff24a, 32'sh3f2fb263, 32'sh3f2f7273, 32'sh3f2f3279, 32'sh3f2ef276, 32'sh3f2eb269, 32'sh3f2e7252, 32'sh3f2e3231, 
               32'sh3f2df206, 32'sh3f2db1d2, 32'sh3f2d7194, 32'sh3f2d314c, 32'sh3f2cf0fb, 32'sh3f2cb09f, 32'sh3f2c703a, 32'sh3f2c2fcc, 
               32'sh3f2bef53, 32'sh3f2baed1, 32'sh3f2b6e45, 32'sh3f2b2daf, 32'sh3f2aed10, 32'sh3f2aac67, 32'sh3f2a6bb4, 32'sh3f2a2af7, 
               32'sh3f29ea31, 32'sh3f29a961, 32'sh3f296887, 32'sh3f2927a3, 32'sh3f28e6b6, 32'sh3f28a5bf, 32'sh3f2864be, 32'sh3f2823b3, 
               32'sh3f27e29f, 32'sh3f27a181, 32'sh3f276059, 32'sh3f271f28, 32'sh3f26ddec, 32'sh3f269ca7, 32'sh3f265b59, 32'sh3f261a00, 
               32'sh3f25d89e, 32'sh3f259732, 32'sh3f2555bc, 32'sh3f25143d, 32'sh3f24d2b4, 32'sh3f249121, 32'sh3f244f84, 32'sh3f240dde, 
               32'sh3f23cc2e, 32'sh3f238a74, 32'sh3f2348b0, 32'sh3f2306e3, 32'sh3f22c50c, 32'sh3f22832b, 32'sh3f224140, 32'sh3f21ff4c, 
               32'sh3f21bd4e, 32'sh3f217b46, 32'sh3f213935, 32'sh3f20f71a, 32'sh3f20b4f5, 32'sh3f2072c6, 32'sh3f20308d, 32'sh3f1fee4b, 
               32'sh3f1fabff, 32'sh3f1f69aa, 32'sh3f1f274a, 32'sh3f1ee4e1, 32'sh3f1ea26e, 32'sh3f1e5ff2, 32'sh3f1e1d6c, 32'sh3f1ddadb, 
               32'sh3f1d9842, 32'sh3f1d559e, 32'sh3f1d12f1, 32'sh3f1cd03a, 32'sh3f1c8d79, 32'sh3f1c4aaf, 32'sh3f1c07db, 32'sh3f1bc4fd, 
               32'sh3f1b8215, 32'sh3f1b3f24, 32'sh3f1afc29, 32'sh3f1ab924, 32'sh3f1a7615, 32'sh3f1a32fd, 32'sh3f19efdb, 32'sh3f19acaf, 
               32'sh3f19697a, 32'sh3f19263b, 32'sh3f18e2f2, 32'sh3f189f9f, 32'sh3f185c43, 32'sh3f1818dc, 32'sh3f17d56d, 32'sh3f1791f3, 
               32'sh3f174e70, 32'sh3f170ae3, 32'sh3f16c74c, 32'sh3f1683ab, 32'sh3f164001, 32'sh3f15fc4d, 32'sh3f15b88f, 32'sh3f1574c8, 
               32'sh3f1530f7, 32'sh3f14ed1c, 32'sh3f14a937, 32'sh3f146549, 32'sh3f142151, 32'sh3f13dd4f, 32'sh3f139944, 32'sh3f13552e, 
               32'sh3f13110f, 32'sh3f12cce7, 32'sh3f1288b4, 32'sh3f124478, 32'sh3f120032, 32'sh3f11bbe2, 32'sh3f117789, 32'sh3f113326, 
               32'sh3f10eeb9, 32'sh3f10aa43, 32'sh3f1065c3, 32'sh3f102139, 32'sh3f0fdca5, 32'sh3f0f9807, 32'sh3f0f5360, 32'sh3f0f0eaf, 
               32'sh3f0ec9f5, 32'sh3f0e8531, 32'sh3f0e4063, 32'sh3f0dfb8b, 32'sh3f0db6a9, 32'sh3f0d71be, 32'sh3f0d2cc9, 32'sh3f0ce7ca, 
               32'sh3f0ca2c2, 32'sh3f0c5db0, 32'sh3f0c1894, 32'sh3f0bd36f, 32'sh3f0b8e3f, 32'sh3f0b4906, 32'sh3f0b03c4, 32'sh3f0abe77, 
               32'sh3f0a7921, 32'sh3f0a33c1, 32'sh3f09ee58, 32'sh3f09a8e4, 32'sh3f096367, 32'sh3f091de0, 32'sh3f08d850, 32'sh3f0892b6, 
               32'sh3f084d12, 32'sh3f080764, 32'sh3f07c1ad, 32'sh3f077bec, 32'sh3f073621, 32'sh3f06f04c, 32'sh3f06aa6e, 32'sh3f066486, 
               32'sh3f061e95, 32'sh3f05d899, 32'sh3f059294, 32'sh3f054c85, 32'sh3f05066d, 32'sh3f04c04a, 32'sh3f047a1e, 32'sh3f0433e9, 
               32'sh3f03eda9, 32'sh3f03a760, 32'sh3f03610d, 32'sh3f031ab1, 32'sh3f02d44a, 32'sh3f028dda, 32'sh3f024760, 32'sh3f0200dd, 
               32'sh3f01ba50, 32'sh3f0173b9, 32'sh3f012d18, 32'sh3f00e66e, 32'sh3f009fba, 32'sh3f0058fc, 32'sh3f001235, 32'sh3effcb64, 
               32'sh3eff8489, 32'sh3eff3da4, 32'sh3efef6b6, 32'sh3efeafbe, 32'sh3efe68bc, 32'sh3efe21b0, 32'sh3efdda9b, 32'sh3efd937c, 
               32'sh3efd4c54, 32'sh3efd0521, 32'sh3efcbde5, 32'sh3efc76a0, 32'sh3efc2f50, 32'sh3efbe7f7, 32'sh3efba094, 32'sh3efb5928, 
               32'sh3efb11b1, 32'sh3efaca31, 32'sh3efa82a7, 32'sh3efa3b14, 32'sh3ef9f377, 32'sh3ef9abd0, 32'sh3ef9641f, 32'sh3ef91c65, 
               32'sh3ef8d4a1, 32'sh3ef88cd3, 32'sh3ef844fc, 32'sh3ef7fd1b, 32'sh3ef7b530, 32'sh3ef76d3b, 32'sh3ef7253d, 32'sh3ef6dd35, 
               32'sh3ef69523, 32'sh3ef64d08, 32'sh3ef604e3, 32'sh3ef5bcb4, 32'sh3ef5747b, 32'sh3ef52c39, 32'sh3ef4e3ed, 32'sh3ef49b98, 
               32'sh3ef45338, 32'sh3ef40acf, 32'sh3ef3c25c, 32'sh3ef379e0, 32'sh3ef3315a, 32'sh3ef2e8ca, 32'sh3ef2a030, 32'sh3ef2578d, 
               32'sh3ef20ee0, 32'sh3ef1c629, 32'sh3ef17d69, 32'sh3ef1349e, 32'sh3ef0ebcb, 32'sh3ef0a2ed, 32'sh3ef05a06, 32'sh3ef01115, 
               32'sh3eefc81a, 32'sh3eef7f16, 32'sh3eef3608, 32'sh3eeeecf0, 32'sh3eeea3ce, 32'sh3eee5aa3, 32'sh3eee116e, 32'sh3eedc830, 
               32'sh3eed7ee7, 32'sh3eed3595, 32'sh3eecec39, 32'sh3eeca2d4, 32'sh3eec5965, 32'sh3eec0fec, 32'sh3eebc669, 32'sh3eeb7cdd, 
               32'sh3eeb3347, 32'sh3eeae9a8, 32'sh3eea9ffe, 32'sh3eea564b, 32'sh3eea0c8e, 32'sh3ee9c2c8, 32'sh3ee978f8, 32'sh3ee92f1e, 
               32'sh3ee8e53a, 32'sh3ee89b4d, 32'sh3ee85156, 32'sh3ee80755, 32'sh3ee7bd4b, 32'sh3ee77337, 32'sh3ee72919, 32'sh3ee6def2, 
               32'sh3ee694c1, 32'sh3ee64a86, 32'sh3ee60041, 32'sh3ee5b5f3, 32'sh3ee56b9b, 32'sh3ee52139, 32'sh3ee4d6ce, 32'sh3ee48c59, 
               32'sh3ee441da, 32'sh3ee3f751, 32'sh3ee3acbf, 32'sh3ee36223, 32'sh3ee3177e, 32'sh3ee2cccf, 32'sh3ee28216, 32'sh3ee23753, 
               32'sh3ee1ec87, 32'sh3ee1a1b1, 32'sh3ee156d1, 32'sh3ee10be7, 32'sh3ee0c0f4, 32'sh3ee075f7, 32'sh3ee02af1, 32'sh3edfdfe1, 
               32'sh3edf94c7, 32'sh3edf49a3, 32'sh3edefe76, 32'sh3edeb33f, 32'sh3ede67fe, 32'sh3ede1cb4, 32'sh3eddd15f, 32'sh3edd8602, 
               32'sh3edd3a9a, 32'sh3edcef29, 32'sh3edca3ae, 32'sh3edc5829, 32'sh3edc0c9b, 32'sh3edbc103, 32'sh3edb7562, 32'sh3edb29b6, 
               32'sh3edade01, 32'sh3eda9242, 32'sh3eda467a, 32'sh3ed9faa8, 32'sh3ed9aecc, 32'sh3ed962e7, 32'sh3ed916f7, 32'sh3ed8caff, 
               32'sh3ed87efc, 32'sh3ed832f0, 32'sh3ed7e6da, 32'sh3ed79aba, 32'sh3ed74e91, 32'sh3ed7025e, 32'sh3ed6b621, 32'sh3ed669da, 
               32'sh3ed61d8a, 32'sh3ed5d131, 32'sh3ed584cd, 32'sh3ed53860, 32'sh3ed4ebe9, 32'sh3ed49f68, 32'sh3ed452de, 32'sh3ed4064a, 
               32'sh3ed3b9ad, 32'sh3ed36d05, 32'sh3ed32054, 32'sh3ed2d39a, 32'sh3ed286d5, 32'sh3ed23a07, 32'sh3ed1ed2f, 32'sh3ed1a04e, 
               32'sh3ed15363, 32'sh3ed1066e, 32'sh3ed0b970, 32'sh3ed06c67, 32'sh3ed01f55, 32'sh3ecfd23a, 32'sh3ecf8515, 32'sh3ecf37e6, 
               32'sh3eceeaad, 32'sh3ece9d6b, 32'sh3ece501f, 32'sh3ece02c9, 32'sh3ecdb56a, 32'sh3ecd6801, 32'sh3ecd1a8e, 32'sh3ecccd11, 
               32'sh3ecc7f8b, 32'sh3ecc31fc, 32'sh3ecbe462, 32'sh3ecb96bf, 32'sh3ecb4912, 32'sh3ecafb5c, 32'sh3ecaad9b, 32'sh3eca5fd1, 
               32'sh3eca11fe, 32'sh3ec9c421, 32'sh3ec9763a, 32'sh3ec92849, 32'sh3ec8da4f, 32'sh3ec88c4b, 32'sh3ec83e3d, 32'sh3ec7f026, 
               32'sh3ec7a205, 32'sh3ec753da, 32'sh3ec705a6, 32'sh3ec6b768, 32'sh3ec66920, 32'sh3ec61ace, 32'sh3ec5cc73, 32'sh3ec57e0e, 
               32'sh3ec52fa0, 32'sh3ec4e128, 32'sh3ec492a6, 32'sh3ec4441a, 32'sh3ec3f585, 32'sh3ec3a6e6, 32'sh3ec3583e, 32'sh3ec3098c, 
               32'sh3ec2bad0, 32'sh3ec26c0a, 32'sh3ec21d3b, 32'sh3ec1ce62, 32'sh3ec17f7f, 32'sh3ec13093, 32'sh3ec0e19d, 32'sh3ec0929d, 
               32'sh3ec04394, 32'sh3ebff481, 32'sh3ebfa564, 32'sh3ebf563e, 32'sh3ebf070e, 32'sh3ebeb7d4, 32'sh3ebe6891, 32'sh3ebe1944, 
               32'sh3ebdc9ed, 32'sh3ebd7a8c, 32'sh3ebd2b22, 32'sh3ebcdbaf, 32'sh3ebc8c31, 32'sh3ebc3caa, 32'sh3ebbed19, 32'sh3ebb9d7f, 
               32'sh3ebb4ddb, 32'sh3ebafe2d, 32'sh3ebaae75, 32'sh3eba5eb4, 32'sh3eba0ee9, 32'sh3eb9bf15, 32'sh3eb96f36, 32'sh3eb91f4f, 
               32'sh3eb8cf5d, 32'sh3eb87f62, 32'sh3eb82f5d, 32'sh3eb7df4e, 32'sh3eb78f36, 32'sh3eb73f14, 32'sh3eb6eee9, 32'sh3eb69eb4, 
               32'sh3eb64e75, 32'sh3eb5fe2c, 32'sh3eb5adda, 32'sh3eb55d7e, 32'sh3eb50d18, 32'sh3eb4bca9, 32'sh3eb46c30, 32'sh3eb41bad, 
               32'sh3eb3cb21, 32'sh3eb37a8b, 32'sh3eb329ec, 32'sh3eb2d942, 32'sh3eb2888f, 32'sh3eb237d3, 32'sh3eb1e70d, 32'sh3eb1963d, 
               32'sh3eb14563, 32'sh3eb0f480, 32'sh3eb0a393, 32'sh3eb0529c, 32'sh3eb0019c, 32'sh3eafb092, 32'sh3eaf5f7e, 32'sh3eaf0e61, 
               32'sh3eaebd3a, 32'sh3eae6c09, 32'sh3eae1acf, 32'sh3eadc98b, 32'sh3ead783d, 32'sh3ead26e6, 32'sh3eacd585, 32'sh3eac841b, 
               32'sh3eac32a6, 32'sh3eabe128, 32'sh3eab8fa1, 32'sh3eab3e0f, 32'sh3eaaec74, 32'sh3eaa9ad0, 32'sh3eaa4922, 32'sh3ea9f76a, 
               32'sh3ea9a5a8, 32'sh3ea953dd, 32'sh3ea90208, 32'sh3ea8b029, 32'sh3ea85e41, 32'sh3ea80c4f, 32'sh3ea7ba54, 32'sh3ea7684e, 
               32'sh3ea7163f, 32'sh3ea6c427, 32'sh3ea67205, 32'sh3ea61fd9, 32'sh3ea5cda3, 32'sh3ea57b64, 32'sh3ea5291b, 32'sh3ea4d6c9, 
               32'sh3ea4846c, 32'sh3ea43206, 32'sh3ea3df97, 32'sh3ea38d1e, 32'sh3ea33a9b, 32'sh3ea2e80e, 32'sh3ea29578, 32'sh3ea242d9, 
               32'sh3ea1f02f, 32'sh3ea19d7c, 32'sh3ea14abf, 32'sh3ea0f7f9, 32'sh3ea0a529, 32'sh3ea0524f, 32'sh3e9fff6b, 32'sh3e9fac7e, 
               32'sh3e9f5988, 32'sh3e9f0687, 32'sh3e9eb37d, 32'sh3e9e6069, 32'sh3e9e0d4c, 32'sh3e9dba25, 32'sh3e9d66f4, 32'sh3e9d13ba, 
               32'sh3e9cc076, 32'sh3e9c6d28, 32'sh3e9c19d1, 32'sh3e9bc670, 32'sh3e9b7306, 32'sh3e9b1f91, 32'sh3e9acc13, 32'sh3e9a788c, 
               32'sh3e9a24fb, 32'sh3e99d160, 32'sh3e997dbb, 32'sh3e992a0d, 32'sh3e98d655, 32'sh3e988294, 32'sh3e982ec9, 32'sh3e97daf4, 
               32'sh3e978715, 32'sh3e97332d, 32'sh3e96df3b, 32'sh3e968b40, 32'sh3e96373b, 32'sh3e95e32c, 32'sh3e958f14, 32'sh3e953af2, 
               32'sh3e94e6c6, 32'sh3e949291, 32'sh3e943e52, 32'sh3e93ea09, 32'sh3e9395b7, 32'sh3e93415b, 32'sh3e92ecf6, 32'sh3e929886, 
               32'sh3e92440d, 32'sh3e91ef8b, 32'sh3e919aff, 32'sh3e914669, 32'sh3e90f1ca, 32'sh3e909d20, 32'sh3e90486e, 32'sh3e8ff3b1, 
               32'sh3e8f9eeb, 32'sh3e8f4a1b, 32'sh3e8ef542, 32'sh3e8ea05f, 32'sh3e8e4b72, 32'sh3e8df67c, 32'sh3e8da17c, 32'sh3e8d4c73, 
               32'sh3e8cf75f, 32'sh3e8ca243, 32'sh3e8c4d1c, 32'sh3e8bf7ec, 32'sh3e8ba2b2, 32'sh3e8b4d6f, 32'sh3e8af821, 32'sh3e8aa2cb, 
               32'sh3e8a4d6a, 32'sh3e89f800, 32'sh3e89a28d, 32'sh3e894d0f, 32'sh3e88f788, 32'sh3e88a1f8, 32'sh3e884c5d, 32'sh3e87f6ba, 
               32'sh3e87a10c, 32'sh3e874b55, 32'sh3e86f594, 32'sh3e869fca, 32'sh3e8649f5, 32'sh3e85f418, 32'sh3e859e30, 32'sh3e85483f, 
               32'sh3e84f245, 32'sh3e849c40, 32'sh3e844632, 32'sh3e83f01b, 32'sh3e8399f9, 32'sh3e8343ce, 32'sh3e82ed9a, 32'sh3e82975c, 
               32'sh3e824114, 32'sh3e81eac3, 32'sh3e819467, 32'sh3e813e03, 32'sh3e80e794, 32'sh3e80911c, 32'sh3e803a9b, 32'sh3e7fe40f, 
               32'sh3e7f8d7b, 32'sh3e7f36dc, 32'sh3e7ee034, 32'sh3e7e8982, 32'sh3e7e32c6, 32'sh3e7ddc01, 32'sh3e7d8533, 32'sh3e7d2e5a, 
               32'sh3e7cd778, 32'sh3e7c808d, 32'sh3e7c2997, 32'sh3e7bd298, 32'sh3e7b7b90, 32'sh3e7b247e, 32'sh3e7acd62, 32'sh3e7a763c, 
               32'sh3e7a1f0d, 32'sh3e79c7d4, 32'sh3e797092, 32'sh3e791946, 32'sh3e78c1f0, 32'sh3e786a91, 32'sh3e781328, 32'sh3e77bbb6, 
               32'sh3e77643a, 32'sh3e770cb4, 32'sh3e76b524, 32'sh3e765d8b, 32'sh3e7605e9, 32'sh3e75ae3c, 32'sh3e755686, 32'sh3e74fec7, 
               32'sh3e74a6fd, 32'sh3e744f2b, 32'sh3e73f74e, 32'sh3e739f68, 32'sh3e734778, 32'sh3e72ef7f, 32'sh3e72977c, 32'sh3e723f6f, 
               32'sh3e71e759, 32'sh3e718f39, 32'sh3e71370f, 32'sh3e70dedc, 32'sh3e70869f, 32'sh3e702e59, 32'sh3e6fd609, 32'sh3e6f7daf, 
               32'sh3e6f254c, 32'sh3e6eccdf, 32'sh3e6e7468, 32'sh3e6e1be8, 32'sh3e6dc35e, 32'sh3e6d6acb, 32'sh3e6d122e, 32'sh3e6cb987, 
               32'sh3e6c60d7, 32'sh3e6c081d, 32'sh3e6baf59, 32'sh3e6b568c, 32'sh3e6afdb5, 32'sh3e6aa4d5, 32'sh3e6a4beb, 32'sh3e69f2f7, 
               32'sh3e6999fa, 32'sh3e6940f3, 32'sh3e68e7e2, 32'sh3e688ec8, 32'sh3e6835a4, 32'sh3e67dc77, 32'sh3e67833f, 32'sh3e6729ff, 
               32'sh3e66d0b4, 32'sh3e667761, 32'sh3e661e03, 32'sh3e65c49c, 32'sh3e656b2b, 32'sh3e6511b0, 32'sh3e64b82c, 32'sh3e645e9f, 
               32'sh3e640507, 32'sh3e63ab66, 32'sh3e6351bc, 32'sh3e62f808, 32'sh3e629e4a, 32'sh3e624483, 32'sh3e61eab2, 32'sh3e6190d7, 
               32'sh3e6136f3, 32'sh3e60dd05, 32'sh3e60830d, 32'sh3e60290c, 32'sh3e5fcf01, 32'sh3e5f74ed, 32'sh3e5f1acf, 32'sh3e5ec0a7, 
               32'sh3e5e6676, 32'sh3e5e0c3b, 32'sh3e5db1f7, 32'sh3e5d57a9, 32'sh3e5cfd51, 32'sh3e5ca2f0, 32'sh3e5c4885, 32'sh3e5bee10, 
               32'sh3e5b9392, 32'sh3e5b390a, 32'sh3e5ade79, 32'sh3e5a83de, 32'sh3e5a2939, 32'sh3e59ce8b, 32'sh3e5973d3, 32'sh3e591912, 
               32'sh3e58be47, 32'sh3e586372, 32'sh3e580894, 32'sh3e57adac, 32'sh3e5752ba, 32'sh3e56f7bf, 32'sh3e569cba, 32'sh3e5641ac, 
               32'sh3e55e694, 32'sh3e558b72, 32'sh3e553047, 32'sh3e54d512, 32'sh3e5479d4, 32'sh3e541e8c, 32'sh3e53c33a, 32'sh3e5367df, 
               32'sh3e530c7a, 32'sh3e52b10b, 32'sh3e525593, 32'sh3e51fa11, 32'sh3e519e86, 32'sh3e5142f1, 32'sh3e50e752, 32'sh3e508baa, 
               32'sh3e502ff9, 32'sh3e4fd43d, 32'sh3e4f7878, 32'sh3e4f1caa, 32'sh3e4ec0d1, 32'sh3e4e64f0, 32'sh3e4e0904, 32'sh3e4dad0f, 
               32'sh3e4d5110, 32'sh3e4cf508, 32'sh3e4c98f6, 32'sh3e4c3cdb, 32'sh3e4be0b6, 32'sh3e4b8487, 32'sh3e4b284f, 32'sh3e4acc0d, 
               32'sh3e4a6fc1, 32'sh3e4a136c, 32'sh3e49b70d, 32'sh3e495aa5, 32'sh3e48fe33, 32'sh3e48a1b8, 32'sh3e484533, 32'sh3e47e8a4, 
               32'sh3e478c0b, 32'sh3e472f69, 32'sh3e46d2be, 32'sh3e467609, 32'sh3e46194a, 32'sh3e45bc82, 32'sh3e455fb0, 32'sh3e4502d4, 
               32'sh3e44a5ef, 32'sh3e444900, 32'sh3e43ec08, 32'sh3e438f06, 32'sh3e4331fa, 32'sh3e42d4e5, 32'sh3e4277c6, 32'sh3e421a9e, 
               32'sh3e41bd6c, 32'sh3e416030, 32'sh3e4102eb, 32'sh3e40a59c, 32'sh3e404844, 32'sh3e3feae2, 32'sh3e3f8d76, 32'sh3e3f3001, 
               32'sh3e3ed282, 32'sh3e3e74fa, 32'sh3e3e1768, 32'sh3e3db9cc, 32'sh3e3d5c27, 32'sh3e3cfe78, 32'sh3e3ca0c0, 32'sh3e3c42fe, 
               32'sh3e3be532, 32'sh3e3b875d, 32'sh3e3b297e, 32'sh3e3acb96, 32'sh3e3a6da4, 32'sh3e3a0fa9, 32'sh3e39b1a3, 32'sh3e395395, 
               32'sh3e38f57c, 32'sh3e38975a, 32'sh3e38392f, 32'sh3e37dafa, 32'sh3e377cbb, 32'sh3e371e73, 32'sh3e36c021, 32'sh3e3661c5, 
               32'sh3e360360, 32'sh3e35a4f1, 32'sh3e354679, 32'sh3e34e7f7, 32'sh3e34896c, 32'sh3e342ad7, 32'sh3e33cc38, 32'sh3e336d90, 
               32'sh3e330ede, 32'sh3e32b022, 32'sh3e32515d, 32'sh3e31f28f, 32'sh3e3193b7, 32'sh3e3134d5, 32'sh3e30d5e9, 32'sh3e3076f4, 
               32'sh3e3017f6, 32'sh3e2fb8ee, 32'sh3e2f59dc, 32'sh3e2efac1, 32'sh3e2e9b9c, 32'sh3e2e3c6d, 32'sh3e2ddd35, 32'sh3e2d7df3, 
               32'sh3e2d1ea8, 32'sh3e2cbf53, 32'sh3e2c5ff5, 32'sh3e2c008d, 32'sh3e2ba11b, 32'sh3e2b41a0, 32'sh3e2ae21b, 32'sh3e2a828c, 
               32'sh3e2a22f4, 32'sh3e29c353, 32'sh3e2963a8, 32'sh3e2903f3, 32'sh3e28a435, 32'sh3e28446d, 32'sh3e27e49b, 32'sh3e2784c0, 
               32'sh3e2724db, 32'sh3e26c4ed, 32'sh3e2664f5, 32'sh3e2604f4, 32'sh3e25a4e9, 32'sh3e2544d4, 32'sh3e24e4b6, 32'sh3e24848e, 
               32'sh3e24245d, 32'sh3e23c422, 32'sh3e2363dd, 32'sh3e23038f, 32'sh3e22a338, 32'sh3e2242d6, 32'sh3e21e26c, 32'sh3e2181f7, 
               32'sh3e212179, 32'sh3e20c0f1, 32'sh3e206060, 32'sh3e1fffc6, 32'sh3e1f9f21, 32'sh3e1f3e73, 32'sh3e1eddbc, 32'sh3e1e7cfb, 
               32'sh3e1e1c30, 32'sh3e1dbb5c, 32'sh3e1d5a7e, 32'sh3e1cf997, 32'sh3e1c98a6, 32'sh3e1c37ab, 32'sh3e1bd6a7, 32'sh3e1b7599, 
               32'sh3e1b1482, 32'sh3e1ab361, 32'sh3e1a5237, 32'sh3e19f103, 32'sh3e198fc5, 32'sh3e192e7e, 32'sh3e18cd2d, 32'sh3e186bd3, 
               32'sh3e180a6f, 32'sh3e17a902, 32'sh3e17478a, 32'sh3e16e60a, 32'sh3e168480, 32'sh3e1622ec, 32'sh3e15c14f, 32'sh3e155fa8, 
               32'sh3e14fdf7, 32'sh3e149c3d, 32'sh3e143a79, 32'sh3e13d8ac, 32'sh3e1376d5, 32'sh3e1314f5, 32'sh3e12b30b, 32'sh3e125118, 
               32'sh3e11ef1b, 32'sh3e118d14, 32'sh3e112b04, 32'sh3e10c8ea, 32'sh3e1066c7, 32'sh3e10049a, 32'sh3e0fa263, 32'sh3e0f4023, 
               32'sh3e0eddd9, 32'sh3e0e7b86, 32'sh3e0e1929, 32'sh3e0db6c3, 32'sh3e0d5453, 32'sh3e0cf1da, 32'sh3e0c8f57, 32'sh3e0c2cca, 
               32'sh3e0bca34, 32'sh3e0b6794, 32'sh3e0b04eb, 32'sh3e0aa238, 32'sh3e0a3f7b, 32'sh3e09dcb5, 32'sh3e0979e6, 32'sh3e09170c, 
               32'sh3e08b42a, 32'sh3e08513d, 32'sh3e07ee47, 32'sh3e078b48, 32'sh3e07283f, 32'sh3e06c52c, 32'sh3e066210, 32'sh3e05feeb, 
               32'sh3e059bbb, 32'sh3e053882, 32'sh3e04d540, 32'sh3e0471f4, 32'sh3e040e9f, 32'sh3e03ab40, 32'sh3e0347d7, 32'sh3e02e465, 
               32'sh3e0280e9, 32'sh3e021d64, 32'sh3e01b9d5, 32'sh3e01563c, 32'sh3e00f29a, 32'sh3e008eef, 32'sh3e002b39, 32'sh3dffc77b, 
               32'sh3dff63b2, 32'sh3dfeffe1, 32'sh3dfe9c05, 32'sh3dfe3820, 32'sh3dfdd432, 32'sh3dfd703a, 32'sh3dfd0c38, 32'sh3dfca82d, 
               32'sh3dfc4418, 32'sh3dfbdffa, 32'sh3dfb7bd2, 32'sh3dfb17a0, 32'sh3dfab365, 32'sh3dfa4f21, 32'sh3df9ead3, 32'sh3df9867b, 
               32'sh3df9221a, 32'sh3df8bdaf, 32'sh3df8593b, 32'sh3df7f4bd, 32'sh3df79036, 32'sh3df72ba5, 32'sh3df6c70a, 32'sh3df66266, 
               32'sh3df5fdb8, 32'sh3df59901, 32'sh3df53440, 32'sh3df4cf76, 32'sh3df46aa2, 32'sh3df405c5, 32'sh3df3a0de, 32'sh3df33bed, 
               32'sh3df2d6f3, 32'sh3df271ef, 32'sh3df20ce2, 32'sh3df1a7cb, 32'sh3df142ab, 32'sh3df0dd81, 32'sh3df0784e, 32'sh3df01311, 
               32'sh3defadca, 32'sh3def487a, 32'sh3deee321, 32'sh3dee7dbd, 32'sh3dee1851, 32'sh3dedb2da, 32'sh3ded4d5b, 32'sh3dece7d1, 
               32'sh3dec823e, 32'sh3dec1ca2, 32'sh3debb6fc, 32'sh3deb514c, 32'sh3deaeb93, 32'sh3dea85d0, 32'sh3dea2004, 32'sh3de9ba2e, 
               32'sh3de9544f, 32'sh3de8ee66, 32'sh3de88874, 32'sh3de82278, 32'sh3de7bc72, 32'sh3de75663, 32'sh3de6f04b, 32'sh3de68a29, 
               32'sh3de623fd, 32'sh3de5bdc8, 32'sh3de55789, 32'sh3de4f141, 32'sh3de48aef, 32'sh3de42493, 32'sh3de3be2e, 32'sh3de357c0, 
               32'sh3de2f148, 32'sh3de28ac6, 32'sh3de2243b, 32'sh3de1bda6, 32'sh3de15708, 32'sh3de0f060, 32'sh3de089af, 32'sh3de022f4, 
               32'sh3ddfbc30, 32'sh3ddf5562, 32'sh3ddeee8a, 32'sh3dde87a9, 32'sh3dde20bf, 32'sh3dddb9cb, 32'sh3ddd52cd, 32'sh3ddcebc6, 
               32'sh3ddc84b5, 32'sh3ddc1d9b, 32'sh3ddbb677, 32'sh3ddb4f4a, 32'sh3ddae813, 32'sh3dda80d3, 32'sh3dda1989, 32'sh3dd9b235, 
               32'sh3dd94ad8, 32'sh3dd8e372, 32'sh3dd87c02, 32'sh3dd81488, 32'sh3dd7ad05, 32'sh3dd74578, 32'sh3dd6dde2, 32'sh3dd67642, 
               32'sh3dd60e99, 32'sh3dd5a6e6, 32'sh3dd53f29, 32'sh3dd4d763, 32'sh3dd46f94, 32'sh3dd407bb, 32'sh3dd39fd8, 32'sh3dd337ec, 
               32'sh3dd2cff7, 32'sh3dd267f8, 32'sh3dd1ffef, 32'sh3dd197dd, 32'sh3dd12fc1, 32'sh3dd0c79c, 32'sh3dd05f6d, 32'sh3dcff735, 
               32'sh3dcf8ef3, 32'sh3dcf26a7, 32'sh3dcebe52, 32'sh3dce55f4, 32'sh3dcded8c, 32'sh3dcd851a, 32'sh3dcd1c9f, 32'sh3dccb41b, 
               32'sh3dcc4b8d, 32'sh3dcbe2f5, 32'sh3dcb7a54, 32'sh3dcb11a9, 32'sh3dcaa8f5, 32'sh3dca4037, 32'sh3dc9d770, 32'sh3dc96e9f, 
               32'sh3dc905c5, 32'sh3dc89ce1, 32'sh3dc833f3, 32'sh3dc7cafc, 32'sh3dc761fc, 32'sh3dc6f8f2, 32'sh3dc68fdf, 32'sh3dc626c1, 
               32'sh3dc5bd9b, 32'sh3dc5546b, 32'sh3dc4eb31, 32'sh3dc481ee, 32'sh3dc418a1, 32'sh3dc3af4b, 32'sh3dc345eb, 32'sh3dc2dc82, 
               32'sh3dc2730f, 32'sh3dc20993, 32'sh3dc1a00d, 32'sh3dc1367e, 32'sh3dc0cce5, 32'sh3dc06343, 32'sh3dbff997, 32'sh3dbf8fe1, 
               32'sh3dbf2622, 32'sh3dbebc5a, 32'sh3dbe5288, 32'sh3dbde8ac, 32'sh3dbd7ec7, 32'sh3dbd14d9, 32'sh3dbcaae1, 32'sh3dbc40df, 
               32'sh3dbbd6d4, 32'sh3dbb6cbf, 32'sh3dbb02a1, 32'sh3dba987a, 32'sh3dba2e48, 32'sh3db9c40e, 32'sh3db959c9, 32'sh3db8ef7c, 
               32'sh3db88524, 32'sh3db81ac4, 32'sh3db7b059, 32'sh3db745e5, 32'sh3db6db68, 32'sh3db670e1, 32'sh3db60651, 32'sh3db59bb7, 
               32'sh3db53113, 32'sh3db4c667, 32'sh3db45bb0, 32'sh3db3f0f0, 32'sh3db38627, 32'sh3db31b54, 32'sh3db2b077, 32'sh3db24591, 
               32'sh3db1daa2, 32'sh3db16fa9, 32'sh3db104a6, 32'sh3db0999a, 32'sh3db02e84, 32'sh3dafc365, 32'sh3daf583d, 32'sh3daeed0a, 
               32'sh3dae81cf, 32'sh3dae168a, 32'sh3dadab3b, 32'sh3dad3fe3, 32'sh3dacd481, 32'sh3dac6916, 32'sh3dabfda1, 32'sh3dab9223, 
               32'sh3dab269b, 32'sh3daabb0a, 32'sh3daa4f6f, 32'sh3da9e3cb, 32'sh3da9781d, 32'sh3da90c66, 32'sh3da8a0a5, 32'sh3da834db, 
               32'sh3da7c907, 32'sh3da75d2a, 32'sh3da6f143, 32'sh3da68553, 32'sh3da61959, 32'sh3da5ad55, 32'sh3da54149, 32'sh3da4d532, 
               32'sh3da46912, 32'sh3da3fce9, 32'sh3da390b6, 32'sh3da3247a, 32'sh3da2b834, 32'sh3da24be4, 32'sh3da1df8c, 32'sh3da17329, 
               32'sh3da106bd, 32'sh3da09a48, 32'sh3da02dc9, 32'sh3d9fc140, 32'sh3d9f54af, 32'sh3d9ee813, 32'sh3d9e7b6e, 32'sh3d9e0ec0, 
               32'sh3d9da208, 32'sh3d9d3546, 32'sh3d9cc87b, 32'sh3d9c5ba7, 32'sh3d9beec9, 32'sh3d9b81e2, 32'sh3d9b14f1, 32'sh3d9aa7f6, 
               32'sh3d9a3af2, 32'sh3d99cde5, 32'sh3d9960ce, 32'sh3d98f3ae, 32'sh3d988684, 32'sh3d981950, 32'sh3d97ac13, 32'sh3d973ecd, 
               32'sh3d96d17d, 32'sh3d966423, 32'sh3d95f6c1, 32'sh3d958954, 32'sh3d951bde, 32'sh3d94ae5f, 32'sh3d9440d6, 32'sh3d93d343, 
               32'sh3d9365a8, 32'sh3d92f802, 32'sh3d928a53, 32'sh3d921c9b, 32'sh3d91aed9, 32'sh3d91410e, 32'sh3d90d339, 32'sh3d90655a, 
               32'sh3d8ff772, 32'sh3d8f8981, 32'sh3d8f1b86, 32'sh3d8ead82, 32'sh3d8e3f74, 32'sh3d8dd15d, 32'sh3d8d633c, 32'sh3d8cf512, 
               32'sh3d8c86de, 32'sh3d8c18a0, 32'sh3d8baa5a, 32'sh3d8b3c09, 32'sh3d8acdb0, 32'sh3d8a5f4c, 32'sh3d89f0e0, 32'sh3d898269, 
               32'sh3d8913ea, 32'sh3d88a560, 32'sh3d8836ce, 32'sh3d87c832, 32'sh3d87598c, 32'sh3d86eadd, 32'sh3d867c24, 32'sh3d860d62, 
               32'sh3d859e96, 32'sh3d852fc1, 32'sh3d84c0e2, 32'sh3d8451fa, 32'sh3d83e309, 32'sh3d83740e, 32'sh3d830509, 32'sh3d8295fb, 
               32'sh3d8226e4, 32'sh3d81b7c3, 32'sh3d814898, 32'sh3d80d964, 32'sh3d806a27, 32'sh3d7ffae0, 32'sh3d7f8b8f, 32'sh3d7f1c35, 
               32'sh3d7eacd2, 32'sh3d7e3d65, 32'sh3d7dcdef, 32'sh3d7d5e6f, 32'sh3d7ceee5, 32'sh3d7c7f53, 32'sh3d7c0fb6, 32'sh3d7ba010, 
               32'sh3d7b3061, 32'sh3d7ac0a8, 32'sh3d7a50e6, 32'sh3d79e11a, 32'sh3d797145, 32'sh3d790167, 32'sh3d78917e, 32'sh3d78218d, 
               32'sh3d77b192, 32'sh3d77418d, 32'sh3d76d17f, 32'sh3d766168, 32'sh3d75f147, 32'sh3d75811c, 32'sh3d7510e8, 32'sh3d74a0ab, 
               32'sh3d743064, 32'sh3d73c013, 32'sh3d734fb9, 32'sh3d72df56, 32'sh3d726ee9, 32'sh3d71fe73, 32'sh3d718df3, 32'sh3d711d6a, 
               32'sh3d70acd7, 32'sh3d703c3b, 32'sh3d6fcb95, 32'sh3d6f5ae6, 32'sh3d6eea2d, 32'sh3d6e796b, 32'sh3d6e08a0, 32'sh3d6d97cb, 
               32'sh3d6d26ec, 32'sh3d6cb604, 32'sh3d6c4513, 32'sh3d6bd418, 32'sh3d6b6313, 32'sh3d6af205, 32'sh3d6a80ee, 32'sh3d6a0fcd, 
               32'sh3d699ea3, 32'sh3d692d6f, 32'sh3d68bc32, 32'sh3d684aeb, 32'sh3d67d99b, 32'sh3d676841, 32'sh3d66f6de, 32'sh3d668571, 
               32'sh3d6613fb, 32'sh3d65a27c, 32'sh3d6530f3, 32'sh3d64bf60, 32'sh3d644dc4, 32'sh3d63dc1f, 32'sh3d636a70, 32'sh3d62f8b8, 
               32'sh3d6286f6, 32'sh3d62152b, 32'sh3d61a356, 32'sh3d613178, 32'sh3d60bf90, 32'sh3d604d9f, 32'sh3d5fdba4, 32'sh3d5f69a0, 
               32'sh3d5ef793, 32'sh3d5e857c, 32'sh3d5e135b, 32'sh3d5da131, 32'sh3d5d2efe, 32'sh3d5cbcc1, 32'sh3d5c4a7b, 32'sh3d5bd82b, 
               32'sh3d5b65d2, 32'sh3d5af36f, 32'sh3d5a8103, 32'sh3d5a0e8d, 32'sh3d599c0e, 32'sh3d592986, 32'sh3d58b6f4, 32'sh3d584458, 
               32'sh3d57d1b3, 32'sh3d575f05, 32'sh3d56ec4d, 32'sh3d56798c, 32'sh3d5606c1, 32'sh3d5593ed, 32'sh3d55210f, 32'sh3d54ae28, 
               32'sh3d543b37, 32'sh3d53c83d, 32'sh3d53553a, 32'sh3d52e22d, 32'sh3d526f16, 32'sh3d51fbf7, 32'sh3d5188cd, 32'sh3d51159a, 
               32'sh3d50a25e, 32'sh3d502f18, 32'sh3d4fbbc9, 32'sh3d4f4871, 32'sh3d4ed50f, 32'sh3d4e61a3, 32'sh3d4dee2e, 32'sh3d4d7ab0, 
               32'sh3d4d0728, 32'sh3d4c9396, 32'sh3d4c1ffc, 32'sh3d4bac57, 32'sh3d4b38aa, 32'sh3d4ac4f3, 32'sh3d4a5132, 32'sh3d49dd68, 
               32'sh3d496994, 32'sh3d48f5b7, 32'sh3d4881d1, 32'sh3d480de1, 32'sh3d4799e8, 32'sh3d4725e5, 32'sh3d46b1d9, 32'sh3d463dc3, 
               32'sh3d45c9a4, 32'sh3d45557c, 32'sh3d44e14a, 32'sh3d446d0e, 32'sh3d43f8c9, 32'sh3d43847b, 32'sh3d431023, 32'sh3d429bc2, 
               32'sh3d422757, 32'sh3d41b2e3, 32'sh3d413e65, 32'sh3d40c9de, 32'sh3d40554e, 32'sh3d3fe0b4, 32'sh3d3f6c11, 32'sh3d3ef764, 
               32'sh3d3e82ae, 32'sh3d3e0dee, 32'sh3d3d9925, 32'sh3d3d2452, 32'sh3d3caf76, 32'sh3d3c3a91, 32'sh3d3bc5a2, 32'sh3d3b50a9, 
               32'sh3d3adba7, 32'sh3d3a669c, 32'sh3d39f188, 32'sh3d397c69, 32'sh3d390742, 32'sh3d389211, 32'sh3d381cd6, 32'sh3d37a792, 
               32'sh3d373245, 32'sh3d36bcee, 32'sh3d36478e, 32'sh3d35d224, 32'sh3d355cb1, 32'sh3d34e735, 32'sh3d3471af, 32'sh3d33fc1f, 
               32'sh3d338687, 32'sh3d3310e4, 32'sh3d329b39, 32'sh3d322583, 32'sh3d31afc5, 32'sh3d3139fd, 32'sh3d30c42b, 32'sh3d304e50, 
               32'sh3d2fd86c, 32'sh3d2f627e, 32'sh3d2eec87, 32'sh3d2e7686, 32'sh3d2e007c, 32'sh3d2d8a69, 32'sh3d2d144c, 32'sh3d2c9e25, 
               32'sh3d2c27f6, 32'sh3d2bb1bc, 32'sh3d2b3b7a, 32'sh3d2ac52d, 32'sh3d2a4ed8, 32'sh3d29d879, 32'sh3d296210, 32'sh3d28eb9f, 
               32'sh3d287523, 32'sh3d27fe9f, 32'sh3d278810, 32'sh3d271179, 32'sh3d269ad8, 32'sh3d26242d, 32'sh3d25ad7a, 32'sh3d2536bc, 
               32'sh3d24bff6, 32'sh3d244925, 32'sh3d23d24c, 32'sh3d235b69, 32'sh3d22e47c, 32'sh3d226d86, 32'sh3d21f687, 32'sh3d217f7e, 
               32'sh3d21086c, 32'sh3d209151, 32'sh3d201a2c, 32'sh3d1fa2fd, 32'sh3d1f2bc5, 32'sh3d1eb484, 32'sh3d1e3d39, 32'sh3d1dc5e5, 
               32'sh3d1d4e88, 32'sh3d1cd721, 32'sh3d1c5fb0, 32'sh3d1be836, 32'sh3d1b70b3, 32'sh3d1af926, 32'sh3d1a8190, 32'sh3d1a09f1, 
               32'sh3d199248, 32'sh3d191a95, 32'sh3d18a2da, 32'sh3d182b14, 32'sh3d17b346, 32'sh3d173b6e, 32'sh3d16c38c, 32'sh3d164ba1, 
               32'sh3d15d3ad, 32'sh3d155baf, 32'sh3d14e3a8, 32'sh3d146b98, 32'sh3d13f37e, 32'sh3d137b5a, 32'sh3d13032d, 32'sh3d128af7, 
               32'sh3d1212b7, 32'sh3d119a6e, 32'sh3d11221c, 32'sh3d10a9c0, 32'sh3d10315a, 32'sh3d0fb8ec, 32'sh3d0f4074, 32'sh3d0ec7f2, 
               32'sh3d0e4f67, 32'sh3d0dd6d2, 32'sh3d0d5e35, 32'sh3d0ce58d, 32'sh3d0c6cdd, 32'sh3d0bf423, 32'sh3d0b7b5f, 32'sh3d0b0292, 
               32'sh3d0a89bc, 32'sh3d0a10dc, 32'sh3d0997f3, 32'sh3d091f00, 32'sh3d08a604, 32'sh3d082cff, 32'sh3d07b3f0, 32'sh3d073ad8, 
               32'sh3d06c1b6, 32'sh3d06488b, 32'sh3d05cf57, 32'sh3d055619, 32'sh3d04dcd2, 32'sh3d046381, 32'sh3d03ea27, 32'sh3d0370c4, 
               32'sh3d02f757, 32'sh3d027de0, 32'sh3d020461, 32'sh3d018ad7, 32'sh3d011145, 32'sh3d0097a9, 32'sh3d001e04, 32'sh3cffa455, 
               32'sh3cff2a9d, 32'sh3cfeb0db, 32'sh3cfe3710, 32'sh3cfdbd3c, 32'sh3cfd435e, 32'sh3cfcc977, 32'sh3cfc4f86, 32'sh3cfbd58c, 
               32'sh3cfb5b89, 32'sh3cfae17c, 32'sh3cfa6766, 32'sh3cf9ed46, 32'sh3cf9731d, 32'sh3cf8f8eb, 32'sh3cf87eaf, 32'sh3cf80469, 
               32'sh3cf78a1b, 32'sh3cf70fc3, 32'sh3cf69561, 32'sh3cf61af7, 32'sh3cf5a082, 32'sh3cf52605, 32'sh3cf4ab7e, 32'sh3cf430ed, 
               32'sh3cf3b653, 32'sh3cf33bb0, 32'sh3cf2c103, 32'sh3cf2464d, 32'sh3cf1cb8e, 32'sh3cf150c5, 32'sh3cf0d5f3, 32'sh3cf05b17, 
               32'sh3cefe032, 32'sh3cef6544, 32'sh3ceeea4c, 32'sh3cee6f4b, 32'sh3cedf440, 32'sh3ced792c, 32'sh3cecfe0f, 32'sh3cec82e8, 
               32'sh3cec07b8, 32'sh3ceb8c7e, 32'sh3ceb113b, 32'sh3cea95ef, 32'sh3cea1a99, 32'sh3ce99f3a, 32'sh3ce923d1, 32'sh3ce8a85f, 
               32'sh3ce82ce4, 32'sh3ce7b15f, 32'sh3ce735d1, 32'sh3ce6ba39, 32'sh3ce63e98, 32'sh3ce5c2ee, 32'sh3ce5473a, 32'sh3ce4cb7d, 
               32'sh3ce44fb7, 32'sh3ce3d3e7, 32'sh3ce3580e, 32'sh3ce2dc2b, 32'sh3ce2603f, 32'sh3ce1e44a, 32'sh3ce1684b, 32'sh3ce0ec43, 
               32'sh3ce07031, 32'sh3cdff416, 32'sh3cdf77f2, 32'sh3cdefbc4, 32'sh3cde7f8d, 32'sh3cde034c, 32'sh3cdd8702, 32'sh3cdd0aaf, 
               32'sh3cdc8e52, 32'sh3cdc11ec, 32'sh3cdb957d, 32'sh3cdb1904, 32'sh3cda9c81, 32'sh3cda1ff6, 32'sh3cd9a361, 32'sh3cd926c2, 
               32'sh3cd8aa1b, 32'sh3cd82d6a, 32'sh3cd7b0af, 32'sh3cd733eb, 32'sh3cd6b71e, 32'sh3cd63a47, 32'sh3cd5bd67, 32'sh3cd5407e, 
               32'sh3cd4c38b, 32'sh3cd4468f, 32'sh3cd3c989, 32'sh3cd34c7a, 32'sh3cd2cf62, 32'sh3cd25240, 32'sh3cd1d515, 32'sh3cd157e0, 
               32'sh3cd0daa2, 32'sh3cd05d5b, 32'sh3ccfe00b, 32'sh3ccf62b0, 32'sh3ccee54d, 32'sh3cce67e0, 32'sh3ccdea6a, 32'sh3ccd6ceb, 
               32'sh3cccef62, 32'sh3ccc71d0, 32'sh3ccbf434, 32'sh3ccb768f, 32'sh3ccaf8e0, 32'sh3cca7b29, 32'sh3cc9fd68, 32'sh3cc97f9d, 
               32'sh3cc901c9, 32'sh3cc883ec, 32'sh3cc80605, 32'sh3cc78815, 32'sh3cc70a1c, 32'sh3cc68c19, 32'sh3cc60e0d, 32'sh3cc58ff7, 
               32'sh3cc511d9, 32'sh3cc493b0, 32'sh3cc4157f, 32'sh3cc39744, 32'sh3cc318ff, 32'sh3cc29ab2, 32'sh3cc21c5b, 32'sh3cc19dfa, 
               32'sh3cc11f90, 32'sh3cc0a11d, 32'sh3cc022a0, 32'sh3cbfa41a, 32'sh3cbf258b, 32'sh3cbea6f2, 32'sh3cbe2850, 32'sh3cbda9a5, 
               32'sh3cbd2af0, 32'sh3cbcac32, 32'sh3cbc2d6b, 32'sh3cbbae9a, 32'sh3cbb2fbf, 32'sh3cbab0dc, 32'sh3cba31ef, 32'sh3cb9b2f9, 
               32'sh3cb933f9, 32'sh3cb8b4f0, 32'sh3cb835dd, 32'sh3cb7b6c1, 32'sh3cb7379c, 32'sh3cb6b86e, 32'sh3cb63936, 32'sh3cb5b9f5, 
               32'sh3cb53aaa, 32'sh3cb4bb56, 32'sh3cb43bf9, 32'sh3cb3bc92, 32'sh3cb33d22, 32'sh3cb2bda9, 32'sh3cb23e26, 32'sh3cb1be9a, 
               32'sh3cb13f04, 32'sh3cb0bf65, 32'sh3cb03fbd, 32'sh3cafc00b, 32'sh3caf4051, 32'sh3caec08c, 32'sh3cae40bf, 32'sh3cadc0e8, 
               32'sh3cad4107, 32'sh3cacc11d, 32'sh3cac412a, 32'sh3cabc12e, 32'sh3cab4128, 32'sh3caac119, 32'sh3caa4100, 32'sh3ca9c0df, 
               32'sh3ca940b3, 32'sh3ca8c07f, 32'sh3ca84041, 32'sh3ca7bffa, 32'sh3ca73fa9, 32'sh3ca6bf4f, 32'sh3ca63eec, 32'sh3ca5be7f, 
               32'sh3ca53e09, 32'sh3ca4bd89, 32'sh3ca43d01, 32'sh3ca3bc6f, 32'sh3ca33bd3, 32'sh3ca2bb2e, 32'sh3ca23a80, 32'sh3ca1b9c9, 
               32'sh3ca13908, 32'sh3ca0b83e, 32'sh3ca0376a, 32'sh3c9fb68d, 32'sh3c9f35a7, 32'sh3c9eb4b7, 32'sh3c9e33be, 32'sh3c9db2bc, 
               32'sh3c9d31b0, 32'sh3c9cb09b, 32'sh3c9c2f7d, 32'sh3c9bae55, 32'sh3c9b2d24, 32'sh3c9aabea, 32'sh3c9a2aa6, 32'sh3c99a959, 
               32'sh3c992803, 32'sh3c98a6a3, 32'sh3c98253a, 32'sh3c97a3c7, 32'sh3c97224c, 32'sh3c96a0c6, 32'sh3c961f38, 32'sh3c959da0, 
               32'sh3c951bff, 32'sh3c949a55, 32'sh3c9418a1, 32'sh3c9396e3, 32'sh3c93151d, 32'sh3c92934d, 32'sh3c921174, 32'sh3c918f91, 
               32'sh3c910da5, 32'sh3c908bb0, 32'sh3c9009b2, 32'sh3c8f87aa, 32'sh3c8f0598, 32'sh3c8e837e, 32'sh3c8e015a, 32'sh3c8d7f2d, 
               32'sh3c8cfcf6, 32'sh3c8c7ab6, 32'sh3c8bf86d, 32'sh3c8b761a, 32'sh3c8af3be, 32'sh3c8a7159, 32'sh3c89eeea, 32'sh3c896c72, 
               32'sh3c88e9f1, 32'sh3c886766, 32'sh3c87e4d2, 32'sh3c876235, 32'sh3c86df8e, 32'sh3c865cde, 32'sh3c85da25, 32'sh3c855762, 
               32'sh3c84d496, 32'sh3c8451c1, 32'sh3c83cee2, 32'sh3c834bfa, 32'sh3c82c909, 32'sh3c82460e, 32'sh3c81c30a, 32'sh3c813ffd, 
               32'sh3c80bce7, 32'sh3c8039c7, 32'sh3c7fb69d, 32'sh3c7f336b, 32'sh3c7eb02f, 32'sh3c7e2ce9, 32'sh3c7da99b, 32'sh3c7d2643, 
               32'sh3c7ca2e2, 32'sh3c7c1f77, 32'sh3c7b9c03, 32'sh3c7b1886, 32'sh3c7a94ff, 32'sh3c7a116f, 32'sh3c798dd6, 32'sh3c790a34, 
               32'sh3c788688, 32'sh3c7802d2, 32'sh3c777f14, 32'sh3c76fb4c, 32'sh3c76777b, 32'sh3c75f3a0, 32'sh3c756fbd, 32'sh3c74ebcf, 
               32'sh3c7467d9, 32'sh3c73e3d9, 32'sh3c735fd0, 32'sh3c72dbbe, 32'sh3c7257a2, 32'sh3c71d37d, 32'sh3c714f4e, 32'sh3c70cb17, 
               32'sh3c7046d6, 32'sh3c6fc28b, 32'sh3c6f3e37, 32'sh3c6eb9da, 32'sh3c6e3574, 32'sh3c6db104, 32'sh3c6d2c8b, 32'sh3c6ca809, 
               32'sh3c6c237e, 32'sh3c6b9ee9, 32'sh3c6b1a4a, 32'sh3c6a95a3, 32'sh3c6a10f2, 32'sh3c698c38, 32'sh3c690774, 32'sh3c6882a7, 
               32'sh3c67fdd1, 32'sh3c6778f2, 32'sh3c66f409, 32'sh3c666f17, 32'sh3c65ea1c, 32'sh3c656517, 32'sh3c64e009, 32'sh3c645af2, 
               32'sh3c63d5d1, 32'sh3c6350a7, 32'sh3c62cb74, 32'sh3c624637, 32'sh3c61c0f1, 32'sh3c613ba2, 32'sh3c60b649, 32'sh3c6030e8, 
               32'sh3c5fab7c, 32'sh3c5f2608, 32'sh3c5ea08a, 32'sh3c5e1b03, 32'sh3c5d9573, 32'sh3c5d0fd9, 32'sh3c5c8a36, 32'sh3c5c048a, 
               32'sh3c5b7ed4, 32'sh3c5af915, 32'sh3c5a734d, 32'sh3c59ed7b, 32'sh3c5967a1, 32'sh3c58e1bc, 32'sh3c585bcf, 32'sh3c57d5d8, 
               32'sh3c574fd8, 32'sh3c56c9cf, 32'sh3c5643bc, 32'sh3c55bda0, 32'sh3c55377b, 32'sh3c54b14c, 32'sh3c542b14, 32'sh3c53a4d3, 
               32'sh3c531e88, 32'sh3c529835, 32'sh3c5211d8, 32'sh3c518b71, 32'sh3c510501, 32'sh3c507e88, 32'sh3c4ff806, 32'sh3c4f717a, 
               32'sh3c4eeae5, 32'sh3c4e6447, 32'sh3c4ddda0, 32'sh3c4d56ef, 32'sh3c4cd035, 32'sh3c4c4971, 32'sh3c4bc2a5, 32'sh3c4b3bcf, 
               32'sh3c4ab4ef, 32'sh3c4a2e07, 32'sh3c49a715, 32'sh3c49201a, 32'sh3c489915, 32'sh3c481207, 32'sh3c478af0, 32'sh3c4703d0, 
               32'sh3c467ca6, 32'sh3c45f573, 32'sh3c456e37, 32'sh3c44e6f1, 32'sh3c445fa2, 32'sh3c43d84a, 32'sh3c4350e9, 32'sh3c42c97e, 
               32'sh3c42420a, 32'sh3c41ba8d, 32'sh3c413306, 32'sh3c40ab76, 32'sh3c4023dd, 32'sh3c3f9c3a, 32'sh3c3f148f, 32'sh3c3e8cd9, 
               32'sh3c3e051b, 32'sh3c3d7d53, 32'sh3c3cf582, 32'sh3c3c6da8, 32'sh3c3be5c5, 32'sh3c3b5dd8, 32'sh3c3ad5e2, 32'sh3c3a4de2, 
               32'sh3c39c5da, 32'sh3c393dc8, 32'sh3c38b5ac, 32'sh3c382d88, 32'sh3c37a55a, 32'sh3c371d23, 32'sh3c3694e2, 32'sh3c360c99, 
               32'sh3c358446, 32'sh3c34fbea, 32'sh3c347384, 32'sh3c33eb15, 32'sh3c33629d, 32'sh3c32da1c, 32'sh3c325191, 32'sh3c31c8fd, 
               32'sh3c314060, 32'sh3c30b7b9, 32'sh3c302f09, 32'sh3c2fa650, 32'sh3c2f1d8e, 32'sh3c2e94c2, 32'sh3c2e0bed, 32'sh3c2d830f, 
               32'sh3c2cfa28, 32'sh3c2c7137, 32'sh3c2be83d, 32'sh3c2b5f39, 32'sh3c2ad62d, 32'sh3c2a4d17, 32'sh3c29c3f8, 32'sh3c293acf, 
               32'sh3c28b19e, 32'sh3c282863, 32'sh3c279f1e, 32'sh3c2715d1, 32'sh3c268c7a, 32'sh3c26031a, 32'sh3c2579b0, 32'sh3c24f03e, 
               32'sh3c2466c2, 32'sh3c23dd3c, 32'sh3c2353ae, 32'sh3c22ca16, 32'sh3c224075, 32'sh3c21b6cb, 32'sh3c212d17, 32'sh3c20a35a, 
               32'sh3c201994, 32'sh3c1f8fc5, 32'sh3c1f05ec, 32'sh3c1e7c0a, 32'sh3c1df21f, 32'sh3c1d682b, 32'sh3c1cde2d, 32'sh3c1c5426, 
               32'sh3c1bca16, 32'sh3c1b3ffc, 32'sh3c1ab5d9, 32'sh3c1a2bad, 32'sh3c19a178, 32'sh3c191739, 32'sh3c188cf1, 32'sh3c1802a0, 
               32'sh3c177845, 32'sh3c16ede2, 32'sh3c166375, 32'sh3c15d8ff, 32'sh3c154e7f, 32'sh3c14c3f6, 32'sh3c143964, 32'sh3c13aec9, 
               32'sh3c132424, 32'sh3c129977, 32'sh3c120ebf, 32'sh3c1183ff, 32'sh3c10f935, 32'sh3c106e63, 32'sh3c0fe386, 32'sh3c0f58a1, 
               32'sh3c0ecdb2, 32'sh3c0e42ba, 32'sh3c0db7b9, 32'sh3c0d2caf, 32'sh3c0ca19b, 32'sh3c0c167e, 32'sh3c0b8b58, 32'sh3c0b0028, 
               32'sh3c0a74f0, 32'sh3c09e9ae, 32'sh3c095e62, 32'sh3c08d30e, 32'sh3c0847b0, 32'sh3c07bc49, 32'sh3c0730d9, 32'sh3c06a55f, 
               32'sh3c0619dc, 32'sh3c058e50, 32'sh3c0502bb, 32'sh3c04771c, 32'sh3c03eb74, 32'sh3c035fc3, 32'sh3c02d409, 32'sh3c024845, 
               32'sh3c01bc78, 32'sh3c0130a2, 32'sh3c00a4c3, 32'sh3c0018da, 32'sh3bff8ce8, 32'sh3bff00ed, 32'sh3bfe74e9, 32'sh3bfde8db, 
               32'sh3bfd5cc4, 32'sh3bfcd0a4, 32'sh3bfc447b, 32'sh3bfbb848, 32'sh3bfb2c0c, 32'sh3bfa9fc7, 32'sh3bfa1379, 32'sh3bf98721, 
               32'sh3bf8fac0, 32'sh3bf86e56, 32'sh3bf7e1e3, 32'sh3bf75566, 32'sh3bf6c8e0, 32'sh3bf63c51, 32'sh3bf5afb9, 32'sh3bf52317, 
               32'sh3bf4966c, 32'sh3bf409b8, 32'sh3bf37cfb, 32'sh3bf2f034, 32'sh3bf26364, 32'sh3bf1d68b, 32'sh3bf149a9, 32'sh3bf0bcbd, 
               32'sh3bf02fc9, 32'sh3befa2ca, 32'sh3bef15c3, 32'sh3bee88b3, 32'sh3bedfb99, 32'sh3bed6e76, 32'sh3bece149, 32'sh3bec5414, 
               32'sh3bebc6d5, 32'sh3beb398d, 32'sh3beaac3c, 32'sh3bea1ee1, 32'sh3be9917e, 32'sh3be90411, 32'sh3be8769b, 32'sh3be7e91b, 
               32'sh3be75b93, 32'sh3be6ce01, 32'sh3be64065, 32'sh3be5b2c1, 32'sh3be52513, 32'sh3be4975d, 32'sh3be4099c, 32'sh3be37bd3, 
               32'sh3be2ee01, 32'sh3be26025, 32'sh3be1d240, 32'sh3be14451, 32'sh3be0b65a, 32'sh3be02859, 32'sh3bdf9a4f, 32'sh3bdf0c3c, 
               32'sh3bde7e20, 32'sh3bddeffa, 32'sh3bdd61cb, 32'sh3bdcd393, 32'sh3bdc4552, 32'sh3bdbb707, 32'sh3bdb28b3, 32'sh3bda9a56, 
               32'sh3bda0bf0, 32'sh3bd97d80, 32'sh3bd8ef07, 32'sh3bd86085, 32'sh3bd7d1fa, 32'sh3bd74366, 32'sh3bd6b4c8, 32'sh3bd62621, 
               32'sh3bd59771, 32'sh3bd508b8, 32'sh3bd479f5, 32'sh3bd3eb29, 32'sh3bd35c54, 32'sh3bd2cd76, 32'sh3bd23e8f, 32'sh3bd1af9e, 
               32'sh3bd120a4, 32'sh3bd091a1, 32'sh3bd00295, 32'sh3bcf737f, 32'sh3bcee460, 32'sh3bce5538, 32'sh3bcdc607, 32'sh3bcd36cc, 
               32'sh3bcca789, 32'sh3bcc183c, 32'sh3bcb88e5, 32'sh3bcaf986, 32'sh3bca6a1d, 32'sh3bc9daac, 32'sh3bc94b31, 32'sh3bc8bbac, 
               32'sh3bc82c1f, 32'sh3bc79c88, 32'sh3bc70ce8, 32'sh3bc67d3f, 32'sh3bc5ed8d, 32'sh3bc55dd1, 32'sh3bc4ce0c, 32'sh3bc43e3e, 
               32'sh3bc3ae67, 32'sh3bc31e87, 32'sh3bc28e9d, 32'sh3bc1feaa, 32'sh3bc16eae, 32'sh3bc0dea9, 32'sh3bc04e9a, 32'sh3bbfbe83, 
               32'sh3bbf2e62, 32'sh3bbe9e37, 32'sh3bbe0e04, 32'sh3bbd7dc7, 32'sh3bbced82, 32'sh3bbc5d33, 32'sh3bbbccda, 32'sh3bbb3c79, 
               32'sh3bbaac0e, 32'sh3bba1b9a, 32'sh3bb98b1d, 32'sh3bb8fa97, 32'sh3bb86a08, 32'sh3bb7d96f, 32'sh3bb748cd, 32'sh3bb6b822, 
               32'sh3bb6276e, 32'sh3bb596b0, 32'sh3bb505e9, 32'sh3bb47519, 32'sh3bb3e440, 32'sh3bb3535e, 32'sh3bb2c272, 32'sh3bb2317e, 
               32'sh3bb1a080, 32'sh3bb10f78, 32'sh3bb07e68, 32'sh3bafed4e, 32'sh3baf5c2c, 32'sh3baecb00, 32'sh3bae39ca, 32'sh3bada88c, 
               32'sh3bad1744, 32'sh3bac85f3, 32'sh3babf499, 32'sh3bab6336, 32'sh3baad1ca, 32'sh3baa4054, 32'sh3ba9aed5, 32'sh3ba91d4d, 
               32'sh3ba88bbc, 32'sh3ba7fa22, 32'sh3ba7687e, 32'sh3ba6d6d1, 32'sh3ba6451b, 32'sh3ba5b35c, 32'sh3ba52194, 32'sh3ba48fc2, 
               32'sh3ba3fde7, 32'sh3ba36c03, 32'sh3ba2da16, 32'sh3ba2481f, 32'sh3ba1b620, 32'sh3ba12417, 32'sh3ba09205, 32'sh3b9fffea, 
               32'sh3b9f6dc5, 32'sh3b9edb98, 32'sh3b9e4961, 32'sh3b9db721, 32'sh3b9d24d8, 32'sh3b9c9286, 32'sh3b9c002a, 32'sh3b9b6dc5, 
               32'sh3b9adb57, 32'sh3b9a48e0, 32'sh3b99b660, 32'sh3b9923d6, 32'sh3b989144, 32'sh3b97fea8, 32'sh3b976c03, 32'sh3b96d954, 
               32'sh3b96469d, 32'sh3b95b3dc, 32'sh3b952112, 32'sh3b948e3f, 32'sh3b93fb63, 32'sh3b93687e, 32'sh3b92d58f, 32'sh3b924297, 
               32'sh3b91af97, 32'sh3b911c8c, 32'sh3b908979, 32'sh3b8ff65c, 32'sh3b8f6337, 32'sh3b8ed008, 32'sh3b8e3cd0, 32'sh3b8da98f, 
               32'sh3b8d1644, 32'sh3b8c82f0, 32'sh3b8bef94, 32'sh3b8b5c2e, 32'sh3b8ac8bf, 32'sh3b8a3546, 32'sh3b89a1c5, 32'sh3b890e3a, 
               32'sh3b887aa6, 32'sh3b87e709, 32'sh3b875363, 32'sh3b86bfb3, 32'sh3b862bfb, 32'sh3b859839, 32'sh3b85046e, 32'sh3b84709a, 
               32'sh3b83dcbc, 32'sh3b8348d6, 32'sh3b82b4e6, 32'sh3b8220ed, 32'sh3b818ceb, 32'sh3b80f8e0, 32'sh3b8064cc, 32'sh3b7fd0ae, 
               32'sh3b7f3c87, 32'sh3b7ea857, 32'sh3b7e141e, 32'sh3b7d7fdc, 32'sh3b7ceb90, 32'sh3b7c573c, 32'sh3b7bc2de, 32'sh3b7b2e77, 
               32'sh3b7a9a07, 32'sh3b7a058e, 32'sh3b79710b, 32'sh3b78dc7f, 32'sh3b7847eb, 32'sh3b77b34d, 32'sh3b771ea5, 32'sh3b7689f5, 
               32'sh3b75f53c, 32'sh3b756079, 32'sh3b74cbad, 32'sh3b7436d8, 32'sh3b73a1fa, 32'sh3b730d12, 32'sh3b727822, 32'sh3b71e328, 
               32'sh3b714e25, 32'sh3b70b919, 32'sh3b702404, 32'sh3b6f8ee6, 32'sh3b6ef9be, 32'sh3b6e648e, 32'sh3b6dcf54, 32'sh3b6d3a11, 
               32'sh3b6ca4c4, 32'sh3b6c0f6f, 32'sh3b6b7a11, 32'sh3b6ae4a9, 32'sh3b6a4f38, 32'sh3b69b9be, 32'sh3b69243b, 32'sh3b688eaf, 
               32'sh3b67f919, 32'sh3b67637a, 32'sh3b66cdd3, 32'sh3b663822, 32'sh3b65a268, 32'sh3b650ca4, 32'sh3b6476d8, 32'sh3b63e102, 
               32'sh3b634b23, 32'sh3b62b53b, 32'sh3b621f4a, 32'sh3b618950, 32'sh3b60f34d, 32'sh3b605d40, 32'sh3b5fc72a, 32'sh3b5f310c, 
               32'sh3b5e9ae4, 32'sh3b5e04b2, 32'sh3b5d6e78, 32'sh3b5cd835, 32'sh3b5c41e8, 32'sh3b5bab92, 32'sh3b5b1533, 32'sh3b5a7ecb, 
               32'sh3b59e85a, 32'sh3b5951df, 32'sh3b58bb5c, 32'sh3b5824cf, 32'sh3b578e39, 32'sh3b56f79a, 32'sh3b5660f2, 32'sh3b55ca41, 
               32'sh3b553386, 32'sh3b549cc3, 32'sh3b5405f6, 32'sh3b536f20, 32'sh3b52d841, 32'sh3b524159, 32'sh3b51aa67, 32'sh3b51136d, 
               32'sh3b507c69, 32'sh3b4fe55c, 32'sh3b4f4e46, 32'sh3b4eb727, 32'sh3b4e1fff, 32'sh3b4d88ce, 32'sh3b4cf193, 32'sh3b4c5a4f, 
               32'sh3b4bc303, 32'sh3b4b2bad, 32'sh3b4a944d, 32'sh3b49fce5, 32'sh3b496574, 32'sh3b48cdf9, 32'sh3b483676, 32'sh3b479ee9, 
               32'sh3b470753, 32'sh3b466fb4, 32'sh3b45d80b, 32'sh3b45405a, 32'sh3b44a8a0, 32'sh3b4410dc, 32'sh3b43790f, 32'sh3b42e139, 
               32'sh3b42495a, 32'sh3b41b172, 32'sh3b411980, 32'sh3b408186, 32'sh3b3fe982, 32'sh3b3f5175, 32'sh3b3eb960, 32'sh3b3e2140, 
               32'sh3b3d8918, 32'sh3b3cf0e7, 32'sh3b3c58ad, 32'sh3b3bc069, 32'sh3b3b281c, 32'sh3b3a8fc6, 32'sh3b39f767, 32'sh3b395eff, 
               32'sh3b38c68e, 32'sh3b382e14, 32'sh3b379590, 32'sh3b36fd03, 32'sh3b36646e, 32'sh3b35cbcf, 32'sh3b353327, 32'sh3b349a75, 
               32'sh3b3401bb, 32'sh3b3368f8, 32'sh3b32d02b, 32'sh3b323755, 32'sh3b319e77, 32'sh3b31058f, 32'sh3b306c9d, 32'sh3b2fd3a3, 
               32'sh3b2f3aa0, 32'sh3b2ea193, 32'sh3b2e087e, 32'sh3b2d6f5f, 32'sh3b2cd637, 32'sh3b2c3d06, 32'sh3b2ba3cc, 32'sh3b2b0a89, 
               32'sh3b2a713d, 32'sh3b29d7e7, 32'sh3b293e89, 32'sh3b28a521, 32'sh3b280bb0, 32'sh3b277236, 32'sh3b26d8b3, 32'sh3b263f27, 
               32'sh3b25a591, 32'sh3b250bf3, 32'sh3b24724b, 32'sh3b23d89b, 32'sh3b233ee1, 32'sh3b22a51e, 32'sh3b220b52, 32'sh3b21717d, 
               32'sh3b20d79e, 32'sh3b203db7, 32'sh3b1fa3c6, 32'sh3b1f09cd, 32'sh3b1e6fca, 32'sh3b1dd5be, 32'sh3b1d3ba9, 32'sh3b1ca18b, 
               32'sh3b1c0764, 32'sh3b1b6d33, 32'sh3b1ad2fa, 32'sh3b1a38b7, 32'sh3b199e6c, 32'sh3b190417, 32'sh3b1869b9, 32'sh3b17cf52, 
               32'sh3b1734e2, 32'sh3b169a69, 32'sh3b15ffe6, 32'sh3b15655b, 32'sh3b14cac6, 32'sh3b143028, 32'sh3b139582, 32'sh3b12fad2, 
               32'sh3b126019, 32'sh3b11c557, 32'sh3b112a8b, 32'sh3b108fb7, 32'sh3b0ff4d9, 32'sh3b0f59f3, 32'sh3b0ebf03, 32'sh3b0e240a, 
               32'sh3b0d8909, 32'sh3b0cedfe, 32'sh3b0c52e9, 32'sh3b0bb7cc, 32'sh3b0b1ca6, 32'sh3b0a8176, 32'sh3b09e63e, 32'sh3b094afc, 
               32'sh3b08afb2, 32'sh3b08145e, 32'sh3b077901, 32'sh3b06dd9b, 32'sh3b06422c, 32'sh3b05a6b3, 32'sh3b050b32, 32'sh3b046fa7, 
               32'sh3b03d414, 32'sh3b033877, 32'sh3b029cd1, 32'sh3b020123, 32'sh3b01656b, 32'sh3b00c9aa, 32'sh3b002ddf, 32'sh3aff920c, 
               32'sh3afef630, 32'sh3afe5a4a, 32'sh3afdbe5c, 32'sh3afd2264, 32'sh3afc8663, 32'sh3afbea5a, 32'sh3afb4e47, 32'sh3afab22b, 
               32'sh3afa1605, 32'sh3af979d7, 32'sh3af8dda0, 32'sh3af8415f, 32'sh3af7a516, 32'sh3af708c3, 32'sh3af66c68, 32'sh3af5d003, 
               32'sh3af53395, 32'sh3af4971e, 32'sh3af3fa9e, 32'sh3af35e15, 32'sh3af2c183, 32'sh3af224e7, 32'sh3af18843, 32'sh3af0eb95, 
               32'sh3af04edf, 32'sh3aefb21f, 32'sh3aef1556, 32'sh3aee7884, 32'sh3aeddba9, 32'sh3aed3ec5, 32'sh3aeca1d8, 32'sh3aec04e2, 
               32'sh3aeb67e3, 32'sh3aeacada, 32'sh3aea2dc9, 32'sh3ae990ae, 32'sh3ae8f38b, 32'sh3ae8565e, 32'sh3ae7b928, 32'sh3ae71be9, 
               32'sh3ae67ea1, 32'sh3ae5e150, 32'sh3ae543f6, 32'sh3ae4a693, 32'sh3ae40926, 32'sh3ae36bb1, 32'sh3ae2ce32, 32'sh3ae230ab, 
               32'sh3ae1931a, 32'sh3ae0f581, 32'sh3ae057de, 32'sh3adfba32, 32'sh3adf1c7d, 32'sh3ade7ebf, 32'sh3adde0f8, 32'sh3add4327, 
               32'sh3adca54e, 32'sh3adc076c, 32'sh3adb6980, 32'sh3adacb8c, 32'sh3ada2d8e, 32'sh3ad98f88, 32'sh3ad8f178, 32'sh3ad8535f, 
               32'sh3ad7b53d, 32'sh3ad71712, 32'sh3ad678de, 32'sh3ad5daa1, 32'sh3ad53c5b, 32'sh3ad49e0c, 32'sh3ad3ffb3, 32'sh3ad36152, 
               32'sh3ad2c2e8, 32'sh3ad22474, 32'sh3ad185f7, 32'sh3ad0e772, 32'sh3ad048e3, 32'sh3acfaa4b, 32'sh3acf0baa, 32'sh3ace6d00, 
               32'sh3acdce4d, 32'sh3acd2f91, 32'sh3acc90cc, 32'sh3acbf1fe, 32'sh3acb5327, 32'sh3acab446, 32'sh3aca155d, 32'sh3ac9766a, 
               32'sh3ac8d76f, 32'sh3ac8386a, 32'sh3ac7995c, 32'sh3ac6fa46, 32'sh3ac65b26, 32'sh3ac5bbfd, 32'sh3ac51ccb, 32'sh3ac47d90, 
               32'sh3ac3de4c, 32'sh3ac33eff, 32'sh3ac29fa9, 32'sh3ac20049, 32'sh3ac160e1, 32'sh3ac0c170, 32'sh3ac021f5, 32'sh3abf8272, 
               32'sh3abee2e5, 32'sh3abe434f, 32'sh3abda3b1, 32'sh3abd0409, 32'sh3abc6458, 32'sh3abbc49e, 32'sh3abb24db, 32'sh3aba850f, 
               32'sh3ab9e53a, 32'sh3ab9455c, 32'sh3ab8a575, 32'sh3ab80585, 32'sh3ab7658c, 32'sh3ab6c58a, 32'sh3ab6257e, 32'sh3ab5856a, 
               32'sh3ab4e54c, 32'sh3ab44526, 32'sh3ab3a4f6, 32'sh3ab304be, 32'sh3ab2647c, 32'sh3ab1c431, 32'sh3ab123dd, 32'sh3ab08381, 
               32'sh3aafe31b, 32'sh3aaf42ac, 32'sh3aaea234, 32'sh3aae01b3, 32'sh3aad6129, 32'sh3aacc095, 32'sh3aac1ff9, 32'sh3aab7f54, 
               32'sh3aaadea6, 32'sh3aaa3def, 32'sh3aa99d2e, 32'sh3aa8fc65, 32'sh3aa85b92, 32'sh3aa7bab7, 32'sh3aa719d2, 32'sh3aa678e5, 
               32'sh3aa5d7ee, 32'sh3aa536ee, 32'sh3aa495e6, 32'sh3aa3f4d4, 32'sh3aa353b9, 32'sh3aa2b295, 32'sh3aa21168, 32'sh3aa17032, 
               32'sh3aa0cef3, 32'sh3aa02dab, 32'sh3a9f8c5a, 32'sh3a9eeb00, 32'sh3a9e499d, 32'sh3a9da831, 32'sh3a9d06bc, 32'sh3a9c653d, 
               32'sh3a9bc3b6, 32'sh3a9b2226, 32'sh3a9a808c, 32'sh3a99deea, 32'sh3a993d3e, 32'sh3a989b8a, 32'sh3a97f9cc, 32'sh3a975806, 
               32'sh3a96b636, 32'sh3a96145e, 32'sh3a95727c, 32'sh3a94d091, 32'sh3a942e9d, 32'sh3a938ca1, 32'sh3a92ea9b, 32'sh3a92488c, 
               32'sh3a91a674, 32'sh3a910453, 32'sh3a906229, 32'sh3a8fbff6, 32'sh3a8f1dba, 32'sh3a8e7b75, 32'sh3a8dd927, 32'sh3a8d36d0, 
               32'sh3a8c9470, 32'sh3a8bf207, 32'sh3a8b4f95, 32'sh3a8aad1a, 32'sh3a8a0a95, 32'sh3a896808, 32'sh3a88c572, 32'sh3a8822d3, 
               32'sh3a87802a, 32'sh3a86dd79, 32'sh3a863abe, 32'sh3a8597fb, 32'sh3a84f52f, 32'sh3a845259, 32'sh3a83af7b, 32'sh3a830c93, 
               32'sh3a8269a3, 32'sh3a81c6a9, 32'sh3a8123a6, 32'sh3a80809b, 32'sh3a7fdd86, 32'sh3a7f3a69, 32'sh3a7e9742, 32'sh3a7df412, 
               32'sh3a7d50da, 32'sh3a7cad98, 32'sh3a7c0a4d, 32'sh3a7b66f9, 32'sh3a7ac39d, 32'sh3a7a2037, 32'sh3a797cc8, 32'sh3a78d950, 
               32'sh3a7835cf, 32'sh3a779245, 32'sh3a76eeb2, 32'sh3a764b17, 32'sh3a75a772, 32'sh3a7503c4, 32'sh3a74600d, 32'sh3a73bc4d, 
               32'sh3a731884, 32'sh3a7274b2, 32'sh3a71d0d7, 32'sh3a712cf3, 32'sh3a708906, 32'sh3a6fe510, 32'sh3a6f4111, 32'sh3a6e9d09, 
               32'sh3a6df8f8, 32'sh3a6d54de, 32'sh3a6cb0ba, 32'sh3a6c0c8e, 32'sh3a6b6859, 32'sh3a6ac41b, 32'sh3a6a1fd4, 32'sh3a697b84, 
               32'sh3a68d72b, 32'sh3a6832c8, 32'sh3a678e5d, 32'sh3a66e9e9, 32'sh3a66456c, 32'sh3a65a0e6, 32'sh3a64fc57, 32'sh3a6457be, 
               32'sh3a63b31d, 32'sh3a630e73, 32'sh3a6269c0, 32'sh3a61c504, 32'sh3a61203e, 32'sh3a607b70, 32'sh3a5fd699, 32'sh3a5f31b9, 
               32'sh3a5e8cd0, 32'sh3a5de7dd, 32'sh3a5d42e2, 32'sh3a5c9dde, 32'sh3a5bf8d1, 32'sh3a5b53ba, 32'sh3a5aae9b, 32'sh3a5a0973, 
               32'sh3a596442, 32'sh3a58bf08, 32'sh3a5819c4, 32'sh3a577478, 32'sh3a56cf23, 32'sh3a5629c5, 32'sh3a55845d, 32'sh3a54deed, 
               32'sh3a543974, 32'sh3a5393f2, 32'sh3a52ee67, 32'sh3a5248d3, 32'sh3a51a335, 32'sh3a50fd8f, 32'sh3a5057e0, 32'sh3a4fb228, 
               32'sh3a4f0c67, 32'sh3a4e669d, 32'sh3a4dc0c9, 32'sh3a4d1aed, 32'sh3a4c7508, 32'sh3a4bcf1a, 32'sh3a4b2923, 32'sh3a4a8323, 
               32'sh3a49dd1a, 32'sh3a493708, 32'sh3a4890ed, 32'sh3a47eac9, 32'sh3a47449c, 32'sh3a469e66, 32'sh3a45f827, 32'sh3a4551df, 
               32'sh3a44ab8e, 32'sh3a440534, 32'sh3a435ed1, 32'sh3a42b865, 32'sh3a4211f0, 32'sh3a416b72, 32'sh3a40c4eb, 32'sh3a401e5b, 
               32'sh3a3f77c3, 32'sh3a3ed121, 32'sh3a3e2a76, 32'sh3a3d83c2, 32'sh3a3cdd05, 32'sh3a3c3640, 32'sh3a3b8f71, 32'sh3a3ae899, 
               32'sh3a3a41b9, 32'sh3a399acf, 32'sh3a38f3dc, 32'sh3a384ce1, 32'sh3a37a5dc, 32'sh3a36fece, 32'sh3a3657b8, 32'sh3a35b098, 
               32'sh3a350970, 32'sh3a34623e, 32'sh3a33bb04, 32'sh3a3313c0, 32'sh3a326c74, 32'sh3a31c51f, 32'sh3a311dc0, 32'sh3a307659, 
               32'sh3a2fcee8, 32'sh3a2f276f, 32'sh3a2e7fed, 32'sh3a2dd862, 32'sh3a2d30cd, 32'sh3a2c8930, 32'sh3a2be18a, 32'sh3a2b39db, 
               32'sh3a2a9223, 32'sh3a29ea62, 32'sh3a294298, 32'sh3a289ac5, 32'sh3a27f2e9, 32'sh3a274b04, 32'sh3a26a316, 32'sh3a25fb1f, 
               32'sh3a25531f, 32'sh3a24ab17, 32'sh3a240305, 32'sh3a235aea, 32'sh3a22b2c6, 32'sh3a220a9a, 32'sh3a216264, 32'sh3a20ba25, 
               32'sh3a2011de, 32'sh3a1f698d, 32'sh3a1ec134, 32'sh3a1e18d1, 32'sh3a1d7066, 32'sh3a1cc7f2, 32'sh3a1c1f74, 32'sh3a1b76ee, 
               32'sh3a1ace5f, 32'sh3a1a25c6, 32'sh3a197d25, 32'sh3a18d47b, 32'sh3a182bc8, 32'sh3a17830c, 32'sh3a16da47, 32'sh3a163179, 
               32'sh3a1588a2, 32'sh3a14dfc2, 32'sh3a1436d9, 32'sh3a138de8, 32'sh3a12e4ed, 32'sh3a123be9, 32'sh3a1192dc, 32'sh3a10e9c7, 
               32'sh3a1040a8, 32'sh3a0f9781, 32'sh3a0eee50, 32'sh3a0e4517, 32'sh3a0d9bd4, 32'sh3a0cf289, 32'sh3a0c4935, 32'sh3a0b9fd7, 
               32'sh3a0af671, 32'sh3a0a4d02, 32'sh3a09a38a, 32'sh3a08fa09, 32'sh3a08507f, 32'sh3a07a6ec, 32'sh3a06fd50, 32'sh3a0653ab, 
               32'sh3a05a9fd, 32'sh3a050047, 32'sh3a045687, 32'sh3a03acbe, 32'sh3a0302ed, 32'sh3a025912, 32'sh3a01af2f, 32'sh3a010542, 
               32'sh3a005b4d, 32'sh39ffb14f, 32'sh39ff0747, 32'sh39fe5d37, 32'sh39fdb31e, 32'sh39fd08fc, 32'sh39fc5ed1, 32'sh39fbb49d, 
               32'sh39fb0a60, 32'sh39fa601a, 32'sh39f9b5cb, 32'sh39f90b74, 32'sh39f86113, 32'sh39f7b6a9, 32'sh39f70c37, 32'sh39f661bb, 
               32'sh39f5b737, 32'sh39f50ca9, 32'sh39f46213, 32'sh39f3b774, 32'sh39f30ccc, 32'sh39f2621b, 32'sh39f1b761, 32'sh39f10c9e, 
               32'sh39f061d2, 32'sh39efb6fd, 32'sh39ef0c1f, 32'sh39ee6138, 32'sh39edb649, 32'sh39ed0b50, 32'sh39ec604e, 32'sh39ebb544, 
               32'sh39eb0a31, 32'sh39ea5f14, 32'sh39e9b3ef, 32'sh39e908c1, 32'sh39e85d8a, 32'sh39e7b24a, 32'sh39e70701, 32'sh39e65baf, 
               32'sh39e5b054, 32'sh39e504f0, 32'sh39e45983, 32'sh39e3ae0e, 32'sh39e3028f, 32'sh39e25708, 32'sh39e1ab77, 32'sh39e0ffde, 
               32'sh39e0543c, 32'sh39dfa891, 32'sh39defcdd, 32'sh39de511f, 32'sh39dda55a, 32'sh39dcf98b, 32'sh39dc4db3, 32'sh39dba1d2, 
               32'sh39daf5e8, 32'sh39da49f6, 32'sh39d99dfa, 32'sh39d8f1f6, 32'sh39d845e9, 32'sh39d799d2, 32'sh39d6edb3, 32'sh39d6418b, 
               32'sh39d5955a, 32'sh39d4e920, 32'sh39d43cdd, 32'sh39d39092, 32'sh39d2e43d, 32'sh39d237df, 32'sh39d18b79, 32'sh39d0df09, 
               32'sh39d03291, 32'sh39cf8610, 32'sh39ced986, 32'sh39ce2cf2, 32'sh39cd8056, 32'sh39ccd3b2, 32'sh39cc2704, 32'sh39cb7a4d, 
               32'sh39cacd8d, 32'sh39ca20c5, 32'sh39c973f3, 32'sh39c8c719, 32'sh39c81a36, 32'sh39c76d49, 32'sh39c6c054, 32'sh39c61356, 
               32'sh39c5664f, 32'sh39c4b93f, 32'sh39c40c27, 32'sh39c35f05, 32'sh39c2b1da, 32'sh39c204a7, 32'sh39c1576a, 32'sh39c0aa25, 
               32'sh39bffcd7, 32'sh39bf4f80, 32'sh39bea220, 32'sh39bdf4b7, 32'sh39bd4745, 32'sh39bc99ca, 32'sh39bbec47, 32'sh39bb3eba, 
               32'sh39ba9125, 32'sh39b9e386, 32'sh39b935df, 32'sh39b8882f, 32'sh39b7da76, 32'sh39b72cb4, 32'sh39b67ee9, 32'sh39b5d115, 
               32'sh39b52339, 32'sh39b47553, 32'sh39b3c765, 32'sh39b3196d, 32'sh39b26b6d, 32'sh39b1bd64, 32'sh39b10f52, 32'sh39b06137, 
               32'sh39afb313, 32'sh39af04e6, 32'sh39ae56b1, 32'sh39ada872, 32'sh39acfa2b, 32'sh39ac4bda, 32'sh39ab9d81, 32'sh39aaef1f, 
               32'sh39aa40b4, 32'sh39a99240, 32'sh39a8e3c4, 32'sh39a8353e, 32'sh39a786af, 32'sh39a6d818, 32'sh39a62978, 32'sh39a57ace, 
               32'sh39a4cc1c, 32'sh39a41d61, 32'sh39a36e9d, 32'sh39a2bfd0, 32'sh39a210fb, 32'sh39a1621c, 32'sh39a0b335, 32'sh39a00444, 
               32'sh399f554b, 32'sh399ea649, 32'sh399df73e, 32'sh399d482a, 32'sh399c990d, 32'sh399be9e8, 32'sh399b3ab9, 32'sh399a8b82, 
               32'sh3999dc42, 32'sh39992cf8, 32'sh39987da6, 32'sh3997ce4b, 32'sh39971ee7, 32'sh39966f7b, 32'sh3995c005, 32'sh39951087, 
               32'sh399460ff, 32'sh3993b16f, 32'sh399301d6, 32'sh39925234, 32'sh3991a289, 32'sh3990f2d5, 32'sh39904319, 32'sh398f9353, 
               32'sh398ee385, 32'sh398e33ae, 32'sh398d83ce, 32'sh398cd3e5, 32'sh398c23f3, 32'sh398b73f8, 32'sh398ac3f4, 32'sh398a13e8, 
               32'sh398963d2, 32'sh3988b3b4, 32'sh3988038d, 32'sh3987535d, 32'sh3986a324, 32'sh3985f2e2, 32'sh39854298, 32'sh39849244, 
               32'sh3983e1e8, 32'sh39833183, 32'sh39828115, 32'sh3981d09e, 32'sh3981201e, 32'sh39806f95, 32'sh397fbf04, 32'sh397f0e69, 
               32'sh397e5dc6, 32'sh397dad1a, 32'sh397cfc65, 32'sh397c4ba7, 32'sh397b9ae0, 32'sh397aea10, 32'sh397a3938, 32'sh39798857, 
               32'sh3978d76c, 32'sh39782679, 32'sh3977757d, 32'sh3976c479, 32'sh3976136b, 32'sh39756254, 32'sh3974b135, 32'sh3974000d, 
               32'sh39734edc, 32'sh39729da2, 32'sh3971ec5f, 32'sh39713b13, 32'sh397089bf, 32'sh396fd861, 32'sh396f26fb, 32'sh396e758c, 
               32'sh396dc414, 32'sh396d1293, 32'sh396c610a, 32'sh396baf77, 32'sh396afddc, 32'sh396a4c37, 32'sh39699a8a, 32'sh3968e8d4, 
               32'sh39683715, 32'sh3967854e, 32'sh3966d37d, 32'sh396621a4, 32'sh39656fc2, 32'sh3964bdd7, 32'sh39640be3, 32'sh396359e6, 
               32'sh3962a7e0, 32'sh3961f5d2, 32'sh396143bb, 32'sh3960919a, 32'sh395fdf71, 32'sh395f2d40, 32'sh395e7b05, 32'sh395dc8c1, 
               32'sh395d1675, 32'sh395c6420, 32'sh395bb1c2, 32'sh395aff5b, 32'sh395a4ceb, 32'sh39599a72, 32'sh3958e7f1, 32'sh39583566, 
               32'sh395782d3, 32'sh3956d037, 32'sh39561d92, 32'sh39556ae5, 32'sh3954b82e, 32'sh3954056f, 32'sh395352a7, 32'sh39529fd6, 
               32'sh3951ecfc, 32'sh39513a19, 32'sh3950872d, 32'sh394fd439, 32'sh394f213c, 32'sh394e6e36, 32'sh394dbb27, 32'sh394d080f, 
               32'sh394c54ee, 32'sh394ba1c5, 32'sh394aee93, 32'sh394a3b58, 32'sh39498814, 32'sh3948d4c7, 32'sh39482171, 32'sh39476e13, 
               32'sh3946baac, 32'sh3946073b, 32'sh394553c3, 32'sh3944a041, 32'sh3943ecb6, 32'sh39433923, 32'sh39428586, 32'sh3941d1e1, 
               32'sh39411e33, 32'sh39406a7d, 32'sh393fb6bd, 32'sh393f02f5, 32'sh393e4f23, 32'sh393d9b49, 32'sh393ce767, 32'sh393c337b, 
               32'sh393b7f86, 32'sh393acb89, 32'sh393a1783, 32'sh39396374, 32'sh3938af5c, 32'sh3937fb3b, 32'sh39374712, 32'sh393692df, 
               32'sh3935dea4, 32'sh39352a60, 32'sh39347613, 32'sh3933c1be, 32'sh39330d5f, 32'sh393258f8, 32'sh3931a488, 32'sh3930f00f, 
               32'sh39303b8e, 32'sh392f8703, 32'sh392ed270, 32'sh392e1dd3, 32'sh392d692f, 32'sh392cb481, 32'sh392bffca, 32'sh392b4b0b, 
               32'sh392a9642, 32'sh3929e171, 32'sh39292c97, 32'sh392877b5, 32'sh3927c2c9, 32'sh39270dd5, 32'sh392658d8, 32'sh3925a3d2, 
               32'sh3924eec3, 32'sh392439ac, 32'sh3923848b, 32'sh3922cf62, 32'sh39221a30, 32'sh392164f5, 32'sh3920afb1, 32'sh391ffa65, 
               32'sh391f4510, 32'sh391e8fb2, 32'sh391dda4b, 32'sh391d24db, 32'sh391c6f63, 32'sh391bb9e1, 32'sh391b0457, 32'sh391a4ec4, 
               32'sh39199929, 32'sh3918e384, 32'sh39182dd7, 32'sh39177821, 32'sh3916c262, 32'sh39160c9a, 32'sh391556ca, 32'sh3914a0f0, 
               32'sh3913eb0e, 32'sh39133523, 32'sh39127f2f, 32'sh3911c933, 32'sh3911132d, 32'sh39105d1f, 32'sh390fa708, 32'sh390ef0e9, 
               32'sh390e3ac0, 32'sh390d848f, 32'sh390cce55, 32'sh390c1812, 32'sh390b61c6, 32'sh390aab71, 32'sh3909f514, 32'sh39093eae, 
               32'sh3908883f, 32'sh3907d1c7, 32'sh39071b47, 32'sh390664bd, 32'sh3905ae2b, 32'sh3904f790, 32'sh390440ed, 32'sh39038a40, 
               32'sh3902d38b, 32'sh39021ccd, 32'sh39016606, 32'sh3900af36, 32'sh38fff85e, 32'sh38ff417d, 32'sh38fe8a93, 32'sh38fdd3a0, 
               32'sh38fd1ca4, 32'sh38fc65a0, 32'sh38fbae93, 32'sh38faf77d, 32'sh38fa405e, 32'sh38f98936, 32'sh38f8d206, 32'sh38f81acd, 
               32'sh38f7638b, 32'sh38f6ac40, 32'sh38f5f4ed, 32'sh38f53d91, 32'sh38f4862c, 32'sh38f3cebe, 32'sh38f31747, 32'sh38f25fc8, 
               32'sh38f1a840, 32'sh38f0f0af, 32'sh38f03915, 32'sh38ef8173, 32'sh38eec9c7, 32'sh38ee1213, 32'sh38ed5a56, 32'sh38eca291, 
               32'sh38ebeac2, 32'sh38eb32eb, 32'sh38ea7b0b, 32'sh38e9c323, 32'sh38e90b31, 32'sh38e85337, 32'sh38e79b34, 32'sh38e6e328, 
               32'sh38e62b13, 32'sh38e572f6, 32'sh38e4bad0, 32'sh38e402a1, 32'sh38e34a69, 32'sh38e29229, 32'sh38e1d9df, 32'sh38e1218d, 
               32'sh38e06932, 32'sh38dfb0cf, 32'sh38def863, 32'sh38de3fed, 32'sh38dd8770, 32'sh38dccee9, 32'sh38dc165a, 32'sh38db5dc1, 
               32'sh38daa520, 32'sh38d9ec77, 32'sh38d933c4, 32'sh38d87b09, 32'sh38d7c245, 32'sh38d70978, 32'sh38d650a3, 32'sh38d597c4, 
               32'sh38d4dedd, 32'sh38d425ed, 32'sh38d36cf5, 32'sh38d2b3f3, 32'sh38d1fae9, 32'sh38d141d6, 32'sh38d088bb, 32'sh38cfcf96, 
               32'sh38cf1669, 32'sh38ce5d33, 32'sh38cda3f4, 32'sh38cceaad, 32'sh38cc315d, 32'sh38cb7804, 32'sh38cabea2, 32'sh38ca0538, 
               32'sh38c94bc4, 32'sh38c89248, 32'sh38c7d8c3, 32'sh38c71f36, 32'sh38c665a0, 32'sh38c5ac01, 32'sh38c4f259, 32'sh38c438a8, 
               32'sh38c37eef, 32'sh38c2c52d, 32'sh38c20b62, 32'sh38c1518f, 32'sh38c097b2, 32'sh38bfddcd, 32'sh38bf23df, 32'sh38be69e9, 
               32'sh38bdafea, 32'sh38bcf5e1, 32'sh38bc3bd1, 32'sh38bb81b7, 32'sh38bac795, 32'sh38ba0d6a, 32'sh38b95336, 32'sh38b898f9, 
               32'sh38b7deb4, 32'sh38b72466, 32'sh38b66a0f, 32'sh38b5afb0, 32'sh38b4f547, 32'sh38b43ad6, 32'sh38b3805c, 32'sh38b2c5da, 
               32'sh38b20b4f, 32'sh38b150bb, 32'sh38b0961e, 32'sh38afdb78, 32'sh38af20ca, 32'sh38ae6613, 32'sh38adab54, 32'sh38acf08b, 
               32'sh38ac35ba, 32'sh38ab7ae0, 32'sh38aabffd, 32'sh38aa0512, 32'sh38a94a1e, 32'sh38a88f21, 32'sh38a7d41b, 32'sh38a7190d, 
               32'sh38a65df6, 32'sh38a5a2d6, 32'sh38a4e7ad, 32'sh38a42c7c, 32'sh38a37142, 32'sh38a2b5ff, 32'sh38a1fab4, 32'sh38a13f5f, 
               32'sh38a08402, 32'sh389fc89d, 32'sh389f0d2e, 32'sh389e51b7, 32'sh389d9637, 32'sh389cdaae, 32'sh389c1f1d, 32'sh389b6383, 
               32'sh389aa7e0, 32'sh3899ec35, 32'sh38993080, 32'sh389874c3, 32'sh3897b8fe, 32'sh3896fd2f, 32'sh38964158, 32'sh38958578, 
               32'sh3894c98f, 32'sh38940d9e, 32'sh389351a4, 32'sh389295a1, 32'sh3891d995, 32'sh38911d81, 32'sh38906164, 32'sh388fa53e, 
               32'sh388ee910, 32'sh388e2cd9, 32'sh388d7099, 32'sh388cb450, 32'sh388bf7ff, 32'sh388b3ba5, 32'sh388a7f42, 32'sh3889c2d7, 
               32'sh38890663, 32'sh388849e6, 32'sh38878d60, 32'sh3886d0d2, 32'sh3886143b, 32'sh3885579b, 32'sh38849af2, 32'sh3883de41, 
               32'sh38832187, 32'sh388264c4, 32'sh3881a7f9, 32'sh3880eb25, 32'sh38802e48, 32'sh387f7163, 32'sh387eb474, 32'sh387df77d, 
               32'sh387d3a7e, 32'sh387c7d75, 32'sh387bc064, 32'sh387b034b, 32'sh387a4628, 32'sh387988fd, 32'sh3878cbc9, 32'sh38780e8c, 
               32'sh38775147, 32'sh387693f9, 32'sh3875d6a2, 32'sh38751943, 32'sh38745bdb, 32'sh38739e6a, 32'sh3872e0f0, 32'sh3872236e, 
               32'sh387165e3, 32'sh3870a84f, 32'sh386feab3, 32'sh386f2d0e, 32'sh386e6f60, 32'sh386db1aa, 32'sh386cf3ea, 32'sh386c3622, 
               32'sh386b7852, 32'sh386aba79, 32'sh3869fc97, 32'sh38693eac, 32'sh386880b8, 32'sh3867c2bc, 32'sh386704b8, 32'sh386646aa, 
               32'sh38658894, 32'sh3864ca75, 32'sh38640c4d, 32'sh38634e1d, 32'sh38628fe4, 32'sh3861d1a3, 32'sh38611358, 32'sh38605505, 
               32'sh385f96a9, 32'sh385ed845, 32'sh385e19d8, 32'sh385d5b62, 32'sh385c9ce3, 32'sh385bde5c, 32'sh385b1fcc, 32'sh385a6134, 
               32'sh3859a292, 32'sh3858e3e8, 32'sh38582536, 32'sh3857667a, 32'sh3856a7b6, 32'sh3855e8ea, 32'sh38552a14, 32'sh38546b36, 
               32'sh3853ac4f, 32'sh3852ed60, 32'sh38522e68, 32'sh38516f67, 32'sh3850b05d, 32'sh384ff14b, 32'sh384f3230, 32'sh384e730d, 
               32'sh384db3e0, 32'sh384cf4ab, 32'sh384c356e, 32'sh384b7627, 32'sh384ab6d8, 32'sh3849f781, 32'sh38493820, 32'sh384878b7, 
               32'sh3847b946, 32'sh3846f9cb, 32'sh38463a48, 32'sh38457abc, 32'sh3844bb28, 32'sh3843fb8b, 32'sh38433be5, 32'sh38427c36, 
               32'sh3841bc7f, 32'sh3840fcc0, 32'sh38403cf7, 32'sh383f7d26, 32'sh383ebd4c, 32'sh383dfd69, 32'sh383d3d7e, 32'sh383c7d8a, 
               32'sh383bbd8e, 32'sh383afd89, 32'sh383a3d7b, 32'sh38397d64, 32'sh3838bd45, 32'sh3837fd1d, 32'sh38373ced, 32'sh38367cb3, 
               32'sh3835bc71, 32'sh3834fc27, 32'sh38343bd4, 32'sh38337b78, 32'sh3832bb13, 32'sh3831faa6, 32'sh38313a30, 32'sh383079b2, 
               32'sh382fb92a, 32'sh382ef89a, 32'sh382e3802, 32'sh382d7761, 32'sh382cb6b7, 32'sh382bf604, 32'sh382b3549, 32'sh382a7485, 
               32'sh3829b3b9, 32'sh3828f2e3, 32'sh38283205, 32'sh3827711f, 32'sh3826b030, 32'sh3825ef38, 32'sh38252e37, 32'sh38246d2e, 
               32'sh3823ac1d, 32'sh3822eb02, 32'sh382229df, 32'sh382168b3, 32'sh3820a77f, 32'sh381fe642, 32'sh381f24fc, 32'sh381e63ad, 
               32'sh381da256, 32'sh381ce0f7, 32'sh381c1f8e, 32'sh381b5e1d, 32'sh381a9ca4, 32'sh3819db21, 32'sh38191996, 32'sh38185803, 
               32'sh38179666, 32'sh3816d4c2, 32'sh38161314, 32'sh3815515e, 32'sh38148f9f, 32'sh3813cdd7, 32'sh38130c07, 32'sh38124a2e, 
               32'sh3811884d, 32'sh3810c663, 32'sh38100470, 32'sh380f4275, 32'sh380e8071, 32'sh380dbe64, 32'sh380cfc4f, 32'sh380c3a31, 
               32'sh380b780a, 32'sh380ab5db, 32'sh3809f3a3, 32'sh38093162, 32'sh38086f19, 32'sh3807acc7, 32'sh3806ea6d, 32'sh3806280a, 
               32'sh3805659e, 32'sh3804a329, 32'sh3803e0ac, 32'sh38031e27, 32'sh38025b98, 32'sh38019902, 32'sh3800d662, 32'sh380013ba, 
               32'sh37ff5109, 32'sh37fe8e4f, 32'sh37fdcb8d, 32'sh37fd08c3, 32'sh37fc45ef, 32'sh37fb8313, 32'sh37fac02e, 32'sh37f9fd41, 
               32'sh37f93a4b, 32'sh37f8774d, 32'sh37f7b446, 32'sh37f6f136, 32'sh37f62e1d, 32'sh37f56afc, 32'sh37f4a7d2, 32'sh37f3e4a0, 
               32'sh37f32165, 32'sh37f25e22, 32'sh37f19ad5, 32'sh37f0d781, 32'sh37f01423, 32'sh37ef50bd, 32'sh37ee8d4e, 32'sh37edc9d7, 
               32'sh37ed0657, 32'sh37ec42ce, 32'sh37eb7f3d, 32'sh37eabba3, 32'sh37e9f801, 32'sh37e93456, 32'sh37e870a2, 32'sh37e7ace6, 
               32'sh37e6e921, 32'sh37e62553, 32'sh37e5617d, 32'sh37e49d9e, 32'sh37e3d9b7, 32'sh37e315c7, 32'sh37e251ce, 32'sh37e18dcd, 
               32'sh37e0c9c3, 32'sh37e005b0, 32'sh37df4195, 32'sh37de7d71, 32'sh37ddb945, 32'sh37dcf510, 32'sh37dc30d2, 32'sh37db6c8c, 
               32'sh37daa83d, 32'sh37d9e3e6, 32'sh37d91f86, 32'sh37d85b1d, 32'sh37d796ac, 32'sh37d6d232, 32'sh37d60daf, 32'sh37d54924, 
               32'sh37d48490, 32'sh37d3bff4, 32'sh37d2fb4f, 32'sh37d236a2, 32'sh37d171eb, 32'sh37d0ad2d, 32'sh37cfe865, 32'sh37cf2395, 
               32'sh37ce5ebd, 32'sh37cd99db, 32'sh37ccd4f2, 32'sh37cc0fff, 32'sh37cb4b04, 32'sh37ca8601, 32'sh37c9c0f4, 32'sh37c8fbe0, 
               32'sh37c836c2, 32'sh37c7719c, 32'sh37c6ac6d, 32'sh37c5e736, 32'sh37c521f6, 32'sh37c45cae, 32'sh37c3975d, 32'sh37c2d203, 
               32'sh37c20ca1, 32'sh37c14736, 32'sh37c081c3, 32'sh37bfbc47, 32'sh37bef6c2, 32'sh37be3135, 32'sh37bd6b9f, 32'sh37bca601, 
               32'sh37bbe05a, 32'sh37bb1aaa, 32'sh37ba54f2, 32'sh37b98f31, 32'sh37b8c968, 32'sh37b80396, 32'sh37b73dbb, 32'sh37b677d8, 
               32'sh37b5b1ec, 32'sh37b4ebf8, 32'sh37b425fb, 32'sh37b35ff5, 32'sh37b299e7, 32'sh37b1d3d1, 32'sh37b10db1, 32'sh37b04789, 
               32'sh37af8159, 32'sh37aebb20, 32'sh37adf4de, 32'sh37ad2e94, 32'sh37ac6841, 32'sh37aba1e6, 32'sh37aadb82, 32'sh37aa1515, 
               32'sh37a94ea0, 32'sh37a88822, 32'sh37a7c19c, 32'sh37a6fb0d, 32'sh37a63476, 32'sh37a56dd5, 32'sh37a4a72d, 32'sh37a3e07c, 
               32'sh37a319c2, 32'sh37a252ff, 32'sh37a18c34, 32'sh37a0c561, 32'sh379ffe85, 32'sh379f37a0, 32'sh379e70b3, 32'sh379da9bd, 
               32'sh379ce2be, 32'sh379c1bb7, 32'sh379b54a8, 32'sh379a8d90, 32'sh3799c66f, 32'sh3798ff46, 32'sh37983814, 32'sh379770d9, 
               32'sh3796a996, 32'sh3795e24a, 32'sh37951af6, 32'sh3794539a, 32'sh37938c34, 32'sh3792c4c6, 32'sh3791fd50, 32'sh379135d1, 
               32'sh37906e49, 32'sh378fa6b9, 32'sh378edf20, 32'sh378e177f, 32'sh378d4fd5, 32'sh378c8823, 32'sh378bc068, 32'sh378af8a4, 
               32'sh378a30d8, 32'sh37896903, 32'sh3788a126, 32'sh3787d940, 32'sh37871152, 32'sh3786495b, 32'sh3785815b, 32'sh3784b953, 
               32'sh3783f143, 32'sh37832929, 32'sh37826108, 32'sh378198dd, 32'sh3780d0aa, 32'sh3780086f, 32'sh377f402b, 32'sh377e77de, 
               32'sh377daf89, 32'sh377ce72b, 32'sh377c1ec5, 32'sh377b5656, 32'sh377a8ddf, 32'sh3779c55f, 32'sh3778fcd7, 32'sh37783446, 
               32'sh37776bac, 32'sh3776a30a, 32'sh3775da5f, 32'sh377511ac, 32'sh377448f0, 32'sh3773802c, 32'sh3772b75f, 32'sh3771ee8a, 
               32'sh377125ac, 32'sh37705cc5, 32'sh376f93d6, 32'sh376ecade, 32'sh376e01de, 32'sh376d38d5, 32'sh376c6fc4, 32'sh376ba6aa, 
               32'sh376add88, 32'sh376a145d, 32'sh37694b2a, 32'sh376881ee, 32'sh3767b8a9, 32'sh3766ef5c, 32'sh37662606, 32'sh37655ca8, 
               32'sh37649341, 32'sh3763c9d2, 32'sh3763005a, 32'sh376236da, 32'sh37616d51, 32'sh3760a3c0, 32'sh375fda26, 32'sh375f1083, 
               32'sh375e46d8, 32'sh375d7d25, 32'sh375cb368, 32'sh375be9a4, 32'sh375b1fd7, 32'sh375a5601, 32'sh37598c23, 32'sh3758c23c, 
               32'sh3757f84c, 32'sh37572e54, 32'sh37566454, 32'sh37559a4b, 32'sh3754d03a, 32'sh37540620, 32'sh37533bfd, 32'sh375271d2, 
               32'sh3751a79e, 32'sh3750dd62, 32'sh3750131e, 32'sh374f48d0, 32'sh374e7e7b, 32'sh374db41c, 32'sh374ce9b6, 32'sh374c1f46, 
               32'sh374b54ce, 32'sh374a8a4e, 32'sh3749bfc5, 32'sh3748f534, 32'sh37482a9a, 32'sh37475ff7, 32'sh3746954c, 32'sh3745ca99, 
               32'sh3744ffdd, 32'sh37443518, 32'sh37436a4b, 32'sh37429f75, 32'sh3741d497, 32'sh374109b1, 32'sh37403ec1, 32'sh373f73ca, 
               32'sh373ea8ca, 32'sh373dddc1, 32'sh373d12b0, 32'sh373c4796, 32'sh373b7c73, 32'sh373ab149, 32'sh3739e615, 32'sh37391ad9, 
               32'sh37384f95, 32'sh37378448, 32'sh3736b8f3, 32'sh3735ed95, 32'sh3735222f, 32'sh373456c0, 32'sh37338b48, 32'sh3732bfc8, 
               32'sh3731f440, 32'sh373128af, 32'sh37305d15, 32'sh372f9173, 32'sh372ec5c9, 32'sh372dfa16, 32'sh372d2e5a, 32'sh372c6296, 
               32'sh372b96ca, 32'sh372acaf4, 32'sh3729ff17, 32'sh37293331, 32'sh37286742, 32'sh37279b4b, 32'sh3726cf4c, 32'sh37260343, 
               32'sh37253733, 32'sh37246b1a, 32'sh37239ef8, 32'sh3722d2ce, 32'sh3722069b, 32'sh37213a60, 32'sh37206e1d, 32'sh371fa1d1, 
               32'sh371ed57c, 32'sh371e091f, 32'sh371d3cb9, 32'sh371c704b, 32'sh371ba3d4, 32'sh371ad755, 32'sh371a0ace, 32'sh37193e3e, 
               32'sh371871a5, 32'sh3717a504, 32'sh3716d85a, 32'sh37160ba8, 32'sh37153eee, 32'sh3714722a, 32'sh3713a55f, 32'sh3712d88b, 
               32'sh37120bae, 32'sh37113ec9, 32'sh371071dc, 32'sh370fa4e6, 32'sh370ed7e7, 32'sh370e0ae0, 32'sh370d3dd0, 32'sh370c70b8, 
               32'sh370ba398, 32'sh370ad66f, 32'sh370a093d, 32'sh37093c03, 32'sh37086ec1, 32'sh3707a176, 32'sh3706d423, 32'sh370606c7, 
               32'sh37053962, 32'sh37046bf5, 32'sh37039e80, 32'sh3702d102, 32'sh3702037c, 32'sh370135ed, 32'sh37006856, 32'sh36ff9ab6, 
               32'sh36fecd0e, 32'sh36fdff5d, 32'sh36fd31a4, 32'sh36fc63e2, 32'sh36fb9618, 32'sh36fac845, 32'sh36f9fa6a, 32'sh36f92c87, 
               32'sh36f85e9a, 32'sh36f790a6, 32'sh36f6c2a9, 32'sh36f5f4a3, 32'sh36f52695, 32'sh36f4587f, 32'sh36f38a60, 32'sh36f2bc38, 
               32'sh36f1ee09, 32'sh36f11fd0, 32'sh36f0518f, 32'sh36ef8346, 32'sh36eeb4f4, 32'sh36ede69a, 32'sh36ed1837, 32'sh36ec49cc, 
               32'sh36eb7b58, 32'sh36eaacdc, 32'sh36e9de58, 32'sh36e90fcb, 32'sh36e84135, 32'sh36e77297, 32'sh36e6a3f1, 32'sh36e5d542, 
               32'sh36e5068a, 32'sh36e437ca, 32'sh36e36902, 32'sh36e29a31, 32'sh36e1cb58, 32'sh36e0fc76, 32'sh36e02d8c, 32'sh36df5e99, 
               32'sh36de8f9e, 32'sh36ddc09b, 32'sh36dcf18f, 32'sh36dc227a, 32'sh36db535d, 32'sh36da8438, 32'sh36d9b50a, 32'sh36d8e5d3, 
               32'sh36d81695, 32'sh36d7474d, 32'sh36d677fe, 32'sh36d5a8a6, 32'sh36d4d945, 32'sh36d409dc, 32'sh36d33a6a, 32'sh36d26af0, 
               32'sh36d19b6e, 32'sh36d0cbe3, 32'sh36cffc50, 32'sh36cf2cb4, 32'sh36ce5d10, 32'sh36cd8d63, 32'sh36ccbdae, 32'sh36cbedf0, 
               32'sh36cb1e2a, 32'sh36ca4e5b, 32'sh36c97e85, 32'sh36c8aea5, 32'sh36c7debd, 32'sh36c70ecd, 32'sh36c63ed4, 32'sh36c56ed3, 
               32'sh36c49ec9, 32'sh36c3ceb7, 32'sh36c2fe9d, 32'sh36c22e7a, 32'sh36c15e4e, 32'sh36c08e1a, 32'sh36bfbdde, 32'sh36beed99, 
               32'sh36be1d4c, 32'sh36bd4cf6, 32'sh36bc7c98, 32'sh36bbac32, 32'sh36badbc3, 32'sh36ba0b4c, 32'sh36b93acc, 32'sh36b86a43, 
               32'sh36b799b3, 32'sh36b6c919, 32'sh36b5f878, 32'sh36b527ce, 32'sh36b4571b, 32'sh36b38660, 32'sh36b2b59d, 32'sh36b1e4d1, 
               32'sh36b113fd, 32'sh36b04320, 32'sh36af723b, 32'sh36aea14e, 32'sh36add058, 32'sh36acff5a, 32'sh36ac2e53, 32'sh36ab5d44, 
               32'sh36aa8c2c, 32'sh36a9bb0c, 32'sh36a8e9e3, 32'sh36a818b2, 32'sh36a74779, 32'sh36a67637, 32'sh36a5a4ed, 32'sh36a4d39a, 
               32'sh36a4023f, 32'sh36a330db, 32'sh36a25f70, 32'sh36a18dfb, 32'sh36a0bc7e, 32'sh369feaf9, 32'sh369f196b, 32'sh369e47d5, 
               32'sh369d7637, 32'sh369ca490, 32'sh369bd2e1, 32'sh369b0129, 32'sh369a2f69, 32'sh36995da0, 32'sh36988bcf, 32'sh3697b9f6, 
               32'sh3696e814, 32'sh36961629, 32'sh36954437, 32'sh3694723c, 32'sh3693a038, 32'sh3692ce2c, 32'sh3691fc18, 32'sh369129fb, 
               32'sh369057d6, 32'sh368f85a8, 32'sh368eb372, 32'sh368de134, 32'sh368d0eed, 32'sh368c3c9e, 32'sh368b6a46, 32'sh368a97e6, 
               32'sh3689c57d, 32'sh3688f30c, 32'sh36882093, 32'sh36874e11, 32'sh36867b87, 32'sh3685a8f5, 32'sh3684d65a, 32'sh368403b6, 
               32'sh3683310b, 32'sh36825e56, 32'sh36818b9a, 32'sh3680b8d5, 32'sh367fe608, 32'sh367f1332, 32'sh367e4054, 32'sh367d6d6d, 
               32'sh367c9a7e, 32'sh367bc787, 32'sh367af487, 32'sh367a217e, 32'sh36794e6e, 32'sh36787b55, 32'sh3677a833, 32'sh3676d50a, 
               32'sh367601d7, 32'sh36752e9d, 32'sh36745b5a, 32'sh3673880e, 32'sh3672b4bb, 32'sh3671e15e, 32'sh36710dfa, 32'sh36703a8d, 
               32'sh366f6717, 32'sh366e939a, 32'sh366dc013, 32'sh366cec85, 32'sh366c18ee, 32'sh366b454f, 32'sh366a71a7, 32'sh36699df7, 
               32'sh3668ca3e, 32'sh3667f67d, 32'sh366722b4, 32'sh36664ee2, 32'sh36657b08, 32'sh3664a726, 32'sh3663d33b, 32'sh3662ff48, 
               32'sh36622b4c, 32'sh36615748, 32'sh3660833b, 32'sh365faf27, 32'sh365edb09, 32'sh365e06e4, 32'sh365d32b6, 32'sh365c5e80, 
               32'sh365b8a41, 32'sh365ab5fa, 32'sh3659e1aa, 32'sh36590d52, 32'sh365838f2, 32'sh3657648a, 32'sh36569019, 32'sh3655bb9f, 
               32'sh3654e71d, 32'sh36541293, 32'sh36533e01, 32'sh36526966, 32'sh365194c3, 32'sh3650c017, 32'sh364feb63, 32'sh364f16a6, 
               32'sh364e41e2, 32'sh364d6d15, 32'sh364c983f, 32'sh364bc361, 32'sh364aee7b, 32'sh364a198c, 32'sh36494495, 32'sh36486f96, 
               32'sh36479a8e, 32'sh3646c57e, 32'sh3645f065, 32'sh36451b44, 32'sh3644461b, 32'sh364370ea, 32'sh36429bb0, 32'sh3641c66d, 
               32'sh3640f123, 32'sh36401bd0, 32'sh363f4674, 32'sh363e7110, 32'sh363d9ba4, 32'sh363cc630, 32'sh363bf0b3, 32'sh363b1b2d, 
               32'sh363a45a0, 32'sh3639700a, 32'sh36389a6b, 32'sh3637c4c5, 32'sh3636ef16, 32'sh3636195e, 32'sh3635439e, 32'sh36346dd6, 
               32'sh36339806, 32'sh3632c22d, 32'sh3631ec4c, 32'sh36311662, 32'sh36304070, 32'sh362f6a76, 32'sh362e9473, 32'sh362dbe68, 
               32'sh362ce855, 32'sh362c1239, 32'sh362b3c15, 32'sh362a65e8, 32'sh36298fb4, 32'sh3628b976, 32'sh3627e331, 32'sh36270ce3, 
               32'sh3626368d, 32'sh3625602e, 32'sh362489c7, 32'sh3623b358, 32'sh3622dce1, 32'sh36220661, 32'sh36212fd8, 32'sh36205948, 
               32'sh361f82af, 32'sh361eac0d, 32'sh361dd564, 32'sh361cfeb2, 32'sh361c27f7, 32'sh361b5135, 32'sh361a7a6a, 32'sh3619a396, 
               32'sh3618ccba, 32'sh3617f5d6, 32'sh36171eea, 32'sh361647f5, 32'sh361570f8, 32'sh361499f3, 32'sh3613c2e5, 32'sh3612ebcf, 
               32'sh361214b0, 32'sh36113d89, 32'sh3610665a, 32'sh360f8f23, 32'sh360eb7e3, 32'sh360de09b, 32'sh360d094a, 32'sh360c31f1, 
               32'sh360b5a90, 32'sh360a8327, 32'sh3609abb5, 32'sh3608d43b, 32'sh3607fcb8, 32'sh3607252d, 32'sh36064d9a, 32'sh360575ff, 
               32'sh36049e5b, 32'sh3603c6af, 32'sh3602eefa, 32'sh3602173e, 32'sh36013f78, 32'sh360067ab, 32'sh35ff8fd5, 32'sh35feb7f7, 
               32'sh35fde011, 32'sh35fd0822, 32'sh35fc302b, 32'sh35fb582b, 32'sh35fa8023, 32'sh35f9a813, 32'sh35f8cffb, 32'sh35f7f7da, 
               32'sh35f71fb1, 32'sh35f64780, 32'sh35f56f46, 32'sh35f49704, 32'sh35f3beba, 32'sh35f2e667, 32'sh35f20e0c, 32'sh35f135a9, 
               32'sh35f05d3d, 32'sh35ef84c9, 32'sh35eeac4d, 32'sh35edd3c9, 32'sh35ecfb3c, 32'sh35ec22a7, 32'sh35eb4a09, 32'sh35ea7163, 
               32'sh35e998b5, 32'sh35e8bfff, 32'sh35e7e740, 32'sh35e70e79, 32'sh35e635a9, 32'sh35e55cd2, 32'sh35e483f2, 32'sh35e3ab09, 
               32'sh35e2d219, 32'sh35e1f920, 32'sh35e1201e, 32'sh35e04715, 32'sh35df6e03, 32'sh35de94e9, 32'sh35ddbbc6, 32'sh35dce29c, 
               32'sh35dc0968, 32'sh35db302d, 32'sh35da56e9, 32'sh35d97d9d, 32'sh35d8a449, 32'sh35d7caec, 32'sh35d6f187, 32'sh35d6181a, 
               32'sh35d53ea5, 32'sh35d46527, 32'sh35d38ba1, 32'sh35d2b212, 32'sh35d1d87c, 32'sh35d0fedd, 32'sh35d02535, 32'sh35cf4b86, 
               32'sh35ce71ce, 32'sh35cd980d, 32'sh35ccbe45, 32'sh35cbe474, 32'sh35cb0a9b, 32'sh35ca30b9, 32'sh35c956d0, 32'sh35c87cde, 
               32'sh35c7a2e3, 32'sh35c6c8e1, 32'sh35c5eed6, 32'sh35c514c3, 32'sh35c43aa7, 32'sh35c36084, 32'sh35c28658, 32'sh35c1ac23, 
               32'sh35c0d1e7, 32'sh35bff7a2, 32'sh35bf1d54, 32'sh35be42ff, 32'sh35bd68a1, 32'sh35bc8e3b, 32'sh35bbb3cd, 32'sh35bad956, 
               32'sh35b9fed7, 32'sh35b92450, 32'sh35b849c0, 32'sh35b76f29, 32'sh35b69489, 32'sh35b5b9e0, 32'sh35b4df30, 32'sh35b40477, 
               32'sh35b329b5, 32'sh35b24eec, 32'sh35b1741a, 32'sh35b09940, 32'sh35afbe5e, 32'sh35aee373, 32'sh35ae0880, 32'sh35ad2d85, 
               32'sh35ac5282, 32'sh35ab7776, 32'sh35aa9c62, 32'sh35a9c146, 32'sh35a8e621, 32'sh35a80af4, 32'sh35a72fbf, 32'sh35a65482, 
               32'sh35a5793c, 32'sh35a49dee, 32'sh35a3c298, 32'sh35a2e73a, 32'sh35a20bd3, 32'sh35a13064, 32'sh35a054ed, 32'sh359f796d, 
               32'sh359e9de5, 32'sh359dc255, 32'sh359ce6bd, 32'sh359c0b1c, 32'sh359b2f73, 32'sh359a53c2, 32'sh35997809, 32'sh35989c47, 
               32'sh3597c07d, 32'sh3596e4ab, 32'sh359608d1, 32'sh35952cee, 32'sh35945103, 32'sh35937510, 32'sh35929914, 32'sh3591bd10, 
               32'sh3590e104, 32'sh359004f0, 32'sh358f28d3, 32'sh358e4caf, 32'sh358d7081, 32'sh358c944c, 32'sh358bb80e, 32'sh358adbc9, 
               32'sh3589ff7a, 32'sh35892324, 32'sh358846c5, 32'sh35876a5f, 32'sh35868def, 32'sh3585b178, 32'sh3584d4f8, 32'sh3583f871, 
               32'sh35831be0, 32'sh35823f48, 32'sh358162a7, 32'sh358085fe, 32'sh357fa94d, 32'sh357ecc94, 32'sh357defd2, 32'sh357d1308, 
               32'sh357c3636, 32'sh357b595c, 32'sh357a7c79, 32'sh35799f8e, 32'sh3578c29b, 32'sh3577e5a0, 32'sh3577089c, 32'sh35762b90, 
               32'sh35754e7c, 32'sh35747160, 32'sh3573943b, 32'sh3572b70e, 32'sh3571d9d9, 32'sh3570fc9c, 32'sh35701f56, 32'sh356f4208, 
               32'sh356e64b2, 32'sh356d8754, 32'sh356ca9ed, 32'sh356bcc7f, 32'sh356aef08, 32'sh356a1188, 32'sh35693401, 32'sh35685671, 
               32'sh356778d9, 32'sh35669b39, 32'sh3565bd90, 32'sh3564dfe0, 32'sh35640227, 32'sh35632466, 32'sh3562469c, 32'sh356168cb, 
               32'sh35608af1, 32'sh355fad0f, 32'sh355ecf25, 32'sh355df132, 32'sh355d1337, 32'sh355c3534, 32'sh355b5729, 32'sh355a7916, 
               32'sh35599afa, 32'sh3558bcd6, 32'sh3557deaa, 32'sh35570076, 32'sh35562239, 32'sh355543f4, 32'sh355465a7, 32'sh35538752, 
               32'sh3552a8f4, 32'sh3551ca8f, 32'sh3550ec21, 32'sh35500dab, 32'sh354f2f2c, 32'sh354e50a6, 32'sh354d7217, 32'sh354c9380, 
               32'sh354bb4e1, 32'sh354ad639, 32'sh3549f789, 32'sh354918d1, 32'sh35483a11, 32'sh35475b49, 32'sh35467c78, 32'sh35459da0, 
               32'sh3544bebf, 32'sh3543dfd6, 32'sh354300e4, 32'sh354221ea, 32'sh354142e9, 32'sh354063df, 32'sh353f84cc, 32'sh353ea5b2, 
               32'sh353dc68f, 32'sh353ce764, 32'sh353c0831, 32'sh353b28f6, 32'sh353a49b2, 32'sh35396a67, 32'sh35388b13, 32'sh3537abb6, 
               32'sh3536cc52, 32'sh3535ece6, 32'sh35350d71, 32'sh35342df4, 32'sh35334e6f, 32'sh35326ee1, 32'sh35318f4c, 32'sh3530afae, 
               32'sh352fd008, 32'sh352ef05a, 32'sh352e10a3, 32'sh352d30e5, 32'sh352c511e, 32'sh352b714f, 32'sh352a9178, 32'sh3529b198, 
               32'sh3528d1b1, 32'sh3527f1c1, 32'sh352711c9, 32'sh352631c9, 32'sh352551c0, 32'sh352471b0, 32'sh35239197, 32'sh3522b176, 
               32'sh3521d14d, 32'sh3520f11c, 32'sh352010e2, 32'sh351f30a0, 32'sh351e5056, 32'sh351d7004, 32'sh351c8faa, 32'sh351baf47, 
               32'sh351acedd, 32'sh3519ee6a, 32'sh35190def, 32'sh35182d6b, 32'sh35174ce0, 32'sh35166c4c, 32'sh35158bb1, 32'sh3514ab0d, 
               32'sh3513ca60, 32'sh3512e9ac, 32'sh351208ef, 32'sh3511282b, 32'sh3510475e, 32'sh350f6689, 32'sh350e85ab, 32'sh350da4c6, 
               32'sh350cc3d8, 32'sh350be2e2, 32'sh350b01e4, 32'sh350a20de, 32'sh35093fd0, 32'sh35085eb9, 32'sh35077d9a, 32'sh35069c73, 
               32'sh3505bb44, 32'sh3504da0d, 32'sh3503f8ce, 32'sh35031786, 32'sh35023636, 32'sh350154de, 32'sh3500737e, 32'sh34ff9216, 
               32'sh34feb0a5, 32'sh34fdcf2d, 32'sh34fcedac, 32'sh34fc0c23, 32'sh34fb2a92, 32'sh34fa48f8, 32'sh34f96757, 32'sh34f885ad, 
               32'sh34f7a3fb, 32'sh34f6c241, 32'sh34f5e07f, 32'sh34f4feb5, 32'sh34f41ce2, 32'sh34f33b07, 32'sh34f25924, 32'sh34f17739, 
               32'sh34f09546, 32'sh34efb34b, 32'sh34eed147, 32'sh34edef3c, 32'sh34ed0d28, 32'sh34ec2b0c, 32'sh34eb48e8, 32'sh34ea66bb, 
               32'sh34e98487, 32'sh34e8a24a, 32'sh34e7c005, 32'sh34e6ddb8, 32'sh34e5fb63, 32'sh34e51906, 32'sh34e436a1, 32'sh34e35433, 
               32'sh34e271bd, 32'sh34e18f3f, 32'sh34e0acb9, 32'sh34dfca2b, 32'sh34dee795, 32'sh34de04f6, 32'sh34dd224f, 32'sh34dc3fa1, 
               32'sh34db5cea, 32'sh34da7a2b, 32'sh34d99763, 32'sh34d8b494, 32'sh34d7d1bc, 32'sh34d6eedd, 32'sh34d60bf5, 32'sh34d52905, 
               32'sh34d4460c, 32'sh34d3630c, 32'sh34d28004, 32'sh34d19cf3, 32'sh34d0b9da, 32'sh34cfd6b9, 32'sh34cef390, 32'sh34ce105f, 
               32'sh34cd2d26, 32'sh34cc49e4, 32'sh34cb669b, 32'sh34ca8349, 32'sh34c99fef, 32'sh34c8bc8d, 32'sh34c7d923, 32'sh34c6f5b0, 
               32'sh34c61236, 32'sh34c52eb3, 32'sh34c44b29, 32'sh34c36796, 32'sh34c283fb, 32'sh34c1a058, 32'sh34c0bcac, 32'sh34bfd8f9, 
               32'sh34bef53d, 32'sh34be117a, 32'sh34bd2dae, 32'sh34bc49da, 32'sh34bb65fe, 32'sh34ba821a, 32'sh34b99e2d, 32'sh34b8ba39, 
               32'sh34b7d63c, 32'sh34b6f237, 32'sh34b60e2b, 32'sh34b52a16, 32'sh34b445f8, 32'sh34b361d3, 32'sh34b27da6, 32'sh34b19970, 
               32'sh34b0b533, 32'sh34afd0ed, 32'sh34aeec9f, 32'sh34ae0849, 32'sh34ad23eb, 32'sh34ac3f85, 32'sh34ab5b16, 32'sh34aa76a0, 
               32'sh34a99221, 32'sh34a8ad9a, 32'sh34a7c90c, 32'sh34a6e475, 32'sh34a5ffd5, 32'sh34a51b2e, 32'sh34a4367f, 32'sh34a351c7, 
               32'sh34a26d08, 32'sh34a18840, 32'sh34a0a370, 32'sh349fbe98, 32'sh349ed9b8, 32'sh349df4d0, 32'sh349d0fe0, 32'sh349c2ae8, 
               32'sh349b45e7, 32'sh349a60de, 32'sh34997bce, 32'sh349896b5, 32'sh3497b194, 32'sh3496cc6b, 32'sh3495e73a, 32'sh34950200, 
               32'sh34941cbf, 32'sh34933776, 32'sh34925224, 32'sh34916cca, 32'sh34908768, 32'sh348fa1ff, 32'sh348ebc8d, 32'sh348dd712, 
               32'sh348cf190, 32'sh348c0c06, 32'sh348b2673, 32'sh348a40d9, 32'sh34895b36, 32'sh3488758b, 32'sh34878fd9, 32'sh3486aa1e, 
               32'sh3485c45b, 32'sh3484de8f, 32'sh3483f8bc, 32'sh348312e1, 32'sh34822cfd, 32'sh34814712, 32'sh3480611e, 32'sh347f7b22, 
               32'sh347e951f, 32'sh347daf13, 32'sh347cc8ff, 32'sh347be2e3, 32'sh347afcbe, 32'sh347a1692, 32'sh3479305e, 32'sh34784a21, 
               32'sh347763dd, 32'sh34767d90, 32'sh3475973b, 32'sh3474b0de, 32'sh3473ca79, 32'sh3472e40c, 32'sh3471fd97, 32'sh3471171a, 
               32'sh34703095, 32'sh346f4a07, 32'sh346e6372, 32'sh346d7cd4, 32'sh346c962f, 32'sh346baf81, 32'sh346ac8cb, 32'sh3469e20d, 
               32'sh3468fb47, 32'sh34681479, 32'sh34672da3, 32'sh346646c5, 32'sh34655fdf, 32'sh346478f0, 32'sh346391fa, 32'sh3462aafb, 
               32'sh3461c3f5, 32'sh3460dce6, 32'sh345ff5cf, 32'sh345f0eb0, 32'sh345e2789, 32'sh345d405a, 32'sh345c5923, 32'sh345b71e4, 
               32'sh345a8a9d, 32'sh3459a34e, 32'sh3458bbf6, 32'sh3457d497, 32'sh3456ed2f, 32'sh345605c0, 32'sh34551e48, 32'sh345436c8, 
               32'sh34534f41, 32'sh345267b1, 32'sh34518019, 32'sh34509879, 32'sh344fb0d1, 32'sh344ec921, 32'sh344de168, 32'sh344cf9a8, 
               32'sh344c11e0, 32'sh344b2a0f, 32'sh344a4237, 32'sh34495a56, 32'sh3448726e, 32'sh34478a7d, 32'sh3446a284, 32'sh3445ba84, 
               32'sh3444d27b, 32'sh3443ea6a, 32'sh34430251, 32'sh34421a30, 32'sh34413207, 32'sh344049d6, 32'sh343f619c, 32'sh343e795b, 
               32'sh343d9112, 32'sh343ca8c1, 32'sh343bc067, 32'sh343ad806, 32'sh3439ef9c, 32'sh3439072b, 32'sh34381eb1, 32'sh3437362f, 
               32'sh34364da6, 32'sh34356514, 32'sh34347c7a, 32'sh343393d8, 32'sh3432ab2e, 32'sh3431c27c, 32'sh3430d9c2, 32'sh342ff100, 
               32'sh342f0836, 32'sh342e1f64, 32'sh342d3689, 32'sh342c4da7, 32'sh342b64bd, 32'sh342a7bca, 32'sh342992d0, 32'sh3428a9cd, 
               32'sh3427c0c3, 32'sh3426d7b0, 32'sh3425ee96, 32'sh34250573, 32'sh34241c49, 32'sh34233316, 32'sh342249db, 32'sh34216098, 
               32'sh3420774d, 32'sh341f8dfb, 32'sh341ea4a0, 32'sh341dbb3d, 32'sh341cd1d2, 32'sh341be85f, 32'sh341afee4, 32'sh341a1561, 
               32'sh34192bd5, 32'sh34184242, 32'sh341758a7, 32'sh34166f04, 32'sh34158559, 32'sh34149ba5, 32'sh3413b1ea, 32'sh3412c827, 
               32'sh3411de5b, 32'sh3410f488, 32'sh34100aac, 32'sh340f20c9, 32'sh340e36dd, 32'sh340d4cea, 32'sh340c62ee, 32'sh340b78eb, 
               32'sh340a8edf, 32'sh3409a4cc, 32'sh3408bab0, 32'sh3407d08c, 32'sh3406e660, 32'sh3405fc2d, 32'sh340511f1, 32'sh340427ad, 
               32'sh34033d61, 32'sh3402530e, 32'sh340168b2, 32'sh34007e4e, 32'sh33ff93e2, 32'sh33fea96e, 32'sh33fdbef2, 32'sh33fcd46e, 
               32'sh33fbe9e2, 32'sh33faff4e, 32'sh33fa14b2, 32'sh33f92a0e, 32'sh33f83f62, 32'sh33f754ae, 32'sh33f669f2, 32'sh33f57f2e, 
               32'sh33f49462, 32'sh33f3a98e, 32'sh33f2beb2, 32'sh33f1d3ce, 32'sh33f0e8e2, 32'sh33effdee, 32'sh33ef12f2, 32'sh33ee27ed, 
               32'sh33ed3ce1, 32'sh33ec51cd, 32'sh33eb66b1, 32'sh33ea7b8d, 32'sh33e99061, 32'sh33e8a52d, 32'sh33e7b9f0, 32'sh33e6ceac, 
               32'sh33e5e360, 32'sh33e4f80c, 32'sh33e40cb0, 32'sh33e3214b, 32'sh33e235df, 32'sh33e14a6b, 32'sh33e05eef, 32'sh33df736b, 
               32'sh33de87de, 32'sh33dd9c4a, 32'sh33dcb0ae, 32'sh33dbc50a, 32'sh33dad95e, 32'sh33d9eda9, 32'sh33d901ed, 32'sh33d81629, 
               32'sh33d72a5d, 32'sh33d63e89, 32'sh33d552ac, 32'sh33d466c8, 32'sh33d37adc, 32'sh33d28ee8, 32'sh33d1a2ec, 32'sh33d0b6e8, 
               32'sh33cfcadc, 32'sh33cedec7, 32'sh33cdf2ab, 32'sh33cd0687, 32'sh33cc1a5b, 32'sh33cb2e27, 32'sh33ca41eb, 32'sh33c955a7, 
               32'sh33c8695b, 32'sh33c77d07, 32'sh33c690ab, 32'sh33c5a447, 32'sh33c4b7db, 32'sh33c3cb67, 32'sh33c2deeb, 32'sh33c1f267, 
               32'sh33c105db, 32'sh33c01948, 32'sh33bf2cac, 32'sh33be4008, 32'sh33bd535c, 32'sh33bc66a8, 32'sh33bb79ec, 32'sh33ba8d29, 
               32'sh33b9a05d, 32'sh33b8b389, 32'sh33b7c6ae, 32'sh33b6d9ca, 32'sh33b5ecde, 32'sh33b4ffeb, 32'sh33b412ef, 32'sh33b325ec, 
               32'sh33b238e0, 32'sh33b14bcd, 32'sh33b05eb1, 32'sh33af718e, 32'sh33ae8462, 32'sh33ad972f, 32'sh33aca9f4, 32'sh33abbcb0, 
               32'sh33aacf65, 32'sh33a9e212, 32'sh33a8f4b6, 32'sh33a80753, 32'sh33a719e8, 32'sh33a62c75, 32'sh33a53efa, 32'sh33a45177, 
               32'sh33a363ec, 32'sh33a27659, 32'sh33a188be, 32'sh33a09b1b, 32'sh339fad70, 32'sh339ebfbd, 32'sh339dd203, 32'sh339ce440, 
               32'sh339bf675, 32'sh339b08a2, 32'sh339a1ac8, 32'sh33992ce5, 32'sh33983efb, 32'sh33975108, 32'sh3396630e, 32'sh3395750b, 
               32'sh33948701, 32'sh339398ef, 32'sh3392aad4, 32'sh3391bcb2, 32'sh3390ce88, 32'sh338fe056, 32'sh338ef21c, 32'sh338e03da, 
               32'sh338d1590, 32'sh338c273e, 32'sh338b38e4, 32'sh338a4a82, 32'sh33895c18, 32'sh33886da7, 32'sh33877f2d, 32'sh338690ab, 
               32'sh3385a222, 32'sh3384b390, 32'sh3383c4f7, 32'sh3382d656, 32'sh3381e7ac, 32'sh3380f8fb, 32'sh33800a42, 32'sh337f1b81, 
               32'sh337e2cb7, 32'sh337d3de6, 32'sh337c4f0d, 32'sh337b602c, 32'sh337a7144, 32'sh33798253, 32'sh3378935a, 32'sh3377a459, 
               32'sh3376b551, 32'sh3375c640, 32'sh3374d728, 32'sh3373e807, 32'sh3372f8df, 32'sh337209af, 32'sh33711a76, 32'sh33702b36, 
               32'sh336f3bee, 32'sh336e4c9e, 32'sh336d5d46, 32'sh336c6de6, 32'sh336b7e7e, 32'sh336a8f0f, 32'sh33699f97, 32'sh3368b017, 
               32'sh3367c090, 32'sh3366d100, 32'sh3365e169, 32'sh3364f1ca, 32'sh33640223, 32'sh33631273, 32'sh336222bc, 32'sh336132fd, 
               32'sh33604336, 32'sh335f5367, 32'sh335e6391, 32'sh335d73b2, 32'sh335c83cb, 32'sh335b93dd, 32'sh335aa3e6, 32'sh3359b3e8, 
               32'sh3358c3e2, 32'sh3357d3d3, 32'sh3356e3bd, 32'sh3355f39f, 32'sh33550379, 32'sh3354134b, 32'sh33532316, 32'sh335232d8, 
               32'sh33514292, 32'sh33505245, 32'sh334f61ef, 32'sh334e7192, 32'sh334d812d, 32'sh334c90bf, 32'sh334ba04a, 32'sh334aafcd, 
               32'sh3349bf48, 32'sh3348cebc, 32'sh3347de27, 32'sh3346ed8a, 32'sh3345fce6, 32'sh33450c39, 32'sh33441b85, 32'sh33432ac8, 
               32'sh33423a04, 32'sh33414938, 32'sh33405864, 32'sh333f6788, 32'sh333e76a4, 32'sh333d85b9, 32'sh333c94c5, 32'sh333ba3ca, 
               32'sh333ab2c6, 32'sh3339c1bb, 32'sh3338d0a8, 32'sh3337df8d, 32'sh3336ee6a, 32'sh3335fd3f, 32'sh33350c0c, 32'sh33341ad1, 
               32'sh3333298f, 32'sh33323844, 32'sh333146f2, 32'sh33305597, 32'sh332f6435, 32'sh332e72cb, 32'sh332d8159, 32'sh332c8fdf, 
               32'sh332b9e5e, 32'sh332aacd4, 32'sh3329bb43, 32'sh3328c9a9, 32'sh3327d808, 32'sh3326e65f, 32'sh3325f4ae, 32'sh332502f5, 
               32'sh33241134, 32'sh33231f6b, 32'sh33222d9a, 32'sh33213bc2, 32'sh332049e1, 32'sh331f57f9, 32'sh331e6609, 32'sh331d7411, 
               32'sh331c8211, 32'sh331b9009, 32'sh331a9dfa, 32'sh3319abe2, 32'sh3318b9c2, 32'sh3317c79b, 32'sh3316d56c, 32'sh3315e335, 
               32'sh3314f0f6, 32'sh3313feaf, 32'sh33130c60, 32'sh33121a0a, 32'sh331127ab, 32'sh33103545, 32'sh330f42d7, 32'sh330e5061, 
               32'sh330d5de3, 32'sh330c6b5d, 32'sh330b78cf, 32'sh330a8639, 32'sh3309939c, 32'sh3308a0f7, 32'sh3307ae49, 32'sh3306bb94, 
               32'sh3305c8d7, 32'sh3304d613, 32'sh3303e346, 32'sh3302f071, 32'sh3301fd95, 32'sh33010ab1, 32'sh330017c4, 32'sh32ff24d0, 
               32'sh32fe31d5, 32'sh32fd3ed1, 32'sh32fc4bc5, 32'sh32fb58b2, 32'sh32fa6596, 32'sh32f97273, 32'sh32f87f48, 32'sh32f78c15, 
               32'sh32f698db, 32'sh32f5a598, 32'sh32f4b24d, 32'sh32f3befb, 32'sh32f2cba1, 32'sh32f1d83f, 32'sh32f0e4d5, 32'sh32eff163, 
               32'sh32eefdea, 32'sh32ee0a68, 32'sh32ed16df, 32'sh32ec234e, 32'sh32eb2fb5, 32'sh32ea3c14, 32'sh32e9486b, 32'sh32e854ba, 
               32'sh32e76102, 32'sh32e66d42, 32'sh32e57979, 32'sh32e485a9, 32'sh32e391d2, 32'sh32e29df2, 32'sh32e1aa0a, 32'sh32e0b61b, 
               32'sh32dfc224, 32'sh32dece25, 32'sh32ddda1e, 32'sh32dce60f, 32'sh32dbf1f8, 32'sh32dafdda, 32'sh32da09b4, 32'sh32d91585, 
               32'sh32d82150, 32'sh32d72d12, 32'sh32d638cc, 32'sh32d5447f, 32'sh32d45029, 32'sh32d35bcc, 32'sh32d26767, 32'sh32d172fa, 
               32'sh32d07e85, 32'sh32cf8a09, 32'sh32ce9585, 32'sh32cda0f8, 32'sh32ccac64, 32'sh32cbb7c9, 32'sh32cac325, 32'sh32c9ce79, 
               32'sh32c8d9c6, 32'sh32c7e50b, 32'sh32c6f048, 32'sh32c5fb7d, 32'sh32c506aa, 32'sh32c411d0, 32'sh32c31ced, 32'sh32c22803, 
               32'sh32c13311, 32'sh32c03e17, 32'sh32bf4916, 32'sh32be540c, 32'sh32bd5efb, 32'sh32bc69e2, 32'sh32bb74c1, 32'sh32ba7f98, 
               32'sh32b98a67, 32'sh32b8952f, 32'sh32b79fef, 32'sh32b6aaa7, 32'sh32b5b557, 32'sh32b4bfff, 32'sh32b3caa0, 32'sh32b2d538, 
               32'sh32b1dfc9, 32'sh32b0ea52, 32'sh32aff4d3, 32'sh32aeff4d, 32'sh32ae09be, 32'sh32ad1428, 32'sh32ac1e8a, 32'sh32ab28e4, 
               32'sh32aa3336, 32'sh32a93d81, 32'sh32a847c4, 32'sh32a751ff, 32'sh32a65c32, 32'sh32a5665d, 32'sh32a47080, 32'sh32a37a9c, 
               32'sh32a284b0, 32'sh32a18ebc, 32'sh32a098c0, 32'sh329fa2bc, 32'sh329eacb1, 32'sh329db69e, 32'sh329cc083, 32'sh329bca60, 
               32'sh329ad435, 32'sh3299de03, 32'sh3298e7c9, 32'sh3297f187, 32'sh3296fb3d, 32'sh329604eb, 32'sh32950e92, 32'sh32941830, 
               32'sh329321c7, 32'sh32922b57, 32'sh329134de, 32'sh32903e5d, 32'sh328f47d5, 32'sh328e5145, 32'sh328d5aad, 32'sh328c640e, 
               32'sh328b6d66, 32'sh328a76b7, 32'sh32898000, 32'sh32888941, 32'sh3287927b, 32'sh32869bac, 32'sh3285a4d6, 32'sh3284adf8, 
               32'sh3283b712, 32'sh3282c025, 32'sh3281c92f, 32'sh3280d232, 32'sh327fdb2d, 32'sh327ee421, 32'sh327ded0c, 32'sh327cf5f0, 
               32'sh327bfecc, 32'sh327b07a0, 32'sh327a106c, 32'sh32791931, 32'sh327821ee, 32'sh32772aa3, 32'sh32763350, 32'sh32753bf5, 
               32'sh32744493, 32'sh32734d29, 32'sh327255b7, 32'sh32715e3d, 32'sh327066bc, 32'sh326f6f33, 32'sh326e77a2, 32'sh326d8009, 
               32'sh326c8868, 32'sh326b90c0, 32'sh326a9910, 32'sh3269a158, 32'sh3268a998, 32'sh3267b1d1, 32'sh3266ba02, 32'sh3265c22b, 
               32'sh3264ca4c, 32'sh3263d266, 32'sh3262da77, 32'sh3261e281, 32'sh3260ea83, 32'sh325ff27e, 32'sh325efa70, 32'sh325e025b, 
               32'sh325d0a3e, 32'sh325c121a, 32'sh325b19ed, 32'sh325a21b9, 32'sh3259297d, 32'sh32583139, 32'sh325738ee, 32'sh3256409b, 
               32'sh32554840, 32'sh32544fdd, 32'sh32535772, 32'sh32525f00, 32'sh32516686, 32'sh32506e04, 32'sh324f757a, 32'sh324e7ce9, 
               32'sh324d8450, 32'sh324c8baf, 32'sh324b9306, 32'sh324a9a56, 32'sh3249a19e, 32'sh3248a8de, 32'sh3247b016, 32'sh3246b747, 
               32'sh3245be70, 32'sh3244c591, 32'sh3243ccaa, 32'sh3242d3bc, 32'sh3241dac6, 32'sh3240e1c8, 32'sh323fe8c2, 32'sh323eefb5, 
               32'sh323df6a0, 32'sh323cfd83, 32'sh323c045e, 32'sh323b0b32, 32'sh323a11fe, 32'sh323918c2, 32'sh32381f7e, 32'sh32372633, 
               32'sh32362ce0, 32'sh32353385, 32'sh32343a22, 32'sh323340b8, 32'sh32324746, 32'sh32314dcc, 32'sh3230544a, 32'sh322f5ac1, 
               32'sh322e6130, 32'sh322d6797, 32'sh322c6df7, 32'sh322b744e, 32'sh322a7a9e, 32'sh322980e7, 32'sh32288727, 32'sh32278d60, 
               32'sh32269391, 32'sh322599ba, 32'sh32249fdc, 32'sh3223a5f6, 32'sh3222ac08, 32'sh3221b212, 32'sh3220b815, 32'sh321fbe10, 
               32'sh321ec403, 32'sh321dc9ef, 32'sh321ccfd2, 32'sh321bd5ae, 32'sh321adb83, 32'sh3219e14f, 32'sh3218e714, 32'sh3217ecd1, 
               32'sh3216f287, 32'sh3215f834, 32'sh3214fdda, 32'sh32140379, 32'sh3213090f, 32'sh32120e9e, 32'sh32111425, 32'sh321019a4, 
               32'sh320f1f1c, 32'sh320e248c, 32'sh320d29f4, 32'sh320c2f54, 32'sh320b34ad, 32'sh320a39fe, 32'sh32093f47, 32'sh32084489, 
               32'sh320749c3, 32'sh32064ef5, 32'sh3205541f, 32'sh32045942, 32'sh32035e5d, 32'sh32026370, 32'sh3201687c, 32'sh32006d80, 
               32'sh31ff727c, 32'sh31fe7771, 32'sh31fd7c5d, 32'sh31fc8142, 32'sh31fb8620, 32'sh31fa8af5, 32'sh31f98fc3, 32'sh31f89489, 
               32'sh31f79948, 32'sh31f69dff, 32'sh31f5a2ae, 32'sh31f4a755, 32'sh31f3abf5, 32'sh31f2b08d, 32'sh31f1b51d, 32'sh31f0b9a6, 
               32'sh31efbe27, 32'sh31eec2a0, 32'sh31edc711, 32'sh31eccb7b, 32'sh31ebcfdd, 32'sh31ead437, 32'sh31e9d88a, 32'sh31e8dcd5, 
               32'sh31e7e118, 32'sh31e6e554, 32'sh31e5e988, 32'sh31e4edb4, 32'sh31e3f1d8, 32'sh31e2f5f5, 32'sh31e1fa0a, 32'sh31e0fe18, 
               32'sh31e0021e, 32'sh31df061c, 32'sh31de0a12, 32'sh31dd0e01, 32'sh31dc11e8, 32'sh31db15c7, 32'sh31da199e, 32'sh31d91d6e, 
               32'sh31d82137, 32'sh31d724f7, 32'sh31d628b0, 32'sh31d52c61, 32'sh31d4300b, 32'sh31d333ac, 32'sh31d23746, 32'sh31d13ad9, 
               32'sh31d03e64, 32'sh31cf41e7, 32'sh31ce4562, 32'sh31cd48d6, 32'sh31cc4c42, 32'sh31cb4fa6, 32'sh31ca5303, 32'sh31c95658, 
               32'sh31c859a5, 32'sh31c75ceb, 32'sh31c66029, 32'sh31c5635f, 32'sh31c4668d, 32'sh31c369b4, 32'sh31c26cd4, 32'sh31c16feb, 
               32'sh31c072fb, 32'sh31bf7603, 32'sh31be7904, 32'sh31bd7bfd, 32'sh31bc7eee, 32'sh31bb81d8, 32'sh31ba84b9, 32'sh31b98794, 
               32'sh31b88a66, 32'sh31b78d31, 32'sh31b68ff4, 32'sh31b592b0, 32'sh31b49564, 32'sh31b39810, 32'sh31b29ab4, 32'sh31b19d51, 
               32'sh31b09fe7, 32'sh31afa274, 32'sh31aea4fa, 32'sh31ada778, 32'sh31aca9ef, 32'sh31abac5e, 32'sh31aaaec5, 32'sh31a9b124, 
               32'sh31a8b37c, 32'sh31a7b5cd, 32'sh31a6b815, 32'sh31a5ba56, 32'sh31a4bc90, 32'sh31a3bec1, 32'sh31a2c0eb, 32'sh31a1c30e, 
               32'sh31a0c528, 32'sh319fc73b, 32'sh319ec947, 32'sh319dcb4a, 32'sh319ccd46, 32'sh319bcf3b, 32'sh319ad128, 32'sh3199d30d, 
               32'sh3198d4ea, 32'sh3197d6c0, 32'sh3196d88e, 32'sh3195da55, 32'sh3194dc14, 32'sh3193ddcb, 32'sh3192df7a, 32'sh3191e122, 
               32'sh3190e2c3, 32'sh318fe45b, 32'sh318ee5ec, 32'sh318de776, 32'sh318ce8f7, 32'sh318bea72, 32'sh318aebe4, 32'sh3189ed4f, 
               32'sh3188eeb2, 32'sh3187f00d, 32'sh3186f161, 32'sh3185f2ae, 32'sh3184f3f2, 32'sh3183f52f, 32'sh3182f665, 32'sh3181f792, 
               32'sh3180f8b8, 32'sh317ff9d7, 32'sh317efaee, 32'sh317dfbfd, 32'sh317cfd04, 32'sh317bfe04, 32'sh317afefc, 32'sh3179ffed, 
               32'sh317900d6, 32'sh317801b8, 32'sh31770291, 32'sh31760363, 32'sh3175042e, 32'sh317404f1, 32'sh317305ac, 32'sh31720660, 
               32'sh3171070c, 32'sh317007b0, 32'sh316f084d, 32'sh316e08e2, 32'sh316d096f, 32'sh316c09f5, 32'sh316b0a74, 32'sh316a0aea, 
               32'sh31690b59, 32'sh31680bc1, 32'sh31670c20, 32'sh31660c79, 32'sh31650cc9, 32'sh31640d12, 32'sh31630d53, 32'sh31620d8d, 
               32'sh31610dbf, 32'sh31600dea, 32'sh315f0e0c, 32'sh315e0e28, 32'sh315d0e3b, 32'sh315c0e47, 32'sh315b0e4c, 32'sh315a0e49, 
               32'sh31590e3e, 32'sh31580e2b, 32'sh31570e11, 32'sh31560df0, 32'sh31550dc6, 32'sh31540d95, 32'sh31530d5d, 32'sh31520d1d, 
               32'sh31510cd5, 32'sh31500c86, 32'sh314f0c2f, 32'sh314e0bd1, 32'sh314d0b6a, 32'sh314c0afd, 32'sh314b0a87, 32'sh314a0a0b, 
               32'sh31490986, 32'sh314808fa, 32'sh31470866, 32'sh314607cb, 32'sh31450728, 32'sh3144067d, 32'sh314305cb, 32'sh31420512, 
               32'sh31410450, 32'sh31400387, 32'sh313f02b7, 32'sh313e01df, 32'sh313d00ff, 32'sh313c0018, 32'sh313aff29, 32'sh3139fe33, 
               32'sh3138fd35, 32'sh3137fc2f, 32'sh3136fb22, 32'sh3135fa0d, 32'sh3134f8f1, 32'sh3133f7cd, 32'sh3132f6a1, 32'sh3131f56e, 
               32'sh3130f433, 32'sh312ff2f1, 32'sh312ef1a7, 32'sh312df055, 32'sh312ceefc, 32'sh312bed9b, 32'sh312aec33, 32'sh3129eac3, 
               32'sh3128e94c, 32'sh3127e7cd, 32'sh3126e646, 32'sh3125e4b8, 32'sh3124e322, 32'sh3123e185, 32'sh3122dfe0, 32'sh3121de34, 
               32'sh3120dc80, 32'sh311fdac4, 32'sh311ed901, 32'sh311dd736, 32'sh311cd564, 32'sh311bd38a, 32'sh311ad1a8, 32'sh3119cfbf, 
               32'sh3118cdcf, 32'sh3117cbd6, 32'sh3116c9d7, 32'sh3115c7cf, 32'sh3114c5c0, 32'sh3113c3aa, 32'sh3112c18c, 32'sh3111bf66, 
               32'sh3110bd39, 32'sh310fbb04, 32'sh310eb8c8, 32'sh310db684, 32'sh310cb438, 32'sh310bb1e5, 32'sh310aaf8b, 32'sh3109ad29, 
               32'sh3108aabf, 32'sh3107a84e, 32'sh3106a5d5, 32'sh3105a354, 32'sh3104a0cc, 32'sh31039e3d, 32'sh31029ba6, 32'sh31019907, 
               32'sh31009661, 32'sh30ff93b3, 32'sh30fe90fe, 32'sh30fd8e41, 32'sh30fc8b7d, 32'sh30fb88b1, 32'sh30fa85dd, 32'sh30f98302, 
               32'sh30f8801f, 32'sh30f77d35, 32'sh30f67a44, 32'sh30f5774a, 32'sh30f47449, 32'sh30f37141, 32'sh30f26e31, 32'sh30f16b1a, 
               32'sh30f067fb, 32'sh30ef64d4, 32'sh30ee61a6, 32'sh30ed5e70, 32'sh30ec5b33, 32'sh30eb57ee, 32'sh30ea54a2, 32'sh30e9514e, 
               32'sh30e84df3, 32'sh30e74a90, 32'sh30e64725, 32'sh30e543b3, 32'sh30e4403a, 32'sh30e33cb9, 32'sh30e23930, 32'sh30e135a0, 
               32'sh30e03208, 32'sh30df2e69, 32'sh30de2ac2, 32'sh30dd2714, 32'sh30dc235e, 32'sh30db1fa1, 32'sh30da1bdc, 32'sh30d9180f, 
               32'sh30d8143b, 32'sh30d71060, 32'sh30d60c7d, 32'sh30d50892, 32'sh30d404a0, 32'sh30d300a6, 32'sh30d1fca5, 32'sh30d0f89c, 
               32'sh30cff48c, 32'sh30cef074, 32'sh30cdec55, 32'sh30cce82e, 32'sh30cbe400, 32'sh30cadfca, 32'sh30c9db8d, 32'sh30c8d748, 
               32'sh30c7d2fb, 32'sh30c6cea7, 32'sh30c5ca4c, 32'sh30c4c5e9, 32'sh30c3c17e, 32'sh30c2bd0c, 32'sh30c1b893, 32'sh30c0b412, 
               32'sh30bfaf89, 32'sh30beaaf9, 32'sh30bda661, 32'sh30bca1c2, 32'sh30bb9d1c, 32'sh30ba986d, 32'sh30b993b8, 32'sh30b88efb, 
               32'sh30b78a36, 32'sh30b6856a, 32'sh30b58096, 32'sh30b47bbb, 32'sh30b376d8, 32'sh30b271ee, 32'sh30b16cfc, 32'sh30b06802, 
               32'sh30af6302, 32'sh30ae5df9, 32'sh30ad58ea, 32'sh30ac53d2, 32'sh30ab4eb3, 32'sh30aa498d, 32'sh30a9445f, 32'sh30a83f2a, 
               32'sh30a739ed, 32'sh30a634a9, 32'sh30a52f5d, 32'sh30a42a09, 32'sh30a324af, 32'sh30a21f4c, 32'sh30a119e2, 32'sh30a01471, 
               32'sh309f0ef8, 32'sh309e0978, 32'sh309d03f0, 32'sh309bfe61, 32'sh309af8ca, 32'sh3099f32b, 32'sh3098ed86, 32'sh3097e7d8, 
               32'sh3096e223, 32'sh3095dc67, 32'sh3094d6a3, 32'sh3093d0d8, 32'sh3092cb05, 32'sh3091c52b, 32'sh3090bf49, 32'sh308fb960, 
               32'sh308eb36f, 32'sh308dad77, 32'sh308ca777, 32'sh308ba170, 32'sh308a9b61, 32'sh3089954b, 32'sh30888f2d, 32'sh30878908, 
               32'sh308682dc, 32'sh30857ca7, 32'sh3084766c, 32'sh30837029, 32'sh308269de, 32'sh3081638c, 32'sh30805d33, 32'sh307f56d2, 
               32'sh307e5069, 32'sh307d49f9, 32'sh307c4382, 32'sh307b3d03, 32'sh307a367c, 32'sh30792fee, 32'sh30782959, 32'sh307722bc, 
               32'sh30761c18, 32'sh3075156c, 32'sh30740eb9, 32'sh307307fe, 32'sh3072013c, 32'sh3070fa72, 32'sh306ff3a1, 32'sh306eecc9, 
               32'sh306de5e9, 32'sh306cdf01, 32'sh306bd812, 32'sh306ad11c, 32'sh3069ca1e, 32'sh3068c318, 32'sh3067bc0b, 32'sh3066b4f7, 
               32'sh3065addb, 32'sh3064a6b8, 32'sh30639f8d, 32'sh3062985b, 32'sh30619121, 32'sh306089e0, 32'sh305f8298, 32'sh305e7b48, 
               32'sh305d73f0, 32'sh305c6c91, 32'sh305b652b, 32'sh305a5dbd, 32'sh30595648, 32'sh30584ecb, 32'sh30574747, 32'sh30563fbb, 
               32'sh30553828, 32'sh3054308d, 32'sh305328eb, 32'sh30522142, 32'sh30511991, 32'sh305011d8, 32'sh304f0a19, 32'sh304e0251, 
               32'sh304cfa83, 32'sh304bf2ac, 32'sh304aeacf, 32'sh3049e2ea, 32'sh3048dafd, 32'sh3047d309, 32'sh3046cb0e, 32'sh3045c30b, 
               32'sh3044bb00, 32'sh3043b2ef, 32'sh3042aad5, 32'sh3041a2b5, 32'sh30409a8d, 32'sh303f925d, 32'sh303e8a26, 32'sh303d81e8, 
               32'sh303c79a2, 32'sh303b7155, 32'sh303a6900, 32'sh303960a4, 32'sh30385840, 32'sh30374fd5, 32'sh30364763, 32'sh30353ee9, 
               32'sh30343667, 32'sh30332ddf, 32'sh3032254e, 32'sh30311cb7, 32'sh30301418, 32'sh302f0b71, 32'sh302e02c3, 32'sh302cfa0e, 
               32'sh302bf151, 32'sh302ae88d, 32'sh3029dfc1, 32'sh3028d6ee, 32'sh3027ce14, 32'sh3026c532, 32'sh3025bc48, 32'sh3024b358, 
               32'sh3023aa5f, 32'sh3022a160, 32'sh30219859, 32'sh30208f4a, 32'sh301f8634, 32'sh301e7d17, 32'sh301d73f2, 32'sh301c6ac6, 
               32'sh301b6193, 32'sh301a5858, 32'sh30194f15, 32'sh301845cb, 32'sh30173c7a, 32'sh30163321, 32'sh301529c1, 32'sh3014205a, 
               32'sh301316eb, 32'sh30120d75, 32'sh301103f7, 32'sh300ffa72, 32'sh300ef0e5, 32'sh300de751, 32'sh300cddb6, 32'sh300bd413, 
               32'sh300aca69, 32'sh3009c0b7, 32'sh3008b6fe, 32'sh3007ad3e, 32'sh3006a376, 32'sh300599a7, 32'sh30048fd0, 32'sh300385f2, 
               32'sh30027c0c, 32'sh30017220, 32'sh3000682b, 32'sh2fff5e30, 32'sh2ffe542d, 32'sh2ffd4a22, 32'sh2ffc4010, 32'sh2ffb35f7, 
               32'sh2ffa2bd6, 32'sh2ff921ae, 32'sh2ff8177f, 32'sh2ff70d48, 32'sh2ff6030a, 32'sh2ff4f8c4, 32'sh2ff3ee77, 32'sh2ff2e423, 
               32'sh2ff1d9c7, 32'sh2ff0cf63, 32'sh2fefc4f9, 32'sh2feeba87, 32'sh2fedb00d, 32'sh2feca58d, 32'sh2feb9b04, 32'sh2fea9075, 
               32'sh2fe985de, 32'sh2fe87b3f, 32'sh2fe7709a, 32'sh2fe665ed, 32'sh2fe55b38, 32'sh2fe4507c, 32'sh2fe345b9, 32'sh2fe23aee, 
               32'sh2fe1301c, 32'sh2fe02543, 32'sh2fdf1a62, 32'sh2fde0f7a, 32'sh2fdd048a, 32'sh2fdbf993, 32'sh2fdaee95, 32'sh2fd9e38f, 
               32'sh2fd8d882, 32'sh2fd7cd6d, 32'sh2fd6c252, 32'sh2fd5b72e, 32'sh2fd4ac04, 32'sh2fd3a0d2, 32'sh2fd29598, 32'sh2fd18a58, 
               32'sh2fd07f0f, 32'sh2fcf73c0, 32'sh2fce6869, 32'sh2fcd5d0b, 32'sh2fcc51a5, 32'sh2fcb4638, 32'sh2fca3ac4, 32'sh2fc92f48, 
               32'sh2fc823c5, 32'sh2fc7183b, 32'sh2fc60ca9, 32'sh2fc5010f, 32'sh2fc3f56f, 32'sh2fc2e9c7, 32'sh2fc1de18, 32'sh2fc0d261, 
               32'sh2fbfc6a3, 32'sh2fbebade, 32'sh2fbdaf11, 32'sh2fbca33d, 32'sh2fbb9761, 32'sh2fba8b7e, 32'sh2fb97f94, 32'sh2fb873a3, 
               32'sh2fb767aa, 32'sh2fb65ba9, 32'sh2fb54fa2, 32'sh2fb44393, 32'sh2fb3377c, 32'sh2fb22b5f, 32'sh2fb11f3a, 32'sh2fb0130d, 
               32'sh2faf06da, 32'sh2fadfa9e, 32'sh2facee5c, 32'sh2fabe212, 32'sh2faad5c1, 32'sh2fa9c968, 32'sh2fa8bd09, 32'sh2fa7b0a1, 
               32'sh2fa6a433, 32'sh2fa597bd, 32'sh2fa48b40, 32'sh2fa37ebb, 32'sh2fa2722f, 32'sh2fa1659c, 32'sh2fa05901, 32'sh2f9f4c5f, 
               32'sh2f9e3fb6, 32'sh2f9d3305, 32'sh2f9c264d, 32'sh2f9b198d, 32'sh2f9a0cc7, 32'sh2f98fff9, 32'sh2f97f323, 32'sh2f96e647, 
               32'sh2f95d963, 32'sh2f94cc77, 32'sh2f93bf84, 32'sh2f92b28a, 32'sh2f91a589, 32'sh2f909880, 32'sh2f8f8b70, 32'sh2f8e7e59, 
               32'sh2f8d713a, 32'sh2f8c6414, 32'sh2f8b56e6, 32'sh2f8a49b1, 32'sh2f893c75, 32'sh2f882f32, 32'sh2f8721e7, 32'sh2f861495, 
               32'sh2f85073c, 32'sh2f83f9db, 32'sh2f82ec73, 32'sh2f81df04, 32'sh2f80d18d, 32'sh2f7fc40f, 32'sh2f7eb689, 32'sh2f7da8fd, 
               32'sh2f7c9b69, 32'sh2f7b8dcd, 32'sh2f7a802b, 32'sh2f797281, 32'sh2f7864cf, 32'sh2f775717, 32'sh2f764957, 32'sh2f753b90, 
               32'sh2f742dc1, 32'sh2f731feb, 32'sh2f72120e, 32'sh2f710429, 32'sh2f6ff63d, 32'sh2f6ee84a, 32'sh2f6dda50, 32'sh2f6ccc4e, 
               32'sh2f6bbe45, 32'sh2f6ab034, 32'sh2f69a21d, 32'sh2f6893fe, 32'sh2f6785d7, 32'sh2f6677aa, 32'sh2f656975, 32'sh2f645b38, 
               32'sh2f634cf5, 32'sh2f623eaa, 32'sh2f613058, 32'sh2f6021fe, 32'sh2f5f139d, 32'sh2f5e0535, 32'sh2f5cf6c6, 32'sh2f5be84f, 
               32'sh2f5ad9d1, 32'sh2f59cb4c, 32'sh2f58bcbf, 32'sh2f57ae2b, 32'sh2f569f90, 32'sh2f5590ed, 32'sh2f548243, 32'sh2f537392, 
               32'sh2f5264da, 32'sh2f51561a, 32'sh2f504753, 32'sh2f4f3885, 32'sh2f4e29af, 32'sh2f4d1ad2, 32'sh2f4c0bee, 32'sh2f4afd02, 
               32'sh2f49ee0f, 32'sh2f48df15, 32'sh2f47d014, 32'sh2f46c10b, 32'sh2f45b1fb, 32'sh2f44a2e4, 32'sh2f4393c6, 32'sh2f4284a0, 
               32'sh2f417573, 32'sh2f40663e, 32'sh2f3f5702, 32'sh2f3e47bf, 32'sh2f3d3875, 32'sh2f3c2924, 32'sh2f3b19cb, 32'sh2f3a0a6b, 
               32'sh2f38fb03, 32'sh2f37eb94, 32'sh2f36dc1f, 32'sh2f35cca1, 32'sh2f34bd1d, 32'sh2f33ad91, 32'sh2f329dfe, 32'sh2f318e63, 
               32'sh2f307ec2, 32'sh2f2f6f19, 32'sh2f2e5f69, 32'sh2f2d4fb1, 32'sh2f2c3ff2, 32'sh2f2b302c, 32'sh2f2a205f, 32'sh2f29108a, 
               32'sh2f2800af, 32'sh2f26f0cb, 32'sh2f25e0e1, 32'sh2f24d0ef, 32'sh2f23c0f6, 32'sh2f22b0f6, 32'sh2f21a0ef, 32'sh2f2090e0, 
               32'sh2f1f80ca, 32'sh2f1e70ad, 32'sh2f1d6088, 32'sh2f1c505c, 32'sh2f1b4029, 32'sh2f1a2fef, 32'sh2f191fad, 32'sh2f180f65, 
               32'sh2f16ff14, 32'sh2f15eebd, 32'sh2f14de5e, 32'sh2f13cdf8, 32'sh2f12bd8b, 32'sh2f11ad17, 32'sh2f109c9b, 32'sh2f0f8c18, 
               32'sh2f0e7b8e, 32'sh2f0d6afd, 32'sh2f0c5a64, 32'sh2f0b49c4, 32'sh2f0a391d, 32'sh2f09286e, 32'sh2f0817b8, 32'sh2f0706fb, 
               32'sh2f05f637, 32'sh2f04e56c, 32'sh2f03d499, 32'sh2f02c3bf, 32'sh2f01b2de, 32'sh2f00a1f5, 32'sh2eff9105, 32'sh2efe800e, 
               32'sh2efd6f10, 32'sh2efc5e0b, 32'sh2efb4cfe, 32'sh2efa3bea, 32'sh2ef92acf, 32'sh2ef819ac, 32'sh2ef70883, 32'sh2ef5f752, 
               32'sh2ef4e619, 32'sh2ef3d4da, 32'sh2ef2c393, 32'sh2ef1b245, 32'sh2ef0a0f0, 32'sh2eef8f94, 32'sh2eee7e30, 32'sh2eed6cc5, 
               32'sh2eec5b53, 32'sh2eeb49da, 32'sh2eea3859, 32'sh2ee926d2, 32'sh2ee81543, 32'sh2ee703ac, 32'sh2ee5f20f, 32'sh2ee4e06a, 
               32'sh2ee3cebe, 32'sh2ee2bd0b, 32'sh2ee1ab50, 32'sh2ee0998f, 32'sh2edf87c6, 32'sh2ede75f6, 32'sh2edd641e, 32'sh2edc5240, 
               32'sh2edb405a, 32'sh2eda2e6d, 32'sh2ed91c79, 32'sh2ed80a7d, 32'sh2ed6f87a, 32'sh2ed5e671, 32'sh2ed4d45f, 32'sh2ed3c247, 
               32'sh2ed2b027, 32'sh2ed19e01, 32'sh2ed08bd3, 32'sh2ecf799d, 32'sh2ece6761, 32'sh2ecd551d, 32'sh2ecc42d2, 32'sh2ecb3080, 
               32'sh2eca1e27, 32'sh2ec90bc6, 32'sh2ec7f95e, 32'sh2ec6e6ef, 32'sh2ec5d479, 32'sh2ec4c1fc, 32'sh2ec3af77, 32'sh2ec29ceb, 
               32'sh2ec18a58, 32'sh2ec077be, 32'sh2ebf651d, 32'sh2ebe5274, 32'sh2ebd3fc4, 32'sh2ebc2d0d, 32'sh2ebb1a4f, 32'sh2eba0789, 
               32'sh2eb8f4bc, 32'sh2eb7e1e9, 32'sh2eb6cf0d, 32'sh2eb5bc2b, 32'sh2eb4a942, 32'sh2eb39651, 32'sh2eb28359, 32'sh2eb1705a, 
               32'sh2eb05d53, 32'sh2eaf4a46, 32'sh2eae3731, 32'sh2ead2415, 32'sh2eac10f2, 32'sh2eaafdc8, 32'sh2ea9ea96, 32'sh2ea8d75e, 
               32'sh2ea7c41e, 32'sh2ea6b0d7, 32'sh2ea59d88, 32'sh2ea48a33, 32'sh2ea376d6, 32'sh2ea26372, 32'sh2ea15007, 32'sh2ea03c95, 
               32'sh2e9f291b, 32'sh2e9e159b, 32'sh2e9d0213, 32'sh2e9bee84, 32'sh2e9adaee, 32'sh2e99c750, 32'sh2e98b3ac, 32'sh2e97a000, 
               32'sh2e968c4d, 32'sh2e957893, 32'sh2e9464d1, 32'sh2e935109, 32'sh2e923d39, 32'sh2e912962, 32'sh2e901584, 32'sh2e8f019f, 
               32'sh2e8dedb3, 32'sh2e8cd9bf, 32'sh2e8bc5c4, 32'sh2e8ab1c2, 32'sh2e899db9, 32'sh2e8889a9, 32'sh2e877591, 32'sh2e866173, 
               32'sh2e854d4d, 32'sh2e843920, 32'sh2e8324ec, 32'sh2e8210b0, 32'sh2e80fc6e, 32'sh2e7fe824, 32'sh2e7ed3d3, 32'sh2e7dbf7b, 
               32'sh2e7cab1c, 32'sh2e7b96b6, 32'sh2e7a8248, 32'sh2e796dd3, 32'sh2e785958, 32'sh2e7744d5, 32'sh2e76304a, 32'sh2e751bb9, 
               32'sh2e740720, 32'sh2e72f281, 32'sh2e71ddda, 32'sh2e70c92c, 32'sh2e6fb477, 32'sh2e6e9fba, 32'sh2e6d8af7, 32'sh2e6c762c, 
               32'sh2e6b615a, 32'sh2e6a4c81, 32'sh2e6937a1, 32'sh2e6822ba, 32'sh2e670dcb, 32'sh2e65f8d6, 32'sh2e64e3d9, 32'sh2e63ced5, 
               32'sh2e62b9ca, 32'sh2e61a4b8, 32'sh2e608f9e, 32'sh2e5f7a7e, 32'sh2e5e6556, 32'sh2e5d5027, 32'sh2e5c3af1, 32'sh2e5b25b4, 
               32'sh2e5a1070, 32'sh2e58fb24, 32'sh2e57e5d2, 32'sh2e56d078, 32'sh2e55bb17, 32'sh2e54a5af, 32'sh2e539040, 32'sh2e527aca, 
               32'sh2e51654c, 32'sh2e504fc8, 32'sh2e4f3a3c, 32'sh2e4e24a9, 32'sh2e4d0f0f, 32'sh2e4bf96e, 32'sh2e4ae3c6, 32'sh2e49ce16, 
               32'sh2e48b860, 32'sh2e47a2a2, 32'sh2e468cdd, 32'sh2e457711, 32'sh2e44613e, 32'sh2e434b64, 32'sh2e423582, 32'sh2e411f9a, 
               32'sh2e4009aa, 32'sh2e3ef3b3, 32'sh2e3dddb5, 32'sh2e3cc7b0, 32'sh2e3bb1a4, 32'sh2e3a9b91, 32'sh2e398576, 32'sh2e386f55, 
               32'sh2e37592c, 32'sh2e3642fc, 32'sh2e352cc5, 32'sh2e341687, 32'sh2e330042, 32'sh2e31e9f6, 32'sh2e30d3a2, 32'sh2e2fbd48, 
               32'sh2e2ea6e6, 32'sh2e2d907d, 32'sh2e2c7a0d, 32'sh2e2b6396, 32'sh2e2a4d18, 32'sh2e293693, 32'sh2e282006, 32'sh2e270973, 
               32'sh2e25f2d8, 32'sh2e24dc36, 32'sh2e23c58d, 32'sh2e22aedd, 32'sh2e219826, 32'sh2e208168, 32'sh2e1f6aa3, 32'sh2e1e53d6, 
               32'sh2e1d3d03, 32'sh2e1c2628, 32'sh2e1b0f46, 32'sh2e19f85d, 32'sh2e18e16d, 32'sh2e17ca76, 32'sh2e16b378, 32'sh2e159c73, 
               32'sh2e148566, 32'sh2e136e53, 32'sh2e125738, 32'sh2e114016, 32'sh2e1028ed, 32'sh2e0f11bd, 32'sh2e0dfa86, 32'sh2e0ce348, 
               32'sh2e0bcc03, 32'sh2e0ab4b7, 32'sh2e099d63, 32'sh2e088608, 32'sh2e076ea7, 32'sh2e06573e, 32'sh2e053fce, 32'sh2e042857, 
               32'sh2e0310d9, 32'sh2e01f954, 32'sh2e00e1c8, 32'sh2dffca34, 32'sh2dfeb29a, 32'sh2dfd9af8, 32'sh2dfc8350, 32'sh2dfb6ba0, 
               32'sh2dfa53e9, 32'sh2df93c2b, 32'sh2df82466, 32'sh2df70c9a, 32'sh2df5f4c7, 32'sh2df4dced, 32'sh2df3c50c, 32'sh2df2ad23, 
               32'sh2df19534, 32'sh2df07d3d, 32'sh2def653f, 32'sh2dee4d3b, 32'sh2ded352f, 32'sh2dec1d1c, 32'sh2deb0502, 32'sh2de9ece1, 
               32'sh2de8d4b8, 32'sh2de7bc89, 32'sh2de6a453, 32'sh2de58c15, 32'sh2de473d1, 32'sh2de35b85, 32'sh2de24333, 32'sh2de12ad9, 
               32'sh2de01278, 32'sh2ddefa10, 32'sh2ddde1a1, 32'sh2ddcc92b, 32'sh2ddbb0ae, 32'sh2dda982a, 32'sh2dd97f9f, 32'sh2dd8670d, 
               32'sh2dd74e73, 32'sh2dd635d3, 32'sh2dd51d2b, 32'sh2dd4047d, 32'sh2dd2ebc7, 32'sh2dd1d30a, 32'sh2dd0ba47, 32'sh2dcfa17c, 
               32'sh2dce88aa, 32'sh2dcd6fd1, 32'sh2dcc56f1, 32'sh2dcb3e0a, 32'sh2dca251c, 32'sh2dc90c26, 32'sh2dc7f32a, 32'sh2dc6da27, 
               32'sh2dc5c11c, 32'sh2dc4a80b, 32'sh2dc38ef2, 32'sh2dc275d3, 32'sh2dc15cac, 32'sh2dc0437e, 32'sh2dbf2a4a, 32'sh2dbe110e, 
               32'sh2dbcf7cb, 32'sh2dbbde81, 32'sh2dbac530, 32'sh2db9abd8, 32'sh2db89279, 32'sh2db77913, 32'sh2db65fa6, 32'sh2db54632, 
               32'sh2db42cb6, 32'sh2db31334, 32'sh2db1f9ab, 32'sh2db0e01a, 32'sh2dafc683, 32'sh2daeace4, 32'sh2dad933f, 32'sh2dac7992, 
               32'sh2dab5fdf, 32'sh2daa4624, 32'sh2da92c62, 32'sh2da81299, 32'sh2da6f8ca, 32'sh2da5def3, 32'sh2da4c515, 32'sh2da3ab30, 
               32'sh2da29144, 32'sh2da17751, 32'sh2da05d57, 32'sh2d9f4356, 32'sh2d9e294e, 32'sh2d9d0f3f, 32'sh2d9bf529, 32'sh2d9adb0b, 
               32'sh2d99c0e7, 32'sh2d98a6bc, 32'sh2d978c8a, 32'sh2d967250, 32'sh2d955810, 32'sh2d943dc9, 32'sh2d93237a, 32'sh2d920925, 
               32'sh2d90eec8, 32'sh2d8fd465, 32'sh2d8eb9fa, 32'sh2d8d9f89, 32'sh2d8c8510, 32'sh2d8b6a90, 32'sh2d8a500a, 32'sh2d89357c, 
               32'sh2d881ae8, 32'sh2d87004c, 32'sh2d85e5a9, 32'sh2d84caff, 32'sh2d83b04f, 32'sh2d829597, 32'sh2d817ad8, 32'sh2d806012, 
               32'sh2d7f4545, 32'sh2d7e2a72, 32'sh2d7d0f97, 32'sh2d7bf4b5, 32'sh2d7ad9cc, 32'sh2d79bedc, 32'sh2d78a3e5, 32'sh2d7788e7, 
               32'sh2d766de2, 32'sh2d7552d6, 32'sh2d7437c3, 32'sh2d731ca9, 32'sh2d720189, 32'sh2d70e661, 32'sh2d6fcb32, 32'sh2d6eaffc, 
               32'sh2d6d94bf, 32'sh2d6c797b, 32'sh2d6b5e30, 32'sh2d6a42dd, 32'sh2d692784, 32'sh2d680c24, 32'sh2d66f0bd, 32'sh2d65d54f, 
               32'sh2d64b9da, 32'sh2d639e5e, 32'sh2d6282db, 32'sh2d616751, 32'sh2d604bc0, 32'sh2d5f3028, 32'sh2d5e1489, 32'sh2d5cf8e3, 
               32'sh2d5bdd36, 32'sh2d5ac182, 32'sh2d59a5c7, 32'sh2d588a05, 32'sh2d576e3c, 32'sh2d56526c, 32'sh2d553695, 32'sh2d541ab7, 
               32'sh2d52fed2, 32'sh2d51e2e6, 32'sh2d50c6f3, 32'sh2d4faafa, 32'sh2d4e8ef9, 32'sh2d4d72f1, 32'sh2d4c56e2, 32'sh2d4b3acc, 
               32'sh2d4a1eaf, 32'sh2d49028b, 32'sh2d47e661, 32'sh2d46ca2f, 32'sh2d45adf6, 32'sh2d4491b6, 32'sh2d43756f, 32'sh2d425922, 
               32'sh2d413ccd, 32'sh2d402071, 32'sh2d3f040f, 32'sh2d3de7a5, 32'sh2d3ccb34, 32'sh2d3baebd, 32'sh2d3a923e, 32'sh2d3975b9, 
               32'sh2d38592c, 32'sh2d373c99, 32'sh2d361ffe, 32'sh2d35035d, 32'sh2d33e6b4, 32'sh2d32ca05, 32'sh2d31ad4f, 32'sh2d309091, 
               32'sh2d2f73cd, 32'sh2d2e5702, 32'sh2d2d3a30, 32'sh2d2c1d56, 32'sh2d2b0076, 32'sh2d29e38f, 32'sh2d28c6a1, 32'sh2d27a9ac, 
               32'sh2d268cb0, 32'sh2d256fad, 32'sh2d2452a3, 32'sh2d233592, 32'sh2d22187a, 32'sh2d20fb5b, 32'sh2d1fde36, 32'sh2d1ec109, 
               32'sh2d1da3d5, 32'sh2d1c869b, 32'sh2d1b6959, 32'sh2d1a4c10, 32'sh2d192ec1, 32'sh2d18116a, 32'sh2d16f40d, 32'sh2d15d6a9, 
               32'sh2d14b93d, 32'sh2d139bcb, 32'sh2d127e52, 32'sh2d1160d2, 32'sh2d10434a, 32'sh2d0f25bc, 32'sh2d0e0827, 32'sh2d0cea8b, 
               32'sh2d0bcce8, 32'sh2d0aaf3e, 32'sh2d09918e, 32'sh2d0873d6, 32'sh2d075617, 32'sh2d063852, 32'sh2d051a85, 32'sh2d03fcb1, 
               32'sh2d02ded7, 32'sh2d01c0f5, 32'sh2d00a30d, 32'sh2cff851e, 32'sh2cfe6728, 32'sh2cfd492a, 32'sh2cfc2b26, 32'sh2cfb0d1b, 
               32'sh2cf9ef09, 32'sh2cf8d0f0, 32'sh2cf7b2d0, 32'sh2cf694aa, 32'sh2cf5767c, 32'sh2cf45847, 32'sh2cf33a0c, 32'sh2cf21bc9, 
               32'sh2cf0fd80, 32'sh2cefdf2f, 32'sh2ceec0d8, 32'sh2ceda27a, 32'sh2cec8414, 32'sh2ceb65a8, 32'sh2cea4735, 32'sh2ce928bb, 
               32'sh2ce80a3a, 32'sh2ce6ebb2, 32'sh2ce5cd24, 32'sh2ce4ae8e, 32'sh2ce38ff1, 32'sh2ce2714e, 32'sh2ce152a4, 32'sh2ce033f2, 
               32'sh2cdf153a, 32'sh2cddf67b, 32'sh2cdcd7b5, 32'sh2cdbb8e8, 32'sh2cda9a14, 32'sh2cd97b39, 32'sh2cd85c57, 32'sh2cd73d6e, 
               32'sh2cd61e7f, 32'sh2cd4ff88, 32'sh2cd3e08b, 32'sh2cd2c186, 32'sh2cd1a27b, 32'sh2cd08369, 32'sh2ccf6450, 32'sh2cce4530, 
               32'sh2ccd2609, 32'sh2ccc06db, 32'sh2ccae7a6, 32'sh2cc9c86b, 32'sh2cc8a928, 32'sh2cc789df, 32'sh2cc66a8e, 32'sh2cc54b37, 
               32'sh2cc42bd9, 32'sh2cc30c74, 32'sh2cc1ed08, 32'sh2cc0cd95, 32'sh2cbfae1b, 32'sh2cbe8e9b, 32'sh2cbd6f13, 32'sh2cbc4f85, 
               32'sh2cbb2fef, 32'sh2cba1053, 32'sh2cb8f0b0, 32'sh2cb7d106, 32'sh2cb6b155, 32'sh2cb5919d, 32'sh2cb471de, 32'sh2cb35218, 
               32'sh2cb2324c, 32'sh2cb11278, 32'sh2caff29e, 32'sh2caed2bd, 32'sh2cadb2d5, 32'sh2cac92e6, 32'sh2cab72f0, 32'sh2caa52f3, 
               32'sh2ca932ef, 32'sh2ca812e5, 32'sh2ca6f2d4, 32'sh2ca5d2bb, 32'sh2ca4b29c, 32'sh2ca39276, 32'sh2ca27249, 32'sh2ca15215, 
               32'sh2ca031da, 32'sh2c9f1199, 32'sh2c9df150, 32'sh2c9cd101, 32'sh2c9bb0ab, 32'sh2c9a904d, 32'sh2c996fe9, 32'sh2c984f7e, 
               32'sh2c972f0d, 32'sh2c960e94, 32'sh2c94ee15, 32'sh2c93cd8e, 32'sh2c92ad01, 32'sh2c918c6d, 32'sh2c906bd2, 32'sh2c8f4b30, 
               32'sh2c8e2a87, 32'sh2c8d09d7, 32'sh2c8be921, 32'sh2c8ac863, 32'sh2c89a79f, 32'sh2c8886d4, 32'sh2c876602, 32'sh2c864529, 
               32'sh2c85244a, 32'sh2c840363, 32'sh2c82e276, 32'sh2c81c181, 32'sh2c80a086, 32'sh2c7f7f84, 32'sh2c7e5e7b, 32'sh2c7d3d6b, 
               32'sh2c7c1c55, 32'sh2c7afb37, 32'sh2c79da13, 32'sh2c78b8e8, 32'sh2c7797b6, 32'sh2c76767d, 32'sh2c75553d, 32'sh2c7433f6, 
               32'sh2c7312a9, 32'sh2c71f154, 32'sh2c70cff9, 32'sh2c6fae97, 32'sh2c6e8d2e, 32'sh2c6d6bbf, 32'sh2c6c4a48, 32'sh2c6b28cb, 
               32'sh2c6a0746, 32'sh2c68e5bb, 32'sh2c67c429, 32'sh2c66a290, 32'sh2c6580f1, 32'sh2c645f4a, 32'sh2c633d9d, 32'sh2c621be8, 
               32'sh2c60fa2d, 32'sh2c5fd86b, 32'sh2c5eb6a3, 32'sh2c5d94d3, 32'sh2c5c72fd, 32'sh2c5b511f, 32'sh2c5a2f3b, 32'sh2c590d50, 
               32'sh2c57eb5e, 32'sh2c56c966, 32'sh2c55a766, 32'sh2c548560, 32'sh2c536353, 32'sh2c52413f, 32'sh2c511f24, 32'sh2c4ffd02, 
               32'sh2c4edada, 32'sh2c4db8aa, 32'sh2c4c9674, 32'sh2c4b7437, 32'sh2c4a51f3, 32'sh2c492fa9, 32'sh2c480d57, 32'sh2c46eaff, 
               32'sh2c45c8a0, 32'sh2c44a63a, 32'sh2c4383cd, 32'sh2c426159, 32'sh2c413edf, 32'sh2c401c5e, 32'sh2c3ef9d6, 32'sh2c3dd747, 
               32'sh2c3cb4b1, 32'sh2c3b9214, 32'sh2c3a6f71, 32'sh2c394cc7, 32'sh2c382a16, 32'sh2c37075e, 32'sh2c35e49f, 32'sh2c34c1da, 
               32'sh2c339f0e, 32'sh2c327c3a, 32'sh2c315961, 32'sh2c303680, 32'sh2c2f1398, 32'sh2c2df0aa, 32'sh2c2ccdb5, 32'sh2c2baab9, 
               32'sh2c2a87b6, 32'sh2c2964ac, 32'sh2c28419c, 32'sh2c271e85, 32'sh2c25fb66, 32'sh2c24d842, 32'sh2c23b516, 32'sh2c2291e4, 
               32'sh2c216eaa, 32'sh2c204b6a, 32'sh2c1f2823, 32'sh2c1e04d6, 32'sh2c1ce181, 32'sh2c1bbe26, 32'sh2c1a9ac4, 32'sh2c19775b, 
               32'sh2c1853eb, 32'sh2c173075, 32'sh2c160cf7, 32'sh2c14e973, 32'sh2c13c5e8, 32'sh2c12a257, 32'sh2c117ebe, 32'sh2c105b1f, 
               32'sh2c0f3779, 32'sh2c0e13cc, 32'sh2c0cf018, 32'sh2c0bcc5e, 32'sh2c0aa89c, 32'sh2c0984d4, 32'sh2c086106, 32'sh2c073d30, 
               32'sh2c061953, 32'sh2c04f570, 32'sh2c03d186, 32'sh2c02ad96, 32'sh2c01899e, 32'sh2c0065a0, 32'sh2bff419a, 32'sh2bfe1d8f, 
               32'sh2bfcf97c, 32'sh2bfbd562, 32'sh2bfab142, 32'sh2bf98d1b, 32'sh2bf868ed, 32'sh2bf744b8, 32'sh2bf6207d, 32'sh2bf4fc3b, 
               32'sh2bf3d7f2, 32'sh2bf2b3a2, 32'sh2bf18f4c, 32'sh2bf06aee, 32'sh2bef468a, 32'sh2bee221f, 32'sh2becfdae, 32'sh2bebd935, 
               32'sh2beab4b6, 32'sh2be99030, 32'sh2be86ba4, 32'sh2be74710, 32'sh2be62276, 32'sh2be4fdd5, 32'sh2be3d92d, 32'sh2be2b47f, 
               32'sh2be18fc9, 32'sh2be06b0d, 32'sh2bdf464a, 32'sh2bde2181, 32'sh2bdcfcb0, 32'sh2bdbd7d9, 32'sh2bdab2fb, 32'sh2bd98e16, 
               32'sh2bd8692b, 32'sh2bd74439, 32'sh2bd61f40, 32'sh2bd4fa40, 32'sh2bd3d53a, 32'sh2bd2b02c, 32'sh2bd18b18, 32'sh2bd065fe, 
               32'sh2bcf40dc, 32'sh2bce1bb4, 32'sh2bccf685, 32'sh2bcbd14f, 32'sh2bcaac12, 32'sh2bc986cf, 32'sh2bc86185, 32'sh2bc73c34, 
               32'sh2bc616dd, 32'sh2bc4f17f, 32'sh2bc3cc19, 32'sh2bc2a6ae, 32'sh2bc1813b, 32'sh2bc05bc2, 32'sh2bbf3642, 32'sh2bbe10bb, 
               32'sh2bbceb2d, 32'sh2bbbc599, 32'sh2bba9ffe, 32'sh2bb97a5c, 32'sh2bb854b4, 32'sh2bb72f05, 32'sh2bb6094f, 32'sh2bb4e392, 
               32'sh2bb3bdce, 32'sh2bb29804, 32'sh2bb17233, 32'sh2bb04c5c, 32'sh2baf267d, 32'sh2bae0098, 32'sh2bacdaac, 32'sh2babb4ba, 
               32'sh2baa8ec0, 32'sh2ba968c0, 32'sh2ba842b9, 32'sh2ba71cac, 32'sh2ba5f697, 32'sh2ba4d07c, 32'sh2ba3aa5b, 32'sh2ba28432, 
               32'sh2ba15e03, 32'sh2ba037cd, 32'sh2b9f1190, 32'sh2b9deb4d, 32'sh2b9cc503, 32'sh2b9b9eb2, 32'sh2b9a785a, 32'sh2b9951fc, 
               32'sh2b982b97, 32'sh2b97052b, 32'sh2b95deb9, 32'sh2b94b840, 32'sh2b9391c0, 32'sh2b926b39, 32'sh2b9144ac, 32'sh2b901e18, 
               32'sh2b8ef77d, 32'sh2b8dd0db, 32'sh2b8caa33, 32'sh2b8b8384, 32'sh2b8a5cce, 32'sh2b893612, 32'sh2b880f4f, 32'sh2b86e885, 
               32'sh2b85c1b5, 32'sh2b849add, 32'sh2b837400, 32'sh2b824d1b, 32'sh2b812630, 32'sh2b7fff3e, 32'sh2b7ed845, 32'sh2b7db145, 
               32'sh2b7c8a3f, 32'sh2b7b6332, 32'sh2b7a3c1f, 32'sh2b791504, 32'sh2b77ede3, 32'sh2b76c6bc, 32'sh2b759f8d, 32'sh2b747858, 
               32'sh2b73511c, 32'sh2b7229da, 32'sh2b710291, 32'sh2b6fdb41, 32'sh2b6eb3ea, 32'sh2b6d8c8d, 32'sh2b6c6529, 32'sh2b6b3dbe, 
               32'sh2b6a164d, 32'sh2b68eed5, 32'sh2b67c756, 32'sh2b669fd0, 32'sh2b657844, 32'sh2b6450b1, 32'sh2b632918, 32'sh2b620177, 
               32'sh2b60d9d0, 32'sh2b5fb223, 32'sh2b5e8a6f, 32'sh2b5d62b4, 32'sh2b5c3af2, 32'sh2b5b1329, 32'sh2b59eb5a, 32'sh2b58c385, 
               32'sh2b579ba8, 32'sh2b5673c5, 32'sh2b554bdb, 32'sh2b5423eb, 32'sh2b52fbf4, 32'sh2b51d3f6, 32'sh2b50abf1, 32'sh2b4f83e6, 
               32'sh2b4e5bd4, 32'sh2b4d33bc, 32'sh2b4c0b9c, 32'sh2b4ae376, 32'sh2b49bb4a, 32'sh2b489317, 32'sh2b476add, 32'sh2b46429c, 
               32'sh2b451a55, 32'sh2b43f207, 32'sh2b42c9b2, 32'sh2b41a157, 32'sh2b4078f5, 32'sh2b3f508c, 32'sh2b3e281d, 32'sh2b3cffa7, 
               32'sh2b3bd72a, 32'sh2b3aaea7, 32'sh2b39861d, 32'sh2b385d8c, 32'sh2b3734f5, 32'sh2b360c57, 32'sh2b34e3b2, 32'sh2b33bb07, 
               32'sh2b329255, 32'sh2b31699c, 32'sh2b3040dd, 32'sh2b2f1817, 32'sh2b2def4b, 32'sh2b2cc677, 32'sh2b2b9d9d, 32'sh2b2a74bd, 
               32'sh2b294bd5, 32'sh2b2822e8, 32'sh2b26f9f3, 32'sh2b25d0f8, 32'sh2b24a7f6, 32'sh2b237eed, 32'sh2b2255de, 32'sh2b212cc8, 
               32'sh2b2003ac, 32'sh2b1eda89, 32'sh2b1db15f, 32'sh2b1c882f, 32'sh2b1b5ef8, 32'sh2b1a35ba, 32'sh2b190c75, 32'sh2b17e32a, 
               32'sh2b16b9d9, 32'sh2b159080, 32'sh2b146722, 32'sh2b133dbc, 32'sh2b121450, 32'sh2b10eadd, 32'sh2b0fc163, 32'sh2b0e97e3, 
               32'sh2b0d6e5c, 32'sh2b0c44cf, 32'sh2b0b1b3b, 32'sh2b09f1a0, 32'sh2b08c7ff, 32'sh2b079e57, 32'sh2b0674a8, 32'sh2b054af3, 
               32'sh2b042137, 32'sh2b02f774, 32'sh2b01cdab, 32'sh2b00a3dc, 32'sh2aff7a05, 32'sh2afe5028, 32'sh2afd2644, 32'sh2afbfc5a, 
               32'sh2afad269, 32'sh2af9a872, 32'sh2af87e73, 32'sh2af7546f, 32'sh2af62a63, 32'sh2af50051, 32'sh2af3d638, 32'sh2af2ac19, 
               32'sh2af181f3, 32'sh2af057c6, 32'sh2aef2d93, 32'sh2aee0359, 32'sh2aecd919, 32'sh2aebaed2, 32'sh2aea8484, 32'sh2ae95a30, 
               32'sh2ae82fd5, 32'sh2ae70574, 32'sh2ae5db0b, 32'sh2ae4b09d, 32'sh2ae38627, 32'sh2ae25bab, 32'sh2ae13129, 32'sh2ae006a0, 
               32'sh2adedc10, 32'sh2addb179, 32'sh2adc86dc, 32'sh2adb5c39, 32'sh2ada318e, 32'sh2ad906dd, 32'sh2ad7dc26, 32'sh2ad6b168, 
               32'sh2ad586a3, 32'sh2ad45bd8, 32'sh2ad33106, 32'sh2ad2062d, 32'sh2ad0db4e, 32'sh2acfb069, 32'sh2ace857c, 32'sh2acd5a89, 
               32'sh2acc2f90, 32'sh2acb0490, 32'sh2ac9d989, 32'sh2ac8ae7c, 32'sh2ac78368, 32'sh2ac6584d, 32'sh2ac52d2c, 32'sh2ac40205, 
               32'sh2ac2d6d6, 32'sh2ac1aba1, 32'sh2ac08066, 32'sh2abf5524, 32'sh2abe29db, 32'sh2abcfe8c, 32'sh2abbd336, 32'sh2abaa7da, 
               32'sh2ab97c77, 32'sh2ab8510d, 32'sh2ab7259d, 32'sh2ab5fa26, 32'sh2ab4cea9, 32'sh2ab3a325, 32'sh2ab2779a, 32'sh2ab14c09, 
               32'sh2ab02071, 32'sh2aaef4d3, 32'sh2aadc92e, 32'sh2aac9d83, 32'sh2aab71d0, 32'sh2aaa4618, 32'sh2aa91a59, 32'sh2aa7ee93, 
               32'sh2aa6c2c6, 32'sh2aa596f4, 32'sh2aa46b1a, 32'sh2aa33f3a, 32'sh2aa21353, 32'sh2aa0e766, 32'sh2a9fbb72, 32'sh2a9e8f78, 
               32'sh2a9d6377, 32'sh2a9c376f, 32'sh2a9b0b61, 32'sh2a99df4d, 32'sh2a98b331, 32'sh2a97870f, 32'sh2a965ae7, 32'sh2a952eb8, 
               32'sh2a940283, 32'sh2a92d647, 32'sh2a91aa04, 32'sh2a907dbb, 32'sh2a8f516b, 32'sh2a8e2515, 32'sh2a8cf8b8, 32'sh2a8bcc54, 
               32'sh2a8a9fea, 32'sh2a89737a, 32'sh2a884702, 32'sh2a871a85, 32'sh2a85ee00, 32'sh2a84c176, 32'sh2a8394e4, 32'sh2a82684c, 
               32'sh2a813bae, 32'sh2a800f09, 32'sh2a7ee25d, 32'sh2a7db5ab, 32'sh2a7c88f2, 32'sh2a7b5c33, 32'sh2a7a2f6d, 32'sh2a7902a1, 
               32'sh2a77d5ce, 32'sh2a76a8f5, 32'sh2a757c15, 32'sh2a744f2e, 32'sh2a732241, 32'sh2a71f54d, 32'sh2a70c853, 32'sh2a6f9b52, 
               32'sh2a6e6e4b, 32'sh2a6d413d, 32'sh2a6c1429, 32'sh2a6ae70e, 32'sh2a69b9ec, 32'sh2a688cc4, 32'sh2a675f96, 32'sh2a663261, 
               32'sh2a650525, 32'sh2a63d7e3, 32'sh2a62aa9a, 32'sh2a617d4b, 32'sh2a604ff5, 32'sh2a5f2299, 32'sh2a5df536, 32'sh2a5cc7cd, 
               32'sh2a5b9a5d, 32'sh2a5a6ce7, 32'sh2a593f6a, 32'sh2a5811e6, 32'sh2a56e45c, 32'sh2a55b6cc, 32'sh2a548935, 32'sh2a535b97, 
               32'sh2a522df3, 32'sh2a510048, 32'sh2a4fd297, 32'sh2a4ea4df, 32'sh2a4d7721, 32'sh2a4c495c, 32'sh2a4b1b91, 32'sh2a49edbf, 
               32'sh2a48bfe7, 32'sh2a479208, 32'sh2a466423, 32'sh2a453637, 32'sh2a440844, 32'sh2a42da4c, 32'sh2a41ac4c, 32'sh2a407e46, 
               32'sh2a3f503a, 32'sh2a3e2227, 32'sh2a3cf40d, 32'sh2a3bc5ed, 32'sh2a3a97c7, 32'sh2a39699a, 32'sh2a383b66, 32'sh2a370d2c, 
               32'sh2a35deeb, 32'sh2a34b0a4, 32'sh2a338257, 32'sh2a325403, 32'sh2a3125a8, 32'sh2a2ff747, 32'sh2a2ec8df, 32'sh2a2d9a71, 
               32'sh2a2c6bfd, 32'sh2a2b3d82, 32'sh2a2a0f00, 32'sh2a28e078, 32'sh2a27b1e9, 32'sh2a268354, 32'sh2a2554b8, 32'sh2a242616, 
               32'sh2a22f76e, 32'sh2a21c8be, 32'sh2a209a09, 32'sh2a1f6b4d, 32'sh2a1e3c8a, 32'sh2a1d0dc1, 32'sh2a1bdef1, 32'sh2a1ab01b, 
               32'sh2a19813f, 32'sh2a18525c, 32'sh2a172372, 32'sh2a15f482, 32'sh2a14c58b, 32'sh2a13968e, 32'sh2a12678b, 32'sh2a113881, 
               32'sh2a100970, 32'sh2a0eda59, 32'sh2a0dab3c, 32'sh2a0c7c18, 32'sh2a0b4ced, 32'sh2a0a1dbc, 32'sh2a08ee85, 32'sh2a07bf47, 
               32'sh2a069003, 32'sh2a0560b8, 32'sh2a043166, 32'sh2a03020f, 32'sh2a01d2b0, 32'sh2a00a34c, 32'sh29ff73e0, 32'sh29fe446f, 
               32'sh29fd14f6, 32'sh29fbe578, 32'sh29fab5f3, 32'sh29f98667, 32'sh29f856d5, 32'sh29f7273c, 32'sh29f5f79d, 32'sh29f4c7f8, 
               32'sh29f3984c, 32'sh29f26899, 32'sh29f138e0, 32'sh29f00921, 32'sh29eed95b, 32'sh29eda98f, 32'sh29ec79bc, 32'sh29eb49e3, 
               32'sh29ea1a03, 32'sh29e8ea1d, 32'sh29e7ba30, 32'sh29e68a3d, 32'sh29e55a43, 32'sh29e42a43, 32'sh29e2fa3d, 32'sh29e1ca30, 
               32'sh29e09a1c, 32'sh29df6a02, 32'sh29de39e2, 32'sh29dd09bb, 32'sh29dbd98e, 32'sh29daa95a, 32'sh29d97920, 32'sh29d848e0, 
               32'sh29d71899, 32'sh29d5e84b, 32'sh29d4b7f7, 32'sh29d3879d, 32'sh29d2573c, 32'sh29d126d4, 32'sh29cff667, 32'sh29cec5f2, 
               32'sh29cd9578, 32'sh29cc64f7, 32'sh29cb346f, 32'sh29ca03e1, 32'sh29c8d34d, 32'sh29c7a2b2, 32'sh29c67210, 32'sh29c54169, 
               32'sh29c410ba, 32'sh29c2e006, 32'sh29c1af4b, 32'sh29c07e89, 32'sh29bf4dc1, 32'sh29be1cf3, 32'sh29bcec1e, 32'sh29bbbb43, 
               32'sh29ba8a61, 32'sh29b95979, 32'sh29b8288a, 32'sh29b6f795, 32'sh29b5c69a, 32'sh29b49598, 32'sh29b3648f, 32'sh29b23381, 
               32'sh29b1026c, 32'sh29afd150, 32'sh29aea02e, 32'sh29ad6f05, 32'sh29ac3dd7, 32'sh29ab0ca1, 32'sh29a9db65, 32'sh29a8aa23, 
               32'sh29a778db, 32'sh29a6478c, 32'sh29a51636, 32'sh29a3e4da, 32'sh29a2b378, 32'sh29a1820f, 32'sh29a050a0, 32'sh299f1f2b, 
               32'sh299dedaf, 32'sh299cbc2c, 32'sh299b8aa4, 32'sh299a5914, 32'sh2999277f, 32'sh2997f5e3, 32'sh2996c440, 32'sh29959297, 
               32'sh299460e8, 32'sh29932f32, 32'sh2991fd76, 32'sh2990cbb4, 32'sh298f99eb, 32'sh298e681b, 32'sh298d3646, 32'sh298c0469, 
               32'sh298ad287, 32'sh2989a09e, 32'sh29886eaf, 32'sh29873cb9, 32'sh29860abd, 32'sh2984d8ba, 32'sh2983a6b1, 32'sh298274a2, 
               32'sh2981428c, 32'sh29801070, 32'sh297ede4d, 32'sh297dac24, 32'sh297c79f5, 32'sh297b47bf, 32'sh297a1583, 32'sh2978e340, 
               32'sh2977b0f7, 32'sh29767ea8, 32'sh29754c52, 32'sh297419f6, 32'sh2972e793, 32'sh2971b52a, 32'sh297082bb, 32'sh296f5045, 
               32'sh296e1dc9, 32'sh296ceb47, 32'sh296bb8be, 32'sh296a862e, 32'sh29695399, 32'sh296820fd, 32'sh2966ee5a, 32'sh2965bbb1, 
               32'sh29648902, 32'sh2963564d, 32'sh29622391, 32'sh2960f0ce, 32'sh295fbe06, 32'sh295e8b36, 32'sh295d5861, 32'sh295c2585, 
               32'sh295af2a3, 32'sh2959bfba, 32'sh29588ccb, 32'sh295759d6, 32'sh295626da, 32'sh2954f3d8, 32'sh2953c0cf, 32'sh29528dc0, 
               32'sh29515aab, 32'sh29502790, 32'sh294ef46e, 32'sh294dc145, 32'sh294c8e16, 32'sh294b5ae1, 32'sh294a27a6, 32'sh2948f464, 
               32'sh2947c11c, 32'sh29468dcd, 32'sh29455a78, 32'sh2944271d, 32'sh2942f3bb, 32'sh2941c053, 32'sh29408ce5, 32'sh293f5970, 
               32'sh293e25f5, 32'sh293cf274, 32'sh293bbeec, 32'sh293a8b5e, 32'sh293957c9, 32'sh2938242e, 32'sh2936f08d, 32'sh2935bce5, 
               32'sh29348937, 32'sh29335583, 32'sh293221c8, 32'sh2930ee07, 32'sh292fba40, 32'sh292e8672, 32'sh292d529e, 32'sh292c1ec3, 
               32'sh292aeae3, 32'sh2929b6fc, 32'sh2928830e, 32'sh29274f1a, 32'sh29261b20, 32'sh2924e720, 32'sh2923b319, 32'sh29227f0b, 
               32'sh29214af8, 32'sh292016de, 32'sh291ee2be, 32'sh291dae97, 32'sh291c7a6a, 32'sh291b4637, 32'sh291a11fd, 32'sh2918ddbd, 
               32'sh2917a977, 32'sh2916752a, 32'sh291540d8, 32'sh29140c7e, 32'sh2912d81f, 32'sh2911a3b9, 32'sh29106f4c, 32'sh290f3ada, 
               32'sh290e0661, 32'sh290cd1e1, 32'sh290b9d5c, 32'sh290a68d0, 32'sh2909343e, 32'sh2907ffa5, 32'sh2906cb06, 32'sh29059661, 
               32'sh290461b5, 32'sh29032d03, 32'sh2901f84b, 32'sh2900c38d, 32'sh28ff8ec8, 32'sh28fe59fc, 32'sh28fd252b, 32'sh28fbf053, 
               32'sh28fabb75, 32'sh28f98690, 32'sh28f851a6, 32'sh28f71cb4, 32'sh28f5e7bd, 32'sh28f4b2bf, 32'sh28f37dbb, 32'sh28f248b1, 
               32'sh28f113a0, 32'sh28efde89, 32'sh28eea96c, 32'sh28ed7448, 32'sh28ec3f1e, 32'sh28eb09ee, 32'sh28e9d4b7, 32'sh28e89f7a, 
               32'sh28e76a37, 32'sh28e634ee, 32'sh28e4ff9e, 32'sh28e3ca48, 32'sh28e294eb, 32'sh28e15f89, 32'sh28e02a20, 32'sh28def4b0, 
               32'sh28ddbf3b, 32'sh28dc89bf, 32'sh28db543c, 32'sh28da1eb4, 32'sh28d8e925, 32'sh28d7b390, 32'sh28d67df4, 32'sh28d54853, 
               32'sh28d412ab, 32'sh28d2dcfc, 32'sh28d1a748, 32'sh28d0718d, 32'sh28cf3bcc, 32'sh28ce0604, 32'sh28ccd036, 32'sh28cb9a62, 
               32'sh28ca6488, 32'sh28c92ea7, 32'sh28c7f8c0, 32'sh28c6c2d3, 32'sh28c58cdf, 32'sh28c456e6, 32'sh28c320e5, 32'sh28c1eadf, 
               32'sh28c0b4d2, 32'sh28bf7ebf, 32'sh28be48a6, 32'sh28bd1287, 32'sh28bbdc61, 32'sh28baa635, 32'sh28b97002, 32'sh28b839ca, 
               32'sh28b7038b, 32'sh28b5cd45, 32'sh28b496fa, 32'sh28b360a8, 32'sh28b22a50, 32'sh28b0f3f2, 32'sh28afbd8d, 32'sh28ae8722, 
               32'sh28ad50b1, 32'sh28ac1a3a, 32'sh28aae3bc, 32'sh28a9ad38, 32'sh28a876ae, 32'sh28a7401d, 32'sh28a60987, 32'sh28a4d2e9, 
               32'sh28a39c46, 32'sh28a2659d, 32'sh28a12eed, 32'sh289ff837, 32'sh289ec17a, 32'sh289d8ab8, 32'sh289c53ef, 32'sh289b1d20, 
               32'sh2899e64a, 32'sh2898af6e, 32'sh2897788c, 32'sh289641a4, 32'sh28950ab6, 32'sh2893d3c1, 32'sh28929cc6, 32'sh289165c5, 
               32'sh28902ebd, 32'sh288ef7b0, 32'sh288dc09c, 32'sh288c8981, 32'sh288b5261, 32'sh288a1b3a, 32'sh2888e40d, 32'sh2887acda, 
               32'sh288675a0, 32'sh28853e60, 32'sh2884071a, 32'sh2882cfce, 32'sh2881987c, 32'sh28806123, 32'sh287f29c4, 32'sh287df25f, 
               32'sh287cbaf3, 32'sh287b8381, 32'sh287a4c09, 32'sh2879148b, 32'sh2877dd07, 32'sh2876a57c, 32'sh28756deb, 32'sh28743654, 
               32'sh2872feb6, 32'sh2871c713, 32'sh28708f69, 32'sh286f57b9, 32'sh286e2002, 32'sh286ce846, 32'sh286bb083, 32'sh286a78ba, 
               32'sh286940ea, 32'sh28680915, 32'sh2866d139, 32'sh28659957, 32'sh2864616f, 32'sh28632980, 32'sh2861f18c, 32'sh2860b991, 
               32'sh285f8190, 32'sh285e4988, 32'sh285d117b, 32'sh285bd967, 32'sh285aa14d, 32'sh2859692d, 32'sh28583106, 32'sh2856f8d9, 
               32'sh2855c0a6, 32'sh2854886d, 32'sh2853502e, 32'sh285217e8, 32'sh2850df9d, 32'sh284fa74a, 32'sh284e6ef2, 32'sh284d3694, 
               32'sh284bfe2f, 32'sh284ac5c4, 32'sh28498d53, 32'sh284854dc, 32'sh28471c5e, 32'sh2845e3db, 32'sh2844ab51, 32'sh284372c0, 
               32'sh28423a2a, 32'sh2841018e, 32'sh283fc8eb, 32'sh283e9042, 32'sh283d5793, 32'sh283c1edd, 32'sh283ae622, 32'sh2839ad60, 
               32'sh28387498, 32'sh28373bca, 32'sh283602f5, 32'sh2834ca1a, 32'sh2833913a, 32'sh28325853, 32'sh28311f65, 32'sh282fe672, 
               32'sh282ead78, 32'sh282d7479, 32'sh282c3b73, 32'sh282b0266, 32'sh2829c954, 32'sh2828903b, 32'sh2827571d, 32'sh28261df8, 
               32'sh2824e4cc, 32'sh2823ab9b, 32'sh28227264, 32'sh28213926, 32'sh281fffe2, 32'sh281ec698, 32'sh281d8d48, 32'sh281c53f1, 
               32'sh281b1a94, 32'sh2819e132, 32'sh2818a7c8, 32'sh28176e59, 32'sh281634e4, 32'sh2814fb68, 32'sh2813c1e6, 32'sh2812885f, 
               32'sh28114ed0, 32'sh2810153c, 32'sh280edba2, 32'sh280da201, 32'sh280c685a, 32'sh280b2ead, 32'sh2809f4fa, 32'sh2808bb41, 
               32'sh28078181, 32'sh280647bb, 32'sh28050def, 32'sh2803d41d, 32'sh28029a45, 32'sh28016067, 32'sh28002682, 32'sh27feec97, 
               32'sh27fdb2a7, 32'sh27fc78af, 32'sh27fb3eb2, 32'sh27fa04af, 32'sh27f8caa5, 32'sh27f79096, 32'sh27f65680, 32'sh27f51c64, 
               32'sh27f3e241, 32'sh27f2a819, 32'sh27f16dea, 32'sh27f033b6, 32'sh27eef97b, 32'sh27edbf3a, 32'sh27ec84f3, 32'sh27eb4aa5, 
               32'sh27ea1052, 32'sh27e8d5f8, 32'sh27e79b98, 32'sh27e66133, 32'sh27e526c6, 32'sh27e3ec54, 32'sh27e2b1dc, 32'sh27e1775d, 
               32'sh27e03cd8, 32'sh27df024e, 32'sh27ddc7bd, 32'sh27dc8d25, 32'sh27db5288, 32'sh27da17e5, 32'sh27d8dd3b, 32'sh27d7a28b, 
               32'sh27d667d5, 32'sh27d52d19, 32'sh27d3f257, 32'sh27d2b78f, 32'sh27d17cc1, 32'sh27d041ec, 32'sh27cf0711, 32'sh27cdcc30, 
               32'sh27cc9149, 32'sh27cb565c, 32'sh27ca1b69, 32'sh27c8e06f, 32'sh27c7a570, 32'sh27c66a6a, 32'sh27c52f5e, 32'sh27c3f44c, 
               32'sh27c2b934, 32'sh27c17e16, 32'sh27c042f2, 32'sh27bf07c7, 32'sh27bdcc97, 32'sh27bc9160, 32'sh27bb5623, 32'sh27ba1ae0, 
               32'sh27b8df97, 32'sh27b7a448, 32'sh27b668f2, 32'sh27b52d97, 32'sh27b3f235, 32'sh27b2b6cd, 32'sh27b17b60, 32'sh27b03fec, 
               32'sh27af0472, 32'sh27adc8f1, 32'sh27ac8d6b, 32'sh27ab51df, 32'sh27aa164c, 32'sh27a8dab3, 32'sh27a79f14, 32'sh27a6636f, 
               32'sh27a527c4, 32'sh27a3ec13, 32'sh27a2b05c, 32'sh27a1749f, 32'sh27a038db, 32'sh279efd12, 32'sh279dc142, 32'sh279c856c, 
               32'sh279b4990, 32'sh279a0dae, 32'sh2798d1c6, 32'sh279795d8, 32'sh279659e3, 32'sh27951de9, 32'sh2793e1e8, 32'sh2792a5e2, 
               32'sh279169d5, 32'sh27902dc2, 32'sh278ef1a9, 32'sh278db58a, 32'sh278c7965, 32'sh278b3d39, 32'sh278a0108, 32'sh2788c4d1, 
               32'sh27878893, 32'sh27864c4f, 32'sh27851006, 32'sh2783d3b6, 32'sh27829760, 32'sh27815b04, 32'sh27801ea2, 32'sh277ee239, 
               32'sh277da5cb, 32'sh277c6957, 32'sh277b2cdc, 32'sh2779f05c, 32'sh2778b3d5, 32'sh27777748, 32'sh27763ab5, 32'sh2774fe1c, 
               32'sh2773c17d, 32'sh277284d8, 32'sh2771482d, 32'sh27700b7c, 32'sh276ecec5, 32'sh276d9207, 32'sh276c5544, 32'sh276b187a, 
               32'sh2769dbaa, 32'sh27689ed5, 32'sh276761f9, 32'sh27662517, 32'sh2764e82f, 32'sh2763ab41, 32'sh27626e4d, 32'sh27613153, 
               32'sh275ff452, 32'sh275eb74c, 32'sh275d7a40, 32'sh275c3d2d, 32'sh275b0014, 32'sh2759c2f6, 32'sh275885d1, 32'sh275748a6, 
               32'sh27560b76, 32'sh2754ce3f, 32'sh27539102, 32'sh275253bf, 32'sh27511676, 32'sh274fd926, 32'sh274e9bd1, 32'sh274d5e76, 
               32'sh274c2115, 32'sh274ae3ad, 32'sh2749a640, 32'sh274868cc, 32'sh27472b53, 32'sh2745edd3, 32'sh2744b04d, 32'sh274372c2, 
               32'sh27423530, 32'sh2740f798, 32'sh273fb9fa, 32'sh273e7c56, 32'sh273d3eac, 32'sh273c00fc, 32'sh273ac346, 32'sh2739858a, 
               32'sh273847c8, 32'sh273709ff, 32'sh2735cc31, 32'sh27348e5d, 32'sh27335082, 32'sh273212a2, 32'sh2730d4bb, 32'sh272f96cf, 
               32'sh272e58dc, 32'sh272d1ae4, 32'sh272bdce5, 32'sh272a9ee0, 32'sh272960d6, 32'sh272822c5, 32'sh2726e4ae, 32'sh2725a691, 
               32'sh2724686e, 32'sh27232a45, 32'sh2721ec16, 32'sh2720ade1, 32'sh271f6fa6, 32'sh271e3165, 32'sh271cf31e, 32'sh271bb4d1, 
               32'sh271a767e, 32'sh27193825, 32'sh2717f9c6, 32'sh2716bb60, 32'sh27157cf5, 32'sh27143e84, 32'sh2713000c, 32'sh2711c18f, 
               32'sh2710830c, 32'sh270f4482, 32'sh270e05f3, 32'sh270cc75d, 32'sh270b88c2, 32'sh270a4a21, 32'sh27090b79, 32'sh2707cccb, 
               32'sh27068e18, 32'sh27054f5e, 32'sh2704109f, 32'sh2702d1d9, 32'sh2701930e, 32'sh2700543c, 32'sh26ff1564, 32'sh26fdd687, 
               32'sh26fc97a3, 32'sh26fb58b9, 32'sh26fa19ca, 32'sh26f8dad4, 32'sh26f79bd8, 32'sh26f65cd6, 32'sh26f51dcf, 32'sh26f3dec1, 
               32'sh26f29fad, 32'sh26f16093, 32'sh26f02174, 32'sh26eee24e, 32'sh26eda322, 32'sh26ec63f0, 32'sh26eb24b9, 32'sh26e9e57b, 
               32'sh26e8a637, 32'sh26e766ed, 32'sh26e6279d, 32'sh26e4e848, 32'sh26e3a8ec, 32'sh26e2698a, 32'sh26e12a22, 32'sh26dfeab5, 
               32'sh26deab41, 32'sh26dd6bc7, 32'sh26dc2c47, 32'sh26daecc2, 32'sh26d9ad36, 32'sh26d86da4, 32'sh26d72e0c, 32'sh26d5ee6f, 
               32'sh26d4aecb, 32'sh26d36f21, 32'sh26d22f72, 32'sh26d0efbc, 32'sh26cfb000, 32'sh26ce703f, 32'sh26cd3077, 32'sh26cbf0aa, 
               32'sh26cab0d6, 32'sh26c970fc, 32'sh26c8311d, 32'sh26c6f137, 32'sh26c5b14c, 32'sh26c4715a, 32'sh26c33163, 32'sh26c1f165, 
               32'sh26c0b162, 32'sh26bf7159, 32'sh26be3149, 32'sh26bcf134, 32'sh26bbb119, 32'sh26ba70f7, 32'sh26b930d0, 32'sh26b7f0a3, 
               32'sh26b6b070, 32'sh26b57036, 32'sh26b42ff7, 32'sh26b2efb2, 32'sh26b1af67, 32'sh26b06f16, 32'sh26af2ebf, 32'sh26adee62, 
               32'sh26acadff, 32'sh26ab6d96, 32'sh26aa2d27, 32'sh26a8ecb3, 32'sh26a7ac38, 32'sh26a66bb7, 32'sh26a52b30, 32'sh26a3eaa4, 
               32'sh26a2aa11, 32'sh26a16978, 32'sh26a028da, 32'sh269ee835, 32'sh269da78b, 32'sh269c66da, 32'sh269b2624, 32'sh2699e568, 
               32'sh2698a4a6, 32'sh269763dd, 32'sh2696230f, 32'sh2694e23b, 32'sh2693a161, 32'sh26926081, 32'sh26911f9b, 32'sh268fdeaf, 
               32'sh268e9dbd, 32'sh268d5cc5, 32'sh268c1bc8, 32'sh268adac4, 32'sh268999ba, 32'sh268858ab, 32'sh26871795, 32'sh2685d67a, 
               32'sh26849558, 32'sh26835431, 32'sh26821303, 32'sh2680d1d0, 32'sh267f9097, 32'sh267e4f58, 32'sh267d0e13, 32'sh267bccc8, 
               32'sh267a8b77, 32'sh26794a20, 32'sh267808c3, 32'sh2676c761, 32'sh267585f8, 32'sh26744489, 32'sh26730315, 32'sh2671c19a, 
               32'sh2670801a, 32'sh266f3e94, 32'sh266dfd08, 32'sh266cbb75, 32'sh266b79dd, 32'sh266a383f, 32'sh2668f69b, 32'sh2667b4f2, 
               32'sh26667342, 32'sh2665318c, 32'sh2663efd1, 32'sh2662ae0f, 32'sh26616c48, 32'sh26602a7a, 32'sh265ee8a7, 32'sh265da6ce, 
               32'sh265c64ef, 32'sh265b230a, 32'sh2659e11f, 32'sh26589f2e, 32'sh26575d37, 32'sh26561b3a, 32'sh2654d938, 32'sh2653972f, 
               32'sh26525521, 32'sh2651130c, 32'sh264fd0f2, 32'sh264e8ed2, 32'sh264d4cac, 32'sh264c0a80, 32'sh264ac84e, 32'sh26498616, 
               32'sh264843d9, 32'sh26470195, 32'sh2645bf4b, 32'sh26447cfc, 32'sh26433aa7, 32'sh2641f84c, 32'sh2640b5eb, 32'sh263f7384, 
               32'sh263e3117, 32'sh263ceea4, 32'sh263bac2b, 32'sh263a69ad, 32'sh26392728, 32'sh2637e49e, 32'sh2636a20d, 32'sh26355f77, 
               32'sh26341cdb, 32'sh2632da39, 32'sh26319792, 32'sh263054e4, 32'sh262f1230, 32'sh262dcf77, 32'sh262c8cb7, 32'sh262b49f2, 
               32'sh262a0727, 32'sh2628c456, 32'sh2627817f, 32'sh26263ea2, 32'sh2624fbbf, 32'sh2623b8d7, 32'sh262275e8, 32'sh262132f4, 
               32'sh261feffa, 32'sh261eacfa, 32'sh261d69f4, 32'sh261c26e8, 32'sh261ae3d6, 32'sh2619a0be, 32'sh26185da1, 32'sh26171a7e, 
               32'sh2615d754, 32'sh26149425, 32'sh261350f0, 32'sh26120db5, 32'sh2610ca75, 32'sh260f872e, 32'sh260e43e2, 32'sh260d008f, 
               32'sh260bbd37, 32'sh260a79d9, 32'sh26093675, 32'sh2607f30b, 32'sh2606af9c, 32'sh26056c26, 32'sh260428ab, 32'sh2602e52a, 
               32'sh2601a1a2, 32'sh26005e15, 32'sh25ff1a83, 32'sh25fdd6ea, 32'sh25fc934b, 32'sh25fb4fa7, 32'sh25fa0bfd, 32'sh25f8c84d, 
               32'sh25f78497, 32'sh25f640db, 32'sh25f4fd19, 32'sh25f3b951, 32'sh25f27584, 32'sh25f131b1, 32'sh25efedd8, 32'sh25eea9f9, 
               32'sh25ed6614, 32'sh25ec2229, 32'sh25eade39, 32'sh25e99a42, 32'sh25e85646, 32'sh25e71244, 32'sh25e5ce3c, 32'sh25e48a2f, 
               32'sh25e3461b, 32'sh25e20202, 32'sh25e0bde2, 32'sh25df79bd, 32'sh25de3592, 32'sh25dcf162, 32'sh25dbad2b, 32'sh25da68ef, 
               32'sh25d924ac, 32'sh25d7e064, 32'sh25d69c16, 32'sh25d557c2, 32'sh25d41369, 32'sh25d2cf09, 32'sh25d18aa4, 32'sh25d04639, 
               32'sh25cf01c8, 32'sh25cdbd51, 32'sh25cc78d4, 32'sh25cb3452, 32'sh25c9efca, 32'sh25c8ab3c, 32'sh25c766a8, 32'sh25c6220e, 
               32'sh25c4dd6e, 32'sh25c398c9, 32'sh25c2541e, 32'sh25c10f6d, 32'sh25bfcab6, 32'sh25be85f9, 32'sh25bd4136, 32'sh25bbfc6e, 
               32'sh25bab7a0, 32'sh25b972cc, 32'sh25b82df2, 32'sh25b6e913, 32'sh25b5a42d, 32'sh25b45f42, 32'sh25b31a51, 32'sh25b1d55a, 
               32'sh25b0905d, 32'sh25af4b5b, 32'sh25ae0652, 32'sh25acc144, 32'sh25ab7c30, 32'sh25aa3717, 32'sh25a8f1f7, 32'sh25a7acd2, 
               32'sh25a667a7, 32'sh25a52276, 32'sh25a3dd3f, 32'sh25a29802, 32'sh25a152c0, 32'sh25a00d78, 32'sh259ec82a, 32'sh259d82d6, 
               32'sh259c3d7c, 32'sh259af81d, 32'sh2599b2b8, 32'sh25986d4d, 32'sh259727dc, 32'sh2595e265, 32'sh25949ce9, 32'sh25935767, 
               32'sh259211df, 32'sh2590cc51, 32'sh258f86be, 32'sh258e4124, 32'sh258cfb85, 32'sh258bb5e0, 32'sh258a7035, 32'sh25892a85, 
               32'sh2587e4cf, 32'sh25869f13, 32'sh25855951, 32'sh25841389, 32'sh2582cdbc, 32'sh258187e8, 32'sh2580420f, 32'sh257efc31, 
               32'sh257db64c, 32'sh257c7062, 32'sh257b2a71, 32'sh2579e47c, 32'sh25789e80, 32'sh2577587e, 32'sh25761277, 32'sh2574cc6a, 
               32'sh25738657, 32'sh2572403f, 32'sh2570fa20, 32'sh256fb3fc, 32'sh256e6dd2, 32'sh256d27a3, 32'sh256be16d, 32'sh256a9b32, 
               32'sh256954f1, 32'sh25680eaa, 32'sh2566c85e, 32'sh2565820b, 32'sh25643bb3, 32'sh2562f555, 32'sh2561aef2, 32'sh25606888, 
               32'sh255f2219, 32'sh255ddba4, 32'sh255c952a, 32'sh255b4ea9, 32'sh255a0823, 32'sh2558c197, 32'sh25577b06, 32'sh2556346e, 
               32'sh2554edd1, 32'sh2553a72e, 32'sh25526085, 32'sh255119d7, 32'sh254fd323, 32'sh254e8c69, 32'sh254d45a9, 32'sh254bfee3, 
               32'sh254ab818, 32'sh25497147, 32'sh25482a70, 32'sh2546e394, 32'sh25459cb2, 32'sh254455ca, 32'sh25430edc, 32'sh2541c7e8, 
               32'sh254080ef, 32'sh253f39f0, 32'sh253df2eb, 32'sh253cabe1, 32'sh253b64d1, 32'sh253a1dbb, 32'sh2538d69f, 32'sh25378f7e, 
               32'sh25364857, 32'sh2535012a, 32'sh2533b9f7, 32'sh253272bf, 32'sh25312b81, 32'sh252fe43d, 32'sh252e9cf3, 32'sh252d55a4, 
               32'sh252c0e4f, 32'sh252ac6f4, 32'sh25297f93, 32'sh2528382d, 32'sh2526f0c1, 32'sh2525a950, 32'sh252461d8, 32'sh25231a5b, 
               32'sh2521d2d8, 32'sh25208b4f, 32'sh251f43c1, 32'sh251dfc2d, 32'sh251cb493, 32'sh251b6cf4, 32'sh251a254e, 32'sh2518dda4, 
               32'sh251795f3, 32'sh25164e3c, 32'sh25150680, 32'sh2513bebf, 32'sh251276f7, 32'sh25112f2a, 32'sh250fe757, 32'sh250e9f7e, 
               32'sh250d57a0, 32'sh250c0fbb, 32'sh250ac7d2, 32'sh25097fe2, 32'sh250837ed, 32'sh2506eff2, 32'sh2505a7f1, 32'sh25045feb, 
               32'sh250317df, 32'sh2501cfcd, 32'sh250087b5, 32'sh24ff3f98, 32'sh24fdf775, 32'sh24fcaf4c, 32'sh24fb671e, 32'sh24fa1eea, 
               32'sh24f8d6b0, 32'sh24f78e71, 32'sh24f6462c, 32'sh24f4fde1, 32'sh24f3b590, 32'sh24f26d3a, 32'sh24f124de, 32'sh24efdc7d, 
               32'sh24ee9415, 32'sh24ed4ba8, 32'sh24ec0335, 32'sh24eababd, 32'sh24e9723f, 32'sh24e829bb, 32'sh24e6e132, 32'sh24e598a2, 
               32'sh24e4500e, 32'sh24e30773, 32'sh24e1bed3, 32'sh24e0762d, 32'sh24df2d81, 32'sh24dde4d0, 32'sh24dc9c19, 32'sh24db535c, 
               32'sh24da0a9a, 32'sh24d8c1d2, 32'sh24d77904, 32'sh24d63031, 32'sh24d4e757, 32'sh24d39e79, 32'sh24d25594, 32'sh24d10caa, 
               32'sh24cfc3ba, 32'sh24ce7ac5, 32'sh24cd31ca, 32'sh24cbe8c9, 32'sh24ca9fc2, 32'sh24c956b6, 32'sh24c80da4, 32'sh24c6c48d, 
               32'sh24c57b6f, 32'sh24c4324d, 32'sh24c2e924, 32'sh24c19ff6, 32'sh24c056c2, 32'sh24bf0d88, 32'sh24bdc449, 32'sh24bc7b04, 
               32'sh24bb31ba, 32'sh24b9e869, 32'sh24b89f14, 32'sh24b755b8, 32'sh24b60c57, 32'sh24b4c2f0, 32'sh24b37983, 32'sh24b23011, 
               32'sh24b0e699, 32'sh24af9d1c, 32'sh24ae5399, 32'sh24ad0a10, 32'sh24abc082, 32'sh24aa76ed, 32'sh24a92d54, 32'sh24a7e3b4, 
               32'sh24a69a0f, 32'sh24a55064, 32'sh24a406b4, 32'sh24a2bcfe, 32'sh24a17342, 32'sh24a02981, 32'sh249edfba, 32'sh249d95ed, 
               32'sh249c4c1b, 32'sh249b0243, 32'sh2499b865, 32'sh24986e82, 32'sh24972499, 32'sh2495daab, 32'sh249490b7, 32'sh249346bd, 
               32'sh2491fcbe, 32'sh2490b2b8, 32'sh248f68ae, 32'sh248e1e9d, 32'sh248cd487, 32'sh248b8a6c, 32'sh248a404b, 32'sh2488f624, 
               32'sh2487abf7, 32'sh248661c5, 32'sh2485178d, 32'sh2483cd50, 32'sh2482830d, 32'sh248138c4, 32'sh247fee76, 32'sh247ea422, 
               32'sh247d59c8, 32'sh247c0f69, 32'sh247ac504, 32'sh24797a9a, 32'sh2478302a, 32'sh2476e5b4, 32'sh24759b39, 32'sh247450b8, 
               32'sh24730631, 32'sh2471bba5, 32'sh24707113, 32'sh246f267c, 32'sh246ddbdf, 32'sh246c913c, 32'sh246b4694, 32'sh2469fbe6, 
               32'sh2468b132, 32'sh24676679, 32'sh24661bbb, 32'sh2464d0f6, 32'sh2463862c, 32'sh24623b5d, 32'sh2460f088, 32'sh245fa5ad, 
               32'sh245e5acc, 32'sh245d0fe6, 32'sh245bc4fb, 32'sh245a7a09, 32'sh24592f13, 32'sh2457e416, 32'sh24569914, 32'sh24554e0d, 
               32'sh245402ff, 32'sh2452b7ec, 32'sh24516cd4, 32'sh245021b6, 32'sh244ed692, 32'sh244d8b69, 32'sh244c403a, 32'sh244af506, 
               32'sh2449a9cc, 32'sh24485e8c, 32'sh24471347, 32'sh2445c7fc, 32'sh24447cac, 32'sh24433156, 32'sh2441e5fa, 32'sh24409a99, 
               32'sh243f4f32, 32'sh243e03c6, 32'sh243cb854, 32'sh243b6cdc, 32'sh243a215f, 32'sh2438d5dc, 32'sh24378a54, 32'sh24363ec6, 
               32'sh2434f332, 32'sh2433a799, 32'sh24325bfb, 32'sh24311056, 32'sh242fc4ad, 32'sh242e78fd, 32'sh242d2d48, 32'sh242be18e, 
               32'sh242a95ce, 32'sh24294a08, 32'sh2427fe3d, 32'sh2426b26c, 32'sh24256695, 32'sh24241ab9, 32'sh2422ced8, 32'sh242182f0, 
               32'sh24203704, 32'sh241eeb11, 32'sh241d9f1a, 32'sh241c531c, 32'sh241b0719, 32'sh2419bb11, 32'sh24186f02, 32'sh241722ef, 
               32'sh2415d6d5, 32'sh24148ab7, 32'sh24133e92, 32'sh2411f268, 32'sh2410a639, 32'sh240f5a04, 32'sh240e0dc9, 32'sh240cc189, 
               32'sh240b7543, 32'sh240a28f8, 32'sh2408dca7, 32'sh24079050, 32'sh240643f4, 32'sh2404f793, 32'sh2403ab2c, 32'sh24025ebf, 
               32'sh2401124d, 32'sh23ffc5d5, 32'sh23fe7958, 32'sh23fd2cd5, 32'sh23fbe04c, 32'sh23fa93be, 32'sh23f9472b, 32'sh23f7fa92, 
               32'sh23f6adf3, 32'sh23f5614f, 32'sh23f414a5, 32'sh23f2c7f6, 32'sh23f17b41, 32'sh23f02e87, 32'sh23eee1c7, 32'sh23ed9502, 
               32'sh23ec4837, 32'sh23eafb66, 32'sh23e9ae90, 32'sh23e861b4, 32'sh23e714d3, 32'sh23e5c7ed, 32'sh23e47b00, 32'sh23e32e0f, 
               32'sh23e1e117, 32'sh23e0941b, 32'sh23df4718, 32'sh23ddfa10, 32'sh23dcad03, 32'sh23db5ff0, 32'sh23da12d8, 32'sh23d8c5ba, 
               32'sh23d77896, 32'sh23d62b6d, 32'sh23d4de3f, 32'sh23d3910b, 32'sh23d243d1, 32'sh23d0f692, 32'sh23cfa94d, 32'sh23ce5c03, 
               32'sh23cd0eb3, 32'sh23cbc15e, 32'sh23ca7403, 32'sh23c926a3, 32'sh23c7d93d, 32'sh23c68bd2, 32'sh23c53e61, 32'sh23c3f0eb, 
               32'sh23c2a36f, 32'sh23c155ee, 32'sh23c00867, 32'sh23bebada, 32'sh23bd6d48, 32'sh23bc1fb1, 32'sh23bad214, 32'sh23b98472, 
               32'sh23b836ca, 32'sh23b6e91c, 32'sh23b59b69, 32'sh23b44db1, 32'sh23b2fff3, 32'sh23b1b22f, 32'sh23b06466, 32'sh23af1698, 
               32'sh23adc8c4, 32'sh23ac7aea, 32'sh23ab2d0b, 32'sh23a9df27, 32'sh23a8913d, 32'sh23a7434d, 32'sh23a5f558, 32'sh23a4a75e, 
               32'sh23a3595e, 32'sh23a20b59, 32'sh23a0bd4e, 32'sh239f6f3d, 32'sh239e2127, 32'sh239cd30c, 32'sh239b84eb, 32'sh239a36c4, 
               32'sh2398e898, 32'sh23979a67, 32'sh23964c30, 32'sh2394fdf4, 32'sh2393afb2, 32'sh2392616a, 32'sh2391131e, 32'sh238fc4cb, 
               32'sh238e7673, 32'sh238d2816, 32'sh238bd9b3, 32'sh238a8b4b, 32'sh23893cdd, 32'sh2387ee6a, 32'sh23869ff1, 32'sh23855173, 
               32'sh238402ef, 32'sh2382b466, 32'sh238165d8, 32'sh23801744, 32'sh237ec8aa, 32'sh237d7a0b, 32'sh237c2b66, 32'sh237adcbc, 
               32'sh23798e0d, 32'sh23783f58, 32'sh2376f09e, 32'sh2375a1de, 32'sh23745318, 32'sh2373044e, 32'sh2371b57d, 32'sh237066a8, 
               32'sh236f17cc, 32'sh236dc8ec, 32'sh236c7a06, 32'sh236b2b1a, 32'sh2369dc29, 32'sh23688d32, 32'sh23673e36, 32'sh2365ef35, 
               32'sh2364a02e, 32'sh23635122, 32'sh23620210, 32'sh2360b2f9, 32'sh235f63dc, 32'sh235e14ba, 32'sh235cc592, 32'sh235b7665, 
               32'sh235a2733, 32'sh2358d7fb, 32'sh235788bd, 32'sh2356397a, 32'sh2354ea32, 32'sh23539ae4, 32'sh23524b91, 32'sh2350fc38, 
               32'sh234facda, 32'sh234e5d76, 32'sh234d0e0d, 32'sh234bbe9f, 32'sh234a6f2b, 32'sh23491fb2, 32'sh2347d033, 32'sh234680af, 
               32'sh23453125, 32'sh2343e196, 32'sh23429201, 32'sh23414267, 32'sh233ff2c8, 32'sh233ea323, 32'sh233d5379, 32'sh233c03c9, 
               32'sh233ab414, 32'sh23396459, 32'sh23381499, 32'sh2336c4d4, 32'sh23357509, 32'sh23342539, 32'sh2332d563, 32'sh23318588, 
               32'sh233035a7, 32'sh232ee5c1, 32'sh232d95d6, 32'sh232c45e5, 32'sh232af5ee, 32'sh2329a5f3, 32'sh232855f2, 32'sh232705eb, 
               32'sh2325b5df, 32'sh232465ce, 32'sh232315b7, 32'sh2321c59a, 32'sh23207579, 32'sh231f2552, 32'sh231dd525, 32'sh231c84f3, 
               32'sh231b34bc, 32'sh2319e47f, 32'sh2318943d, 32'sh231743f5, 32'sh2315f3a8, 32'sh2314a356, 32'sh231352fe, 32'sh231202a1, 
               32'sh2310b23e, 32'sh230f61d6, 32'sh230e1169, 32'sh230cc0f6, 32'sh230b707e, 32'sh230a2000, 32'sh2308cf7d, 32'sh23077ef5, 
               32'sh23062e67, 32'sh2304ddd4, 32'sh23038d3b, 32'sh23023c9d, 32'sh2300ebf9, 32'sh22ff9b51, 32'sh22fe4aa2, 32'sh22fcf9ef, 
               32'sh22fba936, 32'sh22fa5877, 32'sh22f907b3, 32'sh22f7b6ea, 32'sh22f6661c, 32'sh22f51547, 32'sh22f3c46e, 32'sh22f2738f, 
               32'sh22f122ab, 32'sh22efd1c2, 32'sh22ee80d3, 32'sh22ed2fde, 32'sh22ebdee5, 32'sh22ea8de5, 32'sh22e93ce1, 32'sh22e7ebd7, 
               32'sh22e69ac8, 32'sh22e549b3, 32'sh22e3f899, 32'sh22e2a77a, 32'sh22e15655, 32'sh22e0052b, 32'sh22deb3fb, 32'sh22dd62c6, 
               32'sh22dc118c, 32'sh22dac04c, 32'sh22d96f07, 32'sh22d81dbd, 32'sh22d6cc6d, 32'sh22d57b18, 32'sh22d429bd, 32'sh22d2d85d, 
               32'sh22d186f8, 32'sh22d0358d, 32'sh22cee41d, 32'sh22cd92a8, 32'sh22cc412d, 32'sh22caefad, 32'sh22c99e28, 32'sh22c84c9d, 
               32'sh22c6fb0c, 32'sh22c5a977, 32'sh22c457dc, 32'sh22c3063c, 32'sh22c1b496, 32'sh22c062eb, 32'sh22bf113b, 32'sh22bdbf85, 
               32'sh22bc6dca, 32'sh22bb1c09, 32'sh22b9ca43, 32'sh22b87878, 32'sh22b726a8, 32'sh22b5d4d2, 32'sh22b482f7, 32'sh22b33116, 
               32'sh22b1df30, 32'sh22b08d45, 32'sh22af3b54, 32'sh22ade95e, 32'sh22ac9763, 32'sh22ab4562, 32'sh22a9f35c, 32'sh22a8a151, 
               32'sh22a74f40, 32'sh22a5fd2a, 32'sh22a4ab0f, 32'sh22a358ee, 32'sh22a206c8, 32'sh22a0b49c, 32'sh229f626c, 32'sh229e1035, 
               32'sh229cbdfa, 32'sh229b6bb9, 32'sh229a1973, 32'sh2298c728, 32'sh229774d7, 32'sh22962281, 32'sh2294d025, 32'sh22937dc5, 
               32'sh22922b5e, 32'sh2290d8f3, 32'sh228f8682, 32'sh228e340c, 32'sh228ce191, 32'sh228b8f10, 32'sh228a3c8a, 32'sh2288e9fe, 
               32'sh2287976e, 32'sh228644d7, 32'sh2284f23c, 32'sh22839f9b, 32'sh22824cf5, 32'sh2280fa4a, 32'sh227fa799, 32'sh227e54e3, 
               32'sh227d0228, 32'sh227baf67, 32'sh227a5ca1, 32'sh227909d6, 32'sh2277b705, 32'sh2276642f, 32'sh22751154, 32'sh2273be74, 
               32'sh22726b8e, 32'sh227118a3, 32'sh226fc5b2, 32'sh226e72bc, 32'sh226d1fc1, 32'sh226bccc1, 32'sh226a79bb, 32'sh226926b0, 
               32'sh2267d3a0, 32'sh2266808a, 32'sh22652d6f, 32'sh2263da4f, 32'sh22628729, 32'sh226133ff, 32'sh225fe0ce, 32'sh225e8d99, 
               32'sh225d3a5e, 32'sh225be71e, 32'sh225a93d9, 32'sh2259408e, 32'sh2257ed3e, 32'sh225699e9, 32'sh2255468e, 32'sh2253f32f, 
               32'sh22529fca, 32'sh22514c5f, 32'sh224ff8ef, 32'sh224ea57a, 32'sh224d5200, 32'sh224bfe81, 32'sh224aaafc, 32'sh22495771, 
               32'sh224803e2, 32'sh2246b04d, 32'sh22455cb3, 32'sh22440914, 32'sh2242b56f, 32'sh224161c6, 32'sh22400e16, 32'sh223eba62, 
               32'sh223d66a8, 32'sh223c12e9, 32'sh223abf25, 32'sh22396b5b, 32'sh2238178d, 32'sh2236c3b8, 32'sh22356fdf, 32'sh22341c00, 
               32'sh2232c81c, 32'sh22317433, 32'sh22302045, 32'sh222ecc51, 32'sh222d7858, 32'sh222c245a, 32'sh222ad056, 32'sh22297c4d, 
               32'sh2228283f, 32'sh2226d42c, 32'sh22258013, 32'sh22242bf5, 32'sh2222d7d2, 32'sh222183aa, 32'sh22202f7c, 32'sh221edb49, 
               32'sh221d8711, 32'sh221c32d3, 32'sh221ade91, 32'sh22198a49, 32'sh221835fb, 32'sh2216e1a9, 32'sh22158d51, 32'sh221438f4, 
               32'sh2212e492, 32'sh2211902a, 32'sh22103bbd, 32'sh220ee74b, 32'sh220d92d4, 32'sh220c3e57, 32'sh220ae9d6, 32'sh2209954f, 
               32'sh220840c2, 32'sh2206ec31, 32'sh2205979a, 32'sh220442fe, 32'sh2202ee5d, 32'sh220199b6, 32'sh2200450a, 32'sh21fef059, 
               32'sh21fd9ba3, 32'sh21fc46e7, 32'sh21faf227, 32'sh21f99d61, 32'sh21f84895, 32'sh21f6f3c5, 32'sh21f59eef, 32'sh21f44a14, 
               32'sh21f2f534, 32'sh21f1a04f, 32'sh21f04b64, 32'sh21eef674, 32'sh21eda17f, 32'sh21ec4c85, 32'sh21eaf785, 32'sh21e9a280, 
               32'sh21e84d76, 32'sh21e6f867, 32'sh21e5a353, 32'sh21e44e39, 32'sh21e2f91a, 32'sh21e1a3f6, 32'sh21e04ecc, 32'sh21def99e, 
               32'sh21dda46a, 32'sh21dc4f31, 32'sh21daf9f2, 32'sh21d9a4af, 32'sh21d84f66, 32'sh21d6fa18, 32'sh21d5a4c5, 32'sh21d44f6d, 
               32'sh21d2fa0f, 32'sh21d1a4ac, 32'sh21d04f44, 32'sh21cef9d7, 32'sh21cda465, 32'sh21cc4eed, 32'sh21caf970, 32'sh21c9a3ee, 
               32'sh21c84e67, 32'sh21c6f8da, 32'sh21c5a348, 32'sh21c44db1, 32'sh21c2f815, 32'sh21c1a274, 32'sh21c04ccd, 32'sh21bef722, 
               32'sh21bda171, 32'sh21bc4bba, 32'sh21baf5ff, 32'sh21b9a03e, 32'sh21b84a79, 32'sh21b6f4ae, 32'sh21b59ede, 32'sh21b44908, 
               32'sh21b2f32e, 32'sh21b19d4e, 32'sh21b04769, 32'sh21aef17f, 32'sh21ad9b8f, 32'sh21ac459b, 32'sh21aaefa1, 32'sh21a999a2, 
               32'sh21a8439e, 32'sh21a6ed95, 32'sh21a59786, 32'sh21a44173, 32'sh21a2eb5a, 32'sh21a1953c, 32'sh21a03f18, 32'sh219ee8f0, 
               32'sh219d92c2, 32'sh219c3c8f, 32'sh219ae657, 32'sh2199901a, 32'sh219839d8, 32'sh2196e390, 32'sh21958d44, 32'sh219436f2, 
               32'sh2192e09b, 32'sh21918a3e, 32'sh219033dd, 32'sh218edd76, 32'sh218d870b, 32'sh218c309a, 32'sh218ada24, 32'sh218983a8, 
               32'sh21882d28, 32'sh2186d6a2, 32'sh21858017, 32'sh21842987, 32'sh2182d2f2, 32'sh21817c58, 32'sh218025b8, 32'sh217ecf14, 
               32'sh217d786a, 32'sh217c21bb, 32'sh217acb07, 32'sh2179744e, 32'sh21781d8f, 32'sh2176c6cb, 32'sh21757003, 32'sh21741935, 
               32'sh2172c262, 32'sh21716b89, 32'sh217014ac, 32'sh216ebdc9, 32'sh216d66e2, 32'sh216c0ff5, 32'sh216ab903, 32'sh2169620b, 
               32'sh21680b0f, 32'sh2166b40e, 32'sh21655d07, 32'sh216405fb, 32'sh2162aeea, 32'sh216157d4, 32'sh216000b9, 32'sh215ea998, 
               32'sh215d5273, 32'sh215bfb48, 32'sh215aa418, 32'sh21594ce3, 32'sh2157f5a9, 32'sh21569e6a, 32'sh21554726, 32'sh2153efdc, 
               32'sh2152988d, 32'sh2151413a, 32'sh214fe9e1, 32'sh214e9283, 32'sh214d3b1f, 32'sh214be3b7, 32'sh214a8c49, 32'sh214934d7, 
               32'sh2147dd5f, 32'sh214685e2, 32'sh21452e60, 32'sh2143d6d9, 32'sh21427f4d, 32'sh214127bb, 32'sh213fd025, 32'sh213e7889, 
               32'sh213d20e8, 32'sh213bc942, 32'sh213a7197, 32'sh213919e7, 32'sh2137c232, 32'sh21366a77, 32'sh213512b8, 32'sh2133baf3, 
               32'sh21326329, 32'sh21310b5a, 32'sh212fb386, 32'sh212e5bad, 32'sh212d03cf, 32'sh212babec, 32'sh212a5403, 32'sh2128fc15, 
               32'sh2127a423, 32'sh21264c2b, 32'sh2124f42e, 32'sh21239c2c, 32'sh21224425, 32'sh2120ec18, 32'sh211f9407, 32'sh211e3bf1, 
               32'sh211ce3d5, 32'sh211b8bb4, 32'sh211a338e, 32'sh2118db64, 32'sh21178334, 32'sh21162afe, 32'sh2114d2c4, 32'sh21137a85, 
               32'sh21122240, 32'sh2110c9f7, 32'sh210f71a8, 32'sh210e1955, 32'sh210cc0fc, 32'sh210b689e, 32'sh210a103b, 32'sh2108b7d3, 
               32'sh21075f65, 32'sh210606f3, 32'sh2104ae7c, 32'sh210355ff, 32'sh2101fd7e, 32'sh2100a4f7, 32'sh20ff4c6b, 32'sh20fdf3da, 
               32'sh20fc9b44, 32'sh20fb42a9, 32'sh20f9ea09, 32'sh20f89164, 32'sh20f738ba, 32'sh20f5e00b, 32'sh20f48756, 32'sh20f32e9d, 
               32'sh20f1d5de, 32'sh20f07d1a, 32'sh20ef2451, 32'sh20edcb84, 32'sh20ec72b1, 32'sh20eb19d9, 32'sh20e9c0fc, 32'sh20e86819, 
               32'sh20e70f32, 32'sh20e5b646, 32'sh20e45d55, 32'sh20e3045e, 32'sh20e1ab63, 32'sh20e05262, 32'sh20def95c, 32'sh20dda052, 
               32'sh20dc4742, 32'sh20daee2d, 32'sh20d99513, 32'sh20d83bf4, 32'sh20d6e2d0, 32'sh20d589a7, 32'sh20d43079, 32'sh20d2d745, 
               32'sh20d17e0d, 32'sh20d024d0, 32'sh20cecb8d, 32'sh20cd7246, 32'sh20cc18f9, 32'sh20cabfa8, 32'sh20c96651, 32'sh20c80cf5, 
               32'sh20c6b395, 32'sh20c55a2f, 32'sh20c400c4, 32'sh20c2a754, 32'sh20c14ddf, 32'sh20bff465, 32'sh20be9ae6, 32'sh20bd4162, 
               32'sh20bbe7d8, 32'sh20ba8e4a, 32'sh20b934b7, 32'sh20b7db1f, 32'sh20b68181, 32'sh20b527df, 32'sh20b3ce37, 32'sh20b2748b, 
               32'sh20b11ad9, 32'sh20afc123, 32'sh20ae6767, 32'sh20ad0da6, 32'sh20abb3e1, 32'sh20aa5a16, 32'sh20a90046, 32'sh20a7a671, 
               32'sh20a64c97, 32'sh20a4f2b8, 32'sh20a398d5, 32'sh20a23eec, 32'sh20a0e4fe, 32'sh209f8b0b, 32'sh209e3112, 32'sh209cd715, 
               32'sh209b7d13, 32'sh209a230c, 32'sh2098c900, 32'sh20976eef, 32'sh209614d9, 32'sh2094babd, 32'sh2093609d, 32'sh20920678, 
               32'sh2090ac4d, 32'sh208f521e, 32'sh208df7ea, 32'sh208c9db0, 32'sh208b4372, 32'sh2089e92e, 32'sh20888ee6, 32'sh20873499, 
               32'sh2085da46, 32'sh20847fef, 32'sh20832592, 32'sh2081cb31, 32'sh208070ca, 32'sh207f165e, 32'sh207dbbee, 32'sh207c6178, 
               32'sh207b06fe, 32'sh2079ac7e, 32'sh207851fa, 32'sh2076f770, 32'sh20759ce1, 32'sh2074424e, 32'sh2072e7b5, 32'sh20718d18, 
               32'sh20703275, 32'sh206ed7cd, 32'sh206d7d21, 32'sh206c226f, 32'sh206ac7b8, 32'sh20696cfd, 32'sh2068123c, 32'sh2066b776, 
               32'sh20655cac, 32'sh206401dc, 32'sh2062a708, 32'sh20614c2e, 32'sh205ff14f, 32'sh205e966c, 32'sh205d3b83, 32'sh205be096, 
               32'sh205a85a3, 32'sh20592aac, 32'sh2057cfaf, 32'sh205674ad, 32'sh205519a7, 32'sh2053be9b, 32'sh2052638b, 32'sh20510875, 
               32'sh204fad5b, 32'sh204e523c, 32'sh204cf717, 32'sh204b9bee, 32'sh204a40bf, 32'sh2048e58c, 32'sh20478a54, 32'sh20462f16, 
               32'sh2044d3d4, 32'sh2043788d, 32'sh20421d41, 32'sh2040c1ef, 32'sh203f6699, 32'sh203e0b3e, 32'sh203cafde, 32'sh203b5479, 
               32'sh2039f90f, 32'sh20389da0, 32'sh2037422c, 32'sh2035e6b3, 32'sh20348b35, 32'sh20332fb2, 32'sh2031d42a, 32'sh2030789d, 
               32'sh202f1d0b, 32'sh202dc174, 32'sh202c65d9, 32'sh202b0a38, 32'sh2029ae92, 32'sh202852e8, 32'sh2026f738, 32'sh20259b83, 
               32'sh20243fca, 32'sh2022e40b, 32'sh20218848, 32'sh20202c80, 32'sh201ed0b2, 32'sh201d74e0, 32'sh201c1909, 32'sh201abd2d, 
               32'sh2019614c, 32'sh20180565, 32'sh2016a97a, 32'sh20154d8a, 32'sh2013f196, 32'sh2012959c, 32'sh2011399d, 32'sh200fdd99, 
               32'sh200e8190, 32'sh200d2583, 32'sh200bc970, 32'sh200a6d59, 32'sh2009113c, 32'sh2007b51b, 32'sh200658f4, 32'sh2004fcc9, 
               32'sh2003a099, 32'sh20024464, 32'sh2000e829, 32'sh1fff8bea, 32'sh1ffe2fa6, 32'sh1ffcd35e, 32'sh1ffb7710, 32'sh1ffa1abd, 
               32'sh1ff8be65, 32'sh1ff76209, 32'sh1ff605a7, 32'sh1ff4a941, 32'sh1ff34cd5, 32'sh1ff1f065, 32'sh1ff093ef, 32'sh1fef3775, 
               32'sh1feddaf6, 32'sh1fec7e72, 32'sh1feb21e9, 32'sh1fe9c55b, 32'sh1fe868c8, 32'sh1fe70c31, 32'sh1fe5af94, 32'sh1fe452f2, 
               32'sh1fe2f64c, 32'sh1fe199a0, 32'sh1fe03cf0, 32'sh1fdee03b, 32'sh1fdd8381, 32'sh1fdc26c2, 32'sh1fdac9fe, 32'sh1fd96d35, 
               32'sh1fd81067, 32'sh1fd6b394, 32'sh1fd556bd, 32'sh1fd3f9e0, 32'sh1fd29cff, 32'sh1fd14018, 32'sh1fcfe32d, 32'sh1fce863d, 
               32'sh1fcd2948, 32'sh1fcbcc4e, 32'sh1fca6f4f, 32'sh1fc9124b, 32'sh1fc7b542, 32'sh1fc65835, 32'sh1fc4fb22, 32'sh1fc39e0b, 
               32'sh1fc240ef, 32'sh1fc0e3cd, 32'sh1fbf86a7, 32'sh1fbe297c, 32'sh1fbccc4d, 32'sh1fbb6f18, 32'sh1fba11de, 32'sh1fb8b4a0, 
               32'sh1fb7575c, 32'sh1fb5fa14, 32'sh1fb49cc7, 32'sh1fb33f74, 32'sh1fb1e21d, 32'sh1fb084c2, 32'sh1faf2761, 32'sh1fadc9fb, 
               32'sh1fac6c91, 32'sh1fab0f21, 32'sh1fa9b1ad, 32'sh1fa85434, 32'sh1fa6f6b6, 32'sh1fa59933, 32'sh1fa43bab, 32'sh1fa2de1e, 
               32'sh1fa1808c, 32'sh1fa022f6, 32'sh1f9ec55b, 32'sh1f9d67ba, 32'sh1f9c0a15, 32'sh1f9aac6b, 32'sh1f994ebc, 32'sh1f97f109, 
               32'sh1f969350, 32'sh1f953593, 32'sh1f93d7d0, 32'sh1f927a09, 32'sh1f911c3d, 32'sh1f8fbe6c, 32'sh1f8e6096, 32'sh1f8d02bc, 
               32'sh1f8ba4dc, 32'sh1f8a46f8, 32'sh1f88e90e, 32'sh1f878b20, 32'sh1f862d2d, 32'sh1f84cf35, 32'sh1f837139, 32'sh1f821337, 
               32'sh1f80b531, 32'sh1f7f5725, 32'sh1f7df915, 32'sh1f7c9b00, 32'sh1f7b3ce6, 32'sh1f79dec7, 32'sh1f7880a4, 32'sh1f77227b, 
               32'sh1f75c44e, 32'sh1f74661c, 32'sh1f7307e5, 32'sh1f71a9a9, 32'sh1f704b69, 32'sh1f6eed23, 32'sh1f6d8ed9, 32'sh1f6c3089, 
               32'sh1f6ad235, 32'sh1f6973dc, 32'sh1f68157f, 32'sh1f66b71c, 32'sh1f6558b5, 32'sh1f63fa48, 32'sh1f629bd7, 32'sh1f613d61, 
               32'sh1f5fdee6, 32'sh1f5e8067, 32'sh1f5d21e2, 32'sh1f5bc359, 32'sh1f5a64cb, 32'sh1f590638, 32'sh1f57a7a0, 32'sh1f564903, 
               32'sh1f54ea62, 32'sh1f538bbb, 32'sh1f522d10, 32'sh1f50ce60, 32'sh1f4f6fab, 32'sh1f4e10f2, 32'sh1f4cb233, 32'sh1f4b5370, 
               32'sh1f49f4a8, 32'sh1f4895db, 32'sh1f473709, 32'sh1f45d833, 32'sh1f447957, 32'sh1f431a77, 32'sh1f41bb92, 32'sh1f405ca8, 
               32'sh1f3efdb9, 32'sh1f3d9ec6, 32'sh1f3c3fcd, 32'sh1f3ae0d0, 32'sh1f3981ce, 32'sh1f3822c7, 32'sh1f36c3bc, 32'sh1f3564ab, 
               32'sh1f340596, 32'sh1f32a67c, 32'sh1f31475d, 32'sh1f2fe83a, 32'sh1f2e8911, 32'sh1f2d29e4, 32'sh1f2bcab2, 32'sh1f2a6b7b, 
               32'sh1f290c3f, 32'sh1f27acff, 32'sh1f264db9, 32'sh1f24ee6f, 32'sh1f238f20, 32'sh1f222fcd, 32'sh1f20d074, 32'sh1f1f7117, 
               32'sh1f1e11b5, 32'sh1f1cb24e, 32'sh1f1b52e2, 32'sh1f19f372, 32'sh1f1893fc, 32'sh1f173482, 32'sh1f15d503, 32'sh1f147580, 
               32'sh1f1315f7, 32'sh1f11b66a, 32'sh1f1056d8, 32'sh1f0ef741, 32'sh1f0d97a5, 32'sh1f0c3805, 32'sh1f0ad860, 32'sh1f0978b6, 
               32'sh1f081907, 32'sh1f06b953, 32'sh1f05599b, 32'sh1f03f9de, 32'sh1f029a1c, 32'sh1f013a55, 32'sh1effda89, 32'sh1efe7ab9, 
               32'sh1efd1ae4, 32'sh1efbbb0a, 32'sh1efa5b2c, 32'sh1ef8fb48, 32'sh1ef79b60, 32'sh1ef63b73, 32'sh1ef4db81, 32'sh1ef37b8b, 
               32'sh1ef21b90, 32'sh1ef0bb90, 32'sh1eef5b8b, 32'sh1eedfb81, 32'sh1eec9b73, 32'sh1eeb3b60, 32'sh1ee9db48, 32'sh1ee87b2b, 
               32'sh1ee71b0a, 32'sh1ee5bae4, 32'sh1ee45ab9, 32'sh1ee2fa89, 32'sh1ee19a54, 32'sh1ee03a1b, 32'sh1eded9dd, 32'sh1edd799a, 
               32'sh1edc1953, 32'sh1edab907, 32'sh1ed958b6, 32'sh1ed7f860, 32'sh1ed69805, 32'sh1ed537a6, 32'sh1ed3d742, 32'sh1ed276d9, 
               32'sh1ed1166b, 32'sh1ecfb5f9, 32'sh1ece5582, 32'sh1eccf506, 32'sh1ecb9486, 32'sh1eca3400, 32'sh1ec8d376, 32'sh1ec772e7, 
               32'sh1ec61254, 32'sh1ec4b1bc, 32'sh1ec3511f, 32'sh1ec1f07d, 32'sh1ec08fd6, 32'sh1ebf2f2b, 32'sh1ebdce7b, 32'sh1ebc6dc6, 
               32'sh1ebb0d0d, 32'sh1eb9ac4e, 32'sh1eb84b8b, 32'sh1eb6eac4, 32'sh1eb589f7, 32'sh1eb42926, 32'sh1eb2c850, 32'sh1eb16775, 
               32'sh1eb00696, 32'sh1eaea5b2, 32'sh1ead44c9, 32'sh1eabe3db, 32'sh1eaa82e9, 32'sh1ea921f2, 32'sh1ea7c0f6, 32'sh1ea65ff6, 
               32'sh1ea4fef0, 32'sh1ea39de6, 32'sh1ea23cd8, 32'sh1ea0dbc4, 32'sh1e9f7aac, 32'sh1e9e198f, 32'sh1e9cb86e, 32'sh1e9b5748, 
               32'sh1e99f61d, 32'sh1e9894ed, 32'sh1e9733b8, 32'sh1e95d27f, 32'sh1e947141, 32'sh1e930fff, 32'sh1e91aeb7, 32'sh1e904d6b, 
               32'sh1e8eec1b, 32'sh1e8d8ac5, 32'sh1e8c296b, 32'sh1e8ac80c, 32'sh1e8966a8, 32'sh1e880540, 32'sh1e86a3d3, 32'sh1e854261, 
               32'sh1e83e0eb, 32'sh1e827f70, 32'sh1e811df0, 32'sh1e7fbc6b, 32'sh1e7e5ae2, 32'sh1e7cf954, 32'sh1e7b97c2, 32'sh1e7a362a, 
               32'sh1e78d48e, 32'sh1e7772ed, 32'sh1e761148, 32'sh1e74af9e, 32'sh1e734def, 32'sh1e71ec3c, 32'sh1e708a83, 32'sh1e6f28c6, 
               32'sh1e6dc705, 32'sh1e6c653e, 32'sh1e6b0373, 32'sh1e69a1a4, 32'sh1e683fcf, 32'sh1e66ddf6, 32'sh1e657c19, 32'sh1e641a36, 
               32'sh1e62b84f, 32'sh1e615663, 32'sh1e5ff473, 32'sh1e5e927d, 32'sh1e5d3084, 32'sh1e5bce85, 32'sh1e5a6c82, 32'sh1e590a7a, 
               32'sh1e57a86d, 32'sh1e56465c, 32'sh1e54e446, 32'sh1e53822b, 32'sh1e52200c, 32'sh1e50bde8, 32'sh1e4f5bbf, 32'sh1e4df992, 
               32'sh1e4c9760, 32'sh1e4b3529, 32'sh1e49d2ee, 32'sh1e4870ae, 32'sh1e470e69, 32'sh1e45ac20, 32'sh1e4449d2, 32'sh1e42e77f, 
               32'sh1e418528, 32'sh1e4022cc, 32'sh1e3ec06b, 32'sh1e3d5e06, 32'sh1e3bfb9c, 32'sh1e3a992d, 32'sh1e3936ba, 32'sh1e37d442, 
               32'sh1e3671c5, 32'sh1e350f44, 32'sh1e33acbe, 32'sh1e324a33, 32'sh1e30e7a4, 32'sh1e2f8510, 32'sh1e2e2277, 32'sh1e2cbfda, 
               32'sh1e2b5d38, 32'sh1e29fa91, 32'sh1e2897e6, 32'sh1e273536, 32'sh1e25d282, 32'sh1e246fc9, 32'sh1e230d0b, 32'sh1e21aa48, 
               32'sh1e204781, 32'sh1e1ee4b5, 32'sh1e1d81e5, 32'sh1e1c1f10, 32'sh1e1abc36, 32'sh1e195958, 32'sh1e17f675, 32'sh1e16938d, 
               32'sh1e1530a1, 32'sh1e13cdb0, 32'sh1e126abb, 32'sh1e1107c1, 32'sh1e0fa4c2, 32'sh1e0e41be, 32'sh1e0cdeb6, 32'sh1e0b7ba9, 
               32'sh1e0a1898, 32'sh1e08b582, 32'sh1e075268, 32'sh1e05ef48, 32'sh1e048c24, 32'sh1e0328fc, 32'sh1e01c5cf, 32'sh1e00629d, 
               32'sh1dfeff67, 32'sh1dfd9c2c, 32'sh1dfc38ec, 32'sh1dfad5a8, 32'sh1df9725f, 32'sh1df80f11, 32'sh1df6abbf, 32'sh1df54868, 
               32'sh1df3e50d, 32'sh1df281ad, 32'sh1df11e49, 32'sh1defbadf, 32'sh1dee5771, 32'sh1decf3ff, 32'sh1deb9088, 32'sh1dea2d0c, 
               32'sh1de8c98c, 32'sh1de76607, 32'sh1de6027e, 32'sh1de49eef, 32'sh1de33b5d, 32'sh1de1d7c5, 32'sh1de07429, 32'sh1ddf1089, 
               32'sh1dddace4, 32'sh1ddc493a, 32'sh1ddae58b, 32'sh1dd981d8, 32'sh1dd81e21, 32'sh1dd6ba65, 32'sh1dd556a4, 32'sh1dd3f2df, 
               32'sh1dd28f15, 32'sh1dd12b46, 32'sh1dcfc773, 32'sh1dce639b, 32'sh1dccffbf, 32'sh1dcb9bde, 32'sh1dca37f8, 32'sh1dc8d40e, 
               32'sh1dc7701f, 32'sh1dc60c2c, 32'sh1dc4a834, 32'sh1dc34437, 32'sh1dc1e036, 32'sh1dc07c30, 32'sh1dbf1826, 32'sh1dbdb417, 
               32'sh1dbc5004, 32'sh1dbaebec, 32'sh1db987cf, 32'sh1db823ae, 32'sh1db6bf88, 32'sh1db55b5e, 32'sh1db3f72f, 32'sh1db292fb, 
               32'sh1db12ec3, 32'sh1dafca86, 32'sh1dae6645, 32'sh1dad01ff, 32'sh1dab9db5, 32'sh1daa3965, 32'sh1da8d512, 32'sh1da770ba, 
               32'sh1da60c5d, 32'sh1da4a7fc, 32'sh1da34396, 32'sh1da1df2b, 32'sh1da07abc, 32'sh1d9f1649, 32'sh1d9db1d1, 32'sh1d9c4d54, 
               32'sh1d9ae8d2, 32'sh1d99844d, 32'sh1d981fc2, 32'sh1d96bb33, 32'sh1d9556a0, 32'sh1d93f207, 32'sh1d928d6b, 32'sh1d9128ca, 
               32'sh1d8fc424, 32'sh1d8e5f79, 32'sh1d8cfaca, 32'sh1d8b9617, 32'sh1d8a315f, 32'sh1d88cca2, 32'sh1d8767e1, 32'sh1d86031c, 
               32'sh1d849e51, 32'sh1d833983, 32'sh1d81d4af, 32'sh1d806fd7, 32'sh1d7f0afb, 32'sh1d7da61a, 32'sh1d7c4134, 32'sh1d7adc4a, 
               32'sh1d79775c, 32'sh1d781268, 32'sh1d76ad71, 32'sh1d754874, 32'sh1d73e374, 32'sh1d727e6e, 32'sh1d711964, 32'sh1d6fb456, 
               32'sh1d6e4f43, 32'sh1d6cea2b, 32'sh1d6b850f, 32'sh1d6a1fef, 32'sh1d68baca, 32'sh1d6755a0, 32'sh1d65f072, 32'sh1d648b3f, 
               32'sh1d632608, 32'sh1d61c0cc, 32'sh1d605b8c, 32'sh1d5ef647, 32'sh1d5d90fd, 32'sh1d5c2baf, 32'sh1d5ac65d, 32'sh1d596106, 
               32'sh1d57fbaa, 32'sh1d56964a, 32'sh1d5530e6, 32'sh1d53cb7d, 32'sh1d52660f, 32'sh1d51009d, 32'sh1d4f9b26, 32'sh1d4e35ab, 
               32'sh1d4cd02c, 32'sh1d4b6aa7, 32'sh1d4a051f, 32'sh1d489f92, 32'sh1d473a00, 32'sh1d45d46a, 32'sh1d446ecf, 32'sh1d43092f, 
               32'sh1d41a38c, 32'sh1d403de3, 32'sh1d3ed837, 32'sh1d3d7285, 32'sh1d3c0ccf, 32'sh1d3aa715, 32'sh1d394156, 32'sh1d37db93, 
               32'sh1d3675cb, 32'sh1d350fff, 32'sh1d33aa2e, 32'sh1d324458, 32'sh1d30de7e, 32'sh1d2f78a0, 32'sh1d2e12bd, 32'sh1d2cacd6, 
               32'sh1d2b46ea, 32'sh1d29e0f9, 32'sh1d287b05, 32'sh1d27150b, 32'sh1d25af0d, 32'sh1d24490b, 32'sh1d22e304, 32'sh1d217cf9, 
               32'sh1d2016e9, 32'sh1d1eb0d5, 32'sh1d1d4abc, 32'sh1d1be49e, 32'sh1d1a7e7d, 32'sh1d191856, 32'sh1d17b22c, 32'sh1d164bfc, 
               32'sh1d14e5c9, 32'sh1d137f90, 32'sh1d121954, 32'sh1d10b312, 32'sh1d0f4ccd, 32'sh1d0de682, 32'sh1d0c8034, 32'sh1d0b19e1, 
               32'sh1d09b389, 32'sh1d084d2d, 32'sh1d06e6cc, 32'sh1d058067, 32'sh1d0419fe, 32'sh1d02b390, 32'sh1d014d1d, 32'sh1cffe6a6, 
               32'sh1cfe802b, 32'sh1cfd19ab, 32'sh1cfbb327, 32'sh1cfa4c9e, 32'sh1cf8e611, 32'sh1cf77f7f, 32'sh1cf618e9, 32'sh1cf4b24e, 
               32'sh1cf34baf, 32'sh1cf1e50b, 32'sh1cf07e63, 32'sh1cef17b7, 32'sh1cedb106, 32'sh1cec4a50, 32'sh1ceae396, 32'sh1ce97cd8, 
               32'sh1ce81615, 32'sh1ce6af4e, 32'sh1ce54882, 32'sh1ce3e1b2, 32'sh1ce27add, 32'sh1ce11404, 32'sh1cdfad26, 32'sh1cde4644, 
               32'sh1cdcdf5e, 32'sh1cdb7873, 32'sh1cda1183, 32'sh1cd8aa90, 32'sh1cd74397, 32'sh1cd5dc9b, 32'sh1cd47599, 32'sh1cd30e94, 
               32'sh1cd1a78a, 32'sh1cd0407b, 32'sh1cced968, 32'sh1ccd7251, 32'sh1ccc0b35, 32'sh1ccaa415, 32'sh1cc93cf0, 32'sh1cc7d5c7, 
               32'sh1cc66e99, 32'sh1cc50767, 32'sh1cc3a031, 32'sh1cc238f6, 32'sh1cc0d1b6, 32'sh1cbf6a73, 32'sh1cbe032a, 32'sh1cbc9bde, 
               32'sh1cbb348d, 32'sh1cb9cd37, 32'sh1cb865dd, 32'sh1cb6fe7f, 32'sh1cb5971c, 32'sh1cb42fb5, 32'sh1cb2c849, 32'sh1cb160d9, 
               32'sh1caff965, 32'sh1cae91ec, 32'sh1cad2a6e, 32'sh1cabc2ed, 32'sh1caa5b66, 32'sh1ca8f3dc, 32'sh1ca78c4d, 32'sh1ca624b9, 
               32'sh1ca4bd21, 32'sh1ca35585, 32'sh1ca1ede4, 32'sh1ca0863f, 32'sh1c9f1e96, 32'sh1c9db6e8, 32'sh1c9c4f35, 32'sh1c9ae77f, 
               32'sh1c997fc4, 32'sh1c981804, 32'sh1c96b040, 32'sh1c954878, 32'sh1c93e0ab, 32'sh1c9278d9, 32'sh1c911104, 32'sh1c8fa92a, 
               32'sh1c8e414b, 32'sh1c8cd969, 32'sh1c8b7181, 32'sh1c8a0996, 32'sh1c88a1a6, 32'sh1c8739b1, 32'sh1c85d1b8, 32'sh1c8469bb, 
               32'sh1c8301b9, 32'sh1c8199b3, 32'sh1c8031a9, 32'sh1c7ec99a, 32'sh1c7d6187, 32'sh1c7bf96f, 32'sh1c7a9153, 32'sh1c792933, 
               32'sh1c77c10e, 32'sh1c7658e5, 32'sh1c74f0b7, 32'sh1c738885, 32'sh1c72204f, 32'sh1c70b814, 32'sh1c6f4fd5, 32'sh1c6de791, 
               32'sh1c6c7f4a, 32'sh1c6b16fd, 32'sh1c69aead, 32'sh1c684658, 32'sh1c66ddfe, 32'sh1c6575a0, 32'sh1c640d3e, 32'sh1c62a4d8, 
               32'sh1c613c6d, 32'sh1c5fd3fd, 32'sh1c5e6b8a, 32'sh1c5d0312, 32'sh1c5b9a95, 32'sh1c5a3214, 32'sh1c58c98f, 32'sh1c576106, 
               32'sh1c55f878, 32'sh1c548fe5, 32'sh1c53274f, 32'sh1c51beb4, 32'sh1c505614, 32'sh1c4eed71, 32'sh1c4d84c8, 32'sh1c4c1c1c, 
               32'sh1c4ab36b, 32'sh1c494ab6, 32'sh1c47e1fc, 32'sh1c46793e, 32'sh1c45107c, 32'sh1c43a7b5, 32'sh1c423eea, 32'sh1c40d61b, 
               32'sh1c3f6d47, 32'sh1c3e046f, 32'sh1c3c9b93, 32'sh1c3b32b2, 32'sh1c39c9cd, 32'sh1c3860e3, 32'sh1c36f7f5, 32'sh1c358f03, 
               32'sh1c34260c, 32'sh1c32bd12, 32'sh1c315412, 32'sh1c2feb0f, 32'sh1c2e8207, 32'sh1c2d18fa, 32'sh1c2bafea, 32'sh1c2a46d5, 
               32'sh1c28ddbb, 32'sh1c27749e, 32'sh1c260b7c, 32'sh1c24a255, 32'sh1c23392b, 32'sh1c21cffc, 32'sh1c2066c8, 32'sh1c1efd91, 
               32'sh1c1d9454, 32'sh1c1c2b14, 32'sh1c1ac1cf, 32'sh1c195886, 32'sh1c17ef39, 32'sh1c1685e7, 32'sh1c151c91, 32'sh1c13b337, 
               32'sh1c1249d8, 32'sh1c10e075, 32'sh1c0f770e, 32'sh1c0e0da2, 32'sh1c0ca432, 32'sh1c0b3abe, 32'sh1c09d145, 32'sh1c0867c8, 
               32'sh1c06fe46, 32'sh1c0594c1, 32'sh1c042b37, 32'sh1c02c1a9, 32'sh1c015816, 32'sh1bffee7f, 32'sh1bfe84e4, 32'sh1bfd1b44, 
               32'sh1bfbb1a0, 32'sh1bfa47f8, 32'sh1bf8de4c, 32'sh1bf7749b, 32'sh1bf60ae6, 32'sh1bf4a12c, 32'sh1bf3376f, 32'sh1bf1cdac, 
               32'sh1bf063e6, 32'sh1beefa1b, 32'sh1bed904c, 32'sh1bec2679, 32'sh1beabca1, 32'sh1be952c6, 32'sh1be7e8e5, 32'sh1be67f01, 
               32'sh1be51518, 32'sh1be3ab2b, 32'sh1be24139, 32'sh1be0d744, 32'sh1bdf6d4a, 32'sh1bde034b, 32'sh1bdc9949, 32'sh1bdb2f42, 
               32'sh1bd9c537, 32'sh1bd85b27, 32'sh1bd6f113, 32'sh1bd586fb, 32'sh1bd41cdf, 32'sh1bd2b2be, 32'sh1bd14899, 32'sh1bcfde70, 
               32'sh1bce7442, 32'sh1bcd0a11, 32'sh1bcb9fda, 32'sh1bca35a0, 32'sh1bc8cb61, 32'sh1bc7611e, 32'sh1bc5f6d7, 32'sh1bc48c8c, 
               32'sh1bc3223c, 32'sh1bc1b7e8, 32'sh1bc04d8f, 32'sh1bbee333, 32'sh1bbd78d2, 32'sh1bbc0e6c, 32'sh1bbaa403, 32'sh1bb93995, 
               32'sh1bb7cf23, 32'sh1bb664ad, 32'sh1bb4fa32, 32'sh1bb38fb3, 32'sh1bb22530, 32'sh1bb0baa9, 32'sh1baf501d, 32'sh1bade58d, 
               32'sh1bac7af9, 32'sh1bab1060, 32'sh1ba9a5c4, 32'sh1ba83b22, 32'sh1ba6d07d, 32'sh1ba565d4, 32'sh1ba3fb26, 32'sh1ba29074, 
               32'sh1ba125bd, 32'sh1b9fbb03, 32'sh1b9e5044, 32'sh1b9ce581, 32'sh1b9b7ab9, 32'sh1b9a0fee, 32'sh1b98a51e, 32'sh1b973a4a, 
               32'sh1b95cf71, 32'sh1b946495, 32'sh1b92f9b4, 32'sh1b918ecf, 32'sh1b9023e5, 32'sh1b8eb8f7, 32'sh1b8d4e06, 32'sh1b8be30f, 
               32'sh1b8a7815, 32'sh1b890d16, 32'sh1b87a213, 32'sh1b86370c, 32'sh1b84cc01, 32'sh1b8360f1, 32'sh1b81f5dd, 32'sh1b808ac5, 
               32'sh1b7f1fa9, 32'sh1b7db488, 32'sh1b7c4963, 32'sh1b7ade3a, 32'sh1b79730d, 32'sh1b7807db, 32'sh1b769ca6, 32'sh1b75316c, 
               32'sh1b73c62d, 32'sh1b725aeb, 32'sh1b70efa4, 32'sh1b6f8459, 32'sh1b6e190a, 32'sh1b6cadb7, 32'sh1b6b425f, 32'sh1b69d703, 
               32'sh1b686ba3, 32'sh1b67003f, 32'sh1b6594d6, 32'sh1b642969, 32'sh1b62bdf8, 32'sh1b615283, 32'sh1b5fe709, 32'sh1b5e7b8c, 
               32'sh1b5d100a, 32'sh1b5ba484, 32'sh1b5a38f9, 32'sh1b58cd6b, 32'sh1b5761d8, 32'sh1b55f641, 32'sh1b548aa6, 32'sh1b531f06, 
               32'sh1b51b363, 32'sh1b5047bb, 32'sh1b4edc0f, 32'sh1b4d705f, 32'sh1b4c04aa, 32'sh1b4a98f1, 32'sh1b492d35, 32'sh1b47c173, 
               32'sh1b4655ae, 32'sh1b44e9e5, 32'sh1b437e17, 32'sh1b421245, 32'sh1b40a66f, 32'sh1b3f3a95, 32'sh1b3dceb6, 32'sh1b3c62d3, 
               32'sh1b3af6ec, 32'sh1b398b01, 32'sh1b381f12, 32'sh1b36b31e, 32'sh1b354727, 32'sh1b33db2b, 32'sh1b326f2b, 32'sh1b310326, 
               32'sh1b2f971e, 32'sh1b2e2b11, 32'sh1b2cbf00, 32'sh1b2b52eb, 32'sh1b29e6d2, 32'sh1b287ab4, 32'sh1b270e93, 32'sh1b25a26d, 
               32'sh1b243643, 32'sh1b22ca15, 32'sh1b215de2, 32'sh1b1ff1ac, 32'sh1b1e8571, 32'sh1b1d1932, 32'sh1b1bacef, 32'sh1b1a40a7, 
               32'sh1b18d45c, 32'sh1b17680c, 32'sh1b15fbb8, 32'sh1b148f60, 32'sh1b132304, 32'sh1b11b6a4, 32'sh1b104a3f, 32'sh1b0eddd7, 
               32'sh1b0d716a, 32'sh1b0c04f9, 32'sh1b0a9883, 32'sh1b092c0a, 32'sh1b07bf8c, 32'sh1b06530b, 32'sh1b04e685, 32'sh1b0379fb, 
               32'sh1b020d6c, 32'sh1b00a0da, 32'sh1aff3444, 32'sh1afdc7a9, 32'sh1afc5b0a, 32'sh1afaee67, 32'sh1af981c0, 32'sh1af81514, 
               32'sh1af6a865, 32'sh1af53bb1, 32'sh1af3cef9, 32'sh1af2623d, 32'sh1af0f57d, 32'sh1aef88b9, 32'sh1aee1bf0, 32'sh1aecaf24, 
               32'sh1aeb4253, 32'sh1ae9d57e, 32'sh1ae868a5, 32'sh1ae6fbc8, 32'sh1ae58ee6, 32'sh1ae42201, 32'sh1ae2b517, 32'sh1ae14829, 
               32'sh1adfdb37, 32'sh1ade6e41, 32'sh1add0147, 32'sh1adb9448, 32'sh1ada2746, 32'sh1ad8ba3f, 32'sh1ad74d34, 32'sh1ad5e025, 
               32'sh1ad47312, 32'sh1ad305fb, 32'sh1ad198e0, 32'sh1ad02bc0, 32'sh1acebe9d, 32'sh1acd5175, 32'sh1acbe449, 32'sh1aca7719, 
               32'sh1ac909e5, 32'sh1ac79cac, 32'sh1ac62f70, 32'sh1ac4c22f, 32'sh1ac354eb, 32'sh1ac1e7a2, 32'sh1ac07a55, 32'sh1abf0d04, 
               32'sh1abd9faf, 32'sh1abc3255, 32'sh1abac4f8, 32'sh1ab95796, 32'sh1ab7ea31, 32'sh1ab67cc7, 32'sh1ab50f59, 32'sh1ab3a1e7, 
               32'sh1ab23471, 32'sh1ab0c6f7, 32'sh1aaf5978, 32'sh1aadebf6, 32'sh1aac7e6f, 32'sh1aab10e4, 32'sh1aa9a355, 32'sh1aa835c2, 
               32'sh1aa6c82b, 32'sh1aa55a90, 32'sh1aa3ecf1, 32'sh1aa27f4e, 32'sh1aa111a6, 32'sh1a9fa3fa, 32'sh1a9e364b, 32'sh1a9cc897, 
               32'sh1a9b5adf, 32'sh1a99ed23, 32'sh1a987f63, 32'sh1a97119f, 32'sh1a95a3d6, 32'sh1a94360a, 32'sh1a92c839, 32'sh1a915a65, 
               32'sh1a8fec8c, 32'sh1a8e7eaf, 32'sh1a8d10ce, 32'sh1a8ba2e9, 32'sh1a8a3500, 32'sh1a88c713, 32'sh1a875922, 32'sh1a85eb2c, 
               32'sh1a847d33, 32'sh1a830f35, 32'sh1a81a134, 32'sh1a80332e, 32'sh1a7ec524, 32'sh1a7d5716, 32'sh1a7be904, 32'sh1a7a7aee, 
               32'sh1a790cd4, 32'sh1a779eb6, 32'sh1a763093, 32'sh1a74c26d, 32'sh1a735442, 32'sh1a71e614, 32'sh1a7077e1, 32'sh1a6f09aa, 
               32'sh1a6d9b70, 32'sh1a6c2d31, 32'sh1a6abeee, 32'sh1a6950a7, 32'sh1a67e25c, 32'sh1a66740d, 32'sh1a6505b9, 32'sh1a639762, 
               32'sh1a622907, 32'sh1a60baa7, 32'sh1a5f4c44, 32'sh1a5ddddc, 32'sh1a5c6f70, 32'sh1a5b0101, 32'sh1a59928d, 32'sh1a582415, 
               32'sh1a56b599, 32'sh1a554719, 32'sh1a53d895, 32'sh1a526a0d, 32'sh1a50fb81, 32'sh1a4f8cf1, 32'sh1a4e1e5d, 32'sh1a4cafc4, 
               32'sh1a4b4128, 32'sh1a49d287, 32'sh1a4863e3, 32'sh1a46f53a, 32'sh1a45868e, 32'sh1a4417dd, 32'sh1a42a929, 32'sh1a413a70, 
               32'sh1a3fcbb3, 32'sh1a3e5cf2, 32'sh1a3cee2d, 32'sh1a3b7f64, 32'sh1a3a1097, 32'sh1a38a1c6, 32'sh1a3732f1, 32'sh1a35c418, 
               32'sh1a34553b, 32'sh1a32e65a, 32'sh1a317775, 32'sh1a30088b, 32'sh1a2e999e, 32'sh1a2d2aad, 32'sh1a2bbbb7, 32'sh1a2a4cbe, 
               32'sh1a28ddc0, 32'sh1a276ebf, 32'sh1a25ffb9, 32'sh1a2490b0, 32'sh1a2321a2, 32'sh1a21b291, 32'sh1a20437b, 32'sh1a1ed461, 
               32'sh1a1d6544, 32'sh1a1bf622, 32'sh1a1a86fc, 32'sh1a1917d2, 32'sh1a17a8a5, 32'sh1a163973, 32'sh1a14ca3d, 32'sh1a135b03, 
               32'sh1a11ebc5, 32'sh1a107c83, 32'sh1a0f0d3d, 32'sh1a0d9df3, 32'sh1a0c2ea5, 32'sh1a0abf53, 32'sh1a094ffd, 32'sh1a07e0a3, 
               32'sh1a067145, 32'sh1a0501e3, 32'sh1a03927d, 32'sh1a022313, 32'sh1a00b3a5, 32'sh19ff4433, 32'sh19fdd4bd, 32'sh19fc6543, 
               32'sh19faf5c5, 32'sh19f98643, 32'sh19f816bc, 32'sh19f6a732, 32'sh19f537a4, 32'sh19f3c812, 32'sh19f2587c, 32'sh19f0e8e2, 
               32'sh19ef7944, 32'sh19ee09a2, 32'sh19ec99fb, 32'sh19eb2a51, 32'sh19e9baa3, 32'sh19e84af1, 32'sh19e6db3b, 32'sh19e56b81, 
               32'sh19e3fbc3, 32'sh19e28c01, 32'sh19e11c3a, 32'sh19dfac70, 32'sh19de3ca2, 32'sh19dcccd0, 32'sh19db5cfa, 32'sh19d9ed20, 
               32'sh19d87d42, 32'sh19d70d60, 32'sh19d59d7a, 32'sh19d42d90, 32'sh19d2bda2, 32'sh19d14db0, 32'sh19cfddba, 32'sh19ce6dc0, 
               32'sh19ccfdc2, 32'sh19cb8dc0, 32'sh19ca1dbb, 32'sh19c8adb1, 32'sh19c73da3, 32'sh19c5cd91, 32'sh19c45d7b, 32'sh19c2ed62, 
               32'sh19c17d44, 32'sh19c00d22, 32'sh19be9cfd, 32'sh19bd2cd3, 32'sh19bbbca6, 32'sh19ba4c74, 32'sh19b8dc3e, 32'sh19b76c05, 
               32'sh19b5fbc8, 32'sh19b48b86, 32'sh19b31b41, 32'sh19b1aaf7, 32'sh19b03aaa, 32'sh19aeca59, 32'sh19ad5a04, 32'sh19abe9aa, 
               32'sh19aa794d, 32'sh19a908ec, 32'sh19a79887, 32'sh19a6281e, 32'sh19a4b7b1, 32'sh19a34740, 32'sh19a1d6cb, 32'sh19a06652, 
               32'sh199ef5d6, 32'sh199d8555, 32'sh199c14d0, 32'sh199aa448, 32'sh199933bb, 32'sh1997c32b, 32'sh19965296, 32'sh1994e1fe, 
               32'sh19937161, 32'sh199200c1, 32'sh1990901d, 32'sh198f1f74, 32'sh198daec8, 32'sh198c3e18, 32'sh198acd64, 32'sh19895cac, 
               32'sh1987ebf0, 32'sh19867b31, 32'sh19850a6d, 32'sh198399a5, 32'sh198228d9, 32'sh1980b80a, 32'sh197f4736, 32'sh197dd65f, 
               32'sh197c6584, 32'sh197af4a4, 32'sh197983c1, 32'sh197812da, 32'sh1976a1ef, 32'sh19753100, 32'sh1973c00d, 32'sh19724f16, 
               32'sh1970de1b, 32'sh196f6d1c, 32'sh196dfc1a, 32'sh196c8b13, 32'sh196b1a09, 32'sh1969a8fa, 32'sh196837e8, 32'sh1966c6d2, 
               32'sh196555b8, 32'sh1963e49a, 32'sh19627378, 32'sh19610252, 32'sh195f9128, 32'sh195e1ffa, 32'sh195caec9, 32'sh195b3d93, 
               32'sh1959cc5a, 32'sh19585b1c, 32'sh1956e9db, 32'sh19557896, 32'sh1954074d, 32'sh19529600, 32'sh195124af, 32'sh194fb35a, 
               32'sh194e4201, 32'sh194cd0a5, 32'sh194b5f44, 32'sh1949ede0, 32'sh19487c77, 32'sh19470b0b, 32'sh1945999b, 32'sh19442827, 
               32'sh1942b6af, 32'sh19414533, 32'sh193fd3b4, 32'sh193e6230, 32'sh193cf0a9, 32'sh193b7f1d, 32'sh193a0d8e, 32'sh19389bfb, 
               32'sh19372a64, 32'sh1935b8c9, 32'sh1934472a, 32'sh1932d587, 32'sh193163e1, 32'sh192ff236, 32'sh192e8088, 32'sh192d0ed6, 
               32'sh192b9d1f, 32'sh192a2b65, 32'sh1928b9a8, 32'sh192747e6, 32'sh1925d620, 32'sh19246457, 32'sh1922f289, 32'sh192180b8, 
               32'sh19200ee3, 32'sh191e9d0a, 32'sh191d2b2d, 32'sh191bb94c, 32'sh191a4767, 32'sh1918d57f, 32'sh19176393, 32'sh1915f1a2, 
               32'sh19147fae, 32'sh19130db6, 32'sh19119bba, 32'sh191029bb, 32'sh190eb7b7, 32'sh190d45af, 32'sh190bd3a4, 32'sh190a6195, 
               32'sh1908ef82, 32'sh19077d6b, 32'sh19060b50, 32'sh19049932, 32'sh1903270f, 32'sh1901b4e9, 32'sh190042bf, 32'sh18fed091, 
               32'sh18fd5e5f, 32'sh18fbec29, 32'sh18fa79ef, 32'sh18f907b2, 32'sh18f79571, 32'sh18f6232b, 32'sh18f4b0e2, 32'sh18f33e95, 
               32'sh18f1cc45, 32'sh18f059f0, 32'sh18eee798, 32'sh18ed753c, 32'sh18ec02db, 32'sh18ea9077, 32'sh18e91e10, 32'sh18e7aba4, 
               32'sh18e63935, 32'sh18e4c6c1, 32'sh18e3544a, 32'sh18e1e1cf, 32'sh18e06f50, 32'sh18defcce, 32'sh18dd8a47, 32'sh18dc17bd, 
               32'sh18daa52f, 32'sh18d9329d, 32'sh18d7c007, 32'sh18d64d6d, 32'sh18d4dad0, 32'sh18d3682f, 32'sh18d1f589, 32'sh18d082e0, 
               32'sh18cf1034, 32'sh18cd9d83, 32'sh18cc2acf, 32'sh18cab816, 32'sh18c9455a, 32'sh18c7d29a, 32'sh18c65fd7, 32'sh18c4ed0f, 
               32'sh18c37a44, 32'sh18c20774, 32'sh18c094a1, 32'sh18bf21cb, 32'sh18bdaef0, 32'sh18bc3c11, 32'sh18bac92f, 32'sh18b95649, 
               32'sh18b7e35f, 32'sh18b67071, 32'sh18b4fd80, 32'sh18b38a8b, 32'sh18b21791, 32'sh18b0a495, 32'sh18af3194, 32'sh18adbe8f, 
               32'sh18ac4b87, 32'sh18aad87b, 32'sh18a9656b, 32'sh18a7f257, 32'sh18a67f3f, 32'sh18a50c24, 32'sh18a39905, 32'sh18a225e2, 
               32'sh18a0b2bb, 32'sh189f3f90, 32'sh189dcc62, 32'sh189c5930, 32'sh189ae5fa, 32'sh189972c0, 32'sh1897ff82, 32'sh18968c41, 
               32'sh189518fc, 32'sh1893a5b3, 32'sh18923266, 32'sh1890bf16, 32'sh188f4bc2, 32'sh188dd869, 32'sh188c650e, 32'sh188af1ae, 
               32'sh18897e4a, 32'sh18880ae3, 32'sh18869778, 32'sh18852409, 32'sh1883b097, 32'sh18823d20, 32'sh1880c9a6, 32'sh187f5628, 
               32'sh187de2a7, 32'sh187c6f21, 32'sh187afb98, 32'sh1879880b, 32'sh1878147a, 32'sh1876a0e6, 32'sh18752d4d, 32'sh1873b9b1, 
               32'sh18724611, 32'sh1870d26e, 32'sh186f5ec6, 32'sh186deb1b, 32'sh186c776c, 32'sh186b03b9, 32'sh18699003, 32'sh18681c48, 
               32'sh1866a88a, 32'sh186534c9, 32'sh1863c103, 32'sh18624d3a, 32'sh1860d96d, 32'sh185f659c, 32'sh185df1c7, 32'sh185c7def, 
               32'sh185b0a13, 32'sh18599633, 32'sh1858224f, 32'sh1856ae68, 32'sh18553a7d, 32'sh1853c68e, 32'sh1852529b, 32'sh1850dea5, 
               32'sh184f6aab, 32'sh184df6ad, 32'sh184c82ab, 32'sh184b0ea6, 32'sh18499a9d, 32'sh18482690, 32'sh1846b280, 32'sh18453e6b, 
               32'sh1843ca53, 32'sh18425637, 32'sh1840e218, 32'sh183f6df4, 32'sh183df9cd, 32'sh183c85a2, 32'sh183b1174, 32'sh18399d42, 
               32'sh1838290c, 32'sh1836b4d2, 32'sh18354094, 32'sh1833cc53, 32'sh1832580e, 32'sh1830e3c6, 32'sh182f6f79, 32'sh182dfb29, 
               32'sh182c86d5, 32'sh182b127e, 32'sh18299e22, 32'sh182829c3, 32'sh1826b561, 32'sh182540fa, 32'sh1823cc90, 32'sh18225822, 
               32'sh1820e3b0, 32'sh181f6f3b, 32'sh181dfac2, 32'sh181c8645, 32'sh181b11c4, 32'sh18199d40, 32'sh181828b8, 32'sh1816b42d, 
               32'sh18153f9d, 32'sh1813cb0a, 32'sh18125673, 32'sh1810e1d9, 32'sh180f6d3a, 32'sh180df898, 32'sh180c83f3, 32'sh180b0f49, 
               32'sh18099a9c, 32'sh180825ec, 32'sh1806b137, 32'sh18053c7f, 32'sh1803c7c3, 32'sh18025303, 32'sh1800de40, 32'sh17ff6979, 
               32'sh17fdf4ae, 32'sh17fc7fe0, 32'sh17fb0b0e, 32'sh17f99638, 32'sh17f8215e, 32'sh17f6ac81, 32'sh17f537a0, 32'sh17f3c2bc, 
               32'sh17f24dd3, 32'sh17f0d8e7, 32'sh17ef63f8, 32'sh17edef04, 32'sh17ec7a0d, 32'sh17eb0513, 32'sh17e99014, 32'sh17e81b12, 
               32'sh17e6a60c, 32'sh17e53103, 32'sh17e3bbf6, 32'sh17e246e5, 32'sh17e0d1d0, 32'sh17df5cb8, 32'sh17dde79c, 32'sh17dc727c, 
               32'sh17dafd59, 32'sh17d98832, 32'sh17d81308, 32'sh17d69dd9, 32'sh17d528a7, 32'sh17d3b372, 32'sh17d23e38, 32'sh17d0c8fb, 
               32'sh17cf53bb, 32'sh17cdde76, 32'sh17cc692e, 32'sh17caf3e3, 32'sh17c97e93, 32'sh17c80940, 32'sh17c693ea, 32'sh17c51e8f, 
               32'sh17c3a931, 32'sh17c233cf, 32'sh17c0be6a, 32'sh17bf4901, 32'sh17bdd394, 32'sh17bc5e24, 32'sh17bae8b0, 32'sh17b97338, 
               32'sh17b7fdbd, 32'sh17b6883e, 32'sh17b512bb, 32'sh17b39d35, 32'sh17b227ab, 32'sh17b0b21e, 32'sh17af3c8c, 32'sh17adc6f7, 
               32'sh17ac515f, 32'sh17aadbc3, 32'sh17a96623, 32'sh17a7f07f, 32'sh17a67ad8, 32'sh17a5052d, 32'sh17a38f7f, 32'sh17a219cd, 
               32'sh17a0a417, 32'sh179f2e5e, 32'sh179db8a1, 32'sh179c42e0, 32'sh179acd1c, 32'sh17995754, 32'sh1797e188, 32'sh17966bb9, 
               32'sh1794f5e6, 32'sh17938010, 32'sh17920a35, 32'sh17909458, 32'sh178f1e76, 32'sh178da891, 32'sh178c32a9, 32'sh178abcbc, 
               32'sh178946cc, 32'sh1787d0d9, 32'sh17865ae2, 32'sh1784e4e7, 32'sh17836ee8, 32'sh1781f8e6, 32'sh178082e1, 32'sh177f0cd7, 
               32'sh177d96ca, 32'sh177c20ba, 32'sh177aaaa6, 32'sh1779348e, 32'sh1777be72, 32'sh17764853, 32'sh1774d231, 32'sh17735c0a, 
               32'sh1771e5e0, 32'sh17706fb3, 32'sh176ef982, 32'sh176d834d, 32'sh176c0d15, 32'sh176a96d9, 32'sh17692099, 32'sh1767aa56, 
               32'sh1766340f, 32'sh1764bdc5, 32'sh17634777, 32'sh1761d125, 32'sh17605ad0, 32'sh175ee477, 32'sh175d6e1b, 32'sh175bf7bb, 
               32'sh175a8157, 32'sh17590af0, 32'sh17579485, 32'sh17561e16, 32'sh1754a7a4, 32'sh1753312f, 32'sh1751bab5, 32'sh17504439, 
               32'sh174ecdb8, 32'sh174d5734, 32'sh174be0ad, 32'sh174a6a21, 32'sh1748f393, 32'sh17477d00, 32'sh1746066a, 32'sh17448fd1, 
               32'sh17431933, 32'sh1741a293, 32'sh17402bee, 32'sh173eb546, 32'sh173d3e9b, 32'sh173bc7ec, 32'sh173a5139, 32'sh1738da83, 
               32'sh173763c9, 32'sh1735ed0c, 32'sh1734764b, 32'sh1732ff86, 32'sh173188be, 32'sh173011f2, 32'sh172e9b23, 32'sh172d2450, 
               32'sh172bad7a, 32'sh172a36a0, 32'sh1728bfc2, 32'sh172748e1, 32'sh1725d1fc, 32'sh17245b14, 32'sh1722e428, 32'sh17216d39, 
               32'sh171ff646, 32'sh171e7f4f, 32'sh171d0855, 32'sh171b9157, 32'sh171a1a56, 32'sh1718a351, 32'sh17172c49, 32'sh1715b53d, 
               32'sh17143e2d, 32'sh1712c71a, 32'sh17115003, 32'sh170fd8e9, 32'sh170e61cc, 32'sh170ceaaa, 32'sh170b7385, 32'sh1709fc5d, 
               32'sh17088531, 32'sh17070e01, 32'sh170596ce, 32'sh17041f98, 32'sh1702a85e, 32'sh17013120, 32'sh16ffb9df, 32'sh16fe429a, 
               32'sh16fccb51, 32'sh16fb5406, 32'sh16f9dcb6, 32'sh16f86563, 32'sh16f6ee0d, 32'sh16f576b3, 32'sh16f3ff55, 32'sh16f287f4, 
               32'sh16f1108f, 32'sh16ef9927, 32'sh16ee21bb, 32'sh16ecaa4c, 32'sh16eb32d9, 32'sh16e9bb63, 32'sh16e843e9, 32'sh16e6cc6b, 
               32'sh16e554ea, 32'sh16e3dd66, 32'sh16e265de, 32'sh16e0ee52, 32'sh16df76c3, 32'sh16ddff31, 32'sh16dc879a, 32'sh16db1001, 
               32'sh16d99864, 32'sh16d820c3, 32'sh16d6a91f, 32'sh16d53177, 32'sh16d3b9cc, 32'sh16d2421d, 32'sh16d0ca6a, 32'sh16cf52b5, 
               32'sh16cddafb, 32'sh16cc633e, 32'sh16caeb7e, 32'sh16c973ba, 32'sh16c7fbf3, 32'sh16c68428, 32'sh16c50c59, 32'sh16c39487, 
               32'sh16c21cb2, 32'sh16c0a4d9, 32'sh16bf2cfc, 32'sh16bdb51c, 32'sh16bc3d39, 32'sh16bac552, 32'sh16b94d67, 32'sh16b7d579, 
               32'sh16b65d88, 32'sh16b4e593, 32'sh16b36d9a, 32'sh16b1f59e, 32'sh16b07d9f, 32'sh16af059c, 32'sh16ad8d95, 32'sh16ac158b, 
               32'sh16aa9d7e, 32'sh16a9256d, 32'sh16a7ad58, 32'sh16a63540, 32'sh16a4bd25, 32'sh16a34506, 32'sh16a1cce3, 32'sh16a054bd, 
               32'sh169edc94, 32'sh169d6467, 32'sh169bec37, 32'sh169a7403, 32'sh1698fbcb, 32'sh16978390, 32'sh16960b52, 32'sh16949310, 
               32'sh16931acb, 32'sh1691a282, 32'sh16902a36, 32'sh168eb1e6, 32'sh168d3993, 32'sh168bc13c, 32'sh168a48e2, 32'sh1688d084, 
               32'sh16875823, 32'sh1685dfbe, 32'sh16846756, 32'sh1682eeeb, 32'sh1681767c, 32'sh167ffe09, 32'sh167e8593, 32'sh167d0d1a, 
               32'sh167b949d, 32'sh167a1c1c, 32'sh1678a398, 32'sh16772b11, 32'sh1675b286, 32'sh167439f8, 32'sh1672c166, 32'sh167148d1, 
               32'sh166fd039, 32'sh166e579c, 32'sh166cdefd, 32'sh166b665a, 32'sh1669edb3, 32'sh16687509, 32'sh1666fc5c, 32'sh166583ab, 
               32'sh16640af7, 32'sh1662923f, 32'sh16611984, 32'sh165fa0c5, 32'sh165e2803, 32'sh165caf3e, 32'sh165b3675, 32'sh1659bda8, 
               32'sh165844d8, 32'sh1656cc05, 32'sh1655532e, 32'sh1653da54, 32'sh16526176, 32'sh1650e895, 32'sh164f6fb1, 32'sh164df6c9, 
               32'sh164c7ddd, 32'sh164b04ee, 32'sh16498bfc, 32'sh16481306, 32'sh16469a0d, 32'sh16452111, 32'sh1643a810, 32'sh16422f0d, 
               32'sh1640b606, 32'sh163f3cfc, 32'sh163dc3ee, 32'sh163c4add, 32'sh163ad1c8, 32'sh163958b0, 32'sh1637df95, 32'sh16366676, 
               32'sh1634ed53, 32'sh1633742d, 32'sh1631fb04, 32'sh163081d8, 32'sh162f08a8, 32'sh162d8f74, 32'sh162c163d, 32'sh162a9d03, 
               32'sh162923c5, 32'sh1627aa84, 32'sh16263140, 32'sh1624b7f8, 32'sh16233eac, 32'sh1621c55d, 32'sh16204c0b, 32'sh161ed2b6, 
               32'sh161d595d, 32'sh161be000, 32'sh161a66a0, 32'sh1618ed3d, 32'sh161773d6, 32'sh1615fa6c, 32'sh161480ff, 32'sh1613078e, 
               32'sh16118e1a, 32'sh161014a2, 32'sh160e9b27, 32'sh160d21a8, 32'sh160ba826, 32'sh160a2ea1, 32'sh1608b518, 32'sh16073b8c, 
               32'sh1605c1fd, 32'sh1604486a, 32'sh1602ced4, 32'sh1601553a, 32'sh15ffdb9d, 32'sh15fe61fc, 32'sh15fce859, 32'sh15fb6eb1, 
               32'sh15f9f507, 32'sh15f87b59, 32'sh15f701a7, 32'sh15f587f2, 32'sh15f40e3a, 32'sh15f2947f, 32'sh15f11ac0, 32'sh15efa0fd, 
               32'sh15ee2738, 32'sh15ecad6f, 32'sh15eb33a2, 32'sh15e9b9d2, 32'sh15e83fff, 32'sh15e6c628, 32'sh15e54c4e, 32'sh15e3d271, 
               32'sh15e25890, 32'sh15e0deac, 32'sh15df64c5, 32'sh15ddeada, 32'sh15dc70eb, 32'sh15daf6fa, 32'sh15d97d05, 32'sh15d8030c, 
               32'sh15d68911, 32'sh15d50f12, 32'sh15d3950f, 32'sh15d21b09, 32'sh15d0a100, 32'sh15cf26f4, 32'sh15cdace4, 32'sh15cc32d0, 
               32'sh15cab8ba, 32'sh15c93ea0, 32'sh15c7c482, 32'sh15c64a62, 32'sh15c4d03e, 32'sh15c35616, 32'sh15c1dbeb, 32'sh15c061bd, 
               32'sh15bee78c, 32'sh15bd6d57, 32'sh15bbf31f, 32'sh15ba78e3, 32'sh15b8fea4, 32'sh15b78462, 32'sh15b60a1c, 32'sh15b48fd3, 
               32'sh15b31587, 32'sh15b19b37, 32'sh15b020e4, 32'sh15aea68e, 32'sh15ad2c34, 32'sh15abb1d7, 32'sh15aa3777, 32'sh15a8bd13, 
               32'sh15a742ac, 32'sh15a5c842, 32'sh15a44dd4, 32'sh15a2d363, 32'sh15a158ee, 32'sh159fde77, 32'sh159e63fc, 32'sh159ce97d, 
               32'sh159b6efb, 32'sh1599f476, 32'sh159879ee, 32'sh1596ff62, 32'sh159584d3, 32'sh15940a41, 32'sh15928fab, 32'sh15911512, 
               32'sh158f9a76, 32'sh158e1fd6, 32'sh158ca533, 32'sh158b2a8d, 32'sh1589afe3, 32'sh15883536, 32'sh1586ba86, 32'sh15853fd2, 
               32'sh1583c51b, 32'sh15824a61, 32'sh1580cfa3, 32'sh157f54e2, 32'sh157dda1e, 32'sh157c5f57, 32'sh157ae48c, 32'sh157969be, 
               32'sh1577eeec, 32'sh15767417, 32'sh1574f93f, 32'sh15737e64, 32'sh15720385, 32'sh157088a3, 32'sh156f0dbe, 32'sh156d92d5, 
               32'sh156c17e9, 32'sh156a9cfa, 32'sh15692207, 32'sh1567a712, 32'sh15662c18, 32'sh1564b11c, 32'sh1563361c, 32'sh1561bb19, 
               32'sh15604013, 32'sh155ec509, 32'sh155d49fc, 32'sh155bceec, 32'sh155a53d9, 32'sh1558d8c2, 32'sh15575da8, 32'sh1555e28a, 
               32'sh1554676a, 32'sh1552ec46, 32'sh1551711e, 32'sh154ff5f4, 32'sh154e7ac6, 32'sh154cff95, 32'sh154b8461, 32'sh154a0929, 
               32'sh15488dee, 32'sh154712b0, 32'sh1545976e, 32'sh15441c29, 32'sh1542a0e1, 32'sh15412596, 32'sh153faa47, 32'sh153e2ef5, 
               32'sh153cb3a0, 32'sh153b3848, 32'sh1539bcec, 32'sh1538418d, 32'sh1536c62b, 32'sh15354ac5, 32'sh1533cf5c, 32'sh153253f0, 
               32'sh1530d881, 32'sh152f5d0e, 32'sh152de198, 32'sh152c661f, 32'sh152aeaa3, 32'sh15296f23, 32'sh1527f3a0, 32'sh1526781a, 
               32'sh1524fc90, 32'sh15238103, 32'sh15220573, 32'sh152089e0, 32'sh151f0e4a, 32'sh151d92b0, 32'sh151c1713, 32'sh151a9b72, 
               32'sh15191fcf, 32'sh1517a428, 32'sh1516287e, 32'sh1514acd1, 32'sh15133120, 32'sh1511b56c, 32'sh151039b5, 32'sh150ebdfb, 
               32'sh150d423d, 32'sh150bc67d, 32'sh150a4ab9, 32'sh1508cef1, 32'sh15075327, 32'sh1505d759, 32'sh15045b88, 32'sh1502dfb4, 
               32'sh150163dc, 32'sh14ffe801, 32'sh14fe6c23, 32'sh14fcf042, 32'sh14fb745e, 32'sh14f9f876, 32'sh14f87c8b, 32'sh14f7009d, 
               32'sh14f584ac, 32'sh14f408b7, 32'sh14f28cbf, 32'sh14f110c4, 32'sh14ef94c6, 32'sh14ee18c4, 32'sh14ec9cbf, 32'sh14eb20b7, 
               32'sh14e9a4ac, 32'sh14e8289e, 32'sh14e6ac8c, 32'sh14e53077, 32'sh14e3b45f, 32'sh14e23844, 32'sh14e0bc25, 32'sh14df4003, 
               32'sh14ddc3de, 32'sh14dc47b6, 32'sh14dacb8b, 32'sh14d94f5c, 32'sh14d7d32a, 32'sh14d656f5, 32'sh14d4dabd, 32'sh14d35e81, 
               32'sh14d1e242, 32'sh14d06601, 32'sh14cee9bb, 32'sh14cd6d73, 32'sh14cbf127, 32'sh14ca74d9, 32'sh14c8f887, 32'sh14c77c32, 
               32'sh14c5ffd9, 32'sh14c4837e, 32'sh14c3071f, 32'sh14c18abd, 32'sh14c00e58, 32'sh14be91ef, 32'sh14bd1584, 32'sh14bb9915, 
               32'sh14ba1ca3, 32'sh14b8a02e, 32'sh14b723b5, 32'sh14b5a73a, 32'sh14b42abb, 32'sh14b2ae39, 32'sh14b131b4, 32'sh14afb52c, 
               32'sh14ae38a0, 32'sh14acbc11, 32'sh14ab3f7f, 32'sh14a9c2ea, 32'sh14a84652, 32'sh14a6c9b7, 32'sh14a54d18, 32'sh14a3d076, 
               32'sh14a253d1, 32'sh14a0d729, 32'sh149f5a7e, 32'sh149dddcf, 32'sh149c611d, 32'sh149ae468, 32'sh149967b0, 32'sh1497eaf5, 
               32'sh14966e36, 32'sh1494f175, 32'sh149374b0, 32'sh1491f7e8, 32'sh14907b1d, 32'sh148efe4f, 32'sh148d817d, 32'sh148c04a9, 
               32'sh148a87d1, 32'sh14890af6, 32'sh14878e18, 32'sh14861136, 32'sh14849452, 32'sh1483176a, 32'sh14819a7f, 32'sh14801d91, 
               32'sh147ea0a0, 32'sh147d23ac, 32'sh147ba6b4, 32'sh147a29ba, 32'sh1478acbc, 32'sh14772fbb, 32'sh1475b2b7, 32'sh147435b0, 
               32'sh1472b8a5, 32'sh14713b98, 32'sh146fbe87, 32'sh146e4173, 32'sh146cc45c, 32'sh146b4742, 32'sh1469ca25, 32'sh14684d04, 
               32'sh1466cfe1, 32'sh146552ba, 32'sh1463d590, 32'sh14625863, 32'sh1460db33, 32'sh145f5e00, 32'sh145de0c9, 32'sh145c638f, 
               32'sh145ae653, 32'sh14596913, 32'sh1457ebd0, 32'sh14566e8a, 32'sh1454f140, 32'sh145373f4, 32'sh1451f6a4, 32'sh14507952, 
               32'sh144efbfc, 32'sh144d7ea3, 32'sh144c0147, 32'sh144a83e8, 32'sh14490685, 32'sh14478920, 32'sh14460bb7, 32'sh14448e4b, 
               32'sh144310dd, 32'sh1441936b, 32'sh144015f5, 32'sh143e987d, 32'sh143d1b02, 32'sh143b9d83, 32'sh143a2002, 32'sh1438a27d, 
               32'sh143724f5, 32'sh1435a76a, 32'sh143429dc, 32'sh1432ac4b, 32'sh14312eb7, 32'sh142fb11f, 32'sh142e3385, 32'sh142cb5e7, 
               32'sh142b3846, 32'sh1429baa3, 32'sh14283cfc, 32'sh1426bf52, 32'sh142541a4, 32'sh1423c3f4, 32'sh14224641, 32'sh1420c88a, 
               32'sh141f4ad1, 32'sh141dcd14, 32'sh141c4f54, 32'sh141ad191, 32'sh141953cb, 32'sh1417d602, 32'sh14165836, 32'sh1414da66, 
               32'sh14135c94, 32'sh1411debf, 32'sh141060e6, 32'sh140ee30a, 32'sh140d652c, 32'sh140be74a, 32'sh140a6965, 32'sh1408eb7d, 
               32'sh14076d91, 32'sh1405efa3, 32'sh140471b2, 32'sh1402f3be, 32'sh140175c6, 32'sh13fff7cb, 32'sh13fe79ce, 32'sh13fcfbcd, 
               32'sh13fb7dc9, 32'sh13f9ffc2, 32'sh13f881b8, 32'sh13f703ab, 32'sh13f5859b, 32'sh13f40788, 32'sh13f28972, 32'sh13f10b58, 
               32'sh13ef8d3c, 32'sh13ee0f1c, 32'sh13ec90fa, 32'sh13eb12d4, 32'sh13e994ab, 32'sh13e8167f, 32'sh13e69850, 32'sh13e51a1e, 
               32'sh13e39be9, 32'sh13e21db1, 32'sh13e09f76, 32'sh13df2138, 32'sh13dda2f7, 32'sh13dc24b2, 32'sh13daa66b, 32'sh13d92820, 
               32'sh13d7a9d3, 32'sh13d62b82, 32'sh13d4ad2f, 32'sh13d32ed8, 32'sh13d1b07e, 32'sh13d03221, 32'sh13ceb3c1, 32'sh13cd355e, 
               32'sh13cbb6f8, 32'sh13ca388f, 32'sh13c8ba23, 32'sh13c73bb4, 32'sh13c5bd42, 32'sh13c43ecd, 32'sh13c2c054, 32'sh13c141d9, 
               32'sh13bfc35b, 32'sh13be44d9, 32'sh13bcc655, 32'sh13bb47cd, 32'sh13b9c943, 32'sh13b84ab5, 32'sh13b6cc24, 32'sh13b54d91, 
               32'sh13b3cefa, 32'sh13b25060, 32'sh13b0d1c3, 32'sh13af5324, 32'sh13add481, 32'sh13ac55db, 32'sh13aad732, 32'sh13a95886, 
               32'sh13a7d9d7, 32'sh13a65b25, 32'sh13a4dc70, 32'sh13a35db8, 32'sh13a1defd, 32'sh13a0603e, 32'sh139ee17d, 32'sh139d62b9, 
               32'sh139be3f2, 32'sh139a6527, 32'sh1398e65a, 32'sh1397678a, 32'sh1395e8b7, 32'sh139469e0, 32'sh1392eb07, 32'sh13916c2a, 
               32'sh138fed4b, 32'sh138e6e69, 32'sh138cef83, 32'sh138b709b, 32'sh1389f1af, 32'sh138872c1, 32'sh1386f3cf, 32'sh138574db, 
               32'sh1383f5e3, 32'sh138276e9, 32'sh1380f7eb, 32'sh137f78eb, 32'sh137df9e7, 32'sh137c7ae1, 32'sh137afbd7, 32'sh13797ccb, 
               32'sh1377fdbb, 32'sh13767ea8, 32'sh1374ff93, 32'sh1373807a, 32'sh1372015f, 32'sh13708240, 32'sh136f031f, 32'sh136d83fa, 
               32'sh136c04d2, 32'sh136a85a8, 32'sh1369067a, 32'sh1367874a, 32'sh13660816, 32'sh136488e0, 32'sh136309a6, 32'sh13618a6a, 
               32'sh13600b2a, 32'sh135e8be8, 32'sh135d0ca2, 32'sh135b8d5a, 32'sh135a0e0e, 32'sh13588ec0, 32'sh13570f6f, 32'sh1355901a, 
               32'sh135410c3, 32'sh13529169, 32'sh1351120b, 32'sh134f92ab, 32'sh134e1348, 32'sh134c93e1, 32'sh134b1478, 32'sh1349950c, 
               32'sh1348159d, 32'sh1346962b, 32'sh134516b5, 32'sh1343973d, 32'sh134217c2, 32'sh13409844, 32'sh133f18c3, 32'sh133d993f, 
               32'sh133c19b8, 32'sh133a9a2e, 32'sh13391aa1, 32'sh13379b12, 32'sh13361b7f, 32'sh13349be9, 32'sh13331c50, 32'sh13319cb5, 
               32'sh13301d16, 32'sh132e9d74, 32'sh132d1dd0, 32'sh132b9e28, 32'sh132a1e7e, 32'sh13289ed0, 32'sh13271f20, 32'sh13259f6d, 
               32'sh13241fb6, 32'sh13229ffd, 32'sh13212041, 32'sh131fa082, 32'sh131e20c0, 32'sh131ca0fa, 32'sh131b2132, 32'sh1319a168, 
               32'sh1318219a, 32'sh1316a1c9, 32'sh131521f5, 32'sh1313a21e, 32'sh13122245, 32'sh1310a268, 32'sh130f2288, 32'sh130da2a6, 
               32'sh130c22c1, 32'sh130aa2d8, 32'sh130922ed, 32'sh1307a2ff, 32'sh1306230d, 32'sh1304a319, 32'sh13032322, 32'sh1301a328, 
               32'sh1300232c, 32'sh12fea32c, 32'sh12fd2329, 32'sh12fba323, 32'sh12fa231b, 32'sh12f8a30f, 32'sh12f72301, 32'sh12f5a2ef, 
               32'sh12f422db, 32'sh12f2a2c4, 32'sh12f122aa, 32'sh12efa28c, 32'sh12ee226c, 32'sh12eca24a, 32'sh12eb2224, 32'sh12e9a1fb, 
               32'sh12e821cf, 32'sh12e6a1a1, 32'sh12e5216f, 32'sh12e3a13b, 32'sh12e22103, 32'sh12e0a0c9, 32'sh12df208c, 32'sh12dda04c, 
               32'sh12dc2009, 32'sh12da9fc3, 32'sh12d91f7a, 32'sh12d79f2f, 32'sh12d61ee0, 32'sh12d49e8f, 32'sh12d31e3a, 32'sh12d19de3, 
               32'sh12d01d89, 32'sh12ce9d2c, 32'sh12cd1ccc, 32'sh12cb9c69, 32'sh12ca1c03, 32'sh12c89b9a, 32'sh12c71b2e, 32'sh12c59ac0, 
               32'sh12c41a4f, 32'sh12c299da, 32'sh12c11963, 32'sh12bf98e9, 32'sh12be186c, 32'sh12bc97ec, 32'sh12bb1769, 32'sh12b996e4, 
               32'sh12b8165b, 32'sh12b695d0, 32'sh12b51542, 32'sh12b394b0, 32'sh12b2141c, 32'sh12b09385, 32'sh12af12ec, 32'sh12ad924f, 
               32'sh12ac11af, 32'sh12aa910d, 32'sh12a91067, 32'sh12a78fbf, 32'sh12a60f14, 32'sh12a48e66, 32'sh12a30db5, 32'sh12a18d02, 
               32'sh12a00c4b, 32'sh129e8b91, 32'sh129d0ad5, 32'sh129b8a16, 32'sh129a0954, 32'sh1298888f, 32'sh129707c7, 32'sh129586fc, 
               32'sh1294062f, 32'sh1292855e, 32'sh1291048b, 32'sh128f83b5, 32'sh128e02dc, 32'sh128c8200, 32'sh128b0121, 32'sh12898040, 
               32'sh1287ff5b, 32'sh12867e74, 32'sh1284fd8a, 32'sh12837c9d, 32'sh1281fbad, 32'sh12807aba, 32'sh127ef9c5, 32'sh127d78cc, 
               32'sh127bf7d1, 32'sh127a76d3, 32'sh1278f5d2, 32'sh127774ce, 32'sh1275f3c7, 32'sh127472be, 32'sh1272f1b1, 32'sh127170a2, 
               32'sh126fef90, 32'sh126e6e7b, 32'sh126ced63, 32'sh126b6c49, 32'sh1269eb2b, 32'sh12686a0b, 32'sh1266e8e8, 32'sh126567c2, 
               32'sh1263e699, 32'sh1262656e, 32'sh1260e43f, 32'sh125f630e, 32'sh125de1da, 32'sh125c60a3, 32'sh125adf69, 32'sh12595e2c, 
               32'sh1257dced, 32'sh12565bab, 32'sh1254da66, 32'sh1253591e, 32'sh1251d7d3, 32'sh12505685, 32'sh124ed535, 32'sh124d53e2, 
               32'sh124bd28c, 32'sh124a5133, 32'sh1248cfd7, 32'sh12474e79, 32'sh1245cd17, 32'sh12444bb3, 32'sh1242ca4c, 32'sh124148e2, 
               32'sh123fc776, 32'sh123e4606, 32'sh123cc494, 32'sh123b431f, 32'sh1239c1a7, 32'sh1238402d, 32'sh1236beaf, 32'sh12353d2f, 
               32'sh1233bbac, 32'sh12323a26, 32'sh1230b89d, 32'sh122f3712, 32'sh122db583, 32'sh122c33f2, 32'sh122ab25e, 32'sh122930c8, 
               32'sh1227af2e, 32'sh12262d92, 32'sh1224abf3, 32'sh12232a51, 32'sh1221a8ac, 32'sh12202705, 32'sh121ea55a, 32'sh121d23ad, 
               32'sh121ba1fd, 32'sh121a204b, 32'sh12189e95, 32'sh12171cdd, 32'sh12159b22, 32'sh12141964, 32'sh121297a3, 32'sh121115e0, 
               32'sh120f941a, 32'sh120e1251, 32'sh120c9085, 32'sh120b0eb6, 32'sh12098ce5, 32'sh12080b11, 32'sh1206893a, 32'sh12050760, 
               32'sh12038584, 32'sh120203a5, 32'sh120081c3, 32'sh11feffde, 32'sh11fd7df6, 32'sh11fbfc0c, 32'sh11fa7a1f, 32'sh11f8f82f, 
               32'sh11f7763c, 32'sh11f5f447, 32'sh11f4724f, 32'sh11f2f054, 32'sh11f16e56, 32'sh11efec55, 32'sh11ee6a52, 32'sh11ece84c, 
               32'sh11eb6643, 32'sh11e9e438, 32'sh11e86229, 32'sh11e6e018, 32'sh11e55e04, 32'sh11e3dbee, 32'sh11e259d4, 32'sh11e0d7b8, 
               32'sh11df5599, 32'sh11ddd378, 32'sh11dc5153, 32'sh11dacf2c, 32'sh11d94d02, 32'sh11d7cad6, 32'sh11d648a6, 32'sh11d4c674, 
               32'sh11d3443f, 32'sh11d1c208, 32'sh11d03fcd, 32'sh11cebd90, 32'sh11cd3b50, 32'sh11cbb90e, 32'sh11ca36c8, 32'sh11c8b480, 
               32'sh11c73235, 32'sh11c5afe8, 32'sh11c42d97, 32'sh11c2ab44, 32'sh11c128ee, 32'sh11bfa696, 32'sh11be243a, 32'sh11bca1dc, 
               32'sh11bb1f7c, 32'sh11b99d18, 32'sh11b81ab2, 32'sh11b69849, 32'sh11b515dd, 32'sh11b3936f, 32'sh11b210fe, 32'sh11b08e8a, 
               32'sh11af0c13, 32'sh11ad899a, 32'sh11ac071e, 32'sh11aa849f, 32'sh11a9021d, 32'sh11a77f99, 32'sh11a5fd12, 32'sh11a47a88, 
               32'sh11a2f7fc, 32'sh11a1756d, 32'sh119ff2db, 32'sh119e7046, 32'sh119cedaf, 32'sh119b6b15, 32'sh1199e878, 32'sh119865d9, 
               32'sh1196e337, 32'sh11956092, 32'sh1193ddea, 32'sh11925b40, 32'sh1190d893, 32'sh118f55e3, 32'sh118dd331, 32'sh118c507c, 
               32'sh118acdc4, 32'sh11894b09, 32'sh1187c84c, 32'sh1186458c, 32'sh1184c2ca, 32'sh11834004, 32'sh1181bd3c, 32'sh11803a71, 
               32'sh117eb7a4, 32'sh117d34d4, 32'sh117bb201, 32'sh117a2f2c, 32'sh1178ac53, 32'sh11772978, 32'sh1175a69b, 32'sh117423ba, 
               32'sh1172a0d7, 32'sh11711df2, 32'sh116f9b09, 32'sh116e181e, 32'sh116c9531, 32'sh116b1240, 32'sh11698f4d, 32'sh11680c57, 
               32'sh1166895f, 32'sh11650663, 32'sh11638366, 32'sh11620065, 32'sh11607d62, 32'sh115efa5c, 32'sh115d7753, 32'sh115bf448, 
               32'sh115a713a, 32'sh1158ee2a, 32'sh11576b16, 32'sh1155e800, 32'sh115464e8, 32'sh1152e1cc, 32'sh11515eae, 32'sh114fdb8e, 
               32'sh114e586a, 32'sh114cd544, 32'sh114b521c, 32'sh1149cef0, 32'sh11484bc2, 32'sh1146c892, 32'sh1145455e, 32'sh1143c228, 
               32'sh11423ef0, 32'sh1140bbb4, 32'sh113f3876, 32'sh113db536, 32'sh113c31f3, 32'sh113aaead, 32'sh11392b64, 32'sh1137a819, 
               32'sh113624cb, 32'sh1134a17a, 32'sh11331e27, 32'sh11319ad1, 32'sh11301779, 32'sh112e941d, 32'sh112d10c0, 32'sh112b8d5f, 
               32'sh112a09fc, 32'sh11288696, 32'sh1127032e, 32'sh11257fc3, 32'sh1123fc55, 32'sh112278e5, 32'sh1120f572, 32'sh111f71fc, 
               32'sh111dee84, 32'sh111c6b09, 32'sh111ae78b, 32'sh1119640b, 32'sh1117e088, 32'sh11165d03, 32'sh1114d97b, 32'sh111355f0, 
               32'sh1111d263, 32'sh11104ed3, 32'sh110ecb40, 32'sh110d47ab, 32'sh110bc413, 32'sh110a4078, 32'sh1108bcdb, 32'sh1107393b, 
               32'sh1105b599, 32'sh110431f4, 32'sh1102ae4c, 32'sh11012aa2, 32'sh10ffa6f5, 32'sh10fe2346, 32'sh10fc9f94, 32'sh10fb1bdf, 
               32'sh10f99827, 32'sh10f8146d, 32'sh10f690b1, 32'sh10f50cf2, 32'sh10f38930, 32'sh10f2056b, 32'sh10f081a4, 32'sh10eefddb, 
               32'sh10ed7a0e, 32'sh10ebf63f, 32'sh10ea726e, 32'sh10e8ee9a, 32'sh10e76ac3, 32'sh10e5e6ea, 32'sh10e4630e, 32'sh10e2df2f, 
               32'sh10e15b4e, 32'sh10dfd76a, 32'sh10de5384, 32'sh10dccf9b, 32'sh10db4baf, 32'sh10d9c7c1, 32'sh10d843d1, 32'sh10d6bfdd, 
               32'sh10d53be7, 32'sh10d3b7ef, 32'sh10d233f4, 32'sh10d0aff6, 32'sh10cf2bf6, 32'sh10cda7f3, 32'sh10cc23ed, 32'sh10ca9fe5, 
               32'sh10c91bda, 32'sh10c797cd, 32'sh10c613bd, 32'sh10c48fab, 32'sh10c30b96, 32'sh10c1877e, 32'sh10c00364, 32'sh10be7f47, 
               32'sh10bcfb28, 32'sh10bb7706, 32'sh10b9f2e1, 32'sh10b86eba, 32'sh10b6ea90, 32'sh10b56664, 32'sh10b3e235, 32'sh10b25e04, 
               32'sh10b0d9d0, 32'sh10af5599, 32'sh10add160, 32'sh10ac4d24, 32'sh10aac8e6, 32'sh10a944a5, 32'sh10a7c062, 32'sh10a63c1c, 
               32'sh10a4b7d3, 32'sh10a33388, 32'sh10a1af3a, 32'sh10a02aea, 32'sh109ea697, 32'sh109d2242, 32'sh109b9dea, 32'sh109a1990, 
               32'sh10989532, 32'sh109710d3, 32'sh10958c71, 32'sh1094080c, 32'sh109283a5, 32'sh1090ff3b, 32'sh108f7ace, 32'sh108df65f, 
               32'sh108c71ee, 32'sh108aed7a, 32'sh10896903, 32'sh1087e48a, 32'sh1086600e, 32'sh1084db90, 32'sh1083570f, 32'sh1081d28c, 
               32'sh10804e06, 32'sh107ec97d, 32'sh107d44f2, 32'sh107bc065, 32'sh107a3bd5, 32'sh1078b742, 32'sh107732ad, 32'sh1075ae15, 
               32'sh1074297b, 32'sh1072a4de, 32'sh1071203f, 32'sh106f9b9d, 32'sh106e16f9, 32'sh106c9252, 32'sh106b0da8, 32'sh106988fc, 
               32'sh1068044e, 32'sh10667f9d, 32'sh1064fae9, 32'sh10637633, 32'sh1061f17b, 32'sh10606cbf, 32'sh105ee802, 32'sh105d6342, 
               32'sh105bde7f, 32'sh105a59ba, 32'sh1058d4f2, 32'sh10575027, 32'sh1055cb5b, 32'sh1054468b, 32'sh1052c1b9, 32'sh10513ce5, 
               32'sh104fb80e, 32'sh104e3335, 32'sh104cae59, 32'sh104b297a, 32'sh1049a49a, 32'sh10481fb6, 32'sh10469ad0, 32'sh104515e8, 
               32'sh104390fd, 32'sh10420c0f, 32'sh1040871f, 32'sh103f022d, 32'sh103d7d38, 32'sh103bf840, 32'sh103a7346, 32'sh1038ee4a, 
               32'sh1037694b, 32'sh1035e449, 32'sh10345f45, 32'sh1032da3f, 32'sh10315535, 32'sh102fd02a, 32'sh102e4b1c, 32'sh102cc60b, 
               32'sh102b40f8, 32'sh1029bbe3, 32'sh102836cb, 32'sh1026b1b0, 32'sh10252c94, 32'sh1023a774, 32'sh10222252, 32'sh10209d2e, 
               32'sh101f1807, 32'sh101d92dd, 32'sh101c0db1, 32'sh101a8883, 32'sh10190352, 32'sh10177e1f, 32'sh1015f8e9, 32'sh101473b1, 
               32'sh1012ee76, 32'sh10116939, 32'sh100fe3f9, 32'sh100e5eb7, 32'sh100cd972, 32'sh100b542b, 32'sh1009cee1, 32'sh10084995, 
               32'sh1006c446, 32'sh10053ef5, 32'sh1003b9a2, 32'sh1002344c, 32'sh1000aef3, 32'sh0fff2998, 32'sh0ffda43b, 32'sh0ffc1edb, 
               32'sh0ffa9979, 32'sh0ff91414, 32'sh0ff78ead, 32'sh0ff60943, 32'sh0ff483d7, 32'sh0ff2fe68, 32'sh0ff178f7, 32'sh0feff383, 
               32'sh0fee6e0d, 32'sh0fece895, 32'sh0feb631a, 32'sh0fe9dd9d, 32'sh0fe8581d, 32'sh0fe6d29a, 32'sh0fe54d16, 32'sh0fe3c78f, 
               32'sh0fe24205, 32'sh0fe0bc79, 32'sh0fdf36ea, 32'sh0fddb159, 32'sh0fdc2bc6, 32'sh0fdaa630, 32'sh0fd92098, 32'sh0fd79afd, 
               32'sh0fd6155f, 32'sh0fd48fc0, 32'sh0fd30a1e, 32'sh0fd18479, 32'sh0fcffed2, 32'sh0fce7929, 32'sh0fccf37d, 32'sh0fcb6dcf, 
               32'sh0fc9e81e, 32'sh0fc8626b, 32'sh0fc6dcb5, 32'sh0fc556fd, 32'sh0fc3d143, 32'sh0fc24b86, 32'sh0fc0c5c6, 32'sh0fbf4005, 
               32'sh0fbdba40, 32'sh0fbc347a, 32'sh0fbaaeb1, 32'sh0fb928e5, 32'sh0fb7a317, 32'sh0fb61d47, 32'sh0fb49774, 32'sh0fb3119f, 
               32'sh0fb18bc8, 32'sh0fb005ee, 32'sh0fae8011, 32'sh0facfa32, 32'sh0fab7451, 32'sh0fa9ee6d, 32'sh0fa86887, 32'sh0fa6e29f, 
               32'sh0fa55cb4, 32'sh0fa3d6c6, 32'sh0fa250d7, 32'sh0fa0cae5, 32'sh0f9f44f0, 32'sh0f9dbef9, 32'sh0f9c3900, 32'sh0f9ab304, 
               32'sh0f992d06, 32'sh0f97a705, 32'sh0f962102, 32'sh0f949afd, 32'sh0f9314f5, 32'sh0f918eeb, 32'sh0f9008de, 32'sh0f8e82cf, 
               32'sh0f8cfcbe, 32'sh0f8b76aa, 32'sh0f89f094, 32'sh0f886a7b, 32'sh0f86e460, 32'sh0f855e43, 32'sh0f83d823, 32'sh0f825201, 
               32'sh0f80cbdc, 32'sh0f7f45b5, 32'sh0f7dbf8c, 32'sh0f7c3960, 32'sh0f7ab332, 32'sh0f792d01, 32'sh0f77a6ce, 32'sh0f762099, 
               32'sh0f749a61, 32'sh0f731427, 32'sh0f718deb, 32'sh0f7007ac, 32'sh0f6e816b, 32'sh0f6cfb27, 32'sh0f6b74e1, 32'sh0f69ee99, 
               32'sh0f68684e, 32'sh0f66e201, 32'sh0f655bb2, 32'sh0f63d560, 32'sh0f624f0c, 32'sh0f60c8b5, 32'sh0f5f425c, 32'sh0f5dbc01, 
               32'sh0f5c35a3, 32'sh0f5aaf43, 32'sh0f5928e1, 32'sh0f57a27c, 32'sh0f561c15, 32'sh0f5495ab, 32'sh0f530f3f, 32'sh0f5188d1, 
               32'sh0f500260, 32'sh0f4e7bed, 32'sh0f4cf578, 32'sh0f4b6f00, 32'sh0f49e886, 32'sh0f48620a, 32'sh0f46db8b, 32'sh0f45550a, 
               32'sh0f43ce86, 32'sh0f424801, 32'sh0f40c178, 32'sh0f3f3aee, 32'sh0f3db461, 32'sh0f3c2dd2, 32'sh0f3aa740, 32'sh0f3920ac, 
               32'sh0f379a16, 32'sh0f36137d, 32'sh0f348ce2, 32'sh0f330645, 32'sh0f317fa5, 32'sh0f2ff903, 32'sh0f2e725f, 32'sh0f2cebb8, 
               32'sh0f2b650f, 32'sh0f29de64, 32'sh0f2857b6, 32'sh0f26d106, 32'sh0f254a53, 32'sh0f23c39f, 32'sh0f223ce8, 32'sh0f20b62e, 
               32'sh0f1f2f73, 32'sh0f1da8b4, 32'sh0f1c21f4, 32'sh0f1a9b31, 32'sh0f19146c, 32'sh0f178da5, 32'sh0f1606db, 32'sh0f14800f, 
               32'sh0f12f941, 32'sh0f117270, 32'sh0f0feb9d, 32'sh0f0e64c8, 32'sh0f0cddf0, 32'sh0f0b5716, 32'sh0f09d03a, 32'sh0f08495b, 
               32'sh0f06c27a, 32'sh0f053b97, 32'sh0f03b4b1, 32'sh0f022dca, 32'sh0f00a6df, 32'sh0eff1ff3, 32'sh0efd9904, 32'sh0efc1213, 
               32'sh0efa8b20, 32'sh0ef9042a, 32'sh0ef77d32, 32'sh0ef5f637, 32'sh0ef46f3b, 32'sh0ef2e83c, 32'sh0ef1613a, 32'sh0eefda37, 
               32'sh0eee5331, 32'sh0eeccc29, 32'sh0eeb451e, 32'sh0ee9be11, 32'sh0ee83702, 32'sh0ee6aff1, 32'sh0ee528dd, 32'sh0ee3a1c7, 
               32'sh0ee21aaf, 32'sh0ee09394, 32'sh0edf0c77, 32'sh0edd8558, 32'sh0edbfe37, 32'sh0eda7713, 32'sh0ed8efed, 32'sh0ed768c5, 
               32'sh0ed5e19a, 32'sh0ed45a6d, 32'sh0ed2d33e, 32'sh0ed14c0c, 32'sh0ecfc4d9, 32'sh0ece3da3, 32'sh0eccb66a, 32'sh0ecb2f30, 
               32'sh0ec9a7f3, 32'sh0ec820b3, 32'sh0ec69972, 32'sh0ec5122e, 32'sh0ec38ae8, 32'sh0ec203a0, 32'sh0ec07c55, 32'sh0ebef508, 
               32'sh0ebd6db9, 32'sh0ebbe668, 32'sh0eba5f14, 32'sh0eb8d7be, 32'sh0eb75066, 32'sh0eb5c90c, 32'sh0eb441af, 32'sh0eb2ba50, 
               32'sh0eb132ef, 32'sh0eafab8b, 32'sh0eae2425, 32'sh0eac9cbd, 32'sh0eab1553, 32'sh0ea98de6, 32'sh0ea80677, 32'sh0ea67f06, 
               32'sh0ea4f793, 32'sh0ea3701d, 32'sh0ea1e8a5, 32'sh0ea0612b, 32'sh0e9ed9af, 32'sh0e9d5230, 32'sh0e9bcaaf, 32'sh0e9a432c, 
               32'sh0e98bba7, 32'sh0e97341f, 32'sh0e95ac95, 32'sh0e942509, 32'sh0e929d7a, 32'sh0e9115ea, 32'sh0e8f8e57, 32'sh0e8e06c2, 
               32'sh0e8c7f2a, 32'sh0e8af791, 32'sh0e896ff5, 32'sh0e87e857, 32'sh0e8660b6, 32'sh0e84d914, 32'sh0e83516f, 32'sh0e81c9c8, 
               32'sh0e80421e, 32'sh0e7eba73, 32'sh0e7d32c5, 32'sh0e7bab15, 32'sh0e7a2363, 32'sh0e789bae, 32'sh0e7713f7, 32'sh0e758c3e, 
               32'sh0e740483, 32'sh0e727cc6, 32'sh0e70f506, 32'sh0e6f6d44, 32'sh0e6de580, 32'sh0e6c5dba, 32'sh0e6ad5f1, 32'sh0e694e27, 
               32'sh0e67c65a, 32'sh0e663e8a, 32'sh0e64b6b9, 32'sh0e632ee5, 32'sh0e61a70f, 32'sh0e601f37, 32'sh0e5e975d, 32'sh0e5d0f80, 
               32'sh0e5b87a2, 32'sh0e59ffc1, 32'sh0e5877de, 32'sh0e56eff8, 32'sh0e556811, 32'sh0e53e027, 32'sh0e52583b, 32'sh0e50d04d, 
               32'sh0e4f485c, 32'sh0e4dc069, 32'sh0e4c3875, 32'sh0e4ab07e, 32'sh0e492884, 32'sh0e47a089, 32'sh0e46188b, 32'sh0e44908b, 
               32'sh0e430889, 32'sh0e418085, 32'sh0e3ff87f, 32'sh0e3e7076, 32'sh0e3ce86b, 32'sh0e3b605e, 32'sh0e39d84f, 32'sh0e38503d, 
               32'sh0e36c82a, 32'sh0e354014, 32'sh0e33b7fc, 32'sh0e322fe2, 32'sh0e30a7c5, 32'sh0e2f1fa7, 32'sh0e2d9786, 32'sh0e2c0f63, 
               32'sh0e2a873e, 32'sh0e28ff16, 32'sh0e2776ed, 32'sh0e25eec1, 32'sh0e246693, 32'sh0e22de63, 32'sh0e215631, 32'sh0e1fcdfd, 
               32'sh0e1e45c6, 32'sh0e1cbd8d, 32'sh0e1b3552, 32'sh0e19ad15, 32'sh0e1824d6, 32'sh0e169c95, 32'sh0e151451, 32'sh0e138c0b, 
               32'sh0e1203c3, 32'sh0e107b79, 32'sh0e0ef32d, 32'sh0e0d6ade, 32'sh0e0be28e, 32'sh0e0a5a3b, 32'sh0e08d1e6, 32'sh0e07498f, 
               32'sh0e05c135, 32'sh0e0438da, 32'sh0e02b07c, 32'sh0e01281c, 32'sh0dff9fba, 32'sh0dfe1756, 32'sh0dfc8ef0, 32'sh0dfb0688, 
               32'sh0df97e1d, 32'sh0df7f5b0, 32'sh0df66d41, 32'sh0df4e4d0, 32'sh0df35c5d, 32'sh0df1d3e8, 32'sh0df04b70, 32'sh0deec2f7, 
               32'sh0ded3a7b, 32'sh0debb1fd, 32'sh0dea297d, 32'sh0de8a0fa, 32'sh0de71876, 32'sh0de58ff0, 32'sh0de40767, 32'sh0de27edc, 
               32'sh0de0f64f, 32'sh0ddf6dc0, 32'sh0ddde52f, 32'sh0ddc5c9b, 32'sh0ddad406, 32'sh0dd94b6e, 32'sh0dd7c2d4, 32'sh0dd63a39, 
               32'sh0dd4b19a, 32'sh0dd328fa, 32'sh0dd1a058, 32'sh0dd017b4, 32'sh0dce8f0d, 32'sh0dcd0664, 32'sh0dcb7db9, 32'sh0dc9f50c, 
               32'sh0dc86c5d, 32'sh0dc6e3ac, 32'sh0dc55af9, 32'sh0dc3d243, 32'sh0dc2498c, 32'sh0dc0c0d2, 32'sh0dbf3816, 32'sh0dbdaf58, 
               32'sh0dbc2698, 32'sh0dba9dd6, 32'sh0db91512, 32'sh0db78c4b, 32'sh0db60383, 32'sh0db47ab8, 32'sh0db2f1eb, 32'sh0db1691c, 
               32'sh0dafe04b, 32'sh0dae5778, 32'sh0daccea3, 32'sh0dab45cc, 32'sh0da9bcf2, 32'sh0da83417, 32'sh0da6ab39, 32'sh0da52259, 
               32'sh0da39978, 32'sh0da21094, 32'sh0da087ae, 32'sh0d9efec5, 32'sh0d9d75db, 32'sh0d9becef, 32'sh0d9a6400, 32'sh0d98db10, 
               32'sh0d97521d, 32'sh0d95c928, 32'sh0d944032, 32'sh0d92b739, 32'sh0d912e3e, 32'sh0d8fa541, 32'sh0d8e1c41, 32'sh0d8c9340, 
               32'sh0d8b0a3d, 32'sh0d898137, 32'sh0d87f830, 32'sh0d866f26, 32'sh0d84e61a, 32'sh0d835d0c, 32'sh0d81d3fc, 32'sh0d804aea, 
               32'sh0d7ec1d6, 32'sh0d7d38c0, 32'sh0d7bafa8, 32'sh0d7a268e, 32'sh0d789d71, 32'sh0d771453, 32'sh0d758b32, 32'sh0d740210, 
               32'sh0d7278eb, 32'sh0d70efc4, 32'sh0d6f669b, 32'sh0d6ddd70, 32'sh0d6c5443, 32'sh0d6acb14, 32'sh0d6941e3, 32'sh0d67b8b0, 
               32'sh0d662f7b, 32'sh0d64a644, 32'sh0d631d0a, 32'sh0d6193cf, 32'sh0d600a91, 32'sh0d5e8152, 32'sh0d5cf810, 32'sh0d5b6ecc, 
               32'sh0d59e586, 32'sh0d585c3f, 32'sh0d56d2f5, 32'sh0d5549a9, 32'sh0d53c05b, 32'sh0d52370b, 32'sh0d50adb9, 32'sh0d4f2465, 
               32'sh0d4d9b0e, 32'sh0d4c11b6, 32'sh0d4a885c, 32'sh0d48feff, 32'sh0d4775a1, 32'sh0d45ec40, 32'sh0d4462de, 32'sh0d42d979, 
               32'sh0d415013, 32'sh0d3fc6aa, 32'sh0d3e3d40, 32'sh0d3cb3d3, 32'sh0d3b2a64, 32'sh0d39a0f3, 32'sh0d381780, 32'sh0d368e0b, 
               32'sh0d350495, 32'sh0d337b1c, 32'sh0d31f1a1, 32'sh0d306824, 32'sh0d2edea5, 32'sh0d2d5523, 32'sh0d2bcba0, 32'sh0d2a421b, 
               32'sh0d28b894, 32'sh0d272f0b, 32'sh0d25a57f, 32'sh0d241bf2, 32'sh0d229263, 32'sh0d2108d2, 32'sh0d1f7f3e, 32'sh0d1df5a9, 
               32'sh0d1c6c11, 32'sh0d1ae278, 32'sh0d1958dd, 32'sh0d17cf3f, 32'sh0d1645a0, 32'sh0d14bbfe, 32'sh0d13325b, 32'sh0d11a8b5, 
               32'sh0d101f0e, 32'sh0d0e9564, 32'sh0d0d0bb8, 32'sh0d0b820b, 32'sh0d09f85b, 32'sh0d086eaa, 32'sh0d06e4f6, 32'sh0d055b40, 
               32'sh0d03d189, 32'sh0d0247cf, 32'sh0d00be13, 32'sh0cff3456, 32'sh0cfdaa96, 32'sh0cfc20d4, 32'sh0cfa9711, 32'sh0cf90d4b, 
               32'sh0cf78383, 32'sh0cf5f9ba, 32'sh0cf46fee, 32'sh0cf2e620, 32'sh0cf15c51, 32'sh0cefd27f, 32'sh0cee48ab, 32'sh0cecbed6, 
               32'sh0ceb34fe, 32'sh0ce9ab25, 32'sh0ce82149, 32'sh0ce6976b, 32'sh0ce50d8c, 32'sh0ce383aa, 32'sh0ce1f9c7, 32'sh0ce06fe1, 
               32'sh0cdee5f9, 32'sh0cdd5c10, 32'sh0cdbd224, 32'sh0cda4837, 32'sh0cd8be47, 32'sh0cd73456, 32'sh0cd5aa62, 32'sh0cd4206d, 
               32'sh0cd29676, 32'sh0cd10c7c, 32'sh0ccf8281, 32'sh0ccdf884, 32'sh0ccc6e84, 32'sh0ccae483, 32'sh0cc95a80, 32'sh0cc7d07a, 
               32'sh0cc64673, 32'sh0cc4bc6a, 32'sh0cc3325f, 32'sh0cc1a852, 32'sh0cc01e43, 32'sh0cbe9432, 32'sh0cbd0a1f, 32'sh0cbb800a, 
               32'sh0cb9f5f3, 32'sh0cb86bda, 32'sh0cb6e1bf, 32'sh0cb557a2, 32'sh0cb3cd84, 32'sh0cb24363, 32'sh0cb0b940, 32'sh0caf2f1b, 
               32'sh0cada4f5, 32'sh0cac1acc, 32'sh0caa90a2, 32'sh0ca90675, 32'sh0ca77c47, 32'sh0ca5f217, 32'sh0ca467e4, 32'sh0ca2ddb0, 
               32'sh0ca1537a, 32'sh0c9fc942, 32'sh0c9e3f07, 32'sh0c9cb4cb, 32'sh0c9b2a8d, 32'sh0c99a04d, 32'sh0c98160c, 32'sh0c968bc8, 
               32'sh0c950182, 32'sh0c93773a, 32'sh0c91ecf1, 32'sh0c9062a5, 32'sh0c8ed857, 32'sh0c8d4e08, 32'sh0c8bc3b7, 32'sh0c8a3963, 
               32'sh0c88af0e, 32'sh0c8724b7, 32'sh0c859a5e, 32'sh0c841002, 32'sh0c8285a5, 32'sh0c80fb47, 32'sh0c7f70e6, 32'sh0c7de683, 
               32'sh0c7c5c1e, 32'sh0c7ad1b8, 32'sh0c79474f, 32'sh0c77bce5, 32'sh0c763278, 32'sh0c74a80a, 32'sh0c731d9a, 32'sh0c719327, 
               32'sh0c7008b3, 32'sh0c6e7e3d, 32'sh0c6cf3c5, 32'sh0c6b694c, 32'sh0c69ded0, 32'sh0c685452, 32'sh0c66c9d3, 32'sh0c653f51, 
               32'sh0c63b4ce, 32'sh0c622a48, 32'sh0c609fc1, 32'sh0c5f1538, 32'sh0c5d8aad, 32'sh0c5c0020, 32'sh0c5a7591, 32'sh0c58eb00, 
               32'sh0c57606e, 32'sh0c55d5d9, 32'sh0c544b43, 32'sh0c52c0aa, 32'sh0c513610, 32'sh0c4fab74, 32'sh0c4e20d6, 32'sh0c4c9636, 
               32'sh0c4b0b94, 32'sh0c4980f0, 32'sh0c47f64a, 32'sh0c466ba3, 32'sh0c44e0f9, 32'sh0c43564e, 32'sh0c41cba1, 32'sh0c4040f2, 
               32'sh0c3eb641, 32'sh0c3d2b8e, 32'sh0c3ba0d9, 32'sh0c3a1622, 32'sh0c388b6a, 32'sh0c3700af, 32'sh0c3575f3, 32'sh0c33eb35, 
               32'sh0c326075, 32'sh0c30d5b3, 32'sh0c2f4aef, 32'sh0c2dc029, 32'sh0c2c3562, 32'sh0c2aaa98, 32'sh0c291fcd, 32'sh0c279500, 
               32'sh0c260a31, 32'sh0c247f60, 32'sh0c22f48d, 32'sh0c2169b8, 32'sh0c1fdee1, 32'sh0c1e5409, 32'sh0c1cc92f, 32'sh0c1b3e52, 
               32'sh0c19b374, 32'sh0c182894, 32'sh0c169db3, 32'sh0c1512cf, 32'sh0c1387e9, 32'sh0c11fd02, 32'sh0c107219, 32'sh0c0ee72e, 
               32'sh0c0d5c41, 32'sh0c0bd152, 32'sh0c0a4661, 32'sh0c08bb6f, 32'sh0c07307a, 32'sh0c05a584, 32'sh0c041a8c, 32'sh0c028f92, 
               32'sh0c010496, 32'sh0bff7998, 32'sh0bfdee99, 32'sh0bfc6398, 32'sh0bfad894, 32'sh0bf94d8f, 32'sh0bf7c288, 32'sh0bf63780, 
               32'sh0bf4ac75, 32'sh0bf32169, 32'sh0bf1965a, 32'sh0bf00b4a, 32'sh0bee8038, 32'sh0becf524, 32'sh0beb6a0f, 32'sh0be9def7, 
               32'sh0be853de, 32'sh0be6c8c3, 32'sh0be53da6, 32'sh0be3b287, 32'sh0be22766, 32'sh0be09c44, 32'sh0bdf111f, 32'sh0bdd85f9, 
               32'sh0bdbfad1, 32'sh0bda6fa8, 32'sh0bd8e47c, 32'sh0bd7594e, 32'sh0bd5ce1f, 32'sh0bd442ee, 32'sh0bd2b7bb, 32'sh0bd12c86, 
               32'sh0bcfa150, 32'sh0bce1617, 32'sh0bcc8add, 32'sh0bcaffa1, 32'sh0bc97463, 32'sh0bc7e923, 32'sh0bc65de2, 32'sh0bc4d29f, 
               32'sh0bc34759, 32'sh0bc1bc13, 32'sh0bc030ca, 32'sh0bbea57f, 32'sh0bbd1a33, 32'sh0bbb8ee5, 32'sh0bba0395, 32'sh0bb87843, 
               32'sh0bb6ecef, 32'sh0bb5619a, 32'sh0bb3d642, 32'sh0bb24ae9, 32'sh0bb0bf8f, 32'sh0baf3432, 32'sh0bada8d4, 32'sh0bac1d73, 
               32'sh0baa9211, 32'sh0ba906ad, 32'sh0ba77b48, 32'sh0ba5efe0, 32'sh0ba46477, 32'sh0ba2d90c, 32'sh0ba14d9f, 32'sh0b9fc231, 
               32'sh0b9e36c0, 32'sh0b9cab4e, 32'sh0b9b1fda, 32'sh0b999464, 32'sh0b9808ed, 32'sh0b967d73, 32'sh0b94f1f8, 32'sh0b93667b, 
               32'sh0b91dafc, 32'sh0b904f7c, 32'sh0b8ec3fa, 32'sh0b8d3876, 32'sh0b8bacf0, 32'sh0b8a2168, 32'sh0b8895df, 32'sh0b870a53, 
               32'sh0b857ec7, 32'sh0b83f338, 32'sh0b8267a7, 32'sh0b80dc15, 32'sh0b7f5081, 32'sh0b7dc4eb, 32'sh0b7c3953, 32'sh0b7aadba, 
               32'sh0b79221f, 32'sh0b779682, 32'sh0b760ae3, 32'sh0b747f43, 32'sh0b72f3a1, 32'sh0b7167fd, 32'sh0b6fdc57, 32'sh0b6e50af, 
               32'sh0b6cc506, 32'sh0b6b395b, 32'sh0b69adae, 32'sh0b682200, 32'sh0b66964f, 32'sh0b650a9d, 32'sh0b637ee9, 32'sh0b61f334, 
               32'sh0b60677c, 32'sh0b5edbc3, 32'sh0b5d5008, 32'sh0b5bc44c, 32'sh0b5a388d, 32'sh0b58accd, 32'sh0b57210b, 32'sh0b559548, 
               32'sh0b540982, 32'sh0b527dbb, 32'sh0b50f1f3, 32'sh0b4f6628, 32'sh0b4dda5c, 32'sh0b4c4e8d, 32'sh0b4ac2be, 32'sh0b4936ec, 
               32'sh0b47ab19, 32'sh0b461f44, 32'sh0b44936d, 32'sh0b430794, 32'sh0b417bba, 32'sh0b3fefde, 32'sh0b3e6400, 32'sh0b3cd821, 
               32'sh0b3b4c40, 32'sh0b39c05d, 32'sh0b383478, 32'sh0b36a892, 32'sh0b351caa, 32'sh0b3390c0, 32'sh0b3204d4, 32'sh0b3078e7, 
               32'sh0b2eecf8, 32'sh0b2d6107, 32'sh0b2bd515, 32'sh0b2a4920, 32'sh0b28bd2a, 32'sh0b273133, 32'sh0b25a539, 32'sh0b24193e, 
               32'sh0b228d42, 32'sh0b210143, 32'sh0b1f7543, 32'sh0b1de941, 32'sh0b1c5d3d, 32'sh0b1ad138, 32'sh0b194531, 32'sh0b17b928, 
               32'sh0b162d1d, 32'sh0b14a111, 32'sh0b131503, 32'sh0b1188f4, 32'sh0b0ffce2, 32'sh0b0e70cf, 32'sh0b0ce4ba, 32'sh0b0b58a4, 
               32'sh0b09cc8c, 32'sh0b084072, 32'sh0b06b456, 32'sh0b052839, 32'sh0b039c1a, 32'sh0b020ff9, 32'sh0b0083d7, 32'sh0afef7b3, 
               32'sh0afd6b8d, 32'sh0afbdf66, 32'sh0afa533d, 32'sh0af8c712, 32'sh0af73ae5, 32'sh0af5aeb7, 32'sh0af42287, 32'sh0af29656, 
               32'sh0af10a22, 32'sh0aef7ded, 32'sh0aedf1b7, 32'sh0aec657e, 32'sh0aead944, 32'sh0ae94d09, 32'sh0ae7c0cb, 32'sh0ae6348c, 
               32'sh0ae4a84b, 32'sh0ae31c09, 32'sh0ae18fc5, 32'sh0ae0037f, 32'sh0ade7737, 32'sh0adceaee, 32'sh0adb5ea3, 32'sh0ad9d257, 
               32'sh0ad84609, 32'sh0ad6b9b9, 32'sh0ad52d67, 32'sh0ad3a114, 32'sh0ad214bf, 32'sh0ad08869, 32'sh0acefc11, 32'sh0acd6fb7, 
               32'sh0acbe35b, 32'sh0aca56fe, 32'sh0ac8ca9f, 32'sh0ac73e3f, 32'sh0ac5b1dc, 32'sh0ac42579, 32'sh0ac29913, 32'sh0ac10cac, 
               32'sh0abf8043, 32'sh0abdf3d9, 32'sh0abc676d, 32'sh0abadaff, 32'sh0ab94e8f, 32'sh0ab7c21e, 32'sh0ab635ab, 32'sh0ab4a937, 
               32'sh0ab31cc1, 32'sh0ab19049, 32'sh0ab003d0, 32'sh0aae7755, 32'sh0aacead8, 32'sh0aab5e5a, 32'sh0aa9d1da, 32'sh0aa84558, 
               32'sh0aa6b8d5, 32'sh0aa52c50, 32'sh0aa39fca, 32'sh0aa21342, 32'sh0aa086b8, 32'sh0a9efa2c, 32'sh0a9d6d9f, 32'sh0a9be111, 
               32'sh0a9a5480, 32'sh0a98c7ee, 32'sh0a973b5b, 32'sh0a95aec5, 32'sh0a94222f, 32'sh0a929596, 32'sh0a9108fc, 32'sh0a8f7c60, 
               32'sh0a8defc3, 32'sh0a8c6324, 32'sh0a8ad683, 32'sh0a8949e1, 32'sh0a87bd3d, 32'sh0a863097, 32'sh0a84a3f0, 32'sh0a831747, 
               32'sh0a818a9d, 32'sh0a7ffdf1, 32'sh0a7e7143, 32'sh0a7ce494, 32'sh0a7b57e3, 32'sh0a79cb31, 32'sh0a783e7d, 32'sh0a76b1c7, 
               32'sh0a752510, 32'sh0a739857, 32'sh0a720b9c, 32'sh0a707ee0, 32'sh0a6ef222, 32'sh0a6d6563, 32'sh0a6bd8a2, 32'sh0a6a4bdf, 
               32'sh0a68bf1b, 32'sh0a673255, 32'sh0a65a58e, 32'sh0a6418c5, 32'sh0a628bfa, 32'sh0a60ff2e, 32'sh0a5f7260, 32'sh0a5de591, 
               32'sh0a5c58c0, 32'sh0a5acbed, 32'sh0a593f19, 32'sh0a57b243, 32'sh0a56256c, 32'sh0a549893, 32'sh0a530bb8, 32'sh0a517edc, 
               32'sh0a4ff1fe, 32'sh0a4e651f, 32'sh0a4cd83e, 32'sh0a4b4b5b, 32'sh0a49be77, 32'sh0a483191, 32'sh0a46a4aa, 32'sh0a4517c1, 
               32'sh0a438ad7, 32'sh0a41fdeb, 32'sh0a4070fd, 32'sh0a3ee40e, 32'sh0a3d571d, 32'sh0a3bca2b, 32'sh0a3a3d37, 32'sh0a38b041, 
               32'sh0a37234a, 32'sh0a359651, 32'sh0a340957, 32'sh0a327c5b, 32'sh0a30ef5e, 32'sh0a2f625f, 32'sh0a2dd55e, 32'sh0a2c485c, 
               32'sh0a2abb59, 32'sh0a292e53, 32'sh0a27a14d, 32'sh0a261444, 32'sh0a24873a, 32'sh0a22fa2f, 32'sh0a216d22, 32'sh0a1fe013, 
               32'sh0a1e5303, 32'sh0a1cc5f1, 32'sh0a1b38de, 32'sh0a19abc9, 32'sh0a181eb2, 32'sh0a16919a, 32'sh0a150481, 32'sh0a137766, 
               32'sh0a11ea49, 32'sh0a105d2b, 32'sh0a0ed00b, 32'sh0a0d42ea, 32'sh0a0bb5c7, 32'sh0a0a28a2, 32'sh0a089b7c, 32'sh0a070e55, 
               32'sh0a05812c, 32'sh0a03f401, 32'sh0a0266d5, 32'sh0a00d9a7, 32'sh09ff4c78, 32'sh09fdbf47, 32'sh09fc3215, 32'sh09faa4e1, 
               32'sh09f917ac, 32'sh09f78a75, 32'sh09f5fd3d, 32'sh09f47003, 32'sh09f2e2c7, 32'sh09f1558a, 32'sh09efc84b, 32'sh09ee3b0b, 
               32'sh09ecadc9, 32'sh09eb2086, 32'sh09e99342, 32'sh09e805fb, 32'sh09e678b4, 32'sh09e4eb6a, 32'sh09e35e1f, 32'sh09e1d0d3, 
               32'sh09e04385, 32'sh09deb636, 32'sh09dd28e5, 32'sh09db9b92, 32'sh09da0e3e, 32'sh09d880e9, 32'sh09d6f392, 32'sh09d56639, 
               32'sh09d3d8df, 32'sh09d24b84, 32'sh09d0be27, 32'sh09cf30c8, 32'sh09cda368, 32'sh09cc1606, 32'sh09ca88a3, 32'sh09c8fb3f, 
               32'sh09c76dd8, 32'sh09c5e071, 32'sh09c45308, 32'sh09c2c59d, 32'sh09c13831, 32'sh09bfaac3, 32'sh09be1d54, 32'sh09bc8fe3, 
               32'sh09bb0271, 32'sh09b974fd, 32'sh09b7e788, 32'sh09b65a11, 32'sh09b4cc99, 32'sh09b33f20, 32'sh09b1b1a4, 32'sh09b02428, 
               32'sh09ae96aa, 32'sh09ad092a, 32'sh09ab7ba9, 32'sh09a9ee26, 32'sh09a860a2, 32'sh09a6d31c, 32'sh09a54595, 32'sh09a3b80d, 
               32'sh09a22a83, 32'sh09a09cf7, 32'sh099f0f6a, 32'sh099d81dc, 32'sh099bf44c, 32'sh099a66ba, 32'sh0998d927, 32'sh09974b93, 
               32'sh0995bdfd, 32'sh09943065, 32'sh0992a2cc, 32'sh09911532, 32'sh098f8796, 32'sh098df9f9, 32'sh098c6c5a, 32'sh098adeba, 
               32'sh09895118, 32'sh0987c375, 32'sh098635d0, 32'sh0984a82a, 32'sh09831a82, 32'sh09818cd9, 32'sh097fff2f, 32'sh097e7183, 
               32'sh097ce3d5, 32'sh097b5626, 32'sh0979c876, 32'sh09783ac4, 32'sh0976ad11, 32'sh09751f5c, 32'sh097391a6, 32'sh097203ee, 
               32'sh09707635, 32'sh096ee87a, 32'sh096d5abe, 32'sh096bcd01, 32'sh096a3f42, 32'sh0968b181, 32'sh096723bf, 32'sh096595fc, 
               32'sh09640837, 32'sh09627a71, 32'sh0960eca9, 32'sh095f5ee0, 32'sh095dd116, 32'sh095c434a, 32'sh095ab57c, 32'sh095927ad, 
               32'sh095799dd, 32'sh09560c0b, 32'sh09547e38, 32'sh0952f063, 32'sh0951628d, 32'sh094fd4b6, 32'sh094e46dd, 32'sh094cb902, 
               32'sh094b2b27, 32'sh09499d49, 32'sh09480f6b, 32'sh0946818a, 32'sh0944f3a9, 32'sh094365c6, 32'sh0941d7e2, 32'sh094049fc, 
               32'sh093ebc14, 32'sh093d2e2c, 32'sh093ba042, 32'sh093a1256, 32'sh09388469, 32'sh0936f67b, 32'sh0935688b, 32'sh0933da9a, 
               32'sh09324ca7, 32'sh0930beb3, 32'sh092f30bd, 32'sh092da2c7, 32'sh092c14ce, 32'sh092a86d4, 32'sh0928f8d9, 32'sh09276add, 
               32'sh0925dcdf, 32'sh09244edf, 32'sh0922c0df, 32'sh092132dc, 32'sh091fa4d9, 32'sh091e16d4, 32'sh091c88cd, 32'sh091afac6, 
               32'sh09196cbc, 32'sh0917deb2, 32'sh091650a6, 32'sh0914c298, 32'sh09133489, 32'sh0911a679, 32'sh09101868, 32'sh090e8a54, 
               32'sh090cfc40, 32'sh090b6e2a, 32'sh0909e013, 32'sh090851fa, 32'sh0906c3e0, 32'sh090535c5, 32'sh0903a7a8, 32'sh0902198a, 
               32'sh09008b6a, 32'sh08fefd4a, 32'sh08fd6f27, 32'sh08fbe103, 32'sh08fa52de, 32'sh08f8c4b8, 32'sh08f73690, 32'sh08f5a867, 
               32'sh08f41a3c, 32'sh08f28c10, 32'sh08f0fde3, 32'sh08ef6fb4, 32'sh08ede184, 32'sh08ec5352, 32'sh08eac51f, 32'sh08e936eb, 
               32'sh08e7a8b5, 32'sh08e61a7e, 32'sh08e48c46, 32'sh08e2fe0c, 32'sh08e16fd1, 32'sh08dfe194, 32'sh08de5356, 32'sh08dcc517, 
               32'sh08db36d6, 32'sh08d9a894, 32'sh08d81a51, 32'sh08d68c0c, 32'sh08d4fdc6, 32'sh08d36f7f, 32'sh08d1e136, 32'sh08d052ec, 
               32'sh08cec4a0, 32'sh08cd3653, 32'sh08cba805, 32'sh08ca19b6, 32'sh08c88b65, 32'sh08c6fd12, 32'sh08c56ebf, 32'sh08c3e06a, 
               32'sh08c25213, 32'sh08c0c3bc, 32'sh08bf3563, 32'sh08bda708, 32'sh08bc18ac, 32'sh08ba8a4f, 32'sh08b8fbf1, 32'sh08b76d91, 
               32'sh08b5df30, 32'sh08b450cd, 32'sh08b2c26a, 32'sh08b13404, 32'sh08afa59e, 32'sh08ae1736, 32'sh08ac88cd, 32'sh08aafa62, 
               32'sh08a96bf6, 32'sh08a7dd89, 32'sh08a64f1b, 32'sh08a4c0ab, 32'sh08a3323a, 32'sh08a1a3c7, 32'sh08a01553, 32'sh089e86de, 
               32'sh089cf867, 32'sh089b69f0, 32'sh0899db76, 32'sh08984cfc, 32'sh0896be80, 32'sh08953003, 32'sh0893a184, 32'sh08921305, 
               32'sh08908483, 32'sh088ef601, 32'sh088d677d, 32'sh088bd8f8, 32'sh088a4a72, 32'sh0888bbea, 32'sh08872d61, 32'sh08859ed7, 
               32'sh0884104b, 32'sh088281be, 32'sh0880f330, 32'sh087f64a0, 32'sh087dd60f, 32'sh087c477d, 32'sh087ab8e9, 32'sh08792a55, 
               32'sh08779bbe, 32'sh08760d27, 32'sh08747e8e, 32'sh0872eff4, 32'sh08716159, 32'sh086fd2bc, 32'sh086e441e, 32'sh086cb57f, 
               32'sh086b26de, 32'sh0869983c, 32'sh08680999, 32'sh08667af5, 32'sh0864ec4f, 32'sh08635da8, 32'sh0861cf00, 32'sh08604056, 
               32'sh085eb1ab, 32'sh085d22ff, 32'sh085b9451, 32'sh085a05a3, 32'sh085876f3, 32'sh0856e841, 32'sh0855598f, 32'sh0853cadb, 
               32'sh08523c25, 32'sh0850ad6f, 32'sh084f1eb7, 32'sh084d8ffe, 32'sh084c0144, 32'sh084a7288, 32'sh0848e3cb, 32'sh0847550d, 
               32'sh0845c64d, 32'sh0844378d, 32'sh0842a8cb, 32'sh08411a07, 32'sh083f8b43, 32'sh083dfc7d, 32'sh083c6db6, 32'sh083adeee, 
               32'sh08395024, 32'sh0837c159, 32'sh0836328d, 32'sh0834a3bf, 32'sh083314f1, 32'sh08318621, 32'sh082ff74f, 32'sh082e687d, 
               32'sh082cd9a9, 32'sh082b4ad4, 32'sh0829bbfe, 32'sh08282d26, 32'sh08269e4d, 32'sh08250f73, 32'sh08238098, 32'sh0821f1bc, 
               32'sh082062de, 32'sh081ed3ff, 32'sh081d451e, 32'sh081bb63d, 32'sh081a275a, 32'sh08189876, 32'sh08170990, 32'sh08157aaa, 
               32'sh0813ebc2, 32'sh08125cd9, 32'sh0810cdef, 32'sh080f3f03, 32'sh080db016, 32'sh080c2128, 32'sh080a9239, 32'sh08090348, 
               32'sh08077457, 32'sh0805e564, 32'sh0804566f, 32'sh0802c77a, 32'sh08013883, 32'sh07ffa98b, 32'sh07fe1a92, 32'sh07fc8b98, 
               32'sh07fafc9c, 32'sh07f96d9f, 32'sh07f7dea1, 32'sh07f64fa2, 32'sh07f4c0a1, 32'sh07f3319f, 32'sh07f1a29c, 32'sh07f01398, 
               32'sh07ee8493, 32'sh07ecf58c, 32'sh07eb6684, 32'sh07e9d77b, 32'sh07e84871, 32'sh07e6b965, 32'sh07e52a58, 32'sh07e39b4a, 
               32'sh07e20c3b, 32'sh07e07d2b, 32'sh07deee19, 32'sh07dd5f06, 32'sh07dbcff2, 32'sh07da40dd, 32'sh07d8b1c6, 32'sh07d722af, 
               32'sh07d59396, 32'sh07d4047c, 32'sh07d27560, 32'sh07d0e644, 32'sh07cf5726, 32'sh07cdc807, 32'sh07cc38e7, 32'sh07caa9c5, 
               32'sh07c91aa3, 32'sh07c78b7f, 32'sh07c5fc5a, 32'sh07c46d34, 32'sh07c2de0d, 32'sh07c14ee4, 32'sh07bfbfba, 32'sh07be308f, 
               32'sh07bca163, 32'sh07bb1236, 32'sh07b98307, 32'sh07b7f3d8, 32'sh07b664a7, 32'sh07b4d575, 32'sh07b34641, 32'sh07b1b70d, 
               32'sh07b027d7, 32'sh07ae98a0, 32'sh07ad0968, 32'sh07ab7a2f, 32'sh07a9eaf5, 32'sh07a85bb9, 32'sh07a6cc7d, 32'sh07a53d3f, 
               32'sh07a3adff, 32'sh07a21ebf, 32'sh07a08f7e, 32'sh079f003b, 32'sh079d70f7, 32'sh079be1b2, 32'sh079a526c, 32'sh0798c325, 
               32'sh079733dc, 32'sh0795a493, 32'sh07941548, 32'sh079285fc, 32'sh0790f6ae, 32'sh078f6760, 32'sh078dd811, 32'sh078c48c0, 
               32'sh078ab96e, 32'sh07892a1b, 32'sh07879ac7, 32'sh07860b72, 32'sh07847c1b, 32'sh0782ecc3, 32'sh07815d6b, 32'sh077fce11, 
               32'sh077e3eb5, 32'sh077caf59, 32'sh077b1ffc, 32'sh0779909d, 32'sh0778013d, 32'sh077671dd, 32'sh0774e27a, 32'sh07735317, 
               32'sh0771c3b3, 32'sh0770344d, 32'sh076ea4e7, 32'sh076d157f, 32'sh076b8616, 32'sh0769f6ac, 32'sh07686741, 32'sh0766d7d4, 
               32'sh07654867, 32'sh0763b8f8, 32'sh07622988, 32'sh07609a18, 32'sh075f0aa5, 32'sh075d7b32, 32'sh075bebbe, 32'sh075a5c48, 
               32'sh0758ccd2, 32'sh07573d5a, 32'sh0755ade1, 32'sh07541e67, 32'sh07528eec, 32'sh0750ff70, 32'sh074f6ff3, 32'sh074de074, 
               32'sh074c50f4, 32'sh074ac174, 32'sh074931f2, 32'sh0747a26f, 32'sh074612eb, 32'sh07448365, 32'sh0742f3df, 32'sh07416457, 
               32'sh073fd4cf, 32'sh073e4545, 32'sh073cb5ba, 32'sh073b262e, 32'sh073996a1, 32'sh07380713, 32'sh07367784, 32'sh0734e7f3, 
               32'sh07335862, 32'sh0731c8cf, 32'sh0730393b, 32'sh072ea9a6, 32'sh072d1a10, 32'sh072b8a79, 32'sh0729fae1, 32'sh07286b48, 
               32'sh0726dbae, 32'sh07254c12, 32'sh0723bc75, 32'sh07222cd8, 32'sh07209d39, 32'sh071f0d99, 32'sh071d7df8, 32'sh071bee56, 
               32'sh071a5eb3, 32'sh0718cf0e, 32'sh07173f69, 32'sh0715afc3, 32'sh0714201b, 32'sh07129072, 32'sh071100c9, 32'sh070f711e, 
               32'sh070de172, 32'sh070c51c5, 32'sh070ac217, 32'sh07093268, 32'sh0707a2b7, 32'sh07061306, 32'sh07048354, 32'sh0702f3a0, 
               32'sh070163eb, 32'sh06ffd436, 32'sh06fe447f, 32'sh06fcb4c7, 32'sh06fb250e, 32'sh06f99554, 32'sh06f80599, 32'sh06f675dd, 
               32'sh06f4e620, 32'sh06f35662, 32'sh06f1c6a2, 32'sh06f036e2, 32'sh06eea720, 32'sh06ed175e, 32'sh06eb879a, 32'sh06e9f7d5, 
               32'sh06e86810, 32'sh06e6d849, 32'sh06e54881, 32'sh06e3b8b8, 32'sh06e228ee, 32'sh06e09923, 32'sh06df0957, 32'sh06dd7989, 
               32'sh06dbe9bb, 32'sh06da59ec, 32'sh06d8ca1b, 32'sh06d73a4a, 32'sh06d5aa77, 32'sh06d41aa4, 32'sh06d28acf, 32'sh06d0fafa, 
               32'sh06cf6b23, 32'sh06cddb4b, 32'sh06cc4b72, 32'sh06cabb98, 32'sh06c92bbe, 32'sh06c79be2, 32'sh06c60c05, 32'sh06c47c27, 
               32'sh06c2ec48, 32'sh06c15c67, 32'sh06bfcc86, 32'sh06be3ca4, 32'sh06bcacc1, 32'sh06bb1cdd, 32'sh06b98cf7, 32'sh06b7fd11, 
               32'sh06b66d29, 32'sh06b4dd41, 32'sh06b34d58, 32'sh06b1bd6d, 32'sh06b02d81, 32'sh06ae9d95, 32'sh06ad0da7, 32'sh06ab7db9, 
               32'sh06a9edc9, 32'sh06a85dd8, 32'sh06a6cde7, 32'sh06a53df4, 32'sh06a3ae00, 32'sh06a21e0b, 32'sh06a08e16, 32'sh069efe1f, 
               32'sh069d6e27, 32'sh069bde2e, 32'sh069a4e34, 32'sh0698be39, 32'sh06972e3d, 32'sh06959e40, 32'sh06940e42, 32'sh06927e44, 
               32'sh0690ee44, 32'sh068f5e43, 32'sh068dce41, 32'sh068c3e3e, 32'sh068aae3a, 32'sh06891e34, 32'sh06878e2e, 32'sh0685fe27, 
               32'sh06846e1f, 32'sh0682de16, 32'sh06814e0c, 32'sh067fbe01, 32'sh067e2df5, 32'sh067c9de8, 32'sh067b0dda, 32'sh06797dcb, 
               32'sh0677edbb, 32'sh06765daa, 32'sh0674cd98, 32'sh06733d85, 32'sh0671ad71, 32'sh06701d5b, 32'sh066e8d45, 32'sh066cfd2e, 
               32'sh066b6d16, 32'sh0669dcfd, 32'sh06684ce3, 32'sh0666bcc8, 32'sh06652cac, 32'sh06639c8f, 32'sh06620c72, 32'sh06607c53, 
               32'sh065eec33, 32'sh065d5c12, 32'sh065bcbf0, 32'sh065a3bcd, 32'sh0658aba9, 32'sh06571b84, 32'sh06558b5f, 32'sh0653fb38, 
               32'sh06526b10, 32'sh0650dae7, 32'sh064f4abe, 32'sh064dba93, 32'sh064c2a67, 32'sh064a9a3b, 32'sh06490a0d, 32'sh064779df, 
               32'sh0645e9af, 32'sh0644597f, 32'sh0642c94d, 32'sh0641391b, 32'sh063fa8e7, 32'sh063e18b3, 32'sh063c887e, 32'sh063af847, 
               32'sh06396810, 32'sh0637d7d8, 32'sh0636479f, 32'sh0634b765, 32'sh0633272a, 32'sh063196ee, 32'sh063006b1, 32'sh062e7673, 
               32'sh062ce634, 32'sh062b55f4, 32'sh0629c5b3, 32'sh06283571, 32'sh0626a52f, 32'sh062514eb, 32'sh062384a6, 32'sh0621f461, 
               32'sh0620641a, 32'sh061ed3d3, 32'sh061d438b, 32'sh061bb341, 32'sh061a22f7, 32'sh061892ac, 32'sh06170260, 32'sh06157213, 
               32'sh0613e1c5, 32'sh06125176, 32'sh0610c126, 32'sh060f30d5, 32'sh060da083, 32'sh060c1031, 32'sh060a7fdd, 32'sh0608ef88, 
               32'sh06075f33, 32'sh0605cedd, 32'sh06043e85, 32'sh0602ae2d, 32'sh06011dd4, 32'sh05ff8d7a, 32'sh05fdfd1f, 32'sh05fc6cc3, 
               32'sh05fadc66, 32'sh05f94c08, 32'sh05f7bba9, 32'sh05f62b49, 32'sh05f49ae9, 32'sh05f30a87, 32'sh05f17a25, 32'sh05efe9c2, 
               32'sh05ee595d, 32'sh05ecc8f8, 32'sh05eb3892, 32'sh05e9a82b, 32'sh05e817c3, 32'sh05e6875a, 32'sh05e4f6f1, 32'sh05e36686, 
               32'sh05e1d61b, 32'sh05e045ae, 32'sh05deb541, 32'sh05dd24d3, 32'sh05db9463, 32'sh05da03f3, 32'sh05d87382, 32'sh05d6e310, 
               32'sh05d5529e, 32'sh05d3c22a, 32'sh05d231b5, 32'sh05d0a140, 32'sh05cf10ca, 32'sh05cd8052, 32'sh05cbefda, 32'sh05ca5f61, 
               32'sh05c8cee7, 32'sh05c73e6c, 32'sh05c5adf1, 32'sh05c41d74, 32'sh05c28cf7, 32'sh05c0fc78, 32'sh05bf6bf9, 32'sh05bddb79, 
               32'sh05bc4af8, 32'sh05baba76, 32'sh05b929f3, 32'sh05b7996f, 32'sh05b608eb, 32'sh05b47865, 32'sh05b2e7df, 32'sh05b15758, 
               32'sh05afc6d0, 32'sh05ae3647, 32'sh05aca5bd, 32'sh05ab1532, 32'sh05a984a6, 32'sh05a7f41a, 32'sh05a6638d, 32'sh05a4d2fe, 
               32'sh05a3426f, 32'sh05a1b1df, 32'sh05a0214f, 32'sh059e90bd, 32'sh059d002a, 32'sh059b6f97, 32'sh0599df03, 32'sh05984e6d, 
               32'sh0596bdd7, 32'sh05952d41, 32'sh05939ca9, 32'sh05920c10, 32'sh05907b77, 32'sh058eeadc, 32'sh058d5a41, 32'sh058bc9a5, 
               32'sh058a3908, 32'sh0588a86b, 32'sh058717cc, 32'sh0585872d, 32'sh0583f68c, 32'sh058265eb, 32'sh0580d549, 32'sh057f44a6, 
               32'sh057db403, 32'sh057c235e, 32'sh057a92b9, 32'sh05790213, 32'sh0577716b, 32'sh0575e0c4, 32'sh0574501b, 32'sh0572bf71, 
               32'sh05712ec7, 32'sh056f9e1b, 32'sh056e0d6f, 32'sh056c7cc2, 32'sh056aec15, 32'sh05695b66, 32'sh0567cab6, 32'sh05663a06, 
               32'sh0564a955, 32'sh056318a3, 32'sh056187f0, 32'sh055ff73d, 32'sh055e6688, 32'sh055cd5d3, 32'sh055b451d, 32'sh0559b466, 
               32'sh055823ae, 32'sh055692f6, 32'sh0555023c, 32'sh05537182, 32'sh0551e0c7, 32'sh0550500b, 32'sh054ebf4e, 32'sh054d2e91, 
               32'sh054b9dd3, 32'sh054a0d13, 32'sh05487c53, 32'sh0546eb93, 32'sh05455ad1, 32'sh0543ca0f, 32'sh0542394c, 32'sh0540a888, 
               32'sh053f17c3, 32'sh053d86fd, 32'sh053bf637, 32'sh053a656f, 32'sh0538d4a7, 32'sh053743de, 32'sh0535b315, 32'sh0534224a, 
               32'sh0532917f, 32'sh053100b3, 32'sh052f6fe6, 32'sh052ddf18, 32'sh052c4e4a, 32'sh052abd7b, 32'sh05292cab, 32'sh05279bda, 
               32'sh05260b08, 32'sh05247a36, 32'sh0522e962, 32'sh0521588e, 32'sh051fc7b9, 32'sh051e36e4, 32'sh051ca60d, 32'sh051b1536, 
               32'sh0519845e, 32'sh0517f386, 32'sh051662ac, 32'sh0514d1d2, 32'sh051340f6, 32'sh0511b01b, 32'sh05101f3e, 32'sh050e8e60, 
               32'sh050cfd82, 32'sh050b6ca3, 32'sh0509dbc3, 32'sh05084ae3, 32'sh0506ba01, 32'sh0505291f, 32'sh0503983c, 32'sh05020759, 
               32'sh05007674, 32'sh04fee58f, 32'sh04fd54a9, 32'sh04fbc3c2, 32'sh04fa32db, 32'sh04f8a1f2, 32'sh04f71109, 32'sh04f5801f, 
               32'sh04f3ef35, 32'sh04f25e4a, 32'sh04f0cd5d, 32'sh04ef3c71, 32'sh04edab83, 32'sh04ec1a94, 32'sh04ea89a5, 32'sh04e8f8b5, 
               32'sh04e767c5, 32'sh04e5d6d3, 32'sh04e445e1, 32'sh04e2b4ee, 32'sh04e123fa, 32'sh04df9306, 32'sh04de0211, 32'sh04dc711b, 
               32'sh04dae024, 32'sh04d94f2d, 32'sh04d7be34, 32'sh04d62d3b, 32'sh04d49c42, 32'sh04d30b47, 32'sh04d17a4c, 32'sh04cfe950, 
               32'sh04ce5854, 32'sh04ccc756, 32'sh04cb3658, 32'sh04c9a559, 32'sh04c81459, 32'sh04c68359, 32'sh04c4f258, 32'sh04c36156, 
               32'sh04c1d054, 32'sh04c03f50, 32'sh04beae4c, 32'sh04bd1d47, 32'sh04bb8c42, 32'sh04b9fb3c, 32'sh04b86a35, 32'sh04b6d92d, 
               32'sh04b54825, 32'sh04b3b71c, 32'sh04b22612, 32'sh04b09507, 32'sh04af03fc, 32'sh04ad72f0, 32'sh04abe1e3, 32'sh04aa50d6, 
               32'sh04a8bfc7, 32'sh04a72eb8, 32'sh04a59da9, 32'sh04a40c98, 32'sh04a27b87, 32'sh04a0ea76, 32'sh049f5963, 32'sh049dc850, 
               32'sh049c373c, 32'sh049aa627, 32'sh04991512, 32'sh049783fc, 32'sh0495f2e5, 32'sh049461ce, 32'sh0492d0b6, 32'sh04913f9d, 
               32'sh048fae83, 32'sh048e1d69, 32'sh048c8c4e, 32'sh048afb32, 32'sh04896a16, 32'sh0487d8f9, 32'sh048647db, 32'sh0484b6bc, 
               32'sh0483259d, 32'sh0481947d, 32'sh0480035d, 32'sh047e723c, 32'sh047ce11a, 32'sh047b4ff7, 32'sh0479bed4, 32'sh04782db0, 
               32'sh04769c8b, 32'sh04750b65, 32'sh04737a3f, 32'sh0471e919, 32'sh047057f1, 32'sh046ec6c9, 32'sh046d35a0, 32'sh046ba477, 
               32'sh046a134c, 32'sh04688221, 32'sh0466f0f6, 32'sh04655fca, 32'sh0463ce9d, 32'sh04623d6f, 32'sh0460ac41, 32'sh045f1b12, 
               32'sh045d89e2, 32'sh045bf8b2, 32'sh045a6781, 32'sh0458d64f, 32'sh0457451d, 32'sh0455b3ea, 32'sh045422b7, 32'sh04529182, 
               32'sh0451004d, 32'sh044f6f18, 32'sh044ddde1, 32'sh044c4caa, 32'sh044abb73, 32'sh04492a3a, 32'sh04479901, 32'sh044607c8, 
               32'sh0444768d, 32'sh0442e553, 32'sh04415417, 32'sh043fc2db, 32'sh043e319e, 32'sh043ca060, 32'sh043b0f22, 32'sh04397de3, 
               32'sh0437eca4, 32'sh04365b63, 32'sh0434ca23, 32'sh043338e1, 32'sh0431a79f, 32'sh0430165c, 32'sh042e8519, 32'sh042cf3d5, 
               32'sh042b6290, 32'sh0429d14b, 32'sh04284005, 32'sh0426aebe, 32'sh04251d77, 32'sh04238c2f, 32'sh0421fae7, 32'sh0420699d, 
               32'sh041ed854, 32'sh041d4709, 32'sh041bb5be, 32'sh041a2472, 32'sh04189326, 32'sh041701d9, 32'sh0415708b, 32'sh0413df3d, 
               32'sh04124dee, 32'sh0410bc9f, 32'sh040f2b4f, 32'sh040d99fe, 32'sh040c08ad, 32'sh040a775b, 32'sh0408e608, 32'sh040754b5, 
               32'sh0405c361, 32'sh0404320c, 32'sh0402a0b7, 32'sh04010f61, 32'sh03ff7e0b, 32'sh03fdecb4, 32'sh03fc5b5d, 32'sh03faca04, 
               32'sh03f938ac, 32'sh03f7a752, 32'sh03f615f8, 32'sh03f4849e, 32'sh03f2f342, 32'sh03f161e6, 32'sh03efd08a, 32'sh03ee3f2d, 
               32'sh03ecadcf, 32'sh03eb1c71, 32'sh03e98b12, 32'sh03e7f9b3, 32'sh03e66852, 32'sh03e4d6f2, 32'sh03e34591, 32'sh03e1b42f, 
               32'sh03e022cc, 32'sh03de9169, 32'sh03dd0005, 32'sh03db6ea1, 32'sh03d9dd3c, 32'sh03d84bd7, 32'sh03d6ba71, 32'sh03d5290a, 
               32'sh03d397a3, 32'sh03d2063b, 32'sh03d074d2, 32'sh03cee369, 32'sh03cd5200, 32'sh03cbc096, 32'sh03ca2f2b, 32'sh03c89dc0, 
               32'sh03c70c54, 32'sh03c57ae7, 32'sh03c3e97a, 32'sh03c2580c, 32'sh03c0c69e, 32'sh03bf352f, 32'sh03bda3c0, 32'sh03bc1250, 
               32'sh03ba80df, 32'sh03b8ef6e, 32'sh03b75dfc, 32'sh03b5cc8a, 32'sh03b43b17, 32'sh03b2a9a4, 32'sh03b11830, 32'sh03af86bb, 
               32'sh03adf546, 32'sh03ac63d0, 32'sh03aad25a, 32'sh03a940e3, 32'sh03a7af6c, 32'sh03a61df4, 32'sh03a48c7b, 32'sh03a2fb02, 
               32'sh03a16988, 32'sh039fd80e, 32'sh039e4693, 32'sh039cb518, 32'sh039b239c, 32'sh03999220, 32'sh039800a3, 32'sh03966f25, 
               32'sh0394dda7, 32'sh03934c28, 32'sh0391baa9, 32'sh03902929, 32'sh038e97a9, 32'sh038d0628, 32'sh038b74a7, 32'sh0389e325, 
               32'sh038851a2, 32'sh0386c01f, 32'sh03852e9c, 32'sh03839d18, 32'sh03820b93, 32'sh03807a0e, 32'sh037ee888, 32'sh037d5702, 
               32'sh037bc57b, 32'sh037a33f3, 32'sh0378a26b, 32'sh037710e3, 32'sh03757f5a, 32'sh0373edd1, 32'sh03725c46, 32'sh0370cabc, 
               32'sh036f3931, 32'sh036da7a5, 32'sh036c1619, 32'sh036a848c, 32'sh0368f2ff, 32'sh03676171, 32'sh0365cfe3, 32'sh03643e54, 
               32'sh0362acc5, 32'sh03611b35, 32'sh035f89a5, 32'sh035df814, 32'sh035c6682, 32'sh035ad4f1, 32'sh0359435e, 32'sh0357b1cb, 
               32'sh03562038, 32'sh03548ea4, 32'sh0352fd0f, 32'sh03516b7a, 32'sh034fd9e5, 32'sh034e484f, 32'sh034cb6b8, 32'sh034b2521, 
               32'sh03499389, 32'sh034801f1, 32'sh03467059, 32'sh0344dec0, 32'sh03434d26, 32'sh0341bb8c, 32'sh034029f2, 32'sh033e9856, 
               32'sh033d06bb, 32'sh033b751f, 32'sh0339e382, 32'sh033851e5, 32'sh0336c047, 32'sh03352ea9, 32'sh03339d0b, 32'sh03320b6c, 
               32'sh033079cc, 32'sh032ee82c, 32'sh032d568c, 32'sh032bc4eb, 32'sh032a3349, 32'sh0328a1a7, 32'sh03271005, 32'sh03257e62, 
               32'sh0323ecbe, 32'sh03225b1a, 32'sh0320c976, 32'sh031f37d1, 32'sh031da62b, 32'sh031c1486, 32'sh031a82df, 32'sh0318f138, 
               32'sh03175f91, 32'sh0315cde9, 32'sh03143c41, 32'sh0312aa98, 32'sh031118ef, 32'sh030f8745, 32'sh030df59b, 32'sh030c63f1, 
               32'sh030ad245, 32'sh0309409a, 32'sh0307aeee, 32'sh03061d41, 32'sh03048b94, 32'sh0302f9e7, 32'sh03016839, 32'sh02ffd68b, 
               32'sh02fe44dc, 32'sh02fcb32d, 32'sh02fb217d, 32'sh02f98fcd, 32'sh02f7fe1c, 32'sh02f66c6b, 32'sh02f4dab9, 32'sh02f34907, 
               32'sh02f1b755, 32'sh02f025a2, 32'sh02ee93ee, 32'sh02ed023a, 32'sh02eb7086, 32'sh02e9ded1, 32'sh02e84d1c, 32'sh02e6bb67, 
               32'sh02e529b0, 32'sh02e397fa, 32'sh02e20643, 32'sh02e0748c, 32'sh02dee2d4, 32'sh02dd511b, 32'sh02dbbf63, 32'sh02da2da9, 
               32'sh02d89bf0, 32'sh02d70a36, 32'sh02d5787b, 32'sh02d3e6c0, 32'sh02d25505, 32'sh02d0c349, 32'sh02cf318d, 32'sh02cd9fd0, 
               32'sh02cc0e13, 32'sh02ca7c55, 32'sh02c8ea97, 32'sh02c758d9, 32'sh02c5c71a, 32'sh02c4355b, 32'sh02c2a39b, 32'sh02c111db, 
               32'sh02bf801a, 32'sh02bdee59, 32'sh02bc5c98, 32'sh02bacad6, 32'sh02b93914, 32'sh02b7a751, 32'sh02b6158e, 32'sh02b483cb, 
               32'sh02b2f207, 32'sh02b16042, 32'sh02afce7e, 32'sh02ae3cb8, 32'sh02acaaf3, 32'sh02ab192d, 32'sh02a98766, 32'sh02a7f5a0, 
               32'sh02a663d8, 32'sh02a4d211, 32'sh02a34049, 32'sh02a1ae80, 32'sh02a01cb8, 32'sh029e8aee, 32'sh029cf925, 32'sh029b675b, 
               32'sh0299d590, 32'sh029843c5, 32'sh0296b1fa, 32'sh0295202e, 32'sh02938e62, 32'sh0291fc96, 32'sh02906ac9, 32'sh028ed8fc, 
               32'sh028d472e, 32'sh028bb560, 32'sh028a2392, 32'sh028891c3, 32'sh0286fff3, 32'sh02856e24, 32'sh0283dc54, 32'sh02824a84, 
               32'sh0280b8b3, 32'sh027f26e2, 32'sh027d9510, 32'sh027c033e, 32'sh027a716c, 32'sh0278df99, 32'sh02774dc6, 32'sh0275bbf3, 
               32'sh02742a1f, 32'sh0272984b, 32'sh02710676, 32'sh026f74a1, 32'sh026de2cc, 32'sh026c50f6, 32'sh026abf20, 32'sh02692d49, 
               32'sh02679b73, 32'sh0266099b, 32'sh026477c4, 32'sh0262e5ec, 32'sh02615414, 32'sh025fc23b, 32'sh025e3062, 32'sh025c9e88, 
               32'sh025b0caf, 32'sh02597ad5, 32'sh0257e8fa, 32'sh0256571f, 32'sh0254c544, 32'sh02533368, 32'sh0251a18c, 32'sh02500fb0, 
               32'sh024e7dd4, 32'sh024cebf7, 32'sh024b5a19, 32'sh0249c83b, 32'sh0248365d, 32'sh0246a47f, 32'sh024512a0, 32'sh024380c1, 
               32'sh0241eee2, 32'sh02405d02, 32'sh023ecb22, 32'sh023d3941, 32'sh023ba760, 32'sh023a157f, 32'sh0238839e, 32'sh0236f1bc, 
               32'sh02355fd9, 32'sh0233cdf7, 32'sh02323c14, 32'sh0230aa31, 32'sh022f184d, 32'sh022d8669, 32'sh022bf485, 32'sh022a62a0, 
               32'sh0228d0bb, 32'sh02273ed6, 32'sh0225acf1, 32'sh02241b0b, 32'sh02228924, 32'sh0220f73e, 32'sh021f6557, 32'sh021dd370, 
               32'sh021c4188, 32'sh021aafa0, 32'sh02191db8, 32'sh02178bcf, 32'sh0215f9e7, 32'sh021467fd, 32'sh0212d614, 32'sh0211442a, 
               32'sh020fb240, 32'sh020e2055, 32'sh020c8e6b, 32'sh020afc80, 32'sh02096a94, 32'sh0207d8a8, 32'sh020646bc, 32'sh0204b4d0, 
               32'sh020322e3, 32'sh020190f6, 32'sh01ffff09, 32'sh01fe6d1c, 32'sh01fcdb2e, 32'sh01fb4940, 32'sh01f9b751, 32'sh01f82562, 
               32'sh01f69373, 32'sh01f50184, 32'sh01f36f94, 32'sh01f1dda4, 32'sh01f04bb4, 32'sh01eeb9c3, 32'sh01ed27d2, 32'sh01eb95e1, 
               32'sh01ea03ef, 32'sh01e871fe, 32'sh01e6e00b, 32'sh01e54e19, 32'sh01e3bc26, 32'sh01e22a33, 32'sh01e09840, 32'sh01df064d, 
               32'sh01dd7459, 32'sh01dbe265, 32'sh01da5070, 32'sh01d8be7c, 32'sh01d72c87, 32'sh01d59a91, 32'sh01d4089c, 32'sh01d276a6, 
               32'sh01d0e4b0, 32'sh01cf52b9, 32'sh01cdc0c3, 32'sh01cc2ecc, 32'sh01ca9cd4, 32'sh01c90add, 32'sh01c778e5, 32'sh01c5e6ed, 
               32'sh01c454f5, 32'sh01c2c2fc, 32'sh01c13103, 32'sh01bf9f0a, 32'sh01be0d11, 32'sh01bc7b17, 32'sh01bae91d, 32'sh01b95723, 
               32'sh01b7c528, 32'sh01b6332e, 32'sh01b4a133, 32'sh01b30f37, 32'sh01b17d3c, 32'sh01afeb40, 32'sh01ae5944, 32'sh01acc748, 
               32'sh01ab354b, 32'sh01a9a34e, 32'sh01a81151, 32'sh01a67f54, 32'sh01a4ed56, 32'sh01a35b58, 32'sh01a1c95a, 32'sh01a0375c, 
               32'sh019ea55d, 32'sh019d135e, 32'sh019b815f, 32'sh0199ef60, 32'sh01985d60, 32'sh0196cb60, 32'sh01953960, 32'sh0193a760, 
               32'sh0192155f, 32'sh0190835f, 32'sh018ef15e, 32'sh018d5f5c, 32'sh018bcd5b, 32'sh018a3b59, 32'sh0188a957, 32'sh01871755, 
               32'sh01858552, 32'sh0183f34f, 32'sh0182614c, 32'sh0180cf49, 32'sh017f3d46, 32'sh017dab42, 32'sh017c193e, 32'sh017a873a, 
               32'sh0178f536, 32'sh01776331, 32'sh0175d12c, 32'sh01743f27, 32'sh0172ad22, 32'sh01711b1d, 32'sh016f8917, 32'sh016df711, 
               32'sh016c650b, 32'sh016ad305, 32'sh016940fe, 32'sh0167aef7, 32'sh01661cf0, 32'sh01648ae9, 32'sh0162f8e2, 32'sh016166da, 
               32'sh015fd4d2, 32'sh015e42ca, 32'sh015cb0c2, 32'sh015b1eb9, 32'sh01598cb1, 32'sh0157faa8, 32'sh0156689f, 32'sh0154d695, 
               32'sh0153448c, 32'sh0151b282, 32'sh01502078, 32'sh014e8e6e, 32'sh014cfc63, 32'sh014b6a59, 32'sh0149d84e, 32'sh01484643, 
               32'sh0146b438, 32'sh0145222d, 32'sh01439021, 32'sh0141fe16, 32'sh01406c0a, 32'sh013ed9fd, 32'sh013d47f1, 32'sh013bb5e5, 
               32'sh013a23d8, 32'sh013891cb, 32'sh0136ffbe, 32'sh01356db1, 32'sh0133dba3, 32'sh01324996, 32'sh0130b788, 32'sh012f257a, 
               32'sh012d936c, 32'sh012c015d, 32'sh012a6f4f, 32'sh0128dd40, 32'sh01274b31, 32'sh0125b922, 32'sh01242713, 32'sh01229503, 
               32'sh012102f4, 32'sh011f70e4, 32'sh011dded4, 32'sh011c4cc4, 32'sh011abab4, 32'sh011928a3, 32'sh01179693, 32'sh01160482, 
               32'sh01147271, 32'sh0112e060, 32'sh01114e4e, 32'sh010fbc3d, 32'sh010e2a2b, 32'sh010c981a, 32'sh010b0608, 32'sh010973f5, 
               32'sh0107e1e3, 32'sh01064fd1, 32'sh0104bdbe, 32'sh01032bab, 32'sh01019998, 32'sh01000785, 32'sh00fe7572, 32'sh00fce35f, 
               32'sh00fb514b, 32'sh00f9bf38, 32'sh00f82d24, 32'sh00f69b10, 32'sh00f508fc, 32'sh00f376e7, 32'sh00f1e4d3, 32'sh00f052bf, 
               32'sh00eec0aa, 32'sh00ed2e95, 32'sh00eb9c80, 32'sh00ea0a6b, 32'sh00e87856, 32'sh00e6e640, 32'sh00e5542b, 32'sh00e3c215, 
               32'sh00e22fff, 32'sh00e09de9, 32'sh00df0bd3, 32'sh00dd79bd, 32'sh00dbe7a6, 32'sh00da5590, 32'sh00d8c379, 32'sh00d73162, 
               32'sh00d59f4c, 32'sh00d40d35, 32'sh00d27b1d, 32'sh00d0e906, 32'sh00cf56ef, 32'sh00cdc4d7, 32'sh00cc32c0, 32'sh00caa0a8, 
               32'sh00c90e90, 32'sh00c77c78, 32'sh00c5ea60, 32'sh00c45847, 32'sh00c2c62f, 32'sh00c13417, 32'sh00bfa1fe, 32'sh00be0fe5, 
               32'sh00bc7dcc, 32'sh00baebb4, 32'sh00b9599a, 32'sh00b7c781, 32'sh00b63568, 32'sh00b4a34f, 32'sh00b31135, 32'sh00b17f1b, 
               32'sh00afed02, 32'sh00ae5ae8, 32'sh00acc8ce, 32'sh00ab36b4, 32'sh00a9a49a, 32'sh00a81280, 32'sh00a68065, 32'sh00a4ee4b, 
               32'sh00a35c30, 32'sh00a1ca16, 32'sh00a037fb, 32'sh009ea5e0, 32'sh009d13c5, 32'sh009b81aa, 32'sh0099ef8f, 32'sh00985d74, 
               32'sh0096cb58, 32'sh0095393d, 32'sh0093a722, 32'sh00921506, 32'sh009082ea, 32'sh008ef0cf, 32'sh008d5eb3, 32'sh008bcc97, 
               32'sh008a3a7b, 32'sh0088a85f, 32'sh00871643, 32'sh00858426, 32'sh0083f20a, 32'sh00825fee, 32'sh0080cdd1, 32'sh007f3bb5, 
               32'sh007da998, 32'sh007c177b, 32'sh007a855e, 32'sh0078f342, 32'sh00776125, 32'sh0075cf08, 32'sh00743cea, 32'sh0072aacd, 
               32'sh007118b0, 32'sh006f8693, 32'sh006df475, 32'sh006c6258, 32'sh006ad03b, 32'sh00693e1d, 32'sh0067abff, 32'sh006619e2, 
               32'sh006487c4, 32'sh0062f5a6, 32'sh00616388, 32'sh005fd16a, 32'sh005e3f4c, 32'sh005cad2e, 32'sh005b1b10, 32'sh005988f2, 
               32'sh0057f6d4, 32'sh005664b6, 32'sh0054d297, 32'sh00534079, 32'sh0051ae5b, 32'sh00501c3c, 32'sh004e8a1e, 32'sh004cf7ff, 
               32'sh004b65e1, 32'sh0049d3c2, 32'sh004841a3, 32'sh0046af84, 32'sh00451d66, 32'sh00438b47, 32'sh0041f928, 32'sh00406709, 
               32'sh003ed4ea, 32'sh003d42cb, 32'sh003bb0ac, 32'sh003a1e8d, 32'sh00388c6e, 32'sh0036fa4f, 32'sh00356830, 32'sh0033d611, 
               32'sh003243f1, 32'sh0030b1d2, 32'sh002f1fb3, 32'sh002d8d94, 32'sh002bfb74, 32'sh002a6955, 32'sh0028d736, 32'sh00274516, 
               32'sh0025b2f7, 32'sh002420d7, 32'sh00228eb8, 32'sh0020fc98, 32'sh001f6a79, 32'sh001dd859, 32'sh001c463a, 32'sh001ab41a, 
               32'sh001921fb, 32'sh00178fdb, 32'sh0015fdbb, 32'sh00146b9c, 32'sh0012d97c, 32'sh0011475d, 32'sh000fb53d, 32'sh000e231d, 
               32'sh000c90fe, 32'sh000afede, 32'sh00096cbe, 32'sh0007da9f, 32'sh0006487f, 32'sh0004b65f, 32'sh0003243f, 32'sh00019220, 
               32'sh00000000, 32'shfffe6de0, 32'shfffcdbc1, 32'shfffb49a1, 32'shfff9b781, 32'shfff82561, 32'shfff69342, 32'shfff50122, 
               32'shfff36f02, 32'shfff1dce3, 32'shfff04ac3, 32'shffeeb8a3, 32'shffed2684, 32'shffeb9464, 32'shffea0245, 32'shffe87025, 
               32'shffe6de05, 32'shffe54be6, 32'shffe3b9c6, 32'shffe227a7, 32'shffe09587, 32'shffdf0368, 32'shffdd7148, 32'shffdbdf29, 
               32'shffda4d09, 32'shffd8baea, 32'shffd728ca, 32'shffd596ab, 32'shffd4048c, 32'shffd2726c, 32'shffd0e04d, 32'shffcf4e2e, 
               32'shffcdbc0f, 32'shffcc29ef, 32'shffca97d0, 32'shffc905b1, 32'shffc77392, 32'shffc5e173, 32'shffc44f54, 32'shffc2bd35, 
               32'shffc12b16, 32'shffbf98f7, 32'shffbe06d8, 32'shffbc74b9, 32'shffbae29a, 32'shffb9507c, 32'shffb7be5d, 32'shffb62c3e, 
               32'shffb49a1f, 32'shffb30801, 32'shffb175e2, 32'shffafe3c4, 32'shffae51a5, 32'shffacbf87, 32'shffab2d69, 32'shffa99b4a, 
               32'shffa8092c, 32'shffa6770e, 32'shffa4e4f0, 32'shffa352d2, 32'shffa1c0b4, 32'shffa02e96, 32'shff9e9c78, 32'shff9d0a5a, 
               32'shff9b783c, 32'shff99e61e, 32'shff985401, 32'shff96c1e3, 32'shff952fc5, 32'shff939da8, 32'shff920b8b, 32'shff90796d, 
               32'shff8ee750, 32'shff8d5533, 32'shff8bc316, 32'shff8a30f8, 32'shff889edb, 32'shff870cbe, 32'shff857aa2, 32'shff83e885, 
               32'shff825668, 32'shff80c44b, 32'shff7f322f, 32'shff7da012, 32'shff7c0df6, 32'shff7a7bda, 32'shff78e9bd, 32'shff7757a1, 
               32'shff75c585, 32'shff743369, 32'shff72a14d, 32'shff710f31, 32'shff6f7d16, 32'shff6deafa, 32'shff6c58de, 32'shff6ac6c3, 
               32'shff6934a8, 32'shff67a28c, 32'shff661071, 32'shff647e56, 32'shff62ec3b, 32'shff615a20, 32'shff5fc805, 32'shff5e35ea, 
               32'shff5ca3d0, 32'shff5b11b5, 32'shff597f9b, 32'shff57ed80, 32'shff565b66, 32'shff54c94c, 32'shff533732, 32'shff51a518, 
               32'shff5012fe, 32'shff4e80e5, 32'shff4ceecb, 32'shff4b5cb1, 32'shff49ca98, 32'shff48387f, 32'shff46a666, 32'shff45144c, 
               32'shff438234, 32'shff41f01b, 32'shff405e02, 32'shff3ecbe9, 32'shff3d39d1, 32'shff3ba7b9, 32'shff3a15a0, 32'shff388388, 
               32'shff36f170, 32'shff355f58, 32'shff33cd40, 32'shff323b29, 32'shff30a911, 32'shff2f16fa, 32'shff2d84e3, 32'shff2bf2cb, 
               32'shff2a60b4, 32'shff28ce9e, 32'shff273c87, 32'shff25aa70, 32'shff24185a, 32'shff228643, 32'shff20f42d, 32'shff1f6217, 
               32'shff1dd001, 32'shff1c3deb, 32'shff1aabd5, 32'shff1919c0, 32'shff1787aa, 32'shff15f595, 32'shff146380, 32'shff12d16b, 
               32'shff113f56, 32'shff0fad41, 32'shff0e1b2d, 32'shff0c8919, 32'shff0af704, 32'shff0964f0, 32'shff07d2dc, 32'shff0640c8, 
               32'shff04aeb5, 32'shff031ca1, 32'shff018a8e, 32'shfefff87b, 32'shfefe6668, 32'shfefcd455, 32'shfefb4242, 32'shfef9b02f, 
               32'shfef81e1d, 32'shfef68c0b, 32'shfef4f9f8, 32'shfef367e6, 32'shfef1d5d5, 32'shfef043c3, 32'shfeeeb1b2, 32'shfeed1fa0, 
               32'shfeeb8d8f, 32'shfee9fb7e, 32'shfee8696d, 32'shfee6d75d, 32'shfee5454c, 32'shfee3b33c, 32'shfee2212c, 32'shfee08f1c, 
               32'shfedefd0c, 32'shfedd6afd, 32'shfedbd8ed, 32'shfeda46de, 32'shfed8b4cf, 32'shfed722c0, 32'shfed590b1, 32'shfed3fea3, 
               32'shfed26c94, 32'shfed0da86, 32'shfecf4878, 32'shfecdb66a, 32'shfecc245d, 32'shfeca924f, 32'shfec90042, 32'shfec76e35, 
               32'shfec5dc28, 32'shfec44a1b, 32'shfec2b80f, 32'shfec12603, 32'shfebf93f6, 32'shfebe01ea, 32'shfebc6fdf, 32'shfebaddd3, 
               32'shfeb94bc8, 32'shfeb7b9bd, 32'shfeb627b2, 32'shfeb495a7, 32'shfeb3039d, 32'shfeb17192, 32'shfeafdf88, 32'shfeae4d7e, 
               32'shfeacbb74, 32'shfeab296b, 32'shfea99761, 32'shfea80558, 32'shfea6734f, 32'shfea4e147, 32'shfea34f3e, 32'shfea1bd36, 
               32'shfea02b2e, 32'shfe9e9926, 32'shfe9d071e, 32'shfe9b7517, 32'shfe99e310, 32'shfe985109, 32'shfe96bf02, 32'shfe952cfb, 
               32'shfe939af5, 32'shfe9208ef, 32'shfe9076e9, 32'shfe8ee4e3, 32'shfe8d52de, 32'shfe8bc0d9, 32'shfe8a2ed4, 32'shfe889ccf, 
               32'shfe870aca, 32'shfe8578c6, 32'shfe83e6c2, 32'shfe8254be, 32'shfe80c2ba, 32'shfe7f30b7, 32'shfe7d9eb4, 32'shfe7c0cb1, 
               32'shfe7a7aae, 32'shfe78e8ab, 32'shfe7756a9, 32'shfe75c4a7, 32'shfe7432a5, 32'shfe72a0a4, 32'shfe710ea2, 32'shfe6f7ca1, 
               32'shfe6deaa1, 32'shfe6c58a0, 32'shfe6ac6a0, 32'shfe6934a0, 32'shfe67a2a0, 32'shfe6610a0, 32'shfe647ea1, 32'shfe62eca2, 
               32'shfe615aa3, 32'shfe5fc8a4, 32'shfe5e36a6, 32'shfe5ca4a8, 32'shfe5b12aa, 32'shfe5980ac, 32'shfe57eeaf, 32'shfe565cb2, 
               32'shfe54cab5, 32'shfe5338b8, 32'shfe51a6bc, 32'shfe5014c0, 32'shfe4e82c4, 32'shfe4cf0c9, 32'shfe4b5ecd, 32'shfe49ccd2, 
               32'shfe483ad8, 32'shfe46a8dd, 32'shfe4516e3, 32'shfe4384e9, 32'shfe41f2ef, 32'shfe4060f6, 32'shfe3ecefd, 32'shfe3d3d04, 
               32'shfe3bab0b, 32'shfe3a1913, 32'shfe38871b, 32'shfe36f523, 32'shfe35632c, 32'shfe33d134, 32'shfe323f3d, 32'shfe30ad47, 
               32'shfe2f1b50, 32'shfe2d895a, 32'shfe2bf764, 32'shfe2a656f, 32'shfe28d379, 32'shfe274184, 32'shfe25af90, 32'shfe241d9b, 
               32'shfe228ba7, 32'shfe20f9b3, 32'shfe1f67c0, 32'shfe1dd5cd, 32'shfe1c43da, 32'shfe1ab1e7, 32'shfe191ff5, 32'shfe178e02, 
               32'shfe15fc11, 32'shfe146a1f, 32'shfe12d82e, 32'shfe11463d, 32'shfe0fb44c, 32'shfe0e225c, 32'shfe0c906c, 32'shfe0afe7c, 
               32'shfe096c8d, 32'shfe07da9e, 32'shfe0648af, 32'shfe04b6c0, 32'shfe0324d2, 32'shfe0192e4, 32'shfe0000f7, 32'shfdfe6f0a, 
               32'shfdfcdd1d, 32'shfdfb4b30, 32'shfdf9b944, 32'shfdf82758, 32'shfdf6956c, 32'shfdf50380, 32'shfdf37195, 32'shfdf1dfab, 
               32'shfdf04dc0, 32'shfdeebbd6, 32'shfded29ec, 32'shfdeb9803, 32'shfdea0619, 32'shfde87431, 32'shfde6e248, 32'shfde55060, 
               32'shfde3be78, 32'shfde22c90, 32'shfde09aa9, 32'shfddf08c2, 32'shfddd76dc, 32'shfddbe4f5, 32'shfdda530f, 32'shfdd8c12a, 
               32'shfdd72f45, 32'shfdd59d60, 32'shfdd40b7b, 32'shfdd27997, 32'shfdd0e7b3, 32'shfdcf55cf, 32'shfdcdc3ec, 32'shfdcc3209, 
               32'shfdcaa027, 32'shfdc90e44, 32'shfdc77c62, 32'shfdc5ea81, 32'shfdc458a0, 32'shfdc2c6bf, 32'shfdc134de, 32'shfdbfa2fe, 
               32'shfdbe111e, 32'shfdbc7f3f, 32'shfdbaed60, 32'shfdb95b81, 32'shfdb7c9a3, 32'shfdb637c5, 32'shfdb4a5e7, 32'shfdb31409, 
               32'shfdb1822c, 32'shfdaff050, 32'shfdae5e74, 32'shfdaccc98, 32'shfdab3abc, 32'shfda9a8e1, 32'shfda81706, 32'shfda6852b, 
               32'shfda4f351, 32'shfda36178, 32'shfda1cf9e, 32'shfda03dc5, 32'shfd9eabec, 32'shfd9d1a14, 32'shfd9b883c, 32'shfd99f665, 
               32'shfd98648d, 32'shfd96d2b7, 32'shfd9540e0, 32'shfd93af0a, 32'shfd921d34, 32'shfd908b5f, 32'shfd8ef98a, 32'shfd8d67b5, 
               32'shfd8bd5e1, 32'shfd8a440d, 32'shfd88b23a, 32'shfd872067, 32'shfd858e94, 32'shfd83fcc2, 32'shfd826af0, 32'shfd80d91e, 
               32'shfd7f474d, 32'shfd7db57c, 32'shfd7c23ac, 32'shfd7a91dc, 32'shfd79000d, 32'shfd776e3d, 32'shfd75dc6e, 32'shfd744aa0, 
               32'shfd72b8d2, 32'shfd712704, 32'shfd6f9537, 32'shfd6e036a, 32'shfd6c719e, 32'shfd6adfd2, 32'shfd694e06, 32'shfd67bc3b, 
               32'shfd662a70, 32'shfd6498a5, 32'shfd6306db, 32'shfd617512, 32'shfd5fe348, 32'shfd5e5180, 32'shfd5cbfb7, 32'shfd5b2def, 
               32'shfd599c28, 32'shfd580a60, 32'shfd56789a, 32'shfd54e6d3, 32'shfd53550d, 32'shfd51c348, 32'shfd503182, 32'shfd4e9fbe, 
               32'shfd4d0df9, 32'shfd4b7c35, 32'shfd49ea72, 32'shfd4858af, 32'shfd46c6ec, 32'shfd45352a, 32'shfd43a368, 32'shfd4211a7, 
               32'shfd407fe6, 32'shfd3eee25, 32'shfd3d5c65, 32'shfd3bcaa5, 32'shfd3a38e6, 32'shfd38a727, 32'shfd371569, 32'shfd3583ab, 
               32'shfd33f1ed, 32'shfd326030, 32'shfd30ce73, 32'shfd2f3cb7, 32'shfd2daafb, 32'shfd2c1940, 32'shfd2a8785, 32'shfd28f5ca, 
               32'shfd276410, 32'shfd25d257, 32'shfd24409d, 32'shfd22aee5, 32'shfd211d2c, 32'shfd1f8b74, 32'shfd1df9bd, 32'shfd1c6806, 
               32'shfd1ad650, 32'shfd194499, 32'shfd17b2e4, 32'shfd16212f, 32'shfd148f7a, 32'shfd12fdc6, 32'shfd116c12, 32'shfd0fda5e, 
               32'shfd0e48ab, 32'shfd0cb6f9, 32'shfd0b2547, 32'shfd099395, 32'shfd0801e4, 32'shfd067033, 32'shfd04de83, 32'shfd034cd3, 
               32'shfd01bb24, 32'shfd002975, 32'shfcfe97c7, 32'shfcfd0619, 32'shfcfb746c, 32'shfcf9e2bf, 32'shfcf85112, 32'shfcf6bf66, 
               32'shfcf52dbb, 32'shfcf39c0f, 32'shfcf20a65, 32'shfcf078bb, 32'shfceee711, 32'shfced5568, 32'shfcebc3bf, 32'shfcea3217, 
               32'shfce8a06f, 32'shfce70ec8, 32'shfce57d21, 32'shfce3eb7a, 32'shfce259d5, 32'shfce0c82f, 32'shfcdf368a, 32'shfcdda4e6, 
               32'shfcdc1342, 32'shfcda819e, 32'shfcd8effb, 32'shfcd75e59, 32'shfcd5ccb7, 32'shfcd43b15, 32'shfcd2a974, 32'shfcd117d4, 
               32'shfccf8634, 32'shfccdf494, 32'shfccc62f5, 32'shfccad157, 32'shfcc93fb9, 32'shfcc7ae1b, 32'shfcc61c7e, 32'shfcc48ae1, 
               32'shfcc2f945, 32'shfcc167aa, 32'shfcbfd60e, 32'shfcbe4474, 32'shfcbcb2da, 32'shfcbb2140, 32'shfcb98fa7, 32'shfcb7fe0f, 
               32'shfcb66c77, 32'shfcb4dadf, 32'shfcb34948, 32'shfcb1b7b1, 32'shfcb0261b, 32'shfcae9486, 32'shfcad02f1, 32'shfcab715c, 
               32'shfca9dfc8, 32'shfca84e35, 32'shfca6bca2, 32'shfca52b0f, 32'shfca3997e, 32'shfca207ec, 32'shfca0765b, 32'shfc9ee4cb, 
               32'shfc9d533b, 32'shfc9bc1ac, 32'shfc9a301d, 32'shfc989e8f, 32'shfc970d01, 32'shfc957b74, 32'shfc93e9e7, 32'shfc92585b, 
               32'shfc90c6cf, 32'shfc8f3544, 32'shfc8da3ba, 32'shfc8c122f, 32'shfc8a80a6, 32'shfc88ef1d, 32'shfc875d95, 32'shfc85cc0d, 
               32'shfc843a85, 32'shfc82a8fe, 32'shfc811778, 32'shfc7f85f2, 32'shfc7df46d, 32'shfc7c62e8, 32'shfc7ad164, 32'shfc793fe1, 
               32'shfc77ae5e, 32'shfc761cdb, 32'shfc748b59, 32'shfc72f9d8, 32'shfc716857, 32'shfc6fd6d7, 32'shfc6e4557, 32'shfc6cb3d8, 
               32'shfc6b2259, 32'shfc6990db, 32'shfc67ff5d, 32'shfc666de0, 32'shfc64dc64, 32'shfc634ae8, 32'shfc61b96d, 32'shfc6027f2, 
               32'shfc5e9678, 32'shfc5d04fe, 32'shfc5b7385, 32'shfc59e20c, 32'shfc585094, 32'shfc56bf1d, 32'shfc552da6, 32'shfc539c30, 
               32'shfc520aba, 32'shfc507945, 32'shfc4ee7d0, 32'shfc4d565c, 32'shfc4bc4e9, 32'shfc4a3376, 32'shfc48a204, 32'shfc471092, 
               32'shfc457f21, 32'shfc43edb0, 32'shfc425c40, 32'shfc40cad1, 32'shfc3f3962, 32'shfc3da7f4, 32'shfc3c1686, 32'shfc3a8519, 
               32'shfc38f3ac, 32'shfc376240, 32'shfc35d0d5, 32'shfc343f6a, 32'shfc32ae00, 32'shfc311c97, 32'shfc2f8b2e, 32'shfc2df9c5, 
               32'shfc2c685d, 32'shfc2ad6f6, 32'shfc29458f, 32'shfc27b429, 32'shfc2622c4, 32'shfc24915f, 32'shfc22fffb, 32'shfc216e97, 
               32'shfc1fdd34, 32'shfc1e4bd1, 32'shfc1cba6f, 32'shfc1b290e, 32'shfc1997ae, 32'shfc18064d, 32'shfc1674ee, 32'shfc14e38f, 
               32'shfc135231, 32'shfc11c0d3, 32'shfc102f76, 32'shfc0e9e1a, 32'shfc0d0cbe, 32'shfc0b7b62, 32'shfc09ea08, 32'shfc0858ae, 
               32'shfc06c754, 32'shfc0535fc, 32'shfc03a4a3, 32'shfc02134c, 32'shfc0081f5, 32'shfbfef09f, 32'shfbfd5f49, 32'shfbfbcdf4, 
               32'shfbfa3c9f, 32'shfbf8ab4b, 32'shfbf719f8, 32'shfbf588a5, 32'shfbf3f753, 32'shfbf26602, 32'shfbf0d4b1, 32'shfbef4361, 
               32'shfbedb212, 32'shfbec20c3, 32'shfbea8f75, 32'shfbe8fe27, 32'shfbe76cda, 32'shfbe5db8e, 32'shfbe44a42, 32'shfbe2b8f7, 
               32'shfbe127ac, 32'shfbdf9663, 32'shfbde0519, 32'shfbdc73d1, 32'shfbdae289, 32'shfbd95142, 32'shfbd7bffb, 32'shfbd62eb5, 
               32'shfbd49d70, 32'shfbd30c2b, 32'shfbd17ae7, 32'shfbcfe9a4, 32'shfbce5861, 32'shfbccc71f, 32'shfbcb35dd, 32'shfbc9a49d, 
               32'shfbc8135c, 32'shfbc6821d, 32'shfbc4f0de, 32'shfbc35fa0, 32'shfbc1ce62, 32'shfbc03d25, 32'shfbbeabe9, 32'shfbbd1aad, 
               32'shfbbb8973, 32'shfbb9f838, 32'shfbb866ff, 32'shfbb6d5c6, 32'shfbb5448d, 32'shfbb3b356, 32'shfbb2221f, 32'shfbb090e8, 
               32'shfbaeffb3, 32'shfbad6e7e, 32'shfbabdd49, 32'shfbaa4c16, 32'shfba8bae3, 32'shfba729b1, 32'shfba5987f, 32'shfba4074e, 
               32'shfba2761e, 32'shfba0e4ee, 32'shfb9f53bf, 32'shfb9dc291, 32'shfb9c3163, 32'shfb9aa036, 32'shfb990f0a, 32'shfb977ddf, 
               32'shfb95ecb4, 32'shfb945b89, 32'shfb92ca60, 32'shfb913937, 32'shfb8fa80f, 32'shfb8e16e7, 32'shfb8c85c1, 32'shfb8af49b, 
               32'shfb896375, 32'shfb87d250, 32'shfb86412c, 32'shfb84b009, 32'shfb831ee6, 32'shfb818dc4, 32'shfb7ffca3, 32'shfb7e6b83, 
               32'shfb7cda63, 32'shfb7b4944, 32'shfb79b825, 32'shfb782707, 32'shfb7695ea, 32'shfb7504ce, 32'shfb7373b2, 32'shfb71e297, 
               32'shfb70517d, 32'shfb6ec063, 32'shfb6d2f4a, 32'shfb6b9e32, 32'shfb6a0d1b, 32'shfb687c04, 32'shfb66eaee, 32'shfb6559d9, 
               32'shfb63c8c4, 32'shfb6237b0, 32'shfb60a69d, 32'shfb5f158a, 32'shfb5d8479, 32'shfb5bf368, 32'shfb5a6257, 32'shfb58d148, 
               32'shfb574039, 32'shfb55af2a, 32'shfb541e1d, 32'shfb528d10, 32'shfb50fc04, 32'shfb4f6af9, 32'shfb4dd9ee, 32'shfb4c48e4, 
               32'shfb4ab7db, 32'shfb4926d3, 32'shfb4795cb, 32'shfb4604c4, 32'shfb4473be, 32'shfb42e2b9, 32'shfb4151b4, 32'shfb3fc0b0, 
               32'shfb3e2fac, 32'shfb3c9eaa, 32'shfb3b0da8, 32'shfb397ca7, 32'shfb37eba7, 32'shfb365aa7, 32'shfb34c9a8, 32'shfb3338aa, 
               32'shfb31a7ac, 32'shfb3016b0, 32'shfb2e85b4, 32'shfb2cf4b9, 32'shfb2b63be, 32'shfb29d2c5, 32'shfb2841cc, 32'shfb26b0d3, 
               32'shfb251fdc, 32'shfb238ee5, 32'shfb21fdef, 32'shfb206cfa, 32'shfb1edc06, 32'shfb1d4b12, 32'shfb1bba1f, 32'shfb1a292d, 
               32'shfb18983b, 32'shfb17074b, 32'shfb15765b, 32'shfb13e56c, 32'shfb12547d, 32'shfb10c38f, 32'shfb0f32a3, 32'shfb0da1b6, 
               32'shfb0c10cb, 32'shfb0a7fe1, 32'shfb08eef7, 32'shfb075e0e, 32'shfb05cd25, 32'shfb043c3e, 32'shfb02ab57, 32'shfb011a71, 
               32'shfaff898c, 32'shfafdf8a7, 32'shfafc67c4, 32'shfafad6e1, 32'shfaf945ff, 32'shfaf7b51d, 32'shfaf6243d, 32'shfaf4935d, 
               32'shfaf3027e, 32'shfaf171a0, 32'shfaefe0c2, 32'shfaee4fe5, 32'shfaecbf0a, 32'shfaeb2e2e, 32'shfae99d54, 32'shfae80c7a, 
               32'shfae67ba2, 32'shfae4eaca, 32'shfae359f3, 32'shfae1c91c, 32'shfae03847, 32'shfadea772, 32'shfadd169e, 32'shfadb85ca, 
               32'shfad9f4f8, 32'shfad86426, 32'shfad6d355, 32'shfad54285, 32'shfad3b1b6, 32'shfad220e8, 32'shfad0901a, 32'shfaceff4d, 
               32'shfacd6e81, 32'shfacbddb6, 32'shfaca4ceb, 32'shfac8bc22, 32'shfac72b59, 32'shfac59a91, 32'shfac409c9, 32'shfac27903, 
               32'shfac0e83d, 32'shfabf5778, 32'shfabdc6b4, 32'shfabc35f1, 32'shfabaa52f, 32'shfab9146d, 32'shfab783ad, 32'shfab5f2ed, 
               32'shfab4622d, 32'shfab2d16f, 32'shfab140b2, 32'shfaafaff5, 32'shfaae1f39, 32'shfaac8e7e, 32'shfaaafdc4, 32'shfaa96d0a, 
               32'shfaa7dc52, 32'shfaa64b9a, 32'shfaa4bae3, 32'shfaa32a2d, 32'shfaa19978, 32'shfaa008c3, 32'shfa9e7810, 32'shfa9ce75d, 
               32'shfa9b56ab, 32'shfa99c5fa, 32'shfa98354a, 32'shfa96a49a, 32'shfa9513eb, 32'shfa93833e, 32'shfa91f291, 32'shfa9061e5, 
               32'shfa8ed139, 32'shfa8d408f, 32'shfa8bafe5, 32'shfa8a1f3c, 32'shfa888e95, 32'shfa86fded, 32'shfa856d47, 32'shfa83dca2, 
               32'shfa824bfd, 32'shfa80bb5a, 32'shfa7f2ab7, 32'shfa7d9a15, 32'shfa7c0974, 32'shfa7a78d3, 32'shfa78e834, 32'shfa775795, 
               32'shfa75c6f8, 32'shfa74365b, 32'shfa72a5bf, 32'shfa711524, 32'shfa6f8489, 32'shfa6df3f0, 32'shfa6c6357, 32'shfa6ad2bf, 
               32'shfa694229, 32'shfa67b193, 32'shfa6620fd, 32'shfa649069, 32'shfa62ffd6, 32'shfa616f43, 32'shfa5fdeb1, 32'shfa5e4e21, 
               32'shfa5cbd91, 32'shfa5b2d02, 32'shfa599c73, 32'shfa580be6, 32'shfa567b5a, 32'shfa54eace, 32'shfa535a43, 32'shfa51c9b9, 
               32'shfa503930, 32'shfa4ea8a8, 32'shfa4d1821, 32'shfa4b879b, 32'shfa49f715, 32'shfa486691, 32'shfa46d60d, 32'shfa45458a, 
               32'shfa43b508, 32'shfa422487, 32'shfa409407, 32'shfa3f0388, 32'shfa3d7309, 32'shfa3be28c, 32'shfa3a520f, 32'shfa38c194, 
               32'shfa373119, 32'shfa35a09f, 32'shfa341026, 32'shfa327fae, 32'shfa30ef36, 32'shfa2f5ec0, 32'shfa2dce4b, 32'shfa2c3dd6, 
               32'shfa2aad62, 32'shfa291cf0, 32'shfa278c7e, 32'shfa25fc0d, 32'shfa246b9d, 32'shfa22db2d, 32'shfa214abf, 32'shfa1fba52, 
               32'shfa1e29e5, 32'shfa1c997a, 32'shfa1b090f, 32'shfa1978a6, 32'shfa17e83d, 32'shfa1657d5, 32'shfa14c76e, 32'shfa133708, 
               32'shfa11a6a3, 32'shfa10163e, 32'shfa0e85db, 32'shfa0cf579, 32'shfa0b6517, 32'shfa09d4b7, 32'shfa084457, 32'shfa06b3f8, 
               32'shfa05239a, 32'shfa03933d, 32'shfa0202e1, 32'shfa007286, 32'shf9fee22c, 32'shf9fd51d3, 32'shf9fbc17b, 32'shf9fa3123, 
               32'shf9f8a0cd, 32'shf9f71078, 32'shf9f58023, 32'shf9f3efcf, 32'shf9f25f7d, 32'shf9f0cf2b, 32'shf9ef3eda, 32'shf9edae8a, 
               32'shf9ec1e3b, 32'shf9ea8ded, 32'shf9e8fda0, 32'shf9e76d54, 32'shf9e5dd09, 32'shf9e44cbf, 32'shf9e2bc75, 32'shf9e12c2d, 
               32'shf9df9be6, 32'shf9de0b9f, 32'shf9dc7b5a, 32'shf9daeb15, 32'shf9d95ad1, 32'shf9d7ca8f, 32'shf9d63a4d, 32'shf9d4aa0c, 
               32'shf9d319cc, 32'shf9d1898d, 32'shf9cff94f, 32'shf9ce6912, 32'shf9ccd8d6, 32'shf9cb489b, 32'shf9c9b861, 32'shf9c82828, 
               32'shf9c697f0, 32'shf9c507b9, 32'shf9c37782, 32'shf9c1e74d, 32'shf9c05719, 32'shf9bec6e5, 32'shf9bd36b3, 32'shf9bba681, 
               32'shf9ba1651, 32'shf9b88621, 32'shf9b6f5f3, 32'shf9b565c5, 32'shf9b3d599, 32'shf9b2456d, 32'shf9b0b542, 32'shf9af2519, 
               32'shf9ad94f0, 32'shf9ac04c8, 32'shf9aa74a1, 32'shf9a8e47c, 32'shf9a75457, 32'shf9a5c433, 32'shf9a43410, 32'shf9a2a3ee, 
               32'shf9a113cd, 32'shf99f83ad, 32'shf99df38e, 32'shf99c6371, 32'shf99ad354, 32'shf9994338, 32'shf997b31d, 32'shf9962303, 
               32'shf99492ea, 32'shf99302d2, 32'shf99172bb, 32'shf98fe2a5, 32'shf98e528f, 32'shf98cc27b, 32'shf98b3268, 32'shf989a256, 
               32'shf9881245, 32'shf9868235, 32'shf984f226, 32'shf9836218, 32'shf981d20b, 32'shf98041ff, 32'shf97eb1f4, 32'shf97d21ea, 
               32'shf97b91e1, 32'shf97a01d9, 32'shf97871d2, 32'shf976e1cc, 32'shf97551c6, 32'shf973c1c2, 32'shf97231bf, 32'shf970a1bd, 
               32'shf96f11bc, 32'shf96d81bc, 32'shf96bf1be, 32'shf96a61c0, 32'shf968d1c3, 32'shf96741c7, 32'shf965b1cc, 32'shf96421d2, 
               32'shf96291d9, 32'shf96101e1, 32'shf95f71ea, 32'shf95de1f5, 32'shf95c5200, 32'shf95ac20c, 32'shf9593219, 32'shf957a228, 
               32'shf9561237, 32'shf9548247, 32'shf952f259, 32'shf951626b, 32'shf94fd27f, 32'shf94e4293, 32'shf94cb2a8, 32'shf94b22bf, 
               32'shf94992d7, 32'shf94802ef, 32'shf9467309, 32'shf944e323, 32'shf943533f, 32'shf941c35c, 32'shf940337a, 32'shf93ea399, 
               32'shf93d13b8, 32'shf93b83d9, 32'shf939f3fb, 32'shf938641e, 32'shf936d442, 32'shf9354468, 32'shf933b48e, 32'shf93224b5, 
               32'shf93094dd, 32'shf92f0506, 32'shf92d7531, 32'shf92be55c, 32'shf92a5589, 32'shf928c5b6, 32'shf92735e5, 32'shf925a614, 
               32'shf9241645, 32'shf9228677, 32'shf920f6a9, 32'shf91f66dd, 32'shf91dd712, 32'shf91c4748, 32'shf91ab77f, 32'shf91927b7, 
               32'shf91797f0, 32'shf916082b, 32'shf9147866, 32'shf912e8a2, 32'shf91158e0, 32'shf90fc91e, 32'shf90e395e, 32'shf90ca99e, 
               32'shf90b19e0, 32'shf9098a23, 32'shf907fa67, 32'shf9066aac, 32'shf904daf2, 32'shf9034b39, 32'shf901bb81, 32'shf9002bca, 
               32'shf8fe9c15, 32'shf8fd0c60, 32'shf8fb7cac, 32'shf8f9ecfa, 32'shf8f85d49, 32'shf8f6cd98, 32'shf8f53de9, 32'shf8f3ae3b, 
               32'shf8f21e8e, 32'shf8f08ee2, 32'shf8eeff37, 32'shf8ed6f8e, 32'shf8ebdfe5, 32'shf8ea503d, 32'shf8e8c097, 32'shf8e730f2, 
               32'shf8e5a14d, 32'shf8e411aa, 32'shf8e28208, 32'shf8e0f267, 32'shf8df62c7, 32'shf8ddd328, 32'shf8dc438b, 32'shf8dab3ee, 
               32'shf8d92452, 32'shf8d794b8, 32'shf8d6051f, 32'shf8d47587, 32'shf8d2e5f0, 32'shf8d1565a, 32'shf8cfc6c5, 32'shf8ce3731, 
               32'shf8cca79e, 32'shf8cb180d, 32'shf8c9887c, 32'shf8c7f8ed, 32'shf8c6695f, 32'shf8c4d9d2, 32'shf8c34a46, 32'shf8c1babb, 
               32'shf8c02b31, 32'shf8be9ba9, 32'shf8bd0c21, 32'shf8bb7c9b, 32'shf8b9ed15, 32'shf8b85d91, 32'shf8b6ce0e, 32'shf8b53e8c, 
               32'shf8b3af0c, 32'shf8b21f8c, 32'shf8b0900d, 32'shf8af0090, 32'shf8ad7114, 32'shf8abe199, 32'shf8aa521f, 32'shf8a8c2a6, 
               32'shf8a7332e, 32'shf8a5a3b8, 32'shf8a41442, 32'shf8a284ce, 32'shf8a0f55b, 32'shf89f65e8, 32'shf89dd678, 32'shf89c4708, 
               32'shf89ab799, 32'shf899282c, 32'shf89798bf, 32'shf8960954, 32'shf89479ea, 32'shf892ea81, 32'shf8915b19, 32'shf88fcbb3, 
               32'shf88e3c4d, 32'shf88cace9, 32'shf88b1d86, 32'shf8898e23, 32'shf887fec3, 32'shf8866f63, 32'shf884e004, 32'shf88350a7, 
               32'shf881c14b, 32'shf88031ef, 32'shf87ea295, 32'shf87d133d, 32'shf87b83e5, 32'shf879f48e, 32'shf8786539, 32'shf876d5e5, 
               32'shf8754692, 32'shf873b740, 32'shf87227ef, 32'shf87098a0, 32'shf86f0952, 32'shf86d7a04, 32'shf86beab8, 32'shf86a5b6d, 
               32'shf868cc24, 32'shf8673cdb, 32'shf865ad94, 32'shf8641e4e, 32'shf8628f09, 32'shf860ffc5, 32'shf85f7082, 32'shf85de141, 
               32'shf85c5201, 32'shf85ac2c1, 32'shf8593383, 32'shf857a447, 32'shf856150b, 32'shf85485d1, 32'shf852f698, 32'shf8516760, 
               32'shf84fd829, 32'shf84e48f3, 32'shf84cb9bf, 32'shf84b2a8b, 32'shf8499b59, 32'shf8480c28, 32'shf8467cf9, 32'shf844edca, 
               32'shf8435e9d, 32'shf841cf71, 32'shf8404046, 32'shf83eb11c, 32'shf83d21f3, 32'shf83b92cc, 32'shf83a03a6, 32'shf8387481, 
               32'shf836e55d, 32'shf835563b, 32'shf833c719, 32'shf83237f9, 32'shf830a8da, 32'shf82f19bc, 32'shf82d8aa0, 32'shf82bfb84, 
               32'shf82a6c6a, 32'shf828dd51, 32'shf8274e3a, 32'shf825bf23, 32'shf824300e, 32'shf822a0fa, 32'shf82111e7, 32'shf81f82d5, 
               32'shf81df3c5, 32'shf81c64b6, 32'shf81ad5a8, 32'shf819469b, 32'shf817b78f, 32'shf8162885, 32'shf814997c, 32'shf8130a74, 
               32'shf8117b6d, 32'shf80fec68, 32'shf80e5d64, 32'shf80cce61, 32'shf80b3f5f, 32'shf809b05e, 32'shf808215f, 32'shf8069261, 
               32'shf8050364, 32'shf8037468, 32'shf801e56e, 32'shf8005675, 32'shf7fec77d, 32'shf7fd3886, 32'shf7fba991, 32'shf7fa1a9c, 
               32'shf7f88ba9, 32'shf7f6fcb8, 32'shf7f56dc7, 32'shf7f3ded8, 32'shf7f24fea, 32'shf7f0c0fd, 32'shf7ef3211, 32'shf7eda327, 
               32'shf7ec143e, 32'shf7ea8556, 32'shf7e8f670, 32'shf7e7678a, 32'shf7e5d8a6, 32'shf7e449c3, 32'shf7e2bae2, 32'shf7e12c01, 
               32'shf7df9d22, 32'shf7de0e44, 32'shf7dc7f68, 32'shf7daf08d, 32'shf7d961b3, 32'shf7d7d2da, 32'shf7d64402, 32'shf7d4b52c, 
               32'shf7d32657, 32'shf7d19783, 32'shf7d008b1, 32'shf7ce79df, 32'shf7cceb0f, 32'shf7cb5c41, 32'shf7c9cd73, 32'shf7c83ea7, 
               32'shf7c6afdc, 32'shf7c52112, 32'shf7c3924a, 32'shf7c20383, 32'shf7c074bd, 32'shf7bee5f9, 32'shf7bd5735, 32'shf7bbc873, 
               32'shf7ba39b3, 32'shf7b8aaf3, 32'shf7b71c35, 32'shf7b58d78, 32'shf7b3febc, 32'shf7b27002, 32'shf7b0e149, 32'shf7af5291, 
               32'shf7adc3db, 32'shf7ac3525, 32'shf7aaa671, 32'shf7a917bf, 32'shf7a7890d, 32'shf7a5fa5d, 32'shf7a46baf, 32'shf7a2dd01, 
               32'shf7a14e55, 32'shf79fbfaa, 32'shf79e3100, 32'shf79ca258, 32'shf79b13b1, 32'shf799850b, 32'shf797f667, 32'shf79667c4, 
               32'shf794d922, 32'shf7934a81, 32'shf791bbe2, 32'shf7902d44, 32'shf78e9ea7, 32'shf78d100c, 32'shf78b8172, 32'shf789f2d9, 
               32'shf7886442, 32'shf786d5ab, 32'shf7854717, 32'shf783b883, 32'shf78229f1, 32'shf7809b60, 32'shf77f0cd0, 32'shf77d7e42, 
               32'shf77befb5, 32'shf77a6129, 32'shf778d29f, 32'shf7774416, 32'shf775b58e, 32'shf7742708, 32'shf7729883, 32'shf77109ff, 
               32'shf76f7b7d, 32'shf76decfb, 32'shf76c5e7c, 32'shf76acffd, 32'shf7694180, 32'shf767b304, 32'shf766248a, 32'shf7649610, 
               32'shf7630799, 32'shf7617922, 32'shf75feaad, 32'shf75e5c39, 32'shf75ccdc6, 32'shf75b3f55, 32'shf759b0e5, 32'shf7582277, 
               32'shf756940a, 32'shf755059e, 32'shf7537733, 32'shf751e8ca, 32'shf7505a62, 32'shf74ecbfc, 32'shf74d3d96, 32'shf74baf33, 
               32'shf74a20d0, 32'shf748926f, 32'shf747040f, 32'shf74575b1, 32'shf743e754, 32'shf74258f8, 32'shf740ca9d, 32'shf73f3c44, 
               32'shf73daded, 32'shf73c1f96, 32'shf73a9141, 32'shf73902ee, 32'shf737749b, 32'shf735e64a, 32'shf73457fb, 32'shf732c9ad, 
               32'shf7313b60, 32'shf72fad14, 32'shf72e1eca, 32'shf72c9081, 32'shf72b023a, 32'shf72973f4, 32'shf727e5af, 32'shf726576c, 
               32'shf724c92a, 32'shf7233ae9, 32'shf721acaa, 32'shf7201e6c, 32'shf71e902f, 32'shf71d01f4, 32'shf71b73ba, 32'shf719e582, 
               32'shf718574b, 32'shf716c915, 32'shf7153ae1, 32'shf713acae, 32'shf7121e7c, 32'shf710904c, 32'shf70f021d, 32'shf70d73f0, 
               32'shf70be5c4, 32'shf70a5799, 32'shf708c970, 32'shf7073b48, 32'shf705ad22, 32'shf7041efd, 32'shf70290d9, 32'shf70102b6, 
               32'shf6ff7496, 32'shf6fde676, 32'shf6fc5858, 32'shf6faca3b, 32'shf6f93c20, 32'shf6f7ae06, 32'shf6f61fed, 32'shf6f491d6, 
               32'shf6f303c0, 32'shf6f175ac, 32'shf6efe798, 32'shf6ee5987, 32'shf6eccb77, 32'shf6eb3d68, 32'shf6e9af5a, 32'shf6e8214e, 
               32'shf6e69344, 32'shf6e5053a, 32'shf6e37733, 32'shf6e1e92c, 32'shf6e05b27, 32'shf6decd24, 32'shf6dd3f21, 32'shf6dbb121, 
               32'shf6da2321, 32'shf6d89523, 32'shf6d70727, 32'shf6d5792c, 32'shf6d3eb32, 32'shf6d25d39, 32'shf6d0cf43, 32'shf6cf414d, 
               32'shf6cdb359, 32'shf6cc2566, 32'shf6ca9775, 32'shf6c90985, 32'shf6c77b97, 32'shf6c5edaa, 32'shf6c45fbe, 32'shf6c2d1d4, 
               32'shf6c143ec, 32'shf6bfb604, 32'shf6be281e, 32'shf6bc9a3a, 32'shf6bb0c57, 32'shf6b97e76, 32'shf6b7f095, 32'shf6b662b7, 
               32'shf6b4d4d9, 32'shf6b346fe, 32'shf6b1b923, 32'shf6b02b4a, 32'shf6ae9d73, 32'shf6ad0f9d, 32'shf6ab81c8, 32'shf6a9f3f5, 
               32'shf6a86623, 32'shf6a6d853, 32'shf6a54a84, 32'shf6a3bcb6, 32'shf6a22eea, 32'shf6a0a120, 32'shf69f1357, 32'shf69d858f, 
               32'shf69bf7c9, 32'shf69a6a04, 32'shf698dc41, 32'shf6974e7f, 32'shf695c0be, 32'shf69432ff, 32'shf692a542, 32'shf6911786, 
               32'shf68f89cb, 32'shf68dfc12, 32'shf68c6e5a, 32'shf68ae0a4, 32'shf68952ef, 32'shf687c53c, 32'shf686378a, 32'shf684a9da, 
               32'shf6831c2b, 32'shf6818e7d, 32'shf68000d1, 32'shf67e7327, 32'shf67ce57e, 32'shf67b57d6, 32'shf679ca30, 32'shf6783c8b, 
               32'shf676aee8, 32'shf6752146, 32'shf67393a6, 32'shf6720607, 32'shf670786a, 32'shf66eeace, 32'shf66d5d34, 32'shf66bcf9b, 
               32'shf66a4203, 32'shf668b46d, 32'shf66726d9, 32'shf6659946, 32'shf6640bb4, 32'shf6627e24, 32'shf660f096, 32'shf65f6309, 
               32'shf65dd57d, 32'shf65c47f3, 32'shf65aba6b, 32'shf6592ce4, 32'shf6579f5e, 32'shf65611da, 32'shf6548457, 32'shf652f6d6, 
               32'shf6516956, 32'shf64fdbd8, 32'shf64e4e5c, 32'shf64cc0e0, 32'shf64b3367, 32'shf649a5ef, 32'shf6481878, 32'shf6468b03, 
               32'shf644fd8f, 32'shf643701d, 32'shf641e2ac, 32'shf640553d, 32'shf63ec7cf, 32'shf63d3a63, 32'shf63bacf8, 32'shf63a1f8f, 
               32'shf6389228, 32'shf63704c1, 32'shf635775d, 32'shf633e9fa, 32'shf6325c98, 32'shf630cf38, 32'shf62f41d9, 32'shf62db47c, 
               32'shf62c2721, 32'shf62a99c7, 32'shf6290c6e, 32'shf6277f17, 32'shf625f1c2, 32'shf624646e, 32'shf622d71b, 32'shf62149ca, 
               32'shf61fbc7b, 32'shf61e2f2d, 32'shf61ca1e1, 32'shf61b1496, 32'shf619874c, 32'shf617fa05, 32'shf6166cbe, 32'shf614df7a, 
               32'shf6135237, 32'shf611c4f5, 32'shf61037b5, 32'shf60eaa76, 32'shf60d1d39, 32'shf60b8ffd, 32'shf60a02c3, 32'shf608758b, 
               32'shf606e854, 32'shf6055b1f, 32'shf603cdeb, 32'shf60240b9, 32'shf600b388, 32'shf5ff2659, 32'shf5fd992b, 32'shf5fc0bff, 
               32'shf5fa7ed4, 32'shf5f8f1ab, 32'shf5f76484, 32'shf5f5d75e, 32'shf5f44a39, 32'shf5f2bd16, 32'shf5f12ff5, 32'shf5efa2d5, 
               32'shf5ee15b7, 32'shf5ec889a, 32'shf5eafb7f, 32'shf5e96e66, 32'shf5e7e14e, 32'shf5e65437, 32'shf5e4c722, 32'shf5e33a0f, 
               32'shf5e1acfd, 32'shf5e01fed, 32'shf5de92de, 32'shf5dd05d1, 32'shf5db78c6, 32'shf5d9ebbc, 32'shf5d85eb3, 32'shf5d6d1ad, 
               32'shf5d544a7, 32'shf5d3b7a4, 32'shf5d22aa2, 32'shf5d09da1, 32'shf5cf10a2, 32'shf5cd83a5, 32'shf5cbf6a9, 32'shf5ca69af, 
               32'shf5c8dcb6, 32'shf5c74fbf, 32'shf5c5c2c9, 32'shf5c435d5, 32'shf5c2a8e3, 32'shf5c11bf2, 32'shf5bf8f03, 32'shf5be0215, 
               32'shf5bc7529, 32'shf5bae83f, 32'shf5b95b56, 32'shf5b7ce6f, 32'shf5b64189, 32'shf5b4b4a5, 32'shf5b327c2, 32'shf5b19ae1, 
               32'shf5b00e02, 32'shf5ae8124, 32'shf5acf448, 32'shf5ab676d, 32'shf5a9da94, 32'shf5a84dbd, 32'shf5a6c0e7, 32'shf5a53413, 
               32'shf5a3a740, 32'shf5a21a6f, 32'shf5a08da0, 32'shf59f00d2, 32'shf59d7406, 32'shf59be73b, 32'shf59a5a72, 32'shf598cdab, 
               32'shf59740e5, 32'shf595b421, 32'shf594275e, 32'shf5929a9d, 32'shf5910dde, 32'shf58f8120, 32'shf58df464, 32'shf58c67a9, 
               32'shf58adaf0, 32'shf5894e39, 32'shf587c183, 32'shf58634cf, 32'shf584a81d, 32'shf5831b6c, 32'shf5818ebd, 32'shf580020f, 
               32'shf57e7563, 32'shf57ce8b9, 32'shf57b5c10, 32'shf579cf69, 32'shf57842c3, 32'shf576b61f, 32'shf575297d, 32'shf5739cdc, 
               32'shf572103d, 32'shf57083a0, 32'shf56ef704, 32'shf56d6a6a, 32'shf56bddd1, 32'shf56a513b, 32'shf568c4a5, 32'shf5673812, 
               32'shf565ab80, 32'shf5641eef, 32'shf5629261, 32'shf56105d4, 32'shf55f7948, 32'shf55decbe, 32'shf55c6036, 32'shf55ad3b0, 
               32'shf559472b, 32'shf557baa8, 32'shf5562e26, 32'shf554a1a6, 32'shf5531528, 32'shf55188ab, 32'shf54ffc30, 32'shf54e6fb7, 
               32'shf54ce33f, 32'shf54b56c9, 32'shf549ca55, 32'shf5483de2, 32'shf546b171, 32'shf5452501, 32'shf5439893, 32'shf5420c27, 
               32'shf5407fbd, 32'shf53ef354, 32'shf53d66ed, 32'shf53bda87, 32'shf53a4e24, 32'shf538c1c1, 32'shf5373561, 32'shf535a902, 
               32'shf5341ca5, 32'shf5329049, 32'shf53103ef, 32'shf52f7797, 32'shf52deb41, 32'shf52c5eec, 32'shf52ad299, 32'shf5294647, 
               32'shf527b9f7, 32'shf5262da9, 32'shf524a15d, 32'shf5231512, 32'shf52188c9, 32'shf51ffc81, 32'shf51e703b, 32'shf51ce3f7, 
               32'shf51b57b5, 32'shf519cb74, 32'shf5183f35, 32'shf516b2f7, 32'shf51526bc, 32'shf5139a82, 32'shf5120e49, 32'shf5108213, 
               32'shf50ef5de, 32'shf50d69aa, 32'shf50bdd79, 32'shf50a5149, 32'shf508c51b, 32'shf50738ee, 32'shf505acc3, 32'shf504209a, 
               32'shf5029473, 32'shf501084d, 32'shf4ff7c29, 32'shf4fdf007, 32'shf4fc63e6, 32'shf4fad7c7, 32'shf4f94baa, 32'shf4f7bf8e, 
               32'shf4f63374, 32'shf4f4a75c, 32'shf4f31b46, 32'shf4f18f31, 32'shf4f0031e, 32'shf4ee770c, 32'shf4eceafd, 32'shf4eb5eef, 
               32'shf4e9d2e3, 32'shf4e846d8, 32'shf4e6bacf, 32'shf4e52ec8, 32'shf4e3a2c3, 32'shf4e216bf, 32'shf4e08abd, 32'shf4defebd, 
               32'shf4dd72be, 32'shf4dbe6c2, 32'shf4da5ac7, 32'shf4d8cecd, 32'shf4d742d6, 32'shf4d5b6e0, 32'shf4d42aeb, 32'shf4d29ef9, 
               32'shf4d11308, 32'shf4cf8719, 32'shf4cdfb2c, 32'shf4cc6f40, 32'shf4cae356, 32'shf4c9576e, 32'shf4c7cb88, 32'shf4c63fa3, 
               32'shf4c4b3c0, 32'shf4c327df, 32'shf4c19c00, 32'shf4c01022, 32'shf4be8446, 32'shf4bcf86c, 32'shf4bb6c93, 32'shf4b9e0bc, 
               32'shf4b854e7, 32'shf4b6c914, 32'shf4b53d42, 32'shf4b3b173, 32'shf4b225a4, 32'shf4b099d8, 32'shf4af0e0d, 32'shf4ad8245, 
               32'shf4abf67e, 32'shf4aa6ab8, 32'shf4a8def5, 32'shf4a75333, 32'shf4a5c773, 32'shf4a43bb4, 32'shf4a2aff8, 32'shf4a1243d, 
               32'shf49f9884, 32'shf49e0ccc, 32'shf49c8117, 32'shf49af563, 32'shf49969b1, 32'shf497de00, 32'shf4965252, 32'shf494c6a5, 
               32'shf4933afa, 32'shf491af51, 32'shf49023a9, 32'shf48e9803, 32'shf48d0c5f, 32'shf48b80bd, 32'shf489f51d, 32'shf488697e, 
               32'shf486dde1, 32'shf4855246, 32'shf483c6ad, 32'shf4823b15, 32'shf480af7f, 32'shf47f23eb, 32'shf47d9859, 32'shf47c0cc8, 
               32'shf47a8139, 32'shf478f5ad, 32'shf4776a21, 32'shf475de98, 32'shf4745310, 32'shf472c78a, 32'shf4713c06, 32'shf46fb084, 
               32'shf46e2504, 32'shf46c9985, 32'shf46b0e08, 32'shf469828d, 32'shf467f713, 32'shf4666b9c, 32'shf464e026, 32'shf46354b2, 
               32'shf461c940, 32'shf4603dcf, 32'shf45eb261, 32'shf45d26f4, 32'shf45b9b89, 32'shf45a1020, 32'shf45884b8, 32'shf456f953, 
               32'shf4556def, 32'shf453e28d, 32'shf452572c, 32'shf450cbce, 32'shf44f4071, 32'shf44db517, 32'shf44c29be, 32'shf44a9e66, 
               32'shf4491311, 32'shf44787bd, 32'shf445fc6b, 32'shf444711b, 32'shf442e5cd, 32'shf4415a81, 32'shf43fcf36, 32'shf43e43ed, 
               32'shf43cb8a7, 32'shf43b2d61, 32'shf439a21e, 32'shf43816dd, 32'shf4368b9d, 32'shf435005f, 32'shf4337523, 32'shf431e9e9, 
               32'shf4305eb0, 32'shf42ed37a, 32'shf42d4845, 32'shf42bbd12, 32'shf42a31e1, 32'shf428a6b2, 32'shf4271b84, 32'shf4259058, 
               32'shf424052f, 32'shf4227a07, 32'shf420eee1, 32'shf41f63bc, 32'shf41dd89a, 32'shf41c4d79, 32'shf41ac25a, 32'shf419373d, 
               32'shf417ac22, 32'shf4162109, 32'shf41495f1, 32'shf4130adc, 32'shf4117fc8, 32'shf40ff4b6, 32'shf40e69a6, 32'shf40cde97, 
               32'shf40b538b, 32'shf409c880, 32'shf4083d78, 32'shf406b271, 32'shf405276c, 32'shf4039c68, 32'shf4021167, 32'shf4008668, 
               32'shf3fefb6a, 32'shf3fd706e, 32'shf3fbe574, 32'shf3fa5a7c, 32'shf3f8cf86, 32'shf3f74491, 32'shf3f5b99f, 32'shf3f42eae, 
               32'shf3f2a3bf, 32'shf3f118d2, 32'shf3ef8de7, 32'shf3ee02fe, 32'shf3ec7817, 32'shf3eaed31, 32'shf3e9624d, 32'shf3e7d76c, 
               32'shf3e64c8c, 32'shf3e4c1ae, 32'shf3e336d1, 32'shf3e1abf7, 32'shf3e0211f, 32'shf3de9648, 32'shf3dd0b73, 32'shf3db80a0, 
               32'shf3d9f5cf, 32'shf3d86b00, 32'shf3d6e033, 32'shf3d55568, 32'shf3d3ca9e, 32'shf3d23fd7, 32'shf3d0b511, 32'shf3cf2a4d, 
               32'shf3cd9f8b, 32'shf3cc14cb, 32'shf3ca8a0d, 32'shf3c8ff51, 32'shf3c77496, 32'shf3c5e9de, 32'shf3c45f27, 32'shf3c2d472, 
               32'shf3c149bf, 32'shf3bfbf0e, 32'shf3be345f, 32'shf3bca9b2, 32'shf3bb1f07, 32'shf3b9945d, 32'shf3b809b6, 32'shf3b67f10, 
               32'shf3b4f46c, 32'shf3b369ca, 32'shf3b1df2a, 32'shf3b0548c, 32'shf3aec9f0, 32'shf3ad3f56, 32'shf3abb4bd, 32'shf3aa2a27, 
               32'shf3a89f92, 32'shf3a71500, 32'shf3a58a6f, 32'shf3a3ffe0, 32'shf3a27553, 32'shf3a0eac8, 32'shf39f603f, 32'shf39dd5b8, 
               32'shf39c4b32, 32'shf39ac0af, 32'shf399362d, 32'shf397abae, 32'shf3962130, 32'shf39496b4, 32'shf3930c3b, 32'shf39181c3, 
               32'shf38ff74d, 32'shf38e6cd9, 32'shf38ce266, 32'shf38b57f6, 32'shf389cd88, 32'shf388431b, 32'shf386b8b1, 32'shf3852e48, 
               32'shf383a3e2, 32'shf382197d, 32'shf3808f1a, 32'shf37f04b9, 32'shf37d7a5b, 32'shf37beffe, 32'shf37a65a2, 32'shf378db49, 
               32'shf37750f2, 32'shf375c69d, 32'shf3743c49, 32'shf372b1f8, 32'shf37127a9, 32'shf36f9d5b, 32'shf36e130f, 32'shf36c88c6, 
               32'shf36afe7e, 32'shf3697438, 32'shf367e9f4, 32'shf3665fb3, 32'shf364d573, 32'shf3634b35, 32'shf361c0f9, 32'shf36036be, 
               32'shf35eac86, 32'shf35d2250, 32'shf35b981c, 32'shf35a0de9, 32'shf35883b9, 32'shf356f98b, 32'shf3556f5e, 32'shf353e534, 
               32'shf3525b0b, 32'shf350d0e5, 32'shf34f46c0, 32'shf34dbc9d, 32'shf34c327c, 32'shf34aa85e, 32'shf3491e41, 32'shf3479426, 
               32'shf3460a0d, 32'shf3447ff6, 32'shf342f5e1, 32'shf3416bce, 32'shf33fe1bd, 32'shf33e57ae, 32'shf33ccda1, 32'shf33b4396, 
               32'shf339b98d, 32'shf3382f86, 32'shf336a580, 32'shf3351b7d, 32'shf333917c, 32'shf332077c, 32'shf3307d7f, 32'shf32ef384, 
               32'shf32d698a, 32'shf32bdf93, 32'shf32a559e, 32'shf328cbaa, 32'shf32741b9, 32'shf325b7c9, 32'shf3242ddc, 32'shf322a3f0, 
               32'shf3211a07, 32'shf31f901f, 32'shf31e0639, 32'shf31c7c56, 32'shf31af274, 32'shf3196895, 32'shf317deb7, 32'shf31654db, 
               32'shf314cb02, 32'shf313412a, 32'shf311b755, 32'shf3102d81, 32'shf30ea3af, 32'shf30d19e0, 32'shf30b9012, 32'shf30a0646, 
               32'shf3087c7d, 32'shf306f2b5, 32'shf30568ef, 32'shf303df2c, 32'shf302556a, 32'shf300cbaa, 32'shf2ff41ed, 32'shf2fdb831, 
               32'shf2fc2e77, 32'shf2faa4c0, 32'shf2f91b0a, 32'shf2f79156, 32'shf2f607a5, 32'shf2f47df5, 32'shf2f2f448, 32'shf2f16a9c, 
               32'shf2efe0f2, 32'shf2ee574b, 32'shf2eccda5, 32'shf2eb4402, 32'shf2e9ba60, 32'shf2e830c1, 32'shf2e6a723, 32'shf2e51d88, 
               32'shf2e393ef, 32'shf2e20a57, 32'shf2e080c2, 32'shf2def72e, 32'shf2dd6d9d, 32'shf2dbe40e, 32'shf2da5a81, 32'shf2d8d0f5, 
               32'shf2d7476c, 32'shf2d5bde5, 32'shf2d43460, 32'shf2d2aadd, 32'shf2d1215b, 32'shf2cf97dc, 32'shf2ce0e5f, 32'shf2cc84e4, 
               32'shf2cafb6b, 32'shf2c971f5, 32'shf2c7e880, 32'shf2c65f0d, 32'shf2c4d59c, 32'shf2c34c2d, 32'shf2c1c2c0, 32'shf2c03956, 
               32'shf2beafed, 32'shf2bd2687, 32'shf2bb9d22, 32'shf2ba13c0, 32'shf2b88a5f, 32'shf2b70101, 32'shf2b577a4, 32'shf2b3ee4a, 
               32'shf2b264f2, 32'shf2b0db9b, 32'shf2af5247, 32'shf2adc8f5, 32'shf2ac3fa5, 32'shf2aab657, 32'shf2a92d0b, 32'shf2a7a3c1, 
               32'shf2a61a7a, 32'shf2a49134, 32'shf2a307f0, 32'shf2a17eae, 32'shf29ff56f, 32'shf29e6c31, 32'shf29ce2f6, 32'shf29b59bc, 
               32'shf299d085, 32'shf2984750, 32'shf296be1d, 32'shf29534ec, 32'shf293abbd, 32'shf2922290, 32'shf2909965, 32'shf28f103c, 
               32'shf28d8715, 32'shf28bfdf0, 32'shf28a74ce, 32'shf288ebad, 32'shf287628f, 32'shf285d972, 32'shf2845058, 32'shf282c740, 
               32'shf2813e2a, 32'shf27fb516, 32'shf27e2c04, 32'shf27ca2f4, 32'shf27b19e6, 32'shf27990da, 32'shf27807d0, 32'shf2767ec9, 
               32'shf274f5c3, 32'shf2736cc0, 32'shf271e3bf, 32'shf2705abf, 32'shf26ed1c2, 32'shf26d48c7, 32'shf26bbfce, 32'shf26a36d8, 
               32'shf268ade3, 32'shf26724f0, 32'shf2659c00, 32'shf2641311, 32'shf2628a25, 32'shf261013b, 32'shf25f7852, 32'shf25def6c, 
               32'shf25c6688, 32'shf25adda7, 32'shf25954c7, 32'shf257cbe9, 32'shf256430e, 32'shf254ba34, 32'shf253315d, 32'shf251a888, 
               32'shf2501fb5, 32'shf24e96e4, 32'shf24d0e15, 32'shf24b8548, 32'shf249fc7d, 32'shf24873b5, 32'shf246eaee, 32'shf245622a, 
               32'shf243d968, 32'shf24250a8, 32'shf240c7ea, 32'shf23f3f2e, 32'shf23db674, 32'shf23c2dbd, 32'shf23aa507, 32'shf2391c54, 
               32'shf23793a3, 32'shf2360af4, 32'shf2348247, 32'shf232f99c, 32'shf23170f3, 32'shf22fe84c, 32'shf22e5fa8, 32'shf22cd706, 
               32'shf22b4e66, 32'shf229c5c7, 32'shf2283d2c, 32'shf226b492, 32'shf2252bfa, 32'shf223a365, 32'shf2221ad1, 32'shf2209240, 
               32'shf21f09b1, 32'shf21d8124, 32'shf21bf899, 32'shf21a7010, 32'shf218e78a, 32'shf2175f06, 32'shf215d683, 32'shf2144e03, 
               32'shf212c585, 32'shf2113d09, 32'shf20fb490, 32'shf20e2c18, 32'shf20ca3a3, 32'shf20b1b30, 32'shf20992bf, 32'shf2080a50, 
               32'shf20681e3, 32'shf204f978, 32'shf2037110, 32'shf201e8aa, 32'shf2006046, 32'shf1fed7e4, 32'shf1fd4f84, 32'shf1fbc726, 
               32'shf1fa3ecb, 32'shf1f8b671, 32'shf1f72e1a, 32'shf1f5a5c5, 32'shf1f41d72, 32'shf1f29522, 32'shf1f10cd3, 32'shf1ef8487, 
               32'shf1edfc3d, 32'shf1ec73f5, 32'shf1eaebaf, 32'shf1e9636b, 32'shf1e7db2a, 32'shf1e652eb, 32'shf1e4caae, 32'shf1e34273, 
               32'shf1e1ba3a, 32'shf1e03203, 32'shf1dea9cf, 32'shf1dd219d, 32'shf1db996d, 32'shf1da113f, 32'shf1d88913, 32'shf1d700ea, 
               32'shf1d578c2, 32'shf1d3f09d, 32'shf1d2687a, 32'shf1d0e059, 32'shf1cf583b, 32'shf1cdd01e, 32'shf1cc4804, 32'shf1cabfec, 
               32'shf1c937d6, 32'shf1c7afc3, 32'shf1c627b1, 32'shf1c49fa2, 32'shf1c31795, 32'shf1c18f8a, 32'shf1c00781, 32'shf1be7f7b, 
               32'shf1bcf777, 32'shf1bb6f75, 32'shf1b9e775, 32'shf1b85f77, 32'shf1b6d77c, 32'shf1b54f82, 32'shf1b3c78b, 32'shf1b23f97, 
               32'shf1b0b7a4, 32'shf1af2fb3, 32'shf1ada7c5, 32'shf1ac1fd9, 32'shf1aa97ef, 32'shf1a91008, 32'shf1a78822, 32'shf1a6003f, 
               32'shf1a4785e, 32'shf1a2f080, 32'shf1a168a3, 32'shf19fe0c9, 32'shf19e58f1, 32'shf19cd11b, 32'shf19b4947, 32'shf199c176, 
               32'shf19839a6, 32'shf196b1d9, 32'shf1952a0f, 32'shf193a246, 32'shf1921a80, 32'shf19092bc, 32'shf18f0afa, 32'shf18d833a, 
               32'shf18bfb7d, 32'shf18a73c2, 32'shf188ec09, 32'shf1876452, 32'shf185dc9d, 32'shf18454eb, 32'shf182cd3b, 32'shf181458d, 
               32'shf17fbde2, 32'shf17e3638, 32'shf17cae91, 32'shf17b26ec, 32'shf1799f4a, 32'shf17817a9, 32'shf176900b, 32'shf175086f, 
               32'shf17380d6, 32'shf171f93e, 32'shf17071a9, 32'shf16eea16, 32'shf16d6286, 32'shf16bdaf7, 32'shf16a536b, 32'shf168cbe1, 
               32'shf1674459, 32'shf165bcd4, 32'shf1643551, 32'shf162add0, 32'shf1612651, 32'shf15f9ed5, 32'shf15e175b, 32'shf15c8fe3, 
               32'shf15b086d, 32'shf15980fa, 32'shf157f989, 32'shf156721a, 32'shf154eaad, 32'shf1536343, 32'shf151dbdb, 32'shf1505475, 
               32'shf14ecd11, 32'shf14d45b0, 32'shf14bbe51, 32'shf14a36f4, 32'shf148af9a, 32'shf1472842, 32'shf145a0ec, 32'shf1441998, 
               32'shf1429247, 32'shf1410af8, 32'shf13f83ab, 32'shf13dfc60, 32'shf13c7518, 32'shf13aedd2, 32'shf139668e, 32'shf137df4d, 
               32'shf136580d, 32'shf134d0d0, 32'shf1334996, 32'shf131c25d, 32'shf1303b27, 32'shf12eb3f4, 32'shf12d2cc2, 32'shf12ba593, 
               32'shf12a1e66, 32'shf128973b, 32'shf1271013, 32'shf12588ed, 32'shf12401c9, 32'shf1227aa8, 32'shf120f389, 32'shf11f6c6c, 
               32'shf11de551, 32'shf11c5e39, 32'shf11ad723, 32'shf119500f, 32'shf117c8fe, 32'shf11641ef, 32'shf114bae2, 32'shf11333d7, 
               32'shf111accf, 32'shf11025c9, 32'shf10e9ec6, 32'shf10d17c4, 32'shf10b90c5, 32'shf10a09c9, 32'shf10882ce, 32'shf106fbd6, 
               32'shf10574e0, 32'shf103eded, 32'shf10266fc, 32'shf100e00d, 32'shf0ff5921, 32'shf0fdd236, 32'shf0fc4b4f, 32'shf0fac469, 
               32'shf0f93d86, 32'shf0f7b6a5, 32'shf0f62fc6, 32'shf0f4a8ea, 32'shf0f32210, 32'shf0f19b38, 32'shf0f01463, 32'shf0ee8d90, 
               32'shf0ed06bf, 32'shf0eb7ff1, 32'shf0e9f925, 32'shf0e8725b, 32'shf0e6eb94, 32'shf0e564cf, 32'shf0e3de0c, 32'shf0e2574c, 
               32'shf0e0d08d, 32'shf0df49d2, 32'shf0ddc318, 32'shf0dc3c61, 32'shf0dab5ad, 32'shf0d92efa, 32'shf0d7a84a, 32'shf0d6219c, 
               32'shf0d49af1, 32'shf0d31448, 32'shf0d18da1, 32'shf0d006fd, 32'shf0ce805b, 32'shf0ccf9bb, 32'shf0cb731e, 32'shf0c9ec83, 
               32'shf0c865ea, 32'shf0c6df54, 32'shf0c558c0, 32'shf0c3d22e, 32'shf0c24b9f, 32'shf0c0c512, 32'shf0bf3e88, 32'shf0bdb7ff, 
               32'shf0bc317a, 32'shf0baaaf6, 32'shf0b92475, 32'shf0b79df6, 32'shf0b6177a, 32'shf0b49100, 32'shf0b30a88, 32'shf0b18413, 
               32'shf0affda0, 32'shf0ae772f, 32'shf0acf0c1, 32'shf0ab6a55, 32'shf0a9e3eb, 32'shf0a85d84, 32'shf0a6d71f, 32'shf0a550bd, 
               32'shf0a3ca5d, 32'shf0a243ff, 32'shf0a0bda4, 32'shf09f374b, 32'shf09db0f4, 32'shf09c2aa0, 32'shf09aa44e, 32'shf0991dff, 
               32'shf09797b2, 32'shf0961167, 32'shf0948b1f, 32'shf09304d9, 32'shf0917e95, 32'shf08ff854, 32'shf08e7215, 32'shf08cebd9, 
               32'shf08b659f, 32'shf089df67, 32'shf0885932, 32'shf086d2ff, 32'shf0854cce, 32'shf083c6a0, 32'shf0824074, 32'shf080ba4b, 
               32'shf07f3424, 32'shf07dadff, 32'shf07c27dd, 32'shf07aa1bd, 32'shf0791ba0, 32'shf0779585, 32'shf0760f6c, 32'shf0748956, 
               32'shf0730342, 32'shf0717d31, 32'shf06ff722, 32'shf06e7115, 32'shf06ceb0b, 32'shf06b6503, 32'shf069defe, 32'shf06858fb, 
               32'shf066d2fa, 32'shf0654cfc, 32'shf063c700, 32'shf0624107, 32'shf060bb10, 32'shf05f351b, 32'shf05daf29, 32'shf05c293a, 
               32'shf05aa34c, 32'shf0591d61, 32'shf0579779, 32'shf0561193, 32'shf0548baf, 32'shf05305ce, 32'shf0517fef, 32'shf04ffa12, 
               32'shf04e7438, 32'shf04cee61, 32'shf04b688c, 32'shf049e2b9, 32'shf0485ce9, 32'shf046d71b, 32'shf045514f, 32'shf043cb86, 
               32'shf04245c0, 32'shf040bffb, 32'shf03f3a3a, 32'shf03db47a, 32'shf03c2ebd, 32'shf03aa903, 32'shf039234b, 32'shf0379d95, 
               32'shf03617e2, 32'shf0349231, 32'shf0330c83, 32'shf03186d7, 32'shf030012e, 32'shf02e7b87, 32'shf02cf5e2, 32'shf02b7040, 
               32'shf029eaa1, 32'shf0286503, 32'shf026df68, 32'shf02559d0, 32'shf023d43a, 32'shf0224ea7, 32'shf020c916, 32'shf01f4387, 
               32'shf01dbdfb, 32'shf01c3871, 32'shf01ab2ea, 32'shf0192d66, 32'shf017a7e3, 32'shf0162263, 32'shf0149ce6, 32'shf013176b, 
               32'shf01191f3, 32'shf0100c7d, 32'shf00e8709, 32'shf00d0198, 32'shf00b7c29, 32'shf009f6bd, 32'shf0087153, 32'shf006ebec, 
               32'shf0056687, 32'shf003e125, 32'shf0025bc5, 32'shf000d668, 32'shefff510d, 32'sheffdcbb4, 32'sheffc465e, 32'sheffac10b, 
               32'sheff93bba, 32'sheff7b66b, 32'sheff6311f, 32'sheff4abd5, 32'sheff3268e, 32'sheff1a149, 32'sheff01c07, 32'shefee96c7, 
               32'shefed118a, 32'shefeb8c4f, 32'shefea0717, 32'shefe881e1, 32'shefe6fcae, 32'shefe5777d, 32'shefe3f24f, 32'shefe26d23, 
               32'shefe0e7f9, 32'shefdf62d2, 32'shefddddae, 32'shefdc588c, 32'shefdad36c, 32'shefd94e50, 32'shefd7c935, 32'shefd6441d, 
               32'shefd4bf08, 32'shefd339f5, 32'shefd1b4e4, 32'shefd02fd6, 32'shefceaacb, 32'shefcd25c1, 32'shefcba0bb, 32'shefca1bb7, 
               32'shefc896b5, 32'shefc711b6, 32'shefc58cba, 32'shefc407c0, 32'shefc282c8, 32'shefc0fdd3, 32'shefbf78e1, 32'shefbdf3f1, 
               32'shefbc6f03, 32'shefbaea18, 32'shefb96530, 32'shefb7e04a, 32'shefb65b66, 32'shefb4d686, 32'shefb351a7, 32'shefb1cccb, 
               32'shefb047f2, 32'shefaec31b, 32'shefad3e47, 32'shefabb975, 32'shefaa34a5, 32'shefa8afd9, 32'shefa72b0e, 32'shefa5a646, 
               32'shefa42181, 32'shefa29cbe, 32'shefa117fe, 32'shef9f9341, 32'shef9e0e85, 32'shef9c89cd, 32'shef9b0517, 32'shef998063, 
               32'shef97fbb2, 32'shef967704, 32'shef94f258, 32'shef936dae, 32'shef91e907, 32'shef906463, 32'shef8edfc1, 32'shef8d5b22, 
               32'shef8bd685, 32'shef8a51eb, 32'shef88cd53, 32'shef8748be, 32'shef85c42b, 32'shef843f9b, 32'shef82bb0e, 32'shef813683, 
               32'shef7fb1fa, 32'shef7e2d74, 32'shef7ca8f1, 32'shef7b2470, 32'shef799ff2, 32'shef781b76, 32'shef7696fd, 32'shef751286, 
               32'shef738e12, 32'shef7209a1, 32'shef708532, 32'shef6f00c5, 32'shef6d7c5b, 32'shef6bf7f4, 32'shef6a738f, 32'shef68ef2d, 
               32'shef676ace, 32'shef65e670, 32'shef646216, 32'shef62ddbe, 32'shef615969, 32'shef5fd516, 32'shef5e50c6, 32'shef5ccc78, 
               32'shef5b482d, 32'shef59c3e4, 32'shef583f9e, 32'shef56bb5b, 32'shef55371a, 32'shef53b2dc, 32'shef522ea0, 32'shef50aa67, 
               32'shef4f2630, 32'shef4da1fc, 32'shef4c1dcb, 32'shef4a999c, 32'shef491570, 32'shef479146, 32'shef460d1f, 32'shef4488fa, 
               32'shef4304d8, 32'shef4180b9, 32'shef3ffc9c, 32'shef3e7882, 32'shef3cf46a, 32'shef3b7055, 32'shef39ec43, 32'shef386833, 
               32'shef36e426, 32'shef35601b, 32'shef33dc13, 32'shef32580d, 32'shef30d40a, 32'shef2f500a, 32'shef2dcc0c, 32'shef2c4811, 
               32'shef2ac419, 32'shef294023, 32'shef27bc2f, 32'shef26383f, 32'shef24b451, 32'shef233065, 32'shef21ac7c, 32'shef202896, 
               32'shef1ea4b2, 32'shef1d20d1, 32'shef1b9cf2, 32'shef1a1916, 32'shef18953d, 32'shef171166, 32'shef158d92, 32'shef1409c1, 
               32'shef1285f2, 32'shef110225, 32'shef0f7e5c, 32'shef0dfa95, 32'shef0c76d0, 32'shef0af30e, 32'shef096f4f, 32'shef07eb93, 
               32'shef0667d9, 32'shef04e421, 32'shef03606c, 32'shef01dcba, 32'shef00590b, 32'sheefed55e, 32'sheefd51b4, 32'sheefbce0c, 
               32'sheefa4a67, 32'sheef8c6c5, 32'sheef74325, 32'sheef5bf88, 32'sheef43bed, 32'sheef2b855, 32'sheef134c0, 32'sheeefb12d, 
               32'sheeee2d9d, 32'sheeecaa10, 32'sheeeb2685, 32'sheee9a2fd, 32'sheee81f78, 32'sheee69bf5, 32'sheee51875, 32'sheee394f7, 
               32'sheee2117c, 32'sheee08e04, 32'sheedf0a8e, 32'sheedd871b, 32'sheedc03ab, 32'sheeda803d, 32'sheed8fcd2, 32'sheed7796a, 
               32'sheed5f604, 32'sheed472a1, 32'sheed2ef40, 32'sheed16be3, 32'sheecfe887, 32'sheece652f, 32'sheecce1d9, 32'sheecb5e86, 
               32'sheec9db35, 32'sheec857e7, 32'sheec6d49c, 32'sheec55153, 32'sheec3ce0d, 32'sheec24aca, 32'sheec0c78a, 32'sheebf444c, 
               32'sheebdc110, 32'sheebc3dd8, 32'sheebabaa2, 32'sheeb9376e, 32'sheeb7b43e, 32'sheeb63110, 32'sheeb4ade4, 32'sheeb32abc, 
               32'sheeb1a796, 32'sheeb02472, 32'sheeaea152, 32'sheead1e34, 32'sheeab9b18, 32'sheeaa1800, 32'sheea894ea, 32'sheea711d6, 
               32'sheea58ec6, 32'sheea40bb8, 32'sheea288ad, 32'sheea105a4, 32'shee9f829e, 32'shee9dff9b, 32'shee9c7c9a, 32'shee9af99d, 
               32'shee9976a1, 32'shee97f3a9, 32'shee9670b3, 32'shee94edc0, 32'shee936acf, 32'shee91e7e2, 32'shee9064f7, 32'shee8ee20e, 
               32'shee8d5f29, 32'shee8bdc46, 32'shee8a5965, 32'shee88d688, 32'shee8753ad, 32'shee85d0d4, 32'shee844dff, 32'shee82cb2c, 
               32'shee81485c, 32'shee7fc58f, 32'shee7e42c4, 32'shee7cbffc, 32'shee7b3d36, 32'shee79ba74, 32'shee7837b4, 32'shee76b4f7, 
               32'shee75323c, 32'shee73af84, 32'shee722ccf, 32'shee70aa1d, 32'shee6f276d, 32'shee6da4c0, 32'shee6c2216, 32'shee6a9f6e, 
               32'shee691cc9, 32'shee679a27, 32'shee661788, 32'shee6494eb, 32'shee631251, 32'shee618fba, 32'shee600d25, 32'shee5e8a93, 
               32'shee5d0804, 32'shee5b8578, 32'shee5a02ee, 32'shee588067, 32'shee56fde3, 32'shee557b61, 32'shee53f8e2, 32'shee527666, 
               32'shee50f3ed, 32'shee4f7176, 32'shee4def02, 32'shee4c6c91, 32'shee4aea23, 32'shee4967b7, 32'shee47e54e, 32'shee4662e8, 
               32'shee44e084, 32'shee435e24, 32'shee41dbc6, 32'shee40596a, 32'shee3ed712, 32'shee3d54bc, 32'shee3bd269, 32'shee3a5018, 
               32'shee38cdcb, 32'shee374b80, 32'shee35c938, 32'shee3446f2, 32'shee32c4b0, 32'shee314270, 32'shee2fc033, 32'shee2e3df8, 
               32'shee2cbbc1, 32'shee2b398c, 32'shee29b75a, 32'shee28352a, 32'shee26b2fe, 32'shee2530d4, 32'shee23aead, 32'shee222c88, 
               32'shee20aa67, 32'shee1f2848, 32'shee1da62c, 32'shee1c2412, 32'shee1aa1fc, 32'shee191fe8, 32'shee179dd7, 32'shee161bc8, 
               32'shee1499bd, 32'shee1317b4, 32'shee1195ae, 32'shee1013ab, 32'shee0e91aa, 32'shee0d0fac, 32'shee0b8db1, 32'shee0a0bb9, 
               32'shee0889c4, 32'shee0707d1, 32'shee0585e1, 32'shee0403f4, 32'shee02820a, 32'shee010022, 32'shedff7e3d, 32'shedfdfc5b, 
               32'shedfc7a7c, 32'shedfaf8a0, 32'shedf976c6, 32'shedf7f4ef, 32'shedf6731b, 32'shedf4f14a, 32'shedf36f7b, 32'shedf1edaf, 
               32'shedf06be6, 32'shedeeea20, 32'sheded685d, 32'shedebe69c, 32'shedea64de, 32'shede8e323, 32'shede7616b, 32'shede5dfb5, 
               32'shede45e03, 32'shede2dc53, 32'shede15aa6, 32'sheddfd8fb, 32'shedde5754, 32'sheddcd5af, 32'sheddb540d, 32'shedd9d26e, 
               32'shedd850d2, 32'shedd6cf38, 32'shedd54da2, 32'shedd3cc0e, 32'shedd24a7d, 32'shedd0c8ee, 32'shedcf4763, 32'shedcdc5da, 
               32'shedcc4454, 32'shedcac2d1, 32'shedc94151, 32'shedc7bfd3, 32'shedc63e59, 32'shedc4bce1, 32'shedc33b6c, 32'shedc1b9fa, 
               32'shedc0388a, 32'shedbeb71e, 32'shedbd35b4, 32'shedbbb44d, 32'shedba32e9, 32'shedb8b187, 32'shedb73029, 32'shedb5aecd, 
               32'shedb42d74, 32'shedb2ac1e, 32'shedb12acb, 32'shedafa97b, 32'shedae282d, 32'shedaca6e2, 32'shedab259a, 32'sheda9a455, 
               32'sheda82313, 32'sheda6a1d4, 32'sheda52097, 32'sheda39f5d, 32'sheda21e26, 32'sheda09cf2, 32'shed9f1bc1, 32'shed9d9a92, 
               32'shed9c1967, 32'shed9a983e, 32'shed991718, 32'shed9795f5, 32'shed9614d5, 32'shed9493b7, 32'shed93129d, 32'shed919185, 
               32'shed901070, 32'shed8e8f5e, 32'shed8d0e4f, 32'shed8b8d42, 32'shed8a0c39, 32'shed888b32, 32'shed870a2e, 32'shed85892d, 
               32'shed84082f, 32'shed828734, 32'shed81063b, 32'shed7f8546, 32'shed7e0453, 32'shed7c8363, 32'shed7b0276, 32'shed79818c, 
               32'shed7800a5, 32'shed767fc0, 32'shed74fedf, 32'shed737e00, 32'shed71fd24, 32'shed707c4b, 32'shed6efb75, 32'shed6d7aa2, 
               32'shed6bf9d1, 32'shed6a7904, 32'shed68f839, 32'shed677771, 32'shed65f6ac, 32'shed6475ea, 32'shed62f52b, 32'shed61746f, 
               32'shed5ff3b5, 32'shed5e72fe, 32'shed5cf24b, 32'shed5b719a, 32'shed59f0ec, 32'shed587041, 32'shed56ef99, 32'shed556ef3, 
               32'shed53ee51, 32'shed526db1, 32'shed50ed14, 32'shed4f6c7b, 32'shed4debe4, 32'shed4c6b50, 32'shed4aeabe, 32'shed496a30, 
               32'shed47e9a5, 32'shed46691c, 32'shed44e897, 32'shed436814, 32'shed41e794, 32'shed406717, 32'shed3ee69d, 32'shed3d6626, 
               32'shed3be5b1, 32'shed3a6540, 32'shed38e4d2, 32'shed376466, 32'shed35e3fd, 32'shed346397, 32'shed32e334, 32'shed3162d4, 
               32'shed2fe277, 32'shed2e621d, 32'shed2ce1c6, 32'shed2b6171, 32'shed29e120, 32'shed2860d1, 32'shed26e086, 32'shed25603d, 
               32'shed23dff7, 32'shed225fb4, 32'shed20df74, 32'shed1f5f37, 32'shed1ddefd, 32'shed1c5ec5, 32'shed1ade91, 32'shed195e5f, 
               32'shed17de31, 32'shed165e05, 32'shed14dddc, 32'shed135db6, 32'shed11dd94, 32'shed105d74, 32'shed0edd56, 32'shed0d5d3c, 
               32'shed0bdd25, 32'shed0a5d11, 32'shed08dcff, 32'shed075cf1, 32'shed05dce5, 32'shed045cdd, 32'shed02dcd7, 32'shed015cd4, 
               32'shecffdcd4, 32'shecfe5cd8, 32'shecfcdcde, 32'shecfb5ce7, 32'shecf9dcf3, 32'shecf85d01, 32'shecf6dd13, 32'shecf55d28, 
               32'shecf3dd3f, 32'shecf25d5a, 32'shecf0dd78, 32'shecef5d98, 32'shecedddbb, 32'shecec5de2, 32'sheceade0b, 32'shece95e37, 
               32'shece7de66, 32'shece65e98, 32'shece4dece, 32'shece35f06, 32'shece1df40, 32'shece05f7e, 32'shecdedfbf, 32'shecdd6003, 
               32'shecdbe04a, 32'shecda6093, 32'shecd8e0e0, 32'shecd76130, 32'shecd5e182, 32'shecd461d8, 32'shecd2e230, 32'shecd1628c, 
               32'sheccfe2ea, 32'shecce634b, 32'sheccce3b0, 32'sheccb6417, 32'shecc9e481, 32'shecc864ee, 32'shecc6e55f, 32'shecc565d2, 
               32'shecc3e648, 32'shecc266c1, 32'shecc0e73d, 32'shecbf67bc, 32'shecbde83e, 32'shecbc68c3, 32'shecbae94b, 32'shecb969d5, 
               32'shecb7ea63, 32'shecb66af4, 32'shecb4eb88, 32'shecb36c1f, 32'shecb1ecb8, 32'shecb06d55, 32'shecaeedf5, 32'shecad6e97, 
               32'shecabef3d, 32'shecaa6fe6, 32'sheca8f091, 32'sheca77140, 32'sheca5f1f2, 32'sheca472a6, 32'sheca2f35e, 32'sheca17418, 
               32'shec9ff4d6, 32'shec9e7596, 32'shec9cf65a, 32'shec9b7720, 32'shec99f7ea, 32'shec9878b6, 32'shec96f986, 32'shec957a58, 
               32'shec93fb2e, 32'shec927c06, 32'shec90fce1, 32'shec8f7dc0, 32'shec8dfea1, 32'shec8c7f86, 32'shec8b006d, 32'shec898158, 
               32'shec880245, 32'shec868335, 32'shec850429, 32'shec83851f, 32'shec820619, 32'shec808715, 32'shec7f0815, 32'shec7d8917, 
               32'shec7c0a1d, 32'shec7a8b25, 32'shec790c31, 32'shec778d3f, 32'shec760e51, 32'shec748f65, 32'shec73107d, 32'shec719197, 
               32'shec7012b5, 32'shec6e93d6, 32'shec6d14f9, 32'shec6b9620, 32'shec6a1749, 32'shec689876, 32'shec6719a6, 32'shec659ad9, 
               32'shec641c0e, 32'shec629d47, 32'shec611e83, 32'shec5f9fc2, 32'shec5e2103, 32'shec5ca248, 32'shec5b2390, 32'shec59a4db, 
               32'shec582629, 32'shec56a77a, 32'shec5528ce, 32'shec53aa25, 32'shec522b7f, 32'shec50acdc, 32'shec4f2e3d, 32'shec4dafa0, 
               32'shec4c3106, 32'shec4ab26f, 32'shec4933dc, 32'shec47b54b, 32'shec4636bd, 32'shec44b833, 32'shec4339ab, 32'shec41bb27, 
               32'shec403ca5, 32'shec3ebe27, 32'shec3d3fac, 32'shec3bc133, 32'shec3a42be, 32'shec38c44c, 32'shec3745dd, 32'shec35c771, 
               32'shec344908, 32'shec32caa2, 32'shec314c3f, 32'shec2fcddf, 32'shec2e4f82, 32'shec2cd128, 32'shec2b52d1, 32'shec29d47e, 
               32'shec28562d, 32'shec26d7e0, 32'shec255995, 32'shec23db4e, 32'shec225d09, 32'shec20dec8, 32'shec1f608a, 32'shec1de24f, 
               32'shec1c6417, 32'shec1ae5e2, 32'shec1967b0, 32'shec17e981, 32'shec166b55, 32'shec14ed2c, 32'shec136f06, 32'shec11f0e4, 
               32'shec1072c4, 32'shec0ef4a8, 32'shec0d768e, 32'shec0bf878, 32'shec0a7a65, 32'shec08fc55, 32'shec077e48, 32'shec06003e, 
               32'shec048237, 32'shec030433, 32'shec018632, 32'shec000835, 32'shebfe8a3a, 32'shebfd0c42, 32'shebfb8e4e, 32'shebfa105d, 
               32'shebf8926f, 32'shebf71483, 32'shebf5969b, 32'shebf418b6, 32'shebf29ad4, 32'shebf11cf6, 32'shebef9f1a, 32'shebee2141, 
               32'shebeca36c, 32'shebeb259a, 32'shebe9a7ca, 32'shebe829fe, 32'shebe6ac35, 32'shebe52e6f, 32'shebe3b0ac, 32'shebe232ec, 
               32'shebe0b52f, 32'shebdf3776, 32'shebddb9bf, 32'shebdc3c0c, 32'shebdabe5c, 32'shebd940ae, 32'shebd7c304, 32'shebd6455d, 
               32'shebd4c7ba, 32'shebd34a19, 32'shebd1cc7b, 32'shebd04ee1, 32'shebced149, 32'shebcd53b5, 32'shebcbd624, 32'shebca5896, 
               32'shebc8db0b, 32'shebc75d83, 32'shebc5dffe, 32'shebc4627d, 32'shebc2e4fe, 32'shebc16783, 32'shebbfea0b, 32'shebbe6c95, 
               32'shebbcef23, 32'shebbb71b5, 32'shebb9f449, 32'shebb876e0, 32'shebb6f97b, 32'shebb57c18, 32'shebb3feb9, 32'shebb2815d, 
               32'shebb10404, 32'shebaf86ae, 32'shebae095c, 32'shebac8c0c, 32'shebab0ec0, 32'sheba99176, 32'sheba81430, 32'sheba696ed, 
               32'sheba519ad, 32'sheba39c71, 32'sheba21f37, 32'sheba0a200, 32'sheb9f24cd, 32'sheb9da79d, 32'sheb9c2a70, 32'sheb9aad46, 
               32'sheb99301f, 32'sheb97b2fc, 32'sheb9635db, 32'sheb94b8be, 32'sheb933ba4, 32'sheb91be8d, 32'sheb904179, 32'sheb8ec468, 
               32'sheb8d475b, 32'sheb8bca50, 32'sheb8a4d49, 32'sheb88d045, 32'sheb875344, 32'sheb85d646, 32'sheb84594c, 32'sheb82dc54, 
               32'sheb815f60, 32'sheb7fe26f, 32'sheb7e6581, 32'sheb7ce896, 32'sheb7b6bae, 32'sheb79eeca, 32'sheb7871e8, 32'sheb76f50a, 
               32'sheb75782f, 32'sheb73fb57, 32'sheb727e83, 32'sheb7101b1, 32'sheb6f84e3, 32'sheb6e0818, 32'sheb6c8b50, 32'sheb6b0e8b, 
               32'sheb6991ca, 32'sheb68150b, 32'sheb669850, 32'sheb651b98, 32'sheb639ee3, 32'sheb622231, 32'sheb60a582, 32'sheb5f28d7, 
               32'sheb5dac2f, 32'sheb5c2f8a, 32'sheb5ab2e8, 32'sheb593649, 32'sheb57b9ae, 32'sheb563d16, 32'sheb54c081, 32'sheb5343ef, 
               32'sheb51c760, 32'sheb504ad4, 32'sheb4ece4c, 32'sheb4d51c7, 32'sheb4bd545, 32'sheb4a58c6, 32'sheb48dc4b, 32'sheb475fd2, 
               32'sheb45e35d, 32'sheb4466eb, 32'sheb42ea7c, 32'sheb416e11, 32'sheb3ff1a8, 32'sheb3e7543, 32'sheb3cf8e1, 32'sheb3b7c82, 
               32'sheb3a0027, 32'sheb3883ce, 32'sheb370779, 32'sheb358b27, 32'sheb340ed9, 32'sheb32928d, 32'sheb311645, 32'sheb2f99ff, 
               32'sheb2e1dbe, 32'sheb2ca17f, 32'sheb2b2543, 32'sheb29a90b, 32'sheb282cd6, 32'sheb26b0a4, 32'sheb253475, 32'sheb23b84a, 
               32'sheb223c22, 32'sheb20bffd, 32'sheb1f43db, 32'sheb1dc7bc, 32'sheb1c4ba1, 32'sheb1acf89, 32'sheb195374, 32'sheb17d762, 
               32'sheb165b54, 32'sheb14df49, 32'sheb136341, 32'sheb11e73c, 32'sheb106b3a, 32'sheb0eef3c, 32'sheb0d7341, 32'sheb0bf749, 
               32'sheb0a7b54, 32'sheb08ff63, 32'sheb078375, 32'sheb06078a, 32'sheb048ba2, 32'sheb030fbe, 32'sheb0193dd, 32'sheb0017ff, 
               32'sheafe9c24, 32'sheafd204c, 32'sheafba478, 32'sheafa28a7, 32'sheaf8acd9, 32'sheaf7310f, 32'sheaf5b547, 32'sheaf43983, 
               32'sheaf2bdc3, 32'sheaf14205, 32'sheaefc64b, 32'sheaee4a94, 32'sheaeccee0, 32'sheaeb532f, 32'sheae9d782, 32'sheae85bd8, 
               32'sheae6e031, 32'sheae5648e, 32'sheae3e8ed, 32'sheae26d50, 32'sheae0f1b6, 32'sheadf7620, 32'sheaddfa8d, 32'sheadc7efd, 
               32'sheadb0370, 32'shead987e6, 32'shead80c60, 32'shead690dd, 32'shead5155d, 32'shead399e1, 32'shead21e68, 32'shead0a2f2, 
               32'sheacf277f, 32'sheacdac10, 32'sheacc30a4, 32'sheacab53b, 32'sheac939d5, 32'sheac7be73, 32'sheac64314, 32'sheac4c7b8, 
               32'sheac34c60, 32'sheac1d10b, 32'sheac055b9, 32'sheabeda6a, 32'sheabd5f1f, 32'sheabbe3d7, 32'sheaba6892, 32'sheab8ed50, 
               32'sheab77212, 32'sheab5f6d7, 32'sheab47b9f, 32'sheab3006b, 32'sheab1853a, 32'sheab00a0c, 32'sheaae8ee2, 32'sheaad13ba, 
               32'sheaab9896, 32'sheaaa1d76, 32'sheaa8a258, 32'sheaa7273e, 32'sheaa5ac27, 32'sheaa43114, 32'sheaa2b604, 32'sheaa13af7, 
               32'shea9fbfed, 32'shea9e44e7, 32'shea9cc9e4, 32'shea9b4ee4, 32'shea99d3e8, 32'shea9858ee, 32'shea96ddf9, 32'shea956306, 
               32'shea93e817, 32'shea926d2b, 32'shea90f242, 32'shea8f775d, 32'shea8dfc7b, 32'shea8c819c, 32'shea8b06c1, 32'shea898be9, 
               32'shea881114, 32'shea869642, 32'shea851b74, 32'shea83a0a9, 32'shea8225e2, 32'shea80ab1e, 32'shea7f305d, 32'shea7db59f, 
               32'shea7c3ae5, 32'shea7ac02e, 32'shea79457a, 32'shea77caca, 32'shea76501d, 32'shea74d573, 32'shea735acd, 32'shea71e02a, 
               32'shea70658a, 32'shea6eeaee, 32'shea6d7055, 32'shea6bf5bf, 32'shea6a7b2d, 32'shea69009e, 32'shea678612, 32'shea660b8a, 
               32'shea649105, 32'shea631683, 32'shea619c04, 32'shea602189, 32'shea5ea712, 32'shea5d2c9d, 32'shea5bb22c, 32'shea5a37be, 
               32'shea58bd54, 32'shea5742ed, 32'shea55c889, 32'shea544e29, 32'shea52d3cc, 32'shea515972, 32'shea4fdf1c, 32'shea4e64c9, 
               32'shea4cea79, 32'shea4b702d, 32'shea49f5e4, 32'shea487b9e, 32'shea47015c, 32'shea45871d, 32'shea440ce1, 32'shea4292a9, 
               32'shea411874, 32'shea3f9e43, 32'shea3e2415, 32'shea3ca9ea, 32'shea3b2fc2, 32'shea39b59e, 32'shea383b7e, 32'shea36c160, 
               32'shea354746, 32'shea33cd30, 32'shea32531c, 32'shea30d90c, 32'shea2f5f00, 32'shea2de4f7, 32'shea2c6af1, 32'shea2af0ee, 
               32'shea2976ef, 32'shea27fcf4, 32'shea2682fb, 32'shea250906, 32'shea238f15, 32'shea221526, 32'shea209b3b, 32'shea1f2154, 
               32'shea1da770, 32'shea1c2d8f, 32'shea1ab3b2, 32'shea1939d8, 32'shea17c001, 32'shea16462e, 32'shea14cc5e, 32'shea135291, 
               32'shea11d8c8, 32'shea105f03, 32'shea0ee540, 32'shea0d6b81, 32'shea0bf1c6, 32'shea0a780e, 32'shea08fe59, 32'shea0784a7, 
               32'shea060af9, 32'shea04914f, 32'shea0317a7, 32'shea019e04, 32'shea002463, 32'she9feaac6, 32'she9fd312c, 32'she9fbb796, 
               32'she9fa3e03, 32'she9f8c474, 32'she9f74ae8, 32'she9f5d15f, 32'she9f457da, 32'she9f2de58, 32'she9f164d9, 32'she9efeb5e, 
               32'she9ee71e6, 32'she9ecf872, 32'she9eb7f01, 32'she9ea0594, 32'she9e88c2a, 32'she9e712c3, 32'she9e59960, 32'she9e42000, 
               32'she9e2a6a3, 32'she9e12d4a, 32'she9dfb3f5, 32'she9de3aa3, 32'she9dcc154, 32'she9db4808, 32'she9d9cec0, 32'she9d8557c, 
               32'she9d6dc3b, 32'she9d562fd, 32'she9d3e9c3, 32'she9d2708c, 32'she9d0f758, 32'she9cf7e28, 32'she9ce04fc, 32'she9cc8bd3, 
               32'she9cb12ad, 32'she9c9998a, 32'she9c8206b, 32'she9c6a750, 32'she9c52e38, 32'she9c3b523, 32'she9c23c12, 32'she9c0c304, 
               32'she9bf49fa, 32'she9bdd0f3, 32'she9bc57f0, 32'she9badeef, 32'she9b965f3, 32'she9b7ecfa, 32'she9b67404, 32'she9b4fb12, 
               32'she9b38223, 32'she9b20937, 32'she9b0904f, 32'she9af176b, 32'she9ad9e8a, 32'she9ac25ac, 32'she9aaacd2, 32'she9a933fb, 
               32'she9a7bb28, 32'she9a64258, 32'she9a4c98b, 32'she9a350c2, 32'she9a1d7fd, 32'she9a05f3b, 32'she99ee67c, 32'she99d6dc1, 
               32'she99bf509, 32'she99a7c55, 32'she99903a4, 32'she9978af7, 32'she996124d, 32'she99499a6, 32'she9932103, 32'she991a864, 
               32'she9902fc7, 32'she98eb72f, 32'she98d3e9a, 32'she98bc608, 32'she98a4d7a, 32'she988d4ef, 32'she9875c68, 32'she985e3e4, 
               32'she9846b63, 32'she982f2e6, 32'she9817a6d, 32'she98001f7, 32'she97e8984, 32'she97d1115, 32'she97b98aa, 32'she97a2042, 
               32'she978a7dd, 32'she9772f7c, 32'she975b71e, 32'she9743ec4, 32'she972c66d, 32'she9714e1a, 32'she96fd5ca, 32'she96e5d7e, 
               32'she96ce535, 32'she96b6cf0, 32'she969f4ae, 32'she9687c70, 32'she9670435, 32'she9658bfd, 32'she96413c9, 32'she9629b99, 
               32'she961236c, 32'she95fab43, 32'she95e331d, 32'she95cbafa, 32'she95b42db, 32'she959cac0, 32'she95852a8, 32'she956da93, 
               32'she9556282, 32'she953ea75, 32'she952726b, 32'she950fa64, 32'she94f8261, 32'she94e0a62, 32'she94c9266, 32'she94b1a6d, 
               32'she949a278, 32'she9482a87, 32'she946b299, 32'she9453aae, 32'she943c2c7, 32'she9424ae4, 32'she940d304, 32'she93f5b27, 
               32'she93de34e, 32'she93c6b79, 32'she93af3a7, 32'she9397bd8, 32'she938040d, 32'she9368c46, 32'she9351482, 32'she9339cc2, 
               32'she9322505, 32'she930ad4b, 32'she92f3596, 32'she92dbde3, 32'she92c4634, 32'she92ace89, 32'she92956e1, 32'she927df3d, 
               32'she926679c, 32'she924efff, 32'she9237866, 32'she92200cf, 32'she920893d, 32'she91f11ae, 32'she91d9a22, 32'she91c229a, 
               32'she91aab16, 32'she9193395, 32'she917bc17, 32'she916449d, 32'she914cd27, 32'she91355b4, 32'she911de45, 32'she91066d9, 
               32'she90eef71, 32'she90d780c, 32'she90c00ab, 32'she90a894d, 32'she90911f3, 32'she9079a9d, 32'she906234a, 32'she904abfa, 
               32'she90334af, 32'she901bd66, 32'she9004621, 32'she8fecee0, 32'she8fd57a2, 32'she8fbe068, 32'she8fa6932, 32'she8f8f1ff, 
               32'she8f77acf, 32'she8f603a3, 32'she8f48c7b, 32'she8f31556, 32'she8f19e34, 32'she8f02717, 32'she8eeaffd, 32'she8ed38e6, 
               32'she8ebc1d3, 32'she8ea4ac3, 32'she8e8d3b7, 32'she8e75caf, 32'she8e5e5aa, 32'she8e46ea9, 32'she8e2f7ab, 32'she8e180b1, 
               32'she8e009ba, 32'she8de92c7, 32'she8dd1bd8, 32'she8dba4ec, 32'she8da2e04, 32'she8d8b71f, 32'she8d7403e, 32'she8d5c960, 
               32'she8d45286, 32'she8d2dbb0, 32'she8d164dd, 32'she8cfee0e, 32'she8ce7742, 32'she8cd007a, 32'she8cb89b5, 32'she8ca12f4, 
               32'she8c89c37, 32'she8c7257d, 32'she8c5aec7, 32'she8c43814, 32'she8c2c165, 32'she8c14aba, 32'she8bfd412, 32'she8be5d6d, 
               32'she8bce6cd, 32'she8bb702f, 32'she8b9f996, 32'she8b88300, 32'she8b70c6d, 32'she8b595df, 32'she8b41f53, 32'she8b2a8cc, 
               32'she8b13248, 32'she8afbbc7, 32'she8ae454b, 32'she8acced1, 32'she8ab585c, 32'she8a9e1ea, 32'she8a86b7b, 32'she8a6f510, 
               32'she8a57ea9, 32'she8a40845, 32'she8a291e5, 32'she8a11b89, 32'she89fa530, 32'she89e2edb, 32'she89cb889, 32'she89b423b, 
               32'she899cbf1, 32'she89855aa, 32'she896df67, 32'she8956927, 32'she893f2eb, 32'she8927cb3, 32'she891067e, 32'she88f904d, 
               32'she88e1a20, 32'she88ca3f6, 32'she88b2dcf, 32'she889b7ad, 32'she888418e, 32'she886cb72, 32'she885555a, 32'she883df46, 
               32'she8826936, 32'she880f329, 32'she87f7d1f, 32'she87e071a, 32'she87c9118, 32'she87b1b19, 32'she879a51e, 32'she8782f27, 
               32'she876b934, 32'she8754344, 32'she873cd57, 32'she872576f, 32'she870e18a, 32'she86f6ba8, 32'she86df5cb, 32'she86c7ff0, 
               32'she86b0a1a, 32'she8699447, 32'she8681e78, 32'she866a8ac, 32'she86532e4, 32'she863bd20, 32'she862475f, 32'she860d1a2, 
               32'she85f5be9, 32'she85de633, 32'she85c7081, 32'she85afad3, 32'she8598528, 32'she8580f81, 32'she85699dd, 32'she855243d, 
               32'she853aea1, 32'she8523909, 32'she850c374, 32'she84f4de2, 32'she84dd855, 32'she84c62cb, 32'she84aed45, 32'she84977c2, 
               32'she8480243, 32'she8468cc8, 32'she8451750, 32'she843a1dc, 32'she8422c6c, 32'she840b6ff, 32'she83f4196, 32'she83dcc31, 
               32'she83c56cf, 32'she83ae171, 32'she8396c16, 32'she837f6c0, 32'she836816d, 32'she8350c1d, 32'she83396d2, 32'she832218a, 
               32'she830ac45, 32'she82f3705, 32'she82dc1c8, 32'she82c4c8e, 32'she82ad759, 32'she8296227, 32'she827ecf8, 32'she82677ce, 
               32'she82502a7, 32'she8238d84, 32'she8221864, 32'she820a348, 32'she81f2e30, 32'she81db91b, 32'she81c440a, 32'she81acefd, 
               32'she81959f4, 32'she817e4ee, 32'she8166fec, 32'she814faed, 32'she81385f3, 32'she81210fc, 32'she8109c08, 32'she80f2719, 
               32'she80db22d, 32'she80c3d44, 32'she80ac860, 32'she809537f, 32'she807dea2, 32'she80669c8, 32'she804f4f2, 32'she8038020, 
               32'she8020b52, 32'she8009687, 32'she7ff21c0, 32'she7fdacfd, 32'she7fc383d, 32'she7fac381, 32'she7f94ec9, 32'she7f7da14, 
               32'she7f66564, 32'she7f4f0b7, 32'she7f37c0d, 32'she7f20768, 32'she7f092c6, 32'she7ef1e27, 32'she7eda98d, 32'she7ec34f6, 
               32'she7eac063, 32'she7e94bd3, 32'she7e7d748, 32'she7e662c0, 32'she7e4ee3c, 32'she7e379bb, 32'she7e2053e, 32'she7e090c5, 
               32'she7df1c50, 32'she7dda7de, 32'she7dc3370, 32'she7dabf06, 32'she7d94a9f, 32'she7d7d63d, 32'she7d661de, 32'she7d4ed82, 
               32'she7d3792b, 32'she7d204d7, 32'she7d09087, 32'she7cf1c3a, 32'she7cda7f2, 32'she7cc33ad, 32'she7cabf6c, 32'she7c94b2e, 
               32'she7c7d6f4, 32'she7c662be, 32'she7c4ee8c, 32'she7c37a5e, 32'she7c20633, 32'she7c0920c, 32'she7bf1de8, 32'she7bda9c9, 
               32'she7bc35ad, 32'she7bac195, 32'she7b94d80, 32'she7b7d970, 32'she7b66563, 32'she7b4f15a, 32'she7b37d55, 32'she7b20953, 
               32'she7b09555, 32'she7af215b, 32'she7adad65, 32'she7ac3972, 32'she7aac583, 32'she7a95198, 32'she7a7ddb1, 32'she7a669cd, 
               32'she7a4f5ed, 32'she7a38211, 32'she7a20e39, 32'she7a09a64, 32'she79f2693, 32'she79db2c6, 32'she79c3efd, 32'she79acb37, 
               32'she7995776, 32'she797e3b8, 32'she7966ffd, 32'she794fc47, 32'she7938894, 32'she79214e5, 32'she790a13a, 32'she78f2d92, 
               32'she78db9ef, 32'she78c464f, 32'she78ad2b3, 32'she7895f1a, 32'she787eb86, 32'she78677f5, 32'she7850468, 32'she78390df, 
               32'she7821d59, 32'she780a9d8, 32'she77f365a, 32'she77dc2e0, 32'she77c4f69, 32'she77adbf7, 32'she7796888, 32'she777f51d, 
               32'she77681b6, 32'she7750e52, 32'she7739af2, 32'she7722797, 32'she770b43e, 32'she76f40ea, 32'she76dcd9a, 32'she76c5a4d, 
               32'she76ae704, 32'she76973bf, 32'she768007e, 32'she7668d40, 32'she7651a06, 32'she763a6d0, 32'she762339e, 32'she760c070, 
               32'she75f4d45, 32'she75dda1e, 32'she75c66fb, 32'she75af3dc, 32'she75980c1, 32'she7580da9, 32'she7569a95, 32'she7552785, 
               32'she753b479, 32'she7524171, 32'she750ce6c, 32'she74f5b6b, 32'she74de86f, 32'she74c7575, 32'she74b0280, 32'she7498f8f, 
               32'she7481ca1, 32'she746a9b7, 32'she74536d1, 32'she743c3ef, 32'she7425110, 32'she740de35, 32'she73f6b5f, 32'she73df88c, 
               32'she73c85bc, 32'she73b12f1, 32'she739a029, 32'she7382d66, 32'she736baa6, 32'she73547ea, 32'she733d531, 32'she732627d, 
               32'she730efcc, 32'she72f7d20, 32'she72e0a77, 32'she72c97d1, 32'she72b2530, 32'she729b293, 32'she7283ff9, 32'she726cd63, 
               32'she7255ad1, 32'she723e843, 32'she72275b9, 32'she7210332, 32'she71f90b0, 32'she71e1e31, 32'she71cabb6, 32'she71b393f, 
               32'she719c6cb, 32'she718545c, 32'she716e1f0, 32'she7156f89, 32'she713fd25, 32'she7128ac4, 32'she7111868, 32'she70fa610, 
               32'she70e33bb, 32'she70cc16b, 32'she70b4f1e, 32'she709dcd5, 32'she7086a8f, 32'she706f84e, 32'she7058611, 32'she70413d7, 
               32'she702a1a1, 32'she7012f6f, 32'she6ffbd41, 32'she6fe4b17, 32'she6fcd8f1, 32'she6fb66ce, 32'she6f9f4b0, 32'she6f88295, 
               32'she6f7107e, 32'she6f59e6b, 32'she6f42c5c, 32'she6f2ba51, 32'she6f14849, 32'she6efd645, 32'she6ee6446, 32'she6ecf24a, 
               32'she6eb8052, 32'she6ea0e5e, 32'she6e89c6d, 32'she6e72a81, 32'she6e5b899, 32'she6e446b4, 32'she6e2d4d3, 32'she6e162f6, 
               32'she6dff11d, 32'she6de7f48, 32'she6dd0d77, 32'she6db9ba9, 32'she6da29e0, 32'she6d8b81a, 32'she6d74658, 32'she6d5d49b, 
               32'she6d462e1, 32'she6d2f12a, 32'she6d17f78, 32'she6d00dca, 32'she6ce9c1f, 32'she6cd2a79, 32'she6cbb8d6, 32'she6ca4737, 
               32'she6c8d59c, 32'she6c76405, 32'she6c5f272, 32'she6c480e3, 32'she6c30f57, 32'she6c19dd0, 32'she6c02c4c, 32'she6bebacd, 
               32'she6bd4951, 32'she6bbd7d9, 32'she6ba6665, 32'she6b8f4f5, 32'she6b78389, 32'she6b61220, 32'she6b4a0bc, 32'she6b32f5b, 
               32'she6b1bdff, 32'she6b04ca6, 32'she6aedb51, 32'she6ad6a00, 32'she6abf8b3, 32'she6aa876a, 32'she6a91625, 32'she6a7a4e4, 
               32'she6a633a6, 32'she6a4c26d, 32'she6a35137, 32'she6a1e006, 32'she6a06ed8, 32'she69efdae, 32'she69d8c88, 32'she69c1b66, 
               32'she69aaa48, 32'she699392e, 32'she697c818, 32'she6965706, 32'she694e5f7, 32'she69374ed, 32'she69203e6, 32'she69092e4, 
               32'she68f21e5, 32'she68db0ea, 32'she68c3ff3, 32'she68acf00, 32'she6895e11, 32'she687ed26, 32'she6867c3f, 32'she6850b5c, 
               32'she6839a7c, 32'she68229a1, 32'she680b8ca, 32'she67f47f6, 32'she67dd727, 32'she67c665b, 32'she67af593, 32'she67984cf, 
               32'she6781410, 32'she676a354, 32'she675329c, 32'she673c1e8, 32'she6725138, 32'she670e08c, 32'she66f6fe3, 32'she66dff3f, 
               32'she66c8e9f, 32'she66b1e02, 32'she669ad6a, 32'she6683cd5, 32'she666cc45, 32'she6655bb8, 32'she663eb30, 32'she6627aab, 
               32'she6610a2a, 32'she65f99ae, 32'she65e2935, 32'she65cb8c0, 32'she65b484f, 32'she659d7e2, 32'she6586779, 32'she656f714, 
               32'she65586b3, 32'she6541656, 32'she652a5fc, 32'she65135a7, 32'she64fc556, 32'she64e5509, 32'she64ce4bf, 32'she64b747a, 
               32'she64a0438, 32'she64893fb, 32'she64723c2, 32'she645b38c, 32'she644435a, 32'she642d32d, 32'she6416303, 32'she63ff2de, 
               32'she63e82bc, 32'she63d129e, 32'she63ba285, 32'she63a326f, 32'she638c25d, 32'she637524f, 32'she635e245, 32'she6347240, 
               32'she633023e, 32'she6319240, 32'she6302246, 32'she62eb250, 32'she62d425e, 32'she62bd270, 32'she62a6286, 32'she628f2a0, 
               32'she62782be, 32'she62612e0, 32'she624a306, 32'she6233330, 32'she621c35e, 32'she6205390, 32'she61ee3c6, 32'she61d73ff, 
               32'she61c043d, 32'she61a947f, 32'she61924c5, 32'she617b50f, 32'she616455d, 32'she614d5af, 32'she6136605, 32'she611f65e, 
               32'she61086bc, 32'she60f171e, 32'she60da784, 32'she60c37ee, 32'she60ac85c, 32'she60958ce, 32'she607e944, 32'she60679bd, 
               32'she6050a3b, 32'she6039abd, 32'she6022b43, 32'she600bbcd, 32'she5ff4c5b, 32'she5fddced, 32'she5fc6d83, 32'she5fafe1d, 
               32'she5f98ebb, 32'she5f81f5d, 32'she5f6b003, 32'she5f540ad, 32'she5f3d15b, 32'she5f2620d, 32'she5f0f2c3, 32'she5ef837d, 
               32'she5ee143b, 32'she5eca4fd, 32'she5eb35c3, 32'she5e9c68d, 32'she5e8575b, 32'she5e6e82e, 32'she5e57904, 32'she5e409de, 
               32'she5e29abc, 32'she5e12b9f, 32'she5dfbc85, 32'she5de4d6f, 32'she5dcde5e, 32'she5db6f50, 32'she5da0047, 32'she5d89141, 
               32'she5d72240, 32'she5d5b342, 32'she5d44449, 32'she5d2d553, 32'she5d16662, 32'she5cff775, 32'she5ce888b, 32'she5cd19a6, 
               32'she5cbaac5, 32'she5ca3be8, 32'she5c8cd0f, 32'she5c75e3a, 32'she5c5ef69, 32'she5c4809c, 32'she5c311d3, 32'she5c1a30e, 
               32'she5c0344d, 32'she5bec590, 32'she5bd56d7, 32'she5bbe823, 32'she5ba7972, 32'she5b90ac6, 32'she5b79c1d, 32'she5b62d79, 
               32'she5b4bed8, 32'she5b3503c, 32'she5b1e1a3, 32'she5b0730f, 32'she5af047f, 32'she5ad95f3, 32'she5ac276b, 32'she5aab8e7, 
               32'she5a94a67, 32'she5a7dbeb, 32'she5a66d73, 32'she5a4feff, 32'she5a39090, 32'she5a22224, 32'she5a0b3bc, 32'she59f4559, 
               32'she59dd6f9, 32'she59c689e, 32'she59afa47, 32'she5998bf3, 32'she5981da4, 32'she596af59, 32'she5954112, 32'she593d2cf, 
               32'she5926490, 32'she590f656, 32'she58f881f, 32'she58e19ec, 32'she58cabbe, 32'she58b3d93, 32'she589cf6d, 32'she588614a, 
               32'she586f32c, 32'she5858512, 32'she58416fc, 32'she582a8ea, 32'she5813adc, 32'she57fccd2, 32'she57e5ecc, 32'she57cf0cb, 
               32'she57b82cd, 32'she57a14d4, 32'she578a6de, 32'she57738ed, 32'she575cb00, 32'she5745d17, 32'she572ef32, 32'she5718151, 
               32'she5701374, 32'she56ea59b, 32'she56d37c7, 32'she56bc9f6, 32'she56a5c2a, 32'she568ee61, 32'she567809d, 32'she56612dd, 
               32'she564a521, 32'she5633769, 32'she561c9b5, 32'she5605c06, 32'she55eee5a, 32'she55d80b2, 32'she55c130f, 32'she55aa570, 
               32'she55937d5, 32'she557ca3e, 32'she5565cab, 32'she554ef1c, 32'she5538191, 32'she552140a, 32'she550a688, 32'she54f3909, 
               32'she54dcb8f, 32'she54c5e19, 32'she54af0a7, 32'she5498339, 32'she54815cf, 32'she546a86a, 32'she5453b08, 32'she543cdab, 
               32'she5426051, 32'she540f2fc, 32'she53f85ab, 32'she53e185e, 32'she53cab15, 32'she53b3dd1, 32'she539d090, 32'she5386354, 
               32'she536f61b, 32'she53588e7, 32'she5341bb7, 32'she532ae8b, 32'she5314163, 32'she52fd440, 32'she52e6720, 32'she52cfa05, 
               32'she52b8cee, 32'she52a1fdb, 32'she528b2cc, 32'she52745c1, 32'she525d8ba, 32'she5246bb8, 32'she522feb9, 32'she52191bf, 
               32'she52024c9, 32'she51eb7d7, 32'she51d4ae9, 32'she51bddff, 32'she51a711a, 32'she5190438, 32'she517975b, 32'she5162a82, 
               32'she514bdad, 32'she51350dc, 32'she511e410, 32'she5107747, 32'she50f0a83, 32'she50d9dc3, 32'she50c3107, 32'she50ac44f, 
               32'she509579b, 32'she507eaec, 32'she5067e40, 32'she5051199, 32'she503a4f6, 32'she5023857, 32'she500cbbc, 32'she4ff5f26, 
               32'she4fdf294, 32'she4fc8605, 32'she4fb197b, 32'she4f9acf5, 32'she4f84074, 32'she4f6d3f6, 32'she4f5677d, 32'she4f3fb07, 
               32'she4f28e96, 32'she4f12229, 32'she4efb5c1, 32'she4ee495c, 32'she4ecdcfc, 32'she4eb70a0, 32'she4ea0448, 32'she4e897f4, 
               32'she4e72ba4, 32'she4e5bf59, 32'she4e45311, 32'she4e2e6ce, 32'she4e17a8f, 32'she4e00e54, 32'she4dea21e, 32'she4dd35eb, 
               32'she4dbc9bd, 32'she4da5d93, 32'she4d8f16d, 32'she4d7854c, 32'she4d6192e, 32'she4d4ad15, 32'she4d34100, 32'she4d1d4ef, 
               32'she4d068e2, 32'she4cefcda, 32'she4cd90d5, 32'she4cc24d5, 32'she4cab8d9, 32'she4c94ce2, 32'she4c7e0ee, 32'she4c674ff, 
               32'she4c50914, 32'she4c39d2d, 32'she4c2314a, 32'she4c0c56b, 32'she4bf5991, 32'she4bdedbb, 32'she4bc81e9, 32'she4bb161b, 
               32'she4b9aa52, 32'she4b83e8d, 32'she4b6d2cb, 32'she4b5670f, 32'she4b3fb56, 32'she4b28fa1, 32'she4b123f1, 32'she4afb845, 
               32'she4ae4c9d, 32'she4ace0fa, 32'she4ab755a, 32'she4aa09bf, 32'she4a89e28, 32'she4a73295, 32'she4a5c707, 32'she4a45b7c, 
               32'she4a2eff6, 32'she4a18474, 32'she4a018f7, 32'she49ead7d, 32'she49d4208, 32'she49bd697, 32'she49a6b2a, 32'she498ffc1, 
               32'she497945d, 32'she49628fd, 32'she494bda1, 32'she4935249, 32'she491e6f6, 32'she4907ba7, 32'she48f105c, 32'she48da515, 
               32'she48c39d3, 32'she48ace94, 32'she489635a, 32'she487f825, 32'she4868cf3, 32'she48521c6, 32'she483b69d, 32'she4824b78, 
               32'she480e057, 32'she47f753b, 32'she47e0a23, 32'she47c9f0f, 32'she47b33ff, 32'she479c8f4, 32'she4785ded, 32'she476f2ea, 
               32'she47587eb, 32'she4741cf1, 32'she472b1fa, 32'she4714709, 32'she46fdc1b, 32'she46e7131, 32'she46d064c, 32'she46b9b6b, 
               32'she46a308f, 32'she468c5b6, 32'she4675ae2, 32'she465f012, 32'she4648547, 32'she4631a7f, 32'she461afbc, 32'she46044fd, 
               32'she45eda43, 32'she45d6f8c, 32'she45c04da, 32'she45a9a2c, 32'she4592f83, 32'she457c4de, 32'she4565a3c, 32'she454efa0, 
               32'she4538507, 32'she4521a73, 32'she450afe3, 32'she44f4557, 32'she44ddad0, 32'she44c704d, 32'she44b05ce, 32'she4499b53, 
               32'she44830dd, 32'she446c66b, 32'she4455bfd, 32'she443f194, 32'she442872e, 32'she4411ccd, 32'she43fb271, 32'she43e4818, 
               32'she43cddc4, 32'she43b7374, 32'she43a0929, 32'she4389ee2, 32'she437349f, 32'she435ca60, 32'she4346026, 32'she432f5ef, 
               32'she4318bbe, 32'she4302190, 32'she42eb767, 32'she42d4d42, 32'she42be321, 32'she42a7905, 32'she4290eed, 32'she427a4d9, 
               32'she4263ac9, 32'she424d0be, 32'she42366b7, 32'she421fcb5, 32'she42092b6, 32'she41f28bc, 32'she41dbec7, 32'she41c54d5, 
               32'she41aeae8, 32'she41980ff, 32'she418171b, 32'she416ad3a, 32'she415435f, 32'she413d987, 32'she4126fb4, 32'she41105e5, 
               32'she40f9c1a, 32'she40e3254, 32'she40cc891, 32'she40b5ed4, 32'she409f51a, 32'she4088b65, 32'she40721b4, 32'she405b808, 
               32'she4044e60, 32'she402e4bc, 32'she4017b1c, 32'she4001181, 32'she3fea7ea, 32'she3fd3e57, 32'she3fbd4c9, 32'she3fa6b3f, 
               32'she3f901ba, 32'she3f79838, 32'she3f62ebb, 32'she3f4c542, 32'she3f35bce, 32'she3f1f25e, 32'she3f088f2, 32'she3ef1f8b, 
               32'she3edb628, 32'she3ec4cc9, 32'she3eae36f, 32'she3e97a19, 32'she3e810c7, 32'she3e6a77a, 32'she3e53e31, 32'she3e3d4ec, 
               32'she3e26bac, 32'she3e1026f, 32'she3df9938, 32'she3de3004, 32'she3dcc6d5, 32'she3db5dab, 32'she3d9f484, 32'she3d88b62, 
               32'she3d72245, 32'she3d5b92b, 32'she3d45016, 32'she3d2e706, 32'she3d17df9, 32'she3d014f1, 32'she3ceabee, 32'she3cd42ee, 
               32'she3cbd9f4, 32'she3ca70fd, 32'she3c9080b, 32'she3c79f1d, 32'she3c63633, 32'she3c4cd4e, 32'she3c3646d, 32'she3c1fb91, 
               32'she3c092b9, 32'she3bf29e5, 32'she3bdc116, 32'she3bc584b, 32'she3baef84, 32'she3b986c2, 32'she3b81e04, 32'she3b6b54a, 
               32'she3b54c95, 32'she3b3e3e4, 32'she3b27b38, 32'she3b1128f, 32'she3afa9ec, 32'she3ae414c, 32'she3acd8b1, 32'she3ab701b, 
               32'she3aa0788, 32'she3a89efa, 32'she3a73671, 32'she3a5cdec, 32'she3a4656b, 32'she3a2fcee, 32'she3a19476, 32'she3a02c03, 
               32'she39ec393, 32'she39d5b28, 32'she39bf2c2, 32'she39a8a60, 32'she3992202, 32'she397b9a8, 32'she3965153, 32'she394e903, 
               32'she39380b6, 32'she392186f, 32'she390b02b, 32'she38f47ec, 32'she38ddfb1, 32'she38c777b, 32'she38b0f49, 32'she389a71b, 
               32'she3883ef2, 32'she386d6cd, 32'she3856ead, 32'she3840691, 32'she3829e79, 32'she3813666, 32'she37fce57, 32'she37e664d, 
               32'she37cfe47, 32'she37b9645, 32'she37a2e48, 32'she378c64f, 32'she3775e5a, 32'she375f66a, 32'she3748e7f, 32'she3732697, 
               32'she371beb5, 32'she37056d6, 32'she36eeefc, 32'she36d8727, 32'she36c1f55, 32'she36ab788, 32'she3694fc0, 32'she367e7fc, 
               32'she366803c, 32'she3651881, 32'she363b0cb, 32'she3624918, 32'she360e16a, 32'she35f79c1, 32'she35e121c, 32'she35caa7b, 
               32'she35b42df, 32'she359db47, 32'she35873b3, 32'she3570c24, 32'she355a49a, 32'she3543d13, 32'she352d592, 32'she3516e14, 
               32'she350069b, 32'she34e9f27, 32'she34d37b7, 32'she34bd04b, 32'she34a68e4, 32'she3490181, 32'she3479a23, 32'she34632c9, 
               32'she344cb73, 32'she3436422, 32'she341fcd6, 32'she340958d, 32'she33f2e4a, 32'she33dc70a, 32'she33c5fcf, 32'she33af899, 
               32'she3399167, 32'she3382a39, 32'she336c310, 32'she3355beb, 32'she333f4cb, 32'she3328daf, 32'she3312698, 32'she32fbf85, 
               32'she32e5876, 32'she32cf16c, 32'she32b8a67, 32'she32a2365, 32'she328bc69, 32'she3275570, 32'she325ee7d, 32'she324878d, 
               32'she32320a2, 32'she321b9bc, 32'she32052da, 32'she31eebfc, 32'she31d8523, 32'she31c1e4e, 32'she31ab77e, 32'she31950b2, 
               32'she317e9eb, 32'she3168328, 32'she3151c6a, 32'she313b5b0, 32'she3124efa, 32'she310e849, 32'she30f819d, 32'she30e1af5, 
               32'she30cb451, 32'she30b4db2, 32'she309e717, 32'she3088081, 32'she30719ef, 32'she305b362, 32'she3044cd9, 32'she302e655, 
               32'she3017fd5, 32'she300195a, 32'she2feb2e3, 32'she2fd4c70, 32'she2fbe602, 32'she2fa7f99, 32'she2f91934, 32'she2f7b2d3, 
               32'she2f64c77, 32'she2f4e61f, 32'she2f37fcc, 32'she2f2197e, 32'she2f0b333, 32'she2ef4cee, 32'she2ede6ac, 32'she2ec8070, 
               32'she2eb1a37, 32'she2e9b404, 32'she2e84dd4, 32'she2e6e7aa, 32'she2e58183, 32'she2e41b62, 32'she2e2b544, 32'she2e14f2b, 
               32'she2dfe917, 32'she2de8307, 32'she2dd1cfc, 32'she2dbb6f5, 32'she2da50f3, 32'she2d8eaf5, 32'she2d784fb, 32'she2d61f07, 
               32'she2d4b916, 32'she2d3532a, 32'she2d1ed43, 32'she2d08760, 32'she2cf2182, 32'she2cdbba8, 32'she2cc55d2, 32'she2caf001, 
               32'she2c98a35, 32'she2c8246d, 32'she2c6beaa, 32'she2c558eb, 32'she2c3f331, 32'she2c28d7b, 32'she2c127c9, 32'she2bfc21d, 
               32'she2be5c74, 32'she2bcf6d1, 32'she2bb9131, 32'she2ba2b96, 32'she2b8c600, 32'she2b7606e, 32'she2b5fae1, 32'she2b49559, 
               32'she2b32fd4, 32'she2b1ca55, 32'she2b064da, 32'she2aeff63, 32'she2ad99f1, 32'she2ac3483, 32'she2aacf1a, 32'she2a969b6, 
               32'she2a80456, 32'she2a69efa, 32'she2a539a3, 32'she2a3d451, 32'she2a26f03, 32'she2a109b9, 32'she29fa474, 32'she29e3f34, 
               32'she29cd9f8, 32'she29b74c1, 32'she29a0f8e, 32'she298aa60, 32'she2974536, 32'she295e011, 32'she2947af1, 32'she29315d5, 
               32'she291b0bd, 32'she2904baa, 32'she28ee69c, 32'she28d8192, 32'she28c1c8c, 32'she28ab78c, 32'she289528f, 32'she287ed98, 
               32'she28688a4, 32'she28523b6, 32'she283becc, 32'she28259e6, 32'she280f505, 32'she27f9029, 32'she27e2b51, 32'she27cc67d, 
               32'she27b61af, 32'she279fce4, 32'she278981f, 32'she277335e, 32'she275cea1, 32'she27469e9, 32'she2730536, 32'she271a087, 
               32'she2703bdc, 32'she26ed736, 32'she26d7295, 32'she26c0df9, 32'she26aa960, 32'she26944cd, 32'she267e03e, 32'she2667bb3, 
               32'she265172e, 32'she263b2ac, 32'she2624e2f, 32'she260e9b7, 32'she25f8544, 32'she25e20d5, 32'she25cbc6a, 32'she25b5804, 
               32'she259f3a3, 32'she2588f46, 32'she2572aee, 32'she255c69b, 32'she254624b, 32'she252fe01, 32'she25199bb, 32'she250357a, 
               32'she24ed13d, 32'she24d6d05, 32'she24c08d1, 32'she24aa4a2, 32'she2494078, 32'she247dc52, 32'she2467831, 32'she2451414, 
               32'she243affc, 32'she2424be9, 32'she240e7da, 32'she23f83d0, 32'she23e1fca, 32'she23cbbc9, 32'she23b57cc, 32'she239f3d4, 
               32'she2388fe1, 32'she2372bf2, 32'she235c808, 32'she2346422, 32'she2330041, 32'she2319c65, 32'she230388d, 32'she22ed4ba, 
               32'she22d70eb, 32'she22c0d21, 32'she22aa95c, 32'she229459b, 32'she227e1df, 32'she2267e28, 32'she2251a75, 32'she223b6c6, 
               32'she222531c, 32'she220ef77, 32'she21f8bd7, 32'she21e283b, 32'she21cc4a3, 32'she21b6111, 32'she219fd82, 32'she21899f9, 
               32'she2173674, 32'she215d2f4, 32'she2146f78, 32'she2130c01, 32'she211a88f, 32'she2104521, 32'she20ee1b7, 32'she20d7e53, 
               32'she20c1af3, 32'she20ab798, 32'she2095441, 32'she207f0ef, 32'she2068da1, 32'she2052a58, 32'she203c714, 32'she20263d4, 
               32'she2010099, 32'she1ff9d63, 32'she1fe3a31, 32'she1fcd704, 32'she1fb73dc, 32'she1fa10b8, 32'she1f8ad98, 32'she1f74a7e, 
               32'she1f5e768, 32'she1f48457, 32'she1f3214a, 32'she1f1be42, 32'she1f05b3e, 32'she1eef83f, 32'she1ed9545, 32'she1ec3250, 
               32'she1eacf5f, 32'she1e96c73, 32'she1e8098b, 32'she1e6a6a8, 32'she1e543ca, 32'she1e3e0f0, 32'she1e27e1b, 32'she1e11b4b, 
               32'she1dfb87f, 32'she1de55b8, 32'she1dcf2f5, 32'she1db9037, 32'she1da2d7e, 32'she1d8caca, 32'she1d7681a, 32'she1d6056f, 
               32'she1d4a2c8, 32'she1d34026, 32'she1d1dd89, 32'she1d07af0, 32'she1cf185c, 32'she1cdb5cd, 32'she1cc5342, 32'she1caf0bc, 
               32'she1c98e3b, 32'she1c82bbe, 32'she1c6c946, 32'she1c566d3, 32'she1c40464, 32'she1c2a1fa, 32'she1c13f95, 32'she1bfdd34, 
               32'she1be7ad8, 32'she1bd1881, 32'she1bbb62e, 32'she1ba53e0, 32'she1b8f197, 32'she1b78f52, 32'she1b62d12, 32'she1b4cad7, 
               32'she1b368a0, 32'she1b2066e, 32'she1b0a441, 32'she1af4218, 32'she1addff4, 32'she1ac7dd5, 32'she1ab1bba, 32'she1a9b9a4, 
               32'she1a85793, 32'she1a6f586, 32'she1a5937e, 32'she1a4317b, 32'she1a2cf7c, 32'she1a16d83, 32'she1a00b8d, 32'she19ea99d, 
               32'she19d47b1, 32'she19be5ca, 32'she19a83e7, 32'she199220a, 32'she197c031, 32'she1965e5c, 32'she194fc8d, 32'she1939ac2, 
               32'she19238fb, 32'she190d73a, 32'she18f757d, 32'she18e13c4, 32'she18cb211, 32'she18b5062, 32'she189eeb8, 32'she1888d13, 
               32'she1872b72, 32'she185c9d6, 32'she184683e, 32'she18306ac, 32'she181a51e, 32'she1804395, 32'she17ee210, 32'she17d8090, 
               32'she17c1f15, 32'she17abd9f, 32'she1795c2d, 32'she177fac0, 32'she1769958, 32'she17537f4, 32'she173d695, 32'she172753b, 
               32'she17113e5, 32'she16fb295, 32'she16e5149, 32'she16cf001, 32'she16b8ebf, 32'she16a2d81, 32'she168cc48, 32'she1676b13, 
               32'she16609e3, 32'she164a8b8, 32'she1634792, 32'she161e671, 32'she1608554, 32'she15f243c, 32'she15dc328, 32'she15c621a, 
               32'she15b0110, 32'she159a00a, 32'she1583f0a, 32'she156de0e, 32'she1557d17, 32'she1541c25, 32'she152bb37, 32'she1515a4e, 
               32'she14ff96a, 32'she14e988b, 32'she14d37b0, 32'she14bd6da, 32'she14a7609, 32'she149153c, 32'she147b475, 32'she14653b2, 
               32'she144f2f3, 32'she143923a, 32'she1423185, 32'she140d0d5, 32'she13f702a, 32'she13e0f83, 32'she13caee1, 32'she13b4e44, 
               32'she139edac, 32'she1388d19, 32'she1372c8a, 32'she135cc00, 32'she1346b7a, 32'she1330afa, 32'she131aa7e, 32'she1304a07, 
               32'she12ee995, 32'she12d8927, 32'she12c28be, 32'she12ac85a, 32'she12967fb, 32'she12807a0, 32'she126a74a, 32'she12546f9, 
               32'she123e6ad, 32'she1228666, 32'she1212623, 32'she11fc5e5, 32'she11e65ac, 32'she11d0577, 32'she11ba547, 32'she11a451c, 
               32'she118e4f6, 32'she11784d5, 32'she11624b8, 32'she114c4a0, 32'she113648d, 32'she112047f, 32'she110a475, 32'she10f4470, 
               32'she10de470, 32'she10c8475, 32'she10b247f, 32'she109c48d, 32'she10864a0, 32'she10704b8, 32'she105a4d4, 32'she10444f6, 
               32'she102e51c, 32'she1018547, 32'she1002577, 32'she0fec5ab, 32'she0fd65e4, 32'she0fc0622, 32'she0faa665, 32'she0f946ad, 
               32'she0f7e6f9, 32'she0f6874a, 32'she0f527a0, 32'she0f3c7fb, 32'she0f2685b, 32'she0f108bf, 32'she0efa928, 32'she0ee4996, 
               32'she0ecea09, 32'she0eb8a80, 32'she0ea2afd, 32'she0e8cb7e, 32'she0e76c04, 32'she0e60c8e, 32'she0e4ad1e, 32'she0e34db2, 
               32'she0e1ee4b, 32'she0e08ee9, 32'she0df2f8c, 32'she0ddd033, 32'she0dc70e0, 32'she0db1191, 32'she0d9b247, 32'she0d85301, 
               32'she0d6f3c1, 32'she0d59485, 32'she0d4354e, 32'she0d2d61c, 32'she0d176ef, 32'she0d017c6, 32'she0ceb8a3, 32'she0cd5984, 
               32'she0cbfa6a, 32'she0ca9b55, 32'she0c93c44, 32'she0c7dd39, 32'she0c67e32, 32'she0c51f30, 32'she0c3c033, 32'she0c2613a, 
               32'she0c10247, 32'she0bfa358, 32'she0be446e, 32'she0bce589, 32'she0bb86a9, 32'she0ba27cd, 32'she0b8c8f7, 32'she0b76a25, 
               32'she0b60b58, 32'she0b4ac90, 32'she0b34dcd, 32'she0b1ef0e, 32'she0b09055, 32'she0af31a0, 32'she0add2f0, 32'she0ac7445, 
               32'she0ab159e, 32'she0a9b6fd, 32'she0a85860, 32'she0a6f9c8, 32'she0a59b35, 32'she0a43ca7, 32'she0a2de1e, 32'she0a17f99, 
               32'she0a0211a, 32'she09ec29f, 32'she09d6429, 32'she09c05b8, 32'she09aa74b, 32'she09948e4, 32'she097ea81, 32'she0968c24, 
               32'she0952dcb, 32'she093cf77, 32'she0927127, 32'she09112dd, 32'she08fb497, 32'she08e5657, 32'she08cf81b, 32'she08b99e4, 
               32'she08a3bb2, 32'she088dd85, 32'she0877f5c, 32'she0862139, 32'she084c31a, 32'she0836500, 32'she08206eb, 32'she080a8db, 
               32'she07f4acf, 32'she07decc9, 32'she07c8ec7, 32'she07b30cb, 32'she079d2d3, 32'she07874e0, 32'she07716f2, 32'she075b908, 
               32'she0745b24, 32'she072fd44, 32'she0719f6a, 32'she0704194, 32'she06ee3c3, 32'she06d85f7, 32'she06c2830, 32'she06aca6d, 
               32'she0696cb0, 32'she0680ef7, 32'she066b144, 32'she0655395, 32'she063f5eb, 32'she0629846, 32'she0613aa5, 32'she05fdd0a, 
               32'she05e7f74, 32'she05d21e2, 32'she05bc455, 32'she05a66cd, 32'she059094a, 32'she057abcc, 32'she0564e53, 32'she054f0df, 
               32'she053936f, 32'she0523605, 32'she050d89f, 32'she04f7b3e, 32'she04e1de3, 32'she04cc08c, 32'she04b6339, 32'she04a05ec, 
               32'she048a8a4, 32'she0474b60, 32'she045ee22, 32'she04490e8, 32'she04333b3, 32'she041d684, 32'she0407959, 32'she03f1c33, 
               32'she03dbf11, 32'she03c61f5, 32'she03b04de, 32'she039a7cb, 32'she0384abe, 32'she036edb5, 32'she03590b1, 32'she03433b2, 
               32'she032d6b8, 32'she03179c3, 32'she0301cd3, 32'she02ebfe8, 32'she02d6301, 32'she02c0620, 32'she02aa943, 32'she0294c6c, 
               32'she027ef99, 32'she02692cb, 32'she0253602, 32'she023d93e, 32'she0227c7f, 32'she0211fc5, 32'she01fc310, 32'she01e6660, 
               32'she01d09b4, 32'she01bad0e, 32'she01a506c, 32'she018f3cf, 32'she0179738, 32'she0163aa5, 32'she014de17, 32'she013818e, 
               32'she012250a, 32'she010c88b, 32'she00f6c11, 32'she00e0f9b, 32'she00cb32b, 32'she00b56bf, 32'she009fa59, 32'she0089df7, 
               32'she007419b, 32'she005e543, 32'she00488f0, 32'she0032ca2, 32'she001d05a, 32'she0007416, 32'shdfff17d7, 32'shdffdbb9c, 
               32'shdffc5f67, 32'shdffb0337, 32'shdff9a70c, 32'shdff84ae5, 32'shdff6eec4, 32'shdff592a7, 32'shdff43690, 32'shdff2da7d, 
               32'shdff17e70, 32'shdff02267, 32'shdfeec663, 32'shdfed6a64, 32'shdfec0e6a, 32'shdfeab276, 32'shdfe95686, 32'shdfe7fa9b, 
               32'shdfe69eb4, 32'shdfe542d3, 32'shdfe3e6f7, 32'shdfe28b20, 32'shdfe12f4e, 32'shdfdfd380, 32'shdfde77b8, 32'shdfdd1bf5, 
               32'shdfdbc036, 32'shdfda647d, 32'shdfd908c8, 32'shdfd7ad18, 32'shdfd6516e, 32'shdfd4f5c8, 32'shdfd39a27, 32'shdfd23e8c, 
               32'shdfd0e2f5, 32'shdfcf8763, 32'shdfce2bd6, 32'shdfccd04e, 32'shdfcb74cb, 32'shdfca194d, 32'shdfc8bdd4, 32'shdfc76260, 
               32'shdfc606f1, 32'shdfc4ab87, 32'shdfc35022, 32'shdfc1f4c2, 32'shdfc09967, 32'shdfbf3e11, 32'shdfbde2bf, 32'shdfbc8773, 
               32'shdfbb2c2c, 32'shdfb9d0ea, 32'shdfb875ac, 32'shdfb71a74, 32'shdfb5bf41, 32'shdfb46412, 32'shdfb308e9, 32'shdfb1adc4, 
               32'shdfb052a5, 32'shdfaef78b, 32'shdfad9c75, 32'shdfac4165, 32'shdfaae659, 32'shdfa98b53, 32'shdfa83051, 32'shdfa6d554, 
               32'shdfa57a5d, 32'shdfa41f6a, 32'shdfa2c47d, 32'shdfa16994, 32'shdfa00eb1, 32'shdf9eb3d2, 32'shdf9d58f8, 32'shdf9bfe24, 
               32'shdf9aa354, 32'shdf99488a, 32'shdf97edc4, 32'shdf969303, 32'shdf953848, 32'shdf93dd91, 32'shdf9282df, 32'shdf912833, 
               32'shdf8fcd8b, 32'shdf8e72e8, 32'shdf8d184b, 32'shdf8bbdb2, 32'shdf8a631f, 32'shdf890890, 32'shdf87ae06, 32'shdf865382, 
               32'shdf84f902, 32'shdf839e88, 32'shdf824412, 32'shdf80e9a2, 32'shdf7f8f36, 32'shdf7e34cf, 32'shdf7cda6e, 32'shdf7b8011, 
               32'shdf7a25ba, 32'shdf78cb67, 32'shdf77711a, 32'shdf7616d2, 32'shdf74bc8e, 32'shdf736250, 32'shdf720816, 32'shdf70ade2, 
               32'shdf6f53b3, 32'shdf6df988, 32'shdf6c9f63, 32'shdf6b4543, 32'shdf69eb27, 32'shdf689111, 32'shdf673700, 32'shdf65dcf4, 
               32'shdf6482ed, 32'shdf6328eb, 32'shdf61ceee, 32'shdf6074f5, 32'shdf5f1b02, 32'shdf5dc114, 32'shdf5c672b, 32'shdf5b0d48, 
               32'shdf59b369, 32'shdf58598f, 32'shdf56ffba, 32'shdf55a5ea, 32'shdf544c1f, 32'shdf52f25a, 32'shdf519899, 32'shdf503edd, 
               32'shdf4ee527, 32'shdf4d8b75, 32'shdf4c31c9, 32'shdf4ad821, 32'shdf497e7f, 32'shdf4824e1, 32'shdf46cb49, 32'shdf4571b6, 
               32'shdf441828, 32'shdf42be9e, 32'shdf41651a, 32'shdf400b9b, 32'shdf3eb221, 32'shdf3d58ac, 32'shdf3bff3c, 32'shdf3aa5d1, 
               32'shdf394c6b, 32'shdf37f30b, 32'shdf3699af, 32'shdf354058, 32'shdf33e707, 32'shdf328dba, 32'shdf313473, 32'shdf2fdb30, 
               32'shdf2e81f3, 32'shdf2d28bb, 32'shdf2bcf87, 32'shdf2a7659, 32'shdf291d30, 32'shdf27c40c, 32'shdf266aed, 32'shdf2511d3, 
               32'shdf23b8be, 32'shdf225fae, 32'shdf2106a4, 32'shdf1fad9e, 32'shdf1e549d, 32'shdf1cfba2, 32'shdf1ba2ab, 32'shdf1a49ba, 
               32'shdf18f0ce, 32'shdf1797e7, 32'shdf163f04, 32'shdf14e627, 32'shdf138d4f, 32'shdf12347c, 32'shdf10dbaf, 32'shdf0f82e6, 
               32'shdf0e2a22, 32'shdf0cd163, 32'shdf0b78aa, 32'shdf0a1ff5, 32'shdf08c746, 32'shdf076e9c, 32'shdf0615f7, 32'shdf04bd57, 
               32'shdf0364bc, 32'shdf020c26, 32'shdf00b395, 32'shdeff5b09, 32'shdefe0282, 32'shdefcaa01, 32'shdefb5184, 32'shdef9f90d, 
               32'shdef8a09b, 32'shdef7482d, 32'shdef5efc5, 32'shdef49762, 32'shdef33f04, 32'shdef1e6ab, 32'shdef08e58, 32'shdeef3609, 
               32'shdeedddc0, 32'shdeec857b, 32'shdeeb2d3c, 32'shdee9d502, 32'shdee87ccc, 32'shdee7249c, 32'shdee5cc72, 32'shdee4744c, 
               32'shdee31c2b, 32'shdee1c40f, 32'shdee06bf9, 32'shdedf13e8, 32'shdeddbbdb, 32'shdedc63d4, 32'shdedb0bd2, 32'shded9b3d5, 
               32'shded85bdd, 32'shded703eb, 32'shded5abfd, 32'shded45414, 32'shded2fc31, 32'shded1a453, 32'shded04c7a, 32'shdecef4a6, 
               32'shdecd9cd7, 32'shdecc450d, 32'shdecaed48, 32'shdec99589, 32'shdec83dce, 32'shdec6e619, 32'shdec58e69, 32'shdec436be, 
               32'shdec2df18, 32'shdec18777, 32'shdec02fdb, 32'shdebed845, 32'shdebd80b3, 32'shdebc2927, 32'shdebad1a0, 32'shdeb97a1e, 
               32'shdeb822a1, 32'shdeb6cb29, 32'shdeb573b7, 32'shdeb41c49, 32'shdeb2c4e1, 32'shdeb16d7d, 32'shdeb0161f, 32'shdeaebec6, 
               32'shdead6773, 32'shdeac1024, 32'shdeaab8da, 32'shdea96196, 32'shdea80a57, 32'shdea6b31d, 32'shdea55be8, 32'shdea404b8, 
               32'shdea2ad8d, 32'shdea15668, 32'shde9fff47, 32'shde9ea82c, 32'shde9d5116, 32'shde9bfa05, 32'shde9aa2f9, 32'shde994bf2, 
               32'shde97f4f1, 32'shde969df5, 32'shde9546fd, 32'shde93f00b, 32'shde92991e, 32'shde914237, 32'shde8feb54, 32'shde8e9477, 
               32'shde8d3d9e, 32'shde8be6cb, 32'shde8a8ffd, 32'shde893935, 32'shde87e271, 32'shde868bb2, 32'shde8534f9, 32'shde83de45, 
               32'shde828796, 32'shde8130ec, 32'shde7fda48, 32'shde7e83a8, 32'shde7d2d0e, 32'shde7bd679, 32'shde7a7fe9, 32'shde79295e, 
               32'shde77d2d8, 32'shde767c58, 32'shde7525dc, 32'shde73cf66, 32'shde7278f5, 32'shde71228a, 32'shde6fcc23, 32'shde6e75c2, 
               32'shde6d1f65, 32'shde6bc90e, 32'shde6a72bc, 32'shde691c70, 32'shde67c628, 32'shde666fe6, 32'shde6519a9, 32'shde63c371, 
               32'shde626d3e, 32'shde611710, 32'shde5fc0e8, 32'shde5e6ac4, 32'shde5d14a6, 32'shde5bbe8d, 32'shde5a687a, 32'shde59126b, 
               32'shde57bc62, 32'shde56665e, 32'shde55105f, 32'shde53ba65, 32'shde526471, 32'shde510e81, 32'shde4fb897, 32'shde4e62b2, 
               32'shde4d0cd2, 32'shde4bb6f8, 32'shde4a6122, 32'shde490b52, 32'shde47b587, 32'shde465fc2, 32'shde450a01, 32'shde43b446, 
               32'shde425e8f, 32'shde4108de, 32'shde3fb333, 32'shde3e5d8c, 32'shde3d07eb, 32'shde3bb24f, 32'shde3a5cb8, 32'shde390726, 
               32'shde37b199, 32'shde365c12, 32'shde350690, 32'shde33b113, 32'shde325b9b, 32'shde310629, 32'shde2fb0bc, 32'shde2e5b54, 
               32'shde2d05f1, 32'shde2bb093, 32'shde2a5b3b, 32'shde2905e8, 32'shde27b09a, 32'shde265b51, 32'shde25060e, 32'shde23b0cf, 
               32'shde225b96, 32'shde210662, 32'shde1fb134, 32'shde1e5c0a, 32'shde1d06e6, 32'shde1bb1c7, 32'shde1a5cad, 32'shde190799, 
               32'shde17b28a, 32'shde165d80, 32'shde15087b, 32'shde13b37b, 32'shde125e81, 32'shde11098c, 32'shde0fb49c, 32'shde0e5fb1, 
               32'shde0d0acc, 32'shde0bb5ec, 32'shde0a6111, 32'shde090c3b, 32'shde07b76b, 32'shde06629f, 32'shde050dd9, 32'shde03b919, 
               32'shde02645d, 32'shde010fa7, 32'shddffbaf6, 32'shddfe664a, 32'shddfd11a3, 32'shddfbbd02, 32'shddfa6866, 32'shddf913cf, 
               32'shddf7bf3e, 32'shddf66ab1, 32'shddf5162a, 32'shddf3c1a9, 32'shddf26d2c, 32'shddf118b5, 32'shddefc443, 32'shddee6fd6, 
               32'shdded1b6e, 32'shddebc70c, 32'shddea72af, 32'shdde91e57, 32'shdde7ca05, 32'shdde675b7, 32'shdde5216f, 32'shdde3cd2d, 
               32'shdde278ef, 32'shdde124b7, 32'shdddfd084, 32'shddde7c56, 32'shdddd282e, 32'shdddbd40b, 32'shddda7fed, 32'shddd92bd4, 
               32'shddd7d7c1, 32'shddd683b3, 32'shddd52faa, 32'shddd3dba6, 32'shddd287a8, 32'shddd133af, 32'shddcfdfbb, 32'shddce8bcd, 
               32'shddcd37e4, 32'shddcbe400, 32'shddca9021, 32'shddc93c48, 32'shddc7e873, 32'shddc694a5, 32'shddc540db, 32'shddc3ed17, 
               32'shddc29958, 32'shddc1459e, 32'shddbff1ea, 32'shddbe9e3a, 32'shddbd4a91, 32'shddbbf6ec, 32'shddbaa34d, 32'shddb94fb3, 
               32'shddb7fc1e, 32'shddb6a88f, 32'shddb55504, 32'shddb4017f, 32'shddb2ae00, 32'shddb15a86, 32'shddb00711, 32'shddaeb3a1, 
               32'shddad6036, 32'shddac0cd1, 32'shddaab972, 32'shdda96617, 32'shdda812c2, 32'shdda6bf72, 32'shdda56c27, 32'shdda418e2, 
               32'shdda2c5a2, 32'shdda17267, 32'shdda01f32, 32'shdd9ecc01, 32'shdd9d78d7, 32'shdd9c25b1, 32'shdd9ad291, 32'shdd997f76, 
               32'shdd982c60, 32'shdd96d950, 32'shdd958645, 32'shdd94333f, 32'shdd92e03f, 32'shdd918d44, 32'shdd903a4e, 32'shdd8ee75d, 
               32'shdd8d9472, 32'shdd8c418c, 32'shdd8aeeac, 32'shdd899bd1, 32'shdd8848fb, 32'shdd86f62a, 32'shdd85a35f, 32'shdd845099, 
               32'shdd82fdd8, 32'shdd81ab1d, 32'shdd805867, 32'shdd7f05b6, 32'shdd7db30b, 32'shdd7c6065, 32'shdd7b0dc4, 32'shdd79bb29, 
               32'shdd786892, 32'shdd771602, 32'shdd75c376, 32'shdd7470f0, 32'shdd731e6f, 32'shdd71cbf4, 32'shdd70797e, 32'shdd6f270d, 
               32'shdd6dd4a2, 32'shdd6c823b, 32'shdd6b2fdb, 32'shdd69dd7f, 32'shdd688b29, 32'shdd6738d8, 32'shdd65e68d, 32'shdd649447, 
               32'shdd634206, 32'shdd61efcb, 32'shdd609d94, 32'shdd5f4b64, 32'shdd5df938, 32'shdd5ca712, 32'shdd5b54f1, 32'shdd5a02d6, 
               32'shdd58b0c0, 32'shdd575eaf, 32'shdd560ca4, 32'shdd54ba9e, 32'shdd53689d, 32'shdd5216a2, 32'shdd50c4ac, 32'shdd4f72bb, 
               32'shdd4e20d0, 32'shdd4cceea, 32'shdd4b7d09, 32'shdd4a2b2e, 32'shdd48d958, 32'shdd478788, 32'shdd4635bd, 32'shdd44e3f7, 
               32'shdd439236, 32'shdd42407b, 32'shdd40eec5, 32'shdd3f9d15, 32'shdd3e4b6a, 32'shdd3cf9c4, 32'shdd3ba824, 32'shdd3a5689, 
               32'shdd3904f4, 32'shdd37b363, 32'shdd3661d8, 32'shdd351053, 32'shdd33bed3, 32'shdd326d58, 32'shdd311be3, 32'shdd2fca73, 
               32'shdd2e7908, 32'shdd2d27a3, 32'shdd2bd643, 32'shdd2a84e8, 32'shdd293393, 32'shdd27e243, 32'shdd2690f9, 32'shdd253fb4, 
               32'shdd23ee74, 32'shdd229d3a, 32'shdd214c05, 32'shdd1ffad5, 32'shdd1ea9ab, 32'shdd1d5886, 32'shdd1c0767, 32'shdd1ab64d, 
               32'shdd196538, 32'shdd181429, 32'shdd16c31f, 32'shdd15721b, 32'shdd14211b, 32'shdd12d022, 32'shdd117f2d, 32'shdd102e3e, 
               32'shdd0edd55, 32'shdd0d8c71, 32'shdd0c3b92, 32'shdd0aeab9, 32'shdd0999e4, 32'shdd084916, 32'shdd06f84d, 32'shdd05a789, 
               32'shdd0456ca, 32'shdd030611, 32'shdd01b55e, 32'shdd0064af, 32'shdcff1407, 32'shdcfdc363, 32'shdcfc72c5, 32'shdcfb222c, 
               32'shdcf9d199, 32'shdcf8810b, 32'shdcf73083, 32'shdcf5e000, 32'shdcf48f82, 32'shdcf33f0a, 32'shdcf1ee97, 32'shdcf09e2a, 
               32'shdcef4dc2, 32'shdcedfd5f, 32'shdcecad02, 32'shdceb5caa, 32'shdcea0c58, 32'shdce8bc0b, 32'shdce76bc3, 32'shdce61b81, 
               32'shdce4cb44, 32'shdce37b0d, 32'shdce22adb, 32'shdce0daae, 32'shdcdf8a87, 32'shdcde3a66, 32'shdcdcea49, 32'shdcdb9a32, 
               32'shdcda4a21, 32'shdcd8fa15, 32'shdcd7aa0e, 32'shdcd65a0d, 32'shdcd50a12, 32'shdcd3ba1b, 32'shdcd26a2a, 32'shdcd11a3f, 
               32'shdccfca59, 32'shdcce7a78, 32'shdccd2a9d, 32'shdccbdac7, 32'shdcca8af7, 32'shdcc93b2c, 32'shdcc7eb67, 32'shdcc69ba7, 
               32'shdcc54bec, 32'shdcc3fc37, 32'shdcc2ac87, 32'shdcc15cdd, 32'shdcc00d38, 32'shdcbebd99, 32'shdcbd6dff, 32'shdcbc1e6a, 
               32'shdcbacedb, 32'shdcb97f51, 32'shdcb82fcd, 32'shdcb6e04e, 32'shdcb590d5, 32'shdcb44161, 32'shdcb2f1f3, 32'shdcb1a28a, 
               32'shdcb05326, 32'shdcaf03c8, 32'shdcadb46f, 32'shdcac651c, 32'shdcab15ce, 32'shdca9c686, 32'shdca87743, 32'shdca72805, 
               32'shdca5d8cd, 32'shdca4899b, 32'shdca33a6e, 32'shdca1eb46, 32'shdca09c24, 32'shdc9f4d07, 32'shdc9dfdf0, 32'shdc9caede, 
               32'shdc9b5fd2, 32'shdc9a10cb, 32'shdc98c1ca, 32'shdc9772ce, 32'shdc9623d7, 32'shdc94d4e6, 32'shdc9385fa, 32'shdc923714, 
               32'shdc90e834, 32'shdc8f9958, 32'shdc8e4a83, 32'shdc8cfbb2, 32'shdc8bace8, 32'shdc8a5e22, 32'shdc890f62, 32'shdc87c0a8, 
               32'shdc8671f3, 32'shdc852344, 32'shdc83d49a, 32'shdc8285f5, 32'shdc813756, 32'shdc7fe8bc, 32'shdc7e9a28, 32'shdc7d4b9a, 
               32'shdc7bfd11, 32'shdc7aae8d, 32'shdc79600f, 32'shdc781196, 32'shdc76c323, 32'shdc7574b5, 32'shdc74264d, 32'shdc72d7ea, 
               32'shdc71898d, 32'shdc703b35, 32'shdc6eece2, 32'shdc6d9e96, 32'shdc6c504e, 32'shdc6b020c, 32'shdc69b3d0, 32'shdc686599, 
               32'shdc671768, 32'shdc65c93c, 32'shdc647b15, 32'shdc632cf4, 32'shdc61ded9, 32'shdc6090c3, 32'shdc5f42b2, 32'shdc5df4a7, 
               32'shdc5ca6a2, 32'shdc5b58a2, 32'shdc5a0aa8, 32'shdc58bcb3, 32'shdc576ec3, 32'shdc5620d9, 32'shdc54d2f5, 32'shdc538516, 
               32'shdc52373c, 32'shdc50e968, 32'shdc4f9b9a, 32'shdc4e4dd1, 32'shdc4d000d, 32'shdc4bb24f, 32'shdc4a6497, 32'shdc4916e4, 
               32'shdc47c936, 32'shdc467b8e, 32'shdc452dec, 32'shdc43e04f, 32'shdc4292b8, 32'shdc414526, 32'shdc3ff799, 32'shdc3eaa12, 
               32'shdc3d5c91, 32'shdc3c0f15, 32'shdc3ac19f, 32'shdc39742e, 32'shdc3826c3, 32'shdc36d95d, 32'shdc358bfd, 32'shdc343ea2, 
               32'shdc32f14d, 32'shdc31a3fd, 32'shdc3056b3, 32'shdc2f096e, 32'shdc2dbc2f, 32'shdc2c6ef5, 32'shdc2b21c1, 32'shdc29d493, 
               32'shdc28876a, 32'shdc273a46, 32'shdc25ed28, 32'shdc24a010, 32'shdc2352fd, 32'shdc2205f0, 32'shdc20b8e8, 32'shdc1f6be5, 
               32'shdc1e1ee9, 32'shdc1cd1f1, 32'shdc1b8500, 32'shdc1a3813, 32'shdc18eb2d, 32'shdc179e4c, 32'shdc165170, 32'shdc15049a, 
               32'shdc13b7c9, 32'shdc126afe, 32'shdc111e39, 32'shdc0fd179, 32'shdc0e84bf, 32'shdc0d380a, 32'shdc0beb5b, 32'shdc0a9eb1, 
               32'shdc09520d, 32'shdc08056e, 32'shdc06b8d5, 32'shdc056c42, 32'shdc041fb4, 32'shdc02d32b, 32'shdc0186a8, 32'shdc003a2b, 
               32'shdbfeedb3, 32'shdbfda141, 32'shdbfc54d4, 32'shdbfb086d, 32'shdbf9bc0c, 32'shdbf86fb0, 32'shdbf72359, 32'shdbf5d708, 
               32'shdbf48abd, 32'shdbf33e77, 32'shdbf1f237, 32'shdbf0a5fc, 32'shdbef59c7, 32'shdbee0d98, 32'shdbecc16e, 32'shdbeb7549, 
               32'shdbea292b, 32'shdbe8dd11, 32'shdbe790fe, 32'shdbe644ef, 32'shdbe4f8e7, 32'shdbe3ace4, 32'shdbe260e6, 32'shdbe114ef, 
               32'shdbdfc8fc, 32'shdbde7d10, 32'shdbdd3128, 32'shdbdbe547, 32'shdbda996b, 32'shdbd94d94, 32'shdbd801c3, 32'shdbd6b5f8, 
               32'shdbd56a32, 32'shdbd41e72, 32'shdbd2d2b8, 32'shdbd18703, 32'shdbd03b53, 32'shdbceefaa, 32'shdbcda405, 32'shdbcc5867, 
               32'shdbcb0cce, 32'shdbc9c13a, 32'shdbc875ac, 32'shdbc72a24, 32'shdbc5dea1, 32'shdbc49324, 32'shdbc347ac, 32'shdbc1fc3a, 
               32'shdbc0b0ce, 32'shdbbf6567, 32'shdbbe1a06, 32'shdbbcceaa, 32'shdbbb8354, 32'shdbba3804, 32'shdbb8ecb9, 32'shdbb7a174, 
               32'shdbb65634, 32'shdbb50afa, 32'shdbb3bfc6, 32'shdbb27497, 32'shdbb1296e, 32'shdbafde4a, 32'shdbae932c, 32'shdbad4814, 
               32'shdbabfd01, 32'shdbaab1f3, 32'shdba966ec, 32'shdba81bea, 32'shdba6d0ed, 32'shdba585f7, 32'shdba43b05, 32'shdba2f01a, 
               32'shdba1a534, 32'shdba05a53, 32'shdb9f0f78, 32'shdb9dc4a3, 32'shdb9c79d4, 32'shdb9b2f0a, 32'shdb99e445, 32'shdb989987, 
               32'shdb974ece, 32'shdb96041a, 32'shdb94b96c, 32'shdb936ec4, 32'shdb922421, 32'shdb90d984, 32'shdb8f8eed, 32'shdb8e445b, 
               32'shdb8cf9cf, 32'shdb8baf48, 32'shdb8a64c7, 32'shdb891a4c, 32'shdb87cfd6, 32'shdb868566, 32'shdb853afc, 32'shdb83f097, 
               32'shdb82a638, 32'shdb815bde, 32'shdb80118a, 32'shdb7ec73c, 32'shdb7d7cf3, 32'shdb7c32b0, 32'shdb7ae873, 32'shdb799e3b, 
               32'shdb785409, 32'shdb7709dc, 32'shdb75bfb5, 32'shdb747594, 32'shdb732b79, 32'shdb71e163, 32'shdb709752, 32'shdb6f4d48, 
               32'shdb6e0342, 32'shdb6cb943, 32'shdb6b6f49, 32'shdb6a2555, 32'shdb68db67, 32'shdb67917e, 32'shdb66479b, 32'shdb64fdbd, 
               32'shdb63b3e5, 32'shdb626a13, 32'shdb612046, 32'shdb5fd67f, 32'shdb5e8cbe, 32'shdb5d4302, 32'shdb5bf94c, 32'shdb5aaf9c, 
               32'shdb5965f1, 32'shdb581c4c, 32'shdb56d2ac, 32'shdb558913, 32'shdb543f7e, 32'shdb52f5f0, 32'shdb51ac67, 32'shdb5062e4, 
               32'shdb4f1967, 32'shdb4dcfef, 32'shdb4c867d, 32'shdb4b3d10, 32'shdb49f3a9, 32'shdb48aa48, 32'shdb4760ec, 32'shdb461797, 
               32'shdb44ce46, 32'shdb4384fc, 32'shdb423bb7, 32'shdb40f278, 32'shdb3fa93e, 32'shdb3e600a, 32'shdb3d16dc, 32'shdb3bcdb3, 
               32'shdb3a8491, 32'shdb393b73, 32'shdb37f25c, 32'shdb36a94a, 32'shdb35603e, 32'shdb341737, 32'shdb32ce36, 32'shdb31853b, 
               32'shdb303c46, 32'shdb2ef356, 32'shdb2daa6c, 32'shdb2c6187, 32'shdb2b18a9, 32'shdb29cfcf, 32'shdb2886fc, 32'shdb273e2e, 
               32'shdb25f566, 32'shdb24aca4, 32'shdb2363e7, 32'shdb221b30, 32'shdb20d27f, 32'shdb1f89d3, 32'shdb1e412d, 32'shdb1cf88d, 
               32'shdb1baff2, 32'shdb1a675e, 32'shdb191ece, 32'shdb17d645, 32'shdb168dc1, 32'shdb154543, 32'shdb13fccb, 32'shdb12b458, 
               32'shdb116beb, 32'shdb102383, 32'shdb0edb22, 32'shdb0d92c6, 32'shdb0c4a70, 32'shdb0b021f, 32'shdb09b9d4, 32'shdb08718f, 
               32'shdb072950, 32'shdb05e116, 32'shdb0498e2, 32'shdb0350b4, 32'shdb02088b, 32'shdb00c068, 32'shdaff784b, 32'shdafe3033, 
               32'shdafce821, 32'shdafba015, 32'shdafa580f, 32'shdaf9100e, 32'shdaf7c813, 32'shdaf6801e, 32'shdaf5382e, 32'shdaf3f045, 
               32'shdaf2a860, 32'shdaf16082, 32'shdaf018a9, 32'shdaeed0d6, 32'shdaed8909, 32'shdaec4141, 32'shdaeaf980, 32'shdae9b1c4, 
               32'shdae86a0d, 32'shdae7225c, 32'shdae5dab2, 32'shdae4930c, 32'shdae34b6d, 32'shdae203d3, 32'shdae0bc3f, 32'shdadf74b1, 
               32'shdade2d28, 32'shdadce5a5, 32'shdadb9e28, 32'shdada56b0, 32'shdad90f3f, 32'shdad7c7d3, 32'shdad6806d, 32'shdad5390c, 
               32'shdad3f1b1, 32'shdad2aa5c, 32'shdad1630d, 32'shdad01bc3, 32'shdaced47f, 32'shdacd8d41, 32'shdacc4609, 32'shdacafed6, 
               32'shdac9b7a9, 32'shdac87082, 32'shdac72961, 32'shdac5e245, 32'shdac49b2f, 32'shdac3541f, 32'shdac20d15, 32'shdac0c610, 
               32'shdabf7f11, 32'shdabe3818, 32'shdabcf124, 32'shdabbaa36, 32'shdaba634e, 32'shdab91c6c, 32'shdab7d590, 32'shdab68eb9, 
               32'shdab547e8, 32'shdab4011d, 32'shdab2ba57, 32'shdab17397, 32'shdab02cdd, 32'shdaaee629, 32'shdaad9f7b, 32'shdaac58d2, 
               32'shdaab122f, 32'shdaa9cb92, 32'shdaa884fa, 32'shdaa73e69, 32'shdaa5f7dd, 32'shdaa4b157, 32'shdaa36ad6, 32'shdaa2245c, 
               32'shdaa0dde7, 32'shda9f9778, 32'shda9e510e, 32'shda9d0aab, 32'shda9bc44d, 32'shda9a7df5, 32'shda9937a2, 32'shda97f156, 
               32'shda96ab0f, 32'shda9564ce, 32'shda941e93, 32'shda92d85d, 32'shda91922e, 32'shda904c04, 32'shda8f05e0, 32'shda8dbfc1, 
               32'shda8c79a9, 32'shda8b3396, 32'shda89ed89, 32'shda88a782, 32'shda876180, 32'shda861b84, 32'shda84d58f, 32'shda838f9e, 
               32'shda8249b4, 32'shda8103cf, 32'shda7fbdf1, 32'shda7e7818, 32'shda7d3244, 32'shda7bec77, 32'shda7aa6af, 32'shda7960ed, 
               32'shda781b31, 32'shda76d57b, 32'shda758fcb, 32'shda744a20, 32'shda73047b, 32'shda71bedc, 32'shda707942, 32'shda6f33af, 
               32'shda6dee21, 32'shda6ca899, 32'shda6b6317, 32'shda6a1d9b, 32'shda68d824, 32'shda6792b3, 32'shda664d48, 32'shda6507e3, 
               32'shda63c284, 32'shda627d2a, 32'shda6137d6, 32'shda5ff288, 32'shda5ead40, 32'shda5d67fe, 32'shda5c22c1, 32'shda5add8a, 
               32'shda599859, 32'shda58532e, 32'shda570e09, 32'shda55c8e9, 32'shda5483d0, 32'shda533ebc, 32'shda51f9ae, 32'shda50b4a5, 
               32'shda4f6fa3, 32'shda4e2aa6, 32'shda4ce5af, 32'shda4ba0be, 32'shda4a5bd3, 32'shda4916ed, 32'shda47d20e, 32'shda468d34, 
               32'shda454860, 32'shda440392, 32'shda42beca, 32'shda417a07, 32'shda40354a, 32'shda3ef093, 32'shda3dabe2, 32'shda3c6737, 
               32'shda3b2292, 32'shda39ddf2, 32'shda389958, 32'shda3754c4, 32'shda361036, 32'shda34cbae, 32'shda33872c, 32'shda3242af, 
               32'shda30fe38, 32'shda2fb9c7, 32'shda2e755c, 32'shda2d30f7, 32'shda2bec97, 32'shda2aa83e, 32'shda2963ea, 32'shda281f9c, 
               32'shda26db54, 32'shda259711, 32'shda2452d5, 32'shda230e9e, 32'shda21ca6e, 32'shda208643, 32'shda1f421e, 32'shda1dfdfe, 
               32'shda1cb9e5, 32'shda1b75d1, 32'shda1a31c4, 32'shda18edbc, 32'shda17a9ba, 32'shda1665be, 32'shda1521c7, 32'shda13ddd7, 
               32'shda1299ec, 32'shda115607, 32'shda101228, 32'shda0ece4f, 32'shda0d8a7c, 32'shda0c46af, 32'shda0b02e7, 32'shda09bf25, 
               32'shda087b69, 32'shda0737b3, 32'shda05f403, 32'shda04b059, 32'shda036cb5, 32'shda022916, 32'shda00e57d, 32'shd9ffa1eb, 
               32'shd9fe5e5e, 32'shd9fd1ad6, 32'shd9fbd755, 32'shd9fa93da, 32'shd9f95064, 32'shd9f80cf5, 32'shd9f6c98b, 32'shd9f58627, 
               32'shd9f442c9, 32'shd9f2ff71, 32'shd9f1bc1e, 32'shd9f078d2, 32'shd9ef358b, 32'shd9edf24b, 32'shd9ecaf10, 32'shd9eb6bdb, 
               32'shd9ea28ac, 32'shd9e8e582, 32'shd9e7a25f, 32'shd9e65f42, 32'shd9e51c2a, 32'shd9e3d918, 32'shd9e2960c, 32'shd9e15306, 
               32'shd9e01006, 32'shd9decd0c, 32'shd9dd8a18, 32'shd9dc4729, 32'shd9db0441, 32'shd9d9c15e, 32'shd9d87e81, 32'shd9d73baa, 
               32'shd9d5f8d9, 32'shd9d4b60e, 32'shd9d37349, 32'shd9d23089, 32'shd9d0edd0, 32'shd9cfab1c, 32'shd9ce686e, 32'shd9cd25c7, 
               32'shd9cbe325, 32'shd9caa089, 32'shd9c95df3, 32'shd9c81b62, 32'shd9c6d8d8, 32'shd9c59653, 32'shd9c453d5, 32'shd9c3115c, 
               32'shd9c1cee9, 32'shd9c08c7c, 32'shd9bf4a15, 32'shd9be07b4, 32'shd9bcc559, 32'shd9bb8304, 32'shd9ba40b5, 32'shd9b8fe6b, 
               32'shd9b7bc27, 32'shd9b679ea, 32'shd9b537b2, 32'shd9b3f580, 32'shd9b2b354, 32'shd9b1712e, 32'shd9b02f0e, 32'shd9aeecf4, 
               32'shd9adaadf, 32'shd9ac68d1, 32'shd9ab26c8, 32'shd9a9e4c6, 32'shd9a8a2c9, 32'shd9a760d2, 32'shd9a61ee1, 32'shd9a4dcf6, 
               32'shd9a39b11, 32'shd9a25932, 32'shd9a11759, 32'shd99fd586, 32'shd99e93b8, 32'shd99d51f1, 32'shd99c102f, 32'shd99ace74, 
               32'shd9998cbe, 32'shd9984b0e, 32'shd9970965, 32'shd995c7c1, 32'shd9948623, 32'shd993448b, 32'shd99202f8, 32'shd990c16c, 
               32'shd98f7fe6, 32'shd98e3e66, 32'shd98cfceb, 32'shd98bbb77, 32'shd98a7a08, 32'shd989389f, 32'shd987f73d, 32'shd986b5e0, 
               32'shd9857489, 32'shd9843338, 32'shd982f1ed, 32'shd981b0a8, 32'shd9806f69, 32'shd97f2e30, 32'shd97decfd, 32'shd97cabcf, 
               32'shd97b6aa8, 32'shd97a2986, 32'shd978e86b, 32'shd977a755, 32'shd9766646, 32'shd975253c, 32'shd973e438, 32'shd972a33b, 
               32'shd9716243, 32'shd9702151, 32'shd96ee065, 32'shd96d9f7f, 32'shd96c5e9f, 32'shd96b1dc5, 32'shd969dcf1, 32'shd9689c23, 
               32'shd9675b5a, 32'shd9661a98, 32'shd964d9dc, 32'shd9639926, 32'shd9625875, 32'shd96117cb, 32'shd95fd726, 32'shd95e9688, 
               32'shd95d55ef, 32'shd95c155c, 32'shd95ad4d0, 32'shd9599449, 32'shd95853c8, 32'shd957134d, 32'shd955d2d9, 32'shd954926a, 
               32'shd9535201, 32'shd952119e, 32'shd950d141, 32'shd94f90ea, 32'shd94e5099, 32'shd94d104e, 32'shd94bd009, 32'shd94a8fca, 
               32'shd9494f90, 32'shd9480f5d, 32'shd946cf30, 32'shd9458f09, 32'shd9444ee7, 32'shd9430ecc, 32'shd941ceb7, 32'shd9408ea7, 
               32'shd93f4e9e, 32'shd93e0e9b, 32'shd93cce9d, 32'shd93b8ea6, 32'shd93a4eb4, 32'shd9390ec9, 32'shd937cee3, 32'shd9368f04, 
               32'shd9354f2a, 32'shd9340f56, 32'shd932cf89, 32'shd9318fc1, 32'shd9305000, 32'shd92f1044, 32'shd92dd08e, 32'shd92c90df, 
               32'shd92b5135, 32'shd92a1191, 32'shd928d1f4, 32'shd927925c, 32'shd92652ca, 32'shd925133e, 32'shd923d3b9, 32'shd9229439, 
               32'shd92154bf, 32'shd920154b, 32'shd91ed5de, 32'shd91d9676, 32'shd91c5714, 32'shd91b17b8, 32'shd919d863, 32'shd9189913, 
               32'shd91759c9, 32'shd9161a85, 32'shd914db47, 32'shd9139c10, 32'shd9125cde, 32'shd9111db2, 32'shd90fde8c, 32'shd90e9f6d, 
               32'shd90d6053, 32'shd90c213f, 32'shd90ae231, 32'shd909a32a, 32'shd9086428, 32'shd907252c, 32'shd905e636, 32'shd904a747, 
               32'shd903685d, 32'shd9022979, 32'shd900ea9c, 32'shd8ffabc4, 32'shd8fe6cf2, 32'shd8fd2e27, 32'shd8fbef61, 32'shd8fab0a2, 
               32'shd8f971e8, 32'shd8f83335, 32'shd8f6f487, 32'shd8f5b5df, 32'shd8f4773e, 32'shd8f338a3, 32'shd8f1fa0d, 32'shd8f0bb7e, 
               32'shd8ef7cf4, 32'shd8ee3e71, 32'shd8ecfff4, 32'shd8ebc17c, 32'shd8ea830b, 32'shd8e944a0, 32'shd8e8063a, 32'shd8e6c7db, 
               32'shd8e58982, 32'shd8e44b2f, 32'shd8e30ce2, 32'shd8e1ce9b, 32'shd8e0905a, 32'shd8df521f, 32'shd8de13ea, 32'shd8dcd5bb, 
               32'shd8db9792, 32'shd8da596f, 32'shd8d91b52, 32'shd8d7dd3b, 32'shd8d69f2a, 32'shd8d56120, 32'shd8d4231b, 32'shd8d2e51c, 
               32'shd8d1a724, 32'shd8d06931, 32'shd8cf2b45, 32'shd8cded5e, 32'shd8ccaf7e, 32'shd8cb71a3, 32'shd8ca33cf, 32'shd8c8f601, 
               32'shd8c7b838, 32'shd8c67a76, 32'shd8c53cba, 32'shd8c3ff04, 32'shd8c2c154, 32'shd8c183aa, 32'shd8c04606, 32'shd8bf0868, 
               32'shd8bdcad0, 32'shd8bc8d3e, 32'shd8bb4fb3, 32'shd8ba122d, 32'shd8b8d4ad, 32'shd8b79734, 32'shd8b659c0, 32'shd8b51c53, 
               32'shd8b3deeb, 32'shd8b2a18a, 32'shd8b1642f, 32'shd8b026da, 32'shd8aee98a, 32'shd8adac41, 32'shd8ac6efe, 32'shd8ab31c1, 
               32'shd8a9f48a, 32'shd8a8b75a, 32'shd8a77a2f, 32'shd8a63d0a, 32'shd8a4ffec, 32'shd8a3c2d3, 32'shd8a285c0, 32'shd8a148b4, 
               32'shd8a00bae, 32'shd89ecead, 32'shd89d91b3, 32'shd89c54bf, 32'shd89b17d1, 32'shd899dae9, 32'shd8989e07, 32'shd897612b, 
               32'shd8962456, 32'shd894e786, 32'shd893aabc, 32'shd8926df9, 32'shd891313b, 32'shd88ff484, 32'shd88eb7d3, 32'shd88d7b28, 
               32'shd88c3e83, 32'shd88b01e4, 32'shd889c54b, 32'shd88888b8, 32'shd8874c2b, 32'shd8860fa4, 32'shd884d324, 32'shd88396a9, 
               32'shd8825a35, 32'shd8811dc7, 32'shd87fe15e, 32'shd87ea4fc, 32'shd87d68a0, 32'shd87c2c4a, 32'shd87aeffa, 32'shd879b3b1, 
               32'shd878776d, 32'shd8773b2f, 32'shd875fef8, 32'shd874c2c7, 32'shd873869b, 32'shd8724a76, 32'shd8710e57, 32'shd86fd23e, 
               32'shd86e962b, 32'shd86d5a1e, 32'shd86c1e18, 32'shd86ae217, 32'shd869a61d, 32'shd8686a28, 32'shd8672e3a, 32'shd865f252, 
               32'shd864b670, 32'shd8637a94, 32'shd8623ebe, 32'shd86102ee, 32'shd85fc725, 32'shd85e8b61, 32'shd85d4fa4, 32'shd85c13ed, 
               32'shd85ad83c, 32'shd8599c91, 32'shd85860ec, 32'shd857254d, 32'shd855e9b4, 32'shd854ae21, 32'shd8537295, 32'shd852370f, 
               32'shd850fb8e, 32'shd84fc014, 32'shd84e84a0, 32'shd84d4933, 32'shd84c0dcb, 32'shd84ad269, 32'shd849970e, 32'shd8485bb8, 
               32'shd8472069, 32'shd845e520, 32'shd844a9dd, 32'shd8436ea0, 32'shd8423369, 32'shd840f839, 32'shd83fbd0e, 32'shd83e81ea, 
               32'shd83d46cc, 32'shd83c0bb4, 32'shd83ad0a2, 32'shd8399596, 32'shd8385a90, 32'shd8371f91, 32'shd835e497, 32'shd834a9a4, 
               32'shd8336eb7, 32'shd83233d0, 32'shd830f8ef, 32'shd82fbe14, 32'shd82e833f, 32'shd82d4871, 32'shd82c0da9, 32'shd82ad2e7, 
               32'shd829982b, 32'shd8285d75, 32'shd82722c5, 32'shd825e81b, 32'shd824ad78, 32'shd82372db, 32'shd8223843, 32'shd820fdb2, 
               32'shd81fc328, 32'shd81e88a3, 32'shd81d4e24, 32'shd81c13ac, 32'shd81ad93a, 32'shd8199ecd, 32'shd8186468, 32'shd8172a08, 
               32'shd815efae, 32'shd814b55b, 32'shd8137b0d, 32'shd81240c6, 32'shd8110685, 32'shd80fcc4a, 32'shd80e9216, 32'shd80d57e7, 
               32'shd80c1dbf, 32'shd80ae39c, 32'shd809a980, 32'shd8086f6a, 32'shd807355b, 32'shd805fb51, 32'shd804c14e, 32'shd8038751, 
               32'shd8024d59, 32'shd8011369, 32'shd7ffd97e, 32'shd7fe9f99, 32'shd7fd65bb, 32'shd7fc2be3, 32'shd7faf211, 32'shd7f9b845, 
               32'shd7f87e7f, 32'shd7f744bf, 32'shd7f60b06, 32'shd7f4d153, 32'shd7f397a6, 32'shd7f25dff, 32'shd7f1245e, 32'shd7efeac4, 
               32'shd7eeb130, 32'shd7ed77a1, 32'shd7ec3e1a, 32'shd7eb0498, 32'shd7e9cb1c, 32'shd7e891a7, 32'shd7e75838, 32'shd7e61ece, 
               32'shd7e4e56c, 32'shd7e3ac0f, 32'shd7e272b8, 32'shd7e13968, 32'shd7e0001e, 32'shd7dec6da, 32'shd7dd8d9c, 32'shd7dc5465, 
               32'shd7db1b34, 32'shd7d9e208, 32'shd7d8a8e3, 32'shd7d76fc5, 32'shd7d636ac, 32'shd7d4fd9a, 32'shd7d3c48d, 32'shd7d28b87, 
               32'shd7d15288, 32'shd7d0198e, 32'shd7cee09b, 32'shd7cda7ad, 32'shd7cc6ec6, 32'shd7cb35e6, 32'shd7c9fd0b, 32'shd7c8c436, 
               32'shd7c78b68, 32'shd7c652a0, 32'shd7c519de, 32'shd7c3e123, 32'shd7c2a86d, 32'shd7c16fbe, 32'shd7c03715, 32'shd7befe72, 
               32'shd7bdc5d6, 32'shd7bc8d40, 32'shd7bb54af, 32'shd7ba1c25, 32'shd7b8e3a2, 32'shd7b7ab24, 32'shd7b672ad, 32'shd7b53a3c, 
               32'shd7b401d1, 32'shd7b2c96c, 32'shd7b1910e, 32'shd7b058b6, 32'shd7af2063, 32'shd7ade818, 32'shd7acafd2, 32'shd7ab7793, 
               32'shd7aa3f5a, 32'shd7a90727, 32'shd7a7cefa, 32'shd7a696d3, 32'shd7a55eb3, 32'shd7a42699, 32'shd7a2ee85, 32'shd7a1b678, 
               32'shd7a07e70, 32'shd79f466f, 32'shd79e0e74, 32'shd79cd680, 32'shd79b9e91, 32'shd79a66a9, 32'shd7992ec7, 32'shd797f6eb, 
               32'shd796bf16, 32'shd7958746, 32'shd7944f7d, 32'shd79317ba, 32'shd791dffe, 32'shd790a847, 32'shd78f7097, 32'shd78e38ed, 
               32'shd78d014a, 32'shd78bc9ac, 32'shd78a9215, 32'shd7895a84, 32'shd78822f9, 32'shd786eb75, 32'shd785b3f7, 32'shd7847c7f, 
               32'shd783450d, 32'shd7820da1, 32'shd780d63c, 32'shd77f9edd, 32'shd77e6784, 32'shd77d3032, 32'shd77bf8e6, 32'shd77ac1a0, 
               32'shd7798a60, 32'shd7785326, 32'shd7771bf3, 32'shd775e4c6, 32'shd774ad9f, 32'shd773767f, 32'shd7723f64, 32'shd7710850, 
               32'shd76fd143, 32'shd76e9a3b, 32'shd76d633a, 32'shd76c2c3f, 32'shd76af54a, 32'shd769be5c, 32'shd7688774, 32'shd7675092, 
               32'shd76619b6, 32'shd764e2e0, 32'shd763ac11, 32'shd7627548, 32'shd7613e86, 32'shd76007c9, 32'shd75ed113, 32'shd75d9a63, 
               32'shd75c63ba, 32'shd75b2d17, 32'shd759f679, 32'shd758bfe3, 32'shd7578952, 32'shd75652c8, 32'shd7551c44, 32'shd753e5c6, 
               32'shd752af4f, 32'shd75178de, 32'shd7504273, 32'shd74f0c0e, 32'shd74dd5b0, 32'shd74c9f58, 32'shd74b6906, 32'shd74a32bb, 
               32'shd748fc75, 32'shd747c636, 32'shd7468ffe, 32'shd74559cb, 32'shd744239f, 32'shd742ed79, 32'shd741b75a, 32'shd7408141, 
               32'shd73f4b2e, 32'shd73e1521, 32'shd73cdf1b, 32'shd73ba91a, 32'shd73a7321, 32'shd7393d2d, 32'shd7380740, 32'shd736d159, 
               32'shd7359b78, 32'shd734659e, 32'shd7332fca, 32'shd731f9fc, 32'shd730c434, 32'shd72f8e73, 32'shd72e58b8, 32'shd72d2304, 
               32'shd72bed55, 32'shd72ab7ad, 32'shd729820c, 32'shd7284c70, 32'shd72716db, 32'shd725e14c, 32'shd724abc4, 32'shd7237641, 
               32'shd72240c5, 32'shd7210b50, 32'shd71fd5e0, 32'shd71ea077, 32'shd71d6b15, 32'shd71c35b8, 32'shd71b0062, 32'shd719cb12, 
               32'shd71895c9, 32'shd7176086, 32'shd7162b49, 32'shd714f612, 32'shd713c0e2, 32'shd7128bb8, 32'shd7115694, 32'shd7102177, 
               32'shd70eec60, 32'shd70db74f, 32'shd70c8245, 32'shd70b4d41, 32'shd70a1843, 32'shd708e34c, 32'shd707ae5a, 32'shd7067970, 
               32'shd705448b, 32'shd7040fad, 32'shd702dad5, 32'shd701a604, 32'shd7007138, 32'shd6ff3c73, 32'shd6fe07b5, 32'shd6fcd2fd, 
               32'shd6fb9e4b, 32'shd6fa699f, 32'shd6f934fa, 32'shd6f8005b, 32'shd6f6cbc2, 32'shd6f59730, 32'shd6f462a4, 32'shd6f32e1f, 
               32'shd6f1f99f, 32'shd6f0c526, 32'shd6ef90b4, 32'shd6ee5c47, 32'shd6ed27e1, 32'shd6ebf382, 32'shd6eabf28, 32'shd6e98ad6, 
               32'shd6e85689, 32'shd6e72243, 32'shd6e5ee03, 32'shd6e4b9c9, 32'shd6e38596, 32'shd6e25169, 32'shd6e11d42, 32'shd6dfe922, 
               32'shd6deb508, 32'shd6dd80f5, 32'shd6dc4ce7, 32'shd6db18e0, 32'shd6d9e4e0, 32'shd6d8b0e6, 32'shd6d77cf2, 32'shd6d64904, 
               32'shd6d5151d, 32'shd6d3e13d, 32'shd6d2ad62, 32'shd6d1798e, 32'shd6d045c0, 32'shd6cf11f9, 32'shd6cdde38, 32'shd6ccaa7d, 
               32'shd6cb76c9, 32'shd6ca431b, 32'shd6c90f73, 32'shd6c7dbd2, 32'shd6c6a837, 32'shd6c574a2, 32'shd6c44114, 32'shd6c30d8c, 
               32'shd6c1da0b, 32'shd6c0a690, 32'shd6bf731b, 32'shd6be3fad, 32'shd6bd0c45, 32'shd6bbd8e3, 32'shd6baa588, 32'shd6b97233, 
               32'shd6b83ee4, 32'shd6b70b9c, 32'shd6b5d85a, 32'shd6b4a51f, 32'shd6b371ea, 32'shd6b23ebb, 32'shd6b10b92, 32'shd6afd870, 
               32'shd6aea555, 32'shd6ad7240, 32'shd6ac3f31, 32'shd6ab0c28, 32'shd6a9d926, 32'shd6a8a62a, 32'shd6a77335, 32'shd6a64046, 
               32'shd6a50d5d, 32'shd6a3da7b, 32'shd6a2a79f, 32'shd6a174ca, 32'shd6a041fa, 32'shd69f0f32, 32'shd69ddc6f, 32'shd69ca9b3, 
               32'shd69b76fe, 32'shd69a444f, 32'shd69911a6, 32'shd697df03, 32'shd696ac67, 32'shd69579d2, 32'shd6944742, 32'shd69314b9, 
               32'shd691e237, 32'shd690afbb, 32'shd68f7d45, 32'shd68e4ad6, 32'shd68d186d, 32'shd68be60a, 32'shd68ab3ae, 32'shd6898158, 
               32'shd6884f09, 32'shd6871cc0, 32'shd685ea7d, 32'shd684b841, 32'shd683860b, 32'shd68253dc, 32'shd68121b3, 32'shd67fef90, 
               32'shd67ebd74, 32'shd67d8b5e, 32'shd67c594f, 32'shd67b2746, 32'shd679f543, 32'shd678c347, 32'shd6779151, 32'shd6765f62, 
               32'shd6752d79, 32'shd673fb97, 32'shd672c9ba, 32'shd67197e5, 32'shd6706615, 32'shd66f344c, 32'shd66e028a, 32'shd66cd0ce, 
               32'shd66b9f18, 32'shd66a6d69, 32'shd6693bc0, 32'shd6680a1d, 32'shd666d881, 32'shd665a6ec, 32'shd664755c, 32'shd66343d4, 
               32'shd6621251, 32'shd660e0d5, 32'shd65faf60, 32'shd65e7df1, 32'shd65d4c88, 32'shd65c1b26, 32'shd65ae9ca, 32'shd659b874, 
               32'shd6588725, 32'shd65755dd, 32'shd656249b, 32'shd654f35f, 32'shd653c229, 32'shd65290fb, 32'shd6515fd2, 32'shd6502eb0, 
               32'shd64efd94, 32'shd64dcc7f, 32'shd64c9b71, 32'shd64b6a68, 32'shd64a3966, 32'shd649086b, 32'shd647d776, 32'shd646a687, 
               32'shd645759f, 32'shd64444bd, 32'shd64313e2, 32'shd641e30d, 32'shd640b23f, 32'shd63f8177, 32'shd63e50b5, 32'shd63d1ffa, 
               32'shd63bef46, 32'shd63abe97, 32'shd6398df0, 32'shd6385d4e, 32'shd6372cb3, 32'shd635fc1f, 32'shd634cb91, 32'shd6339b09, 
               32'shd6326a88, 32'shd6313a0e, 32'shd6300999, 32'shd62ed92c, 32'shd62da8c4, 32'shd62c7863, 32'shd62b4809, 32'shd62a17b5, 
               32'shd628e767, 32'shd627b720, 32'shd62686e0, 32'shd62556a6, 32'shd6242672, 32'shd622f645, 32'shd621c61e, 32'shd62095fe, 
               32'shd61f65e4, 32'shd61e35d0, 32'shd61d05c3, 32'shd61bd5bd, 32'shd61aa5bd, 32'shd61975c3, 32'shd61845d0, 32'shd61715e3, 
               32'shd615e5fd, 32'shd614b61d, 32'shd6138644, 32'shd6125671, 32'shd61126a5, 32'shd60ff6df, 32'shd60ec720, 32'shd60d9767, 
               32'shd60c67b4, 32'shd60b3808, 32'shd60a0863, 32'shd608d8c4, 32'shd607a92b, 32'shd6067999, 32'shd6054a0d, 32'shd6041a88, 
               32'shd602eb0a, 32'shd601bb91, 32'shd6008c20, 32'shd5ff5cb4, 32'shd5fe2d50, 32'shd5fcfdf1, 32'shd5fbce9a, 32'shd5fa9f48, 
               32'shd5f96ffd, 32'shd5f840b9, 32'shd5f7117b, 32'shd5f5e244, 32'shd5f4b313, 32'shd5f383e8, 32'shd5f254c4, 32'shd5f125a7, 
               32'shd5eff690, 32'shd5eec77f, 32'shd5ed9875, 32'shd5ec6972, 32'shd5eb3a75, 32'shd5ea0b7e, 32'shd5e8dc8e, 32'shd5e7ada4, 
               32'shd5e67ec1, 32'shd5e54fe5, 32'shd5e4210f, 32'shd5e2f23f, 32'shd5e1c376, 32'shd5e094b3, 32'shd5df65f7, 32'shd5de3742, 
               32'shd5dd0892, 32'shd5dbd9ea, 32'shd5daab48, 32'shd5d97cac, 32'shd5d84e17, 32'shd5d71f88, 32'shd5d5f100, 32'shd5d4c27e, 
               32'shd5d39403, 32'shd5d2658f, 32'shd5d13721, 32'shd5d008b9, 32'shd5ceda58, 32'shd5cdabfd, 32'shd5cc7da9, 32'shd5cb4f5c, 
               32'shd5ca2115, 32'shd5c8f2d4, 32'shd5c7c49a, 32'shd5c69666, 32'shd5c56839, 32'shd5c43a13, 32'shd5c30bf3, 32'shd5c1ddd9, 
               32'shd5c0afc6, 32'shd5bf81ba, 32'shd5be53b4, 32'shd5bd25b4, 32'shd5bbf7bc, 32'shd5bac9c9, 32'shd5b99bdd, 32'shd5b86df8, 
               32'shd5b74019, 32'shd5b61241, 32'shd5b4e46f, 32'shd5b3b6a4, 32'shd5b288df, 32'shd5b15b21, 32'shd5b02d69, 32'shd5aeffb8, 
               32'shd5add20d, 32'shd5aca469, 32'shd5ab76cb, 32'shd5aa4934, 32'shd5a91ba4, 32'shd5a7ee1a, 32'shd5a6c096, 32'shd5a59319, 
               32'shd5a465a3, 32'shd5a33833, 32'shd5a20aca, 32'shd5a0dd67, 32'shd59fb00b, 32'shd59e82b5, 32'shd59d5566, 32'shd59c281d, 
               32'shd59afadb, 32'shd599cd9f, 32'shd598a06a, 32'shd597733c, 32'shd5964614, 32'shd59518f2, 32'shd593ebd7, 32'shd592bec3, 
               32'shd59191b5, 32'shd59064ae, 32'shd58f37ad, 32'shd58e0ab3, 32'shd58cddbf, 32'shd58bb0d2, 32'shd58a83eb, 32'shd589570b, 
               32'shd5882a32, 32'shd586fd5f, 32'shd585d093, 32'shd584a3cd, 32'shd583770e, 32'shd5824a55, 32'shd5811da3, 32'shd57ff0f7, 
               32'shd57ec452, 32'shd57d97b4, 32'shd57c6b1c, 32'shd57b3e8a, 32'shd57a1200, 32'shd578e57b, 32'shd577b8fe, 32'shd5768c86, 
               32'shd5756016, 32'shd57433ac, 32'shd5730748, 32'shd571daeb, 32'shd570ae95, 32'shd56f8245, 32'shd56e55fc, 32'shd56d29b9, 
               32'shd56bfd7d, 32'shd56ad148, 32'shd569a519, 32'shd56878f1, 32'shd5674ccf, 32'shd56620b3, 32'shd564f49f, 32'shd563c891, 
               32'shd5629c89, 32'shd5617088, 32'shd560448e, 32'shd55f189a, 32'shd55decad, 32'shd55cc0c6, 32'shd55b94e6, 32'shd55a690c, 
               32'shd5593d3a, 32'shd558116d, 32'shd556e5a7, 32'shd555b9e8, 32'shd5548e30, 32'shd553627d, 32'shd55236d2, 32'shd5510b2d, 
               32'shd54fdf8f, 32'shd54eb3f7, 32'shd54d8866, 32'shd54c5cdb, 32'shd54b3157, 32'shd54a05da, 32'shd548da63, 32'shd547aef3, 
               32'shd5468389, 32'shd5455826, 32'shd5442cca, 32'shd5430174, 32'shd541d625, 32'shd540aadc, 32'shd53f7f9a, 32'shd53e545f, 
               32'shd53d292a, 32'shd53bfdfb, 32'shd53ad2d4, 32'shd539a7b3, 32'shd5387c98, 32'shd5375184, 32'shd5362677, 32'shd534fb70, 
               32'shd533d070, 32'shd532a577, 32'shd5317a84, 32'shd5304f97, 32'shd52f24b2, 32'shd52df9d3, 32'shd52ccefa, 32'shd52ba428, 
               32'shd52a795d, 32'shd5294e98, 32'shd52823da, 32'shd526f923, 32'shd525ce72, 32'shd524a3c7, 32'shd5237924, 32'shd5224e87, 
               32'shd52123f0, 32'shd51ff960, 32'shd51eced7, 32'shd51da455, 32'shd51c79d9, 32'shd51b4f63, 32'shd51a24f5, 32'shd518fa8c, 
               32'shd517d02b, 32'shd516a5d0, 32'shd5157b7c, 32'shd514512e, 32'shd51326e7, 32'shd511fca7, 32'shd510d26d, 32'shd50fa83a, 
               32'shd50e7e0d, 32'shd50d53e7, 32'shd50c29c8, 32'shd50affaf, 32'shd509d59d, 32'shd508ab91, 32'shd507818d, 32'shd506578e, 
               32'shd5052d97, 32'shd50403a6, 32'shd502d9bc, 32'shd501afd8, 32'shd50085fb, 32'shd4ff5c24, 32'shd4fe3255, 32'shd4fd088c, 
               32'shd4fbdec9, 32'shd4fab50d, 32'shd4f98b58, 32'shd4f861a9, 32'shd4f73801, 32'shd4f60e60, 32'shd4f4e4c5, 32'shd4f3bb31, 
               32'shd4f291a4, 32'shd4f1681d, 32'shd4f03e9d, 32'shd4ef1523, 32'shd4edebb0, 32'shd4ecc244, 32'shd4eb98de, 32'shd4ea6f80, 
               32'shd4e94627, 32'shd4e81cd6, 32'shd4e6f38b, 32'shd4e5ca46, 32'shd4e4a108, 32'shd4e377d1, 32'shd4e24ea1, 32'shd4e12577, 
               32'shd4dffc54, 32'shd4ded338, 32'shd4ddaa22, 32'shd4dc8113, 32'shd4db580a, 32'shd4da2f08, 32'shd4d9060d, 32'shd4d7dd18, 
               32'shd4d6b42b, 32'shd4d58b43, 32'shd4d46263, 32'shd4d33989, 32'shd4d210b5, 32'shd4d0e7e9, 32'shd4cfbf23, 32'shd4ce9664, 
               32'shd4cd6dab, 32'shd4cc44f9, 32'shd4cb1c4e, 32'shd4c9f3a9, 32'shd4c8cb0b, 32'shd4c7a274, 32'shd4c679e3, 32'shd4c55159, 
               32'shd4c428d6, 32'shd4c30059, 32'shd4c1d7e3, 32'shd4c0af74, 32'shd4bf870b, 32'shd4be5ea9, 32'shd4bd364e, 32'shd4bc0df9, 
               32'shd4bae5ab, 32'shd4b9bd64, 32'shd4b89523, 32'shd4b76ce9, 32'shd4b644b6, 32'shd4b51c8a, 32'shd4b3f464, 32'shd4b2cc44, 
               32'shd4b1a42c, 32'shd4b07c1a, 32'shd4af540f, 32'shd4ae2c0a, 32'shd4ad040c, 32'shd4abdc15, 32'shd4aab425, 32'shd4a98c3b, 
               32'shd4a86458, 32'shd4a73c7b, 32'shd4a614a6, 32'shd4a4ecd7, 32'shd4a3c50e, 32'shd4a29d4c, 32'shd4a17591, 32'shd4a04ddd, 
               32'shd49f2630, 32'shd49dfe89, 32'shd49cd6e8, 32'shd49baf4f, 32'shd49a87bc, 32'shd4996030, 32'shd49838aa, 32'shd497112b, 
               32'shd495e9b3, 32'shd494c242, 32'shd4939ad7, 32'shd4927373, 32'shd4914c16, 32'shd49024bf, 32'shd48efd6f, 32'shd48dd626, 
               32'shd48caee4, 32'shd48b87a8, 32'shd48a6073, 32'shd4893944, 32'shd488121d, 32'shd486eafc, 32'shd485c3e1, 32'shd4849cce, 
               32'shd48375c1, 32'shd4824ebb, 32'shd48127bb, 32'shd48000c2, 32'shd47ed9d0, 32'shd47db2e5, 32'shd47c8c00, 32'shd47b6523, 
               32'shd47a3e4b, 32'shd479177b, 32'shd477f0b1, 32'shd476c9ee, 32'shd475a332, 32'shd4747c7c, 32'shd47355cd, 32'shd4722f25, 
               32'shd4710883, 32'shd46fe1e8, 32'shd46ebb54, 32'shd46d94c7, 32'shd46c6e40, 32'shd46b47c0, 32'shd46a2147, 32'shd468fad5, 
               32'shd467d469, 32'shd466ae04, 32'shd46587a6, 32'shd464614e, 32'shd4633afd, 32'shd46214b3, 32'shd460ee70, 32'shd45fc833, 
               32'shd45ea1fd, 32'shd45d7bce, 32'shd45c55a5, 32'shd45b2f84, 32'shd45a0969, 32'shd458e354, 32'shd457bd47, 32'shd4569740, 
               32'shd4557140, 32'shd4544b46, 32'shd4532554, 32'shd451ff68, 32'shd450d983, 32'shd44fb3a4, 32'shd44e8dcd, 32'shd44d67fc, 
               32'shd44c4232, 32'shd44b1c6e, 32'shd449f6b1, 32'shd448d0fb, 32'shd447ab4c, 32'shd44685a4, 32'shd4456002, 32'shd4443a67, 
               32'shd44314d3, 32'shd441ef45, 32'shd440c9be, 32'shd43fa43e, 32'shd43e7ec5, 32'shd43d5952, 32'shd43c33e7, 32'shd43b0e81, 
               32'shd439e923, 32'shd438c3cc, 32'shd4379e7b, 32'shd4367931, 32'shd43553ee, 32'shd4342eb1, 32'shd433097b, 32'shd431e44c, 
               32'shd430bf24, 32'shd42f9a02, 32'shd42e74e8, 32'shd42d4fd4, 32'shd42c2ac6, 32'shd42b05c0, 32'shd429e0c0, 32'shd428bbc7, 
               32'shd42796d5, 32'shd42671ea, 32'shd4254d05, 32'shd4242827, 32'shd4230350, 32'shd421de7f, 32'shd420b9b6, 32'shd41f94f3, 
               32'shd41e7037, 32'shd41d4b81, 32'shd41c26d3, 32'shd41b022b, 32'shd419dd8a, 32'shd418b8f0, 32'shd417945c, 32'shd4166fd0, 
               32'shd4154b4a, 32'shd41426cb, 32'shd4130252, 32'shd411dde1, 32'shd410b976, 32'shd40f9512, 32'shd40e70b4, 32'shd40d4c5e, 
               32'shd40c280e, 32'shd40b03c5, 32'shd409df83, 32'shd408bb48, 32'shd4079713, 32'shd40672e5, 32'shd4054ebe, 32'shd4042a9e, 
               32'shd4030684, 32'shd401e271, 32'shd400be66, 32'shd3ff9a60, 32'shd3fe7662, 32'shd3fd526a, 32'shd3fc2e7a, 32'shd3fb0a90, 
               32'shd3f9e6ad, 32'shd3f8c2d0, 32'shd3f79efa, 32'shd3f67b2c, 32'shd3f55764, 32'shd3f433a2, 32'shd3f30fe8, 32'shd3f1ec34, 
               32'shd3f0c887, 32'shd3efa4e1, 32'shd3ee8142, 32'shd3ed5da9, 32'shd3ec3a18, 32'shd3eb168d, 32'shd3e9f309, 32'shd3e8cf8b, 
               32'shd3e7ac15, 32'shd3e688a5, 32'shd3e5653c, 32'shd3e441da, 32'shd3e31e7f, 32'shd3e1fb2a, 32'shd3e0d7dd, 32'shd3dfb496, 
               32'shd3de9156, 32'shd3dd6e1c, 32'shd3dc4aea, 32'shd3db27be, 32'shd3da049a, 32'shd3d8e17b, 32'shd3d7be64, 32'shd3d69b54, 
               32'shd3d5784a, 32'shd3d45547, 32'shd3d3324b, 32'shd3d20f56, 32'shd3d0ec68, 32'shd3cfc980, 32'shd3cea69f, 32'shd3cd83c6, 
               32'shd3cc60f2, 32'shd3cb3e26, 32'shd3ca1b61, 32'shd3c8f8a2, 32'shd3c7d5ea, 32'shd3c6b339, 32'shd3c5908f, 32'shd3c46dec, 
               32'shd3c34b4f, 32'shd3c228b9, 32'shd3c1062a, 32'shd3bfe3a2, 32'shd3bec121, 32'shd3bd9ea7, 32'shd3bc7c33, 32'shd3bb59c6, 
               32'shd3ba3760, 32'shd3b91501, 32'shd3b7f2a9, 32'shd3b6d057, 32'shd3b5ae0d, 32'shd3b48bc9, 32'shd3b3698c, 32'shd3b24756, 
               32'shd3b12526, 32'shd3b002fe, 32'shd3aee0dc, 32'shd3adbec1, 32'shd3ac9cad, 32'shd3ab7aa0, 32'shd3aa589a, 32'shd3a9369a, 
               32'shd3a814a2, 32'shd3a6f2b0, 32'shd3a5d0c5, 32'shd3a4aee1, 32'shd3a38d03, 32'shd3a26b2d, 32'shd3a1495d, 32'shd3a02795, 
               32'shd39f05d3, 32'shd39de418, 32'shd39cc263, 32'shd39ba0b6, 32'shd39a7f0f, 32'shd3995d70, 32'shd3983bd7, 32'shd3971a45, 
               32'shd395f8ba, 32'shd394d735, 32'shd393b5b8, 32'shd3929441, 32'shd39172d2, 32'shd3905169, 32'shd38f3007, 32'shd38e0eac, 
               32'shd38ced57, 32'shd38bcc0a, 32'shd38aaac3, 32'shd3898983, 32'shd388684a, 32'shd3874718, 32'shd38625ed, 32'shd38504c9, 
               32'shd383e3ab, 32'shd382c295, 32'shd381a185, 32'shd380807c, 32'shd37f5f7a, 32'shd37e3e7f, 32'shd37d1d8a, 32'shd37bfc9d, 
               32'shd37adbb6, 32'shd379bad7, 32'shd37899fe, 32'shd377792c, 32'shd3765861, 32'shd375379d, 32'shd37416df, 32'shd372f629, 
               32'shd371d579, 32'shd370b4d0, 32'shd36f942e, 32'shd36e7393, 32'shd36d52ff, 32'shd36c3272, 32'shd36b11eb, 32'shd369f16c, 
               32'shd368d0f3, 32'shd367b082, 32'shd3669017, 32'shd3656fb3, 32'shd3644f55, 32'shd3632eff, 32'shd3620eb0, 32'shd360ee67, 
               32'shd35fce26, 32'shd35eadeb, 32'shd35d8db7, 32'shd35c6d8a, 32'shd35b4d64, 32'shd35a2d45, 32'shd3590d2c, 32'shd357ed1b, 
               32'shd356cd11, 32'shd355ad0d, 32'shd3548d10, 32'shd3536d1a, 32'shd3524d2b, 32'shd3512d43, 32'shd3500d62, 32'shd34eed88, 
               32'shd34dcdb4, 32'shd34cade8, 32'shd34b8e22, 32'shd34a6e63, 32'shd3494eab, 32'shd3482efa, 32'shd3470f50, 32'shd345efad, 
               32'shd344d011, 32'shd343b07b, 32'shd34290ed, 32'shd3417165, 32'shd34051e5, 32'shd33f326b, 32'shd33e12f8, 32'shd33cf38c, 
               32'shd33bd427, 32'shd33ab4c9, 32'shd3399572, 32'shd3387621, 32'shd33756d8, 32'shd3363795, 32'shd335185a, 32'shd333f925, 
               32'shd332d9f7, 32'shd331bad0, 32'shd3309bb0, 32'shd32f7c97, 32'shd32e5d85, 32'shd32d3e7a, 32'shd32c1f75, 32'shd32b0078, 
               32'shd329e181, 32'shd328c292, 32'shd327a3a9, 32'shd32684c7, 32'shd32565ec, 32'shd3244718, 32'shd323284b, 32'shd3220985, 
               32'shd320eac6, 32'shd31fcc0e, 32'shd31ead5c, 32'shd31d8eb2, 32'shd31c700f, 32'shd31b5172, 32'shd31a32dc, 32'shd319144e, 
               32'shd317f5c6, 32'shd316d745, 32'shd315b8cb, 32'shd3149a58, 32'shd3137bec, 32'shd3125d86, 32'shd3113f28, 32'shd31020d1, 
               32'shd30f0280, 32'shd30de437, 32'shd30cc5f4, 32'shd30ba7b9, 32'shd30a8984, 32'shd3096b56, 32'shd3084d30, 32'shd3072f10, 
               32'shd30610f7, 32'shd304f2e5, 32'shd303d4da, 32'shd302b6d6, 32'shd30198d8, 32'shd3007ae2, 32'shd2ff5cf3, 32'shd2fe3f0b, 
               32'shd2fd2129, 32'shd2fc034f, 32'shd2fae57b, 32'shd2f9c7ae, 32'shd2f8a9e9, 32'shd2f78c2a, 32'shd2f66e72, 32'shd2f550c2, 
               32'shd2f43318, 32'shd2f31575, 32'shd2f1f7d9, 32'shd2f0da44, 32'shd2efbcb6, 32'shd2ee9f2e, 32'shd2ed81ae, 32'shd2ec6435, 
               32'shd2eb46c3, 32'shd2ea2957, 32'shd2e90bf3, 32'shd2e7ee96, 32'shd2e6d13f, 32'shd2e5b3f0, 32'shd2e496a7, 32'shd2e37965, 
               32'shd2e25c2b, 32'shd2e13ef7, 32'shd2e021ca, 32'shd2df04a5, 32'shd2dde786, 32'shd2dcca6e, 32'shd2dbad5d, 32'shd2da9053, 
               32'shd2d97350, 32'shd2d85654, 32'shd2d7395f, 32'shd2d61c71, 32'shd2d4ff8a, 32'shd2d3e2aa, 32'shd2d2c5d0, 32'shd2d1a8fe, 
               32'shd2d08c33, 32'shd2cf6f6f, 32'shd2ce52b1, 32'shd2cd35fb, 32'shd2cc194c, 32'shd2cafca3, 32'shd2c9e002, 32'shd2c8c367, 
               32'shd2c7a6d4, 32'shd2c68a47, 32'shd2c56dc2, 32'shd2c45143, 32'shd2c334cc, 32'shd2c2185b, 32'shd2c0fbf1, 32'shd2bfdf8f, 
               32'shd2bec333, 32'shd2bda6de, 32'shd2bc8a91, 32'shd2bb6e4a, 32'shd2ba520a, 32'shd2b935d1, 32'shd2b8199f, 32'shd2b6fd75, 
               32'shd2b5e151, 32'shd2b4c534, 32'shd2b3a91e, 32'shd2b28d0f, 32'shd2b17107, 32'shd2b05506, 32'shd2af390d, 32'shd2ae1d1a, 
               32'shd2ad012e, 32'shd2abe549, 32'shd2aac96b, 32'shd2a9ad94, 32'shd2a891c4, 32'shd2a775fb, 32'shd2a65a39, 32'shd2a53e7e, 
               32'shd2a422ca, 32'shd2a3071d, 32'shd2a1eb77, 32'shd2a0cfd8, 32'shd29fb440, 32'shd29e98af, 32'shd29d7d25, 32'shd29c61a2, 
               32'shd29b4626, 32'shd29a2ab1, 32'shd2990f43, 32'shd297f3dc, 32'shd296d87c, 32'shd295bd23, 32'shd294a1d0, 32'shd2938685, 
               32'shd2926b41, 32'shd2915004, 32'shd29034ce, 32'shd28f199f, 32'shd28dfe77, 32'shd28ce357, 32'shd28bc83d, 32'shd28aad2a, 
               32'shd289921e, 32'shd2887719, 32'shd2875c1b, 32'shd2864124, 32'shd2852634, 32'shd2840b4b, 32'shd282f069, 32'shd281d58e, 
               32'shd280babb, 32'shd27f9fee, 32'shd27e8528, 32'shd27d6a69, 32'shd27c4fb1, 32'shd27b3501, 32'shd27a1a57, 32'shd278ffb4, 
               32'shd277e518, 32'shd276ca84, 32'shd275aff6, 32'shd2749570, 32'shd2737af0, 32'shd2726077, 32'shd2714606, 32'shd2702b9b, 
               32'shd26f1138, 32'shd26df6db, 32'shd26cdc86, 32'shd26bc237, 32'shd26aa7f0, 32'shd2698db0, 32'shd2687376, 32'shd2675944, 
               32'shd2663f19, 32'shd26524f5, 32'shd2640ad7, 32'shd262f0c1, 32'shd261d6b2, 32'shd260bcaa, 32'shd25fa2a9, 32'shd25e88af, 
               32'shd25d6ebc, 32'shd25c54d0, 32'shd25b3aeb, 32'shd25a210d, 32'shd2590736, 32'shd257ed67, 32'shd256d39e, 32'shd255b9dc, 
               32'shd254a021, 32'shd253866e, 32'shd2526cc1, 32'shd251531c, 32'shd250397d, 32'shd24f1fe6, 32'shd24e0655, 32'shd24ceccc, 
               32'shd24bd34a, 32'shd24ab9ce, 32'shd249a05a, 32'shd24886ed, 32'shd2476d87, 32'shd2465428, 32'shd2453ad0, 32'shd244217f, 
               32'shd2430835, 32'shd241eef2, 32'shd240d5b6, 32'shd23fbc82, 32'shd23ea354, 32'shd23d8a2d, 32'shd23c710e, 32'shd23b57f5, 
               32'shd23a3ee4, 32'shd23925d9, 32'shd2380cd6, 32'shd236f3da, 32'shd235dae4, 32'shd234c1f6, 32'shd233a90f, 32'shd232902f, 
               32'shd2317756, 32'shd2305e84, 32'shd22f45b9, 32'shd22e2cf6, 32'shd22d1439, 32'shd22bfb83, 32'shd22ae2d5, 32'shd229ca2d, 
               32'shd228b18d, 32'shd22798f3, 32'shd2268061, 32'shd22567d6, 32'shd2244f52, 32'shd22336d5, 32'shd2221e5f, 32'shd22105f0, 
               32'shd21fed88, 32'shd21ed527, 32'shd21dbccd, 32'shd21ca47b, 32'shd21b8c2f, 32'shd21a73eb, 32'shd2195bad, 32'shd2184377, 
               32'shd2172b48, 32'shd216131f, 32'shd214fafe, 32'shd213e2e4, 32'shd212cad1, 32'shd211b2c5, 32'shd2109ac1, 32'shd20f82c3, 
               32'shd20e6acc, 32'shd20d52dd, 32'shd20c3af4, 32'shd20b2313, 32'shd20a0b39, 32'shd208f366, 32'shd207db9a, 32'shd206c3d5, 
               32'shd205ac17, 32'shd2049460, 32'shd2037cb0, 32'shd2026508, 32'shd2014d66, 32'shd20035cc, 32'shd1ff1e38, 32'shd1fe06ac, 
               32'shd1fcef27, 32'shd1fbd7a9, 32'shd1fac032, 32'shd1f9a8c2, 32'shd1f89159, 32'shd1f779f8, 32'shd1f6629d, 32'shd1f54b49, 
               32'shd1f433fd, 32'shd1f31cb8, 32'shd1f2057a, 32'shd1f0ee43, 32'shd1efd713, 32'shd1eebfea, 32'shd1eda8c8, 32'shd1ec91ad, 
               32'shd1eb7a9a, 32'shd1ea638d, 32'shd1e94c88, 32'shd1e8358a, 32'shd1e71e93, 32'shd1e607a3, 32'shd1e4f0ba, 32'shd1e3d9d8, 
               32'shd1e2c2fd, 32'shd1e1ac2a, 32'shd1e0955d, 32'shd1df7e98, 32'shd1de67da, 32'shd1dd5123, 32'shd1dc3a73, 32'shd1db23ca, 
               32'shd1da0d28, 32'shd1d8f68d, 32'shd1d7dffa, 32'shd1d6c96d, 32'shd1d5b2e8, 32'shd1d49c6a, 32'shd1d385f3, 32'shd1d26f83, 
               32'shd1d1591a, 32'shd1d042b8, 32'shd1cf2c5e, 32'shd1ce160a, 32'shd1ccffbe, 32'shd1cbe979, 32'shd1cad33b, 32'shd1c9bd04, 
               32'shd1c8a6d4, 32'shd1c790ab, 32'shd1c67a8a, 32'shd1c5646f, 32'shd1c44e5c, 32'shd1c33850, 32'shd1c2224b, 32'shd1c10c4d, 
               32'shd1bff656, 32'shd1bee066, 32'shd1bdca7e, 32'shd1bcb49c, 32'shd1bb9ec2, 32'shd1ba88ef, 32'shd1b97323, 32'shd1b85d5e, 
               32'shd1b747a0, 32'shd1b631ea, 32'shd1b51c3a, 32'shd1b40692, 32'shd1b2f0f1, 32'shd1b1db57, 32'shd1b0c5c4, 32'shd1afb038, 
               32'shd1ae9ab4, 32'shd1ad8536, 32'shd1ac6fc0, 32'shd1ab5a51, 32'shd1aa44e9, 32'shd1a92f88, 32'shd1a81a2e, 32'shd1a704dc, 
               32'shd1a5ef90, 32'shd1a4da4c, 32'shd1a3c50f, 32'shd1a2afd9, 32'shd1a19aaa, 32'shd1a08582, 32'shd19f7062, 32'shd19e5b48, 
               32'shd19d4636, 32'shd19c312b, 32'shd19b1c27, 32'shd19a072a, 32'shd198f235, 32'shd197dd46, 32'shd196c85f, 32'shd195b37f, 
               32'shd1949ea6, 32'shd19389d4, 32'shd1927509, 32'shd1916046, 32'shd1904b89, 32'shd18f36d4, 32'shd18e2226, 32'shd18d0d7f, 
               32'shd18bf8e0, 32'shd18ae447, 32'shd189cfb6, 32'shd188bb2b, 32'shd187a6a8, 32'shd186922d, 32'shd1857db8, 32'shd184694a, 
               32'shd18354e4, 32'shd1824085, 32'shd1812c2d, 32'shd18017dc, 32'shd17f0392, 32'shd17def50, 32'shd17cdb14, 32'shd17bc6e0, 
               32'shd17ab2b3, 32'shd1799e8d, 32'shd1788a6f, 32'shd1777657, 32'shd1766247, 32'shd1754e3e, 32'shd1743a3c, 32'shd1732641, 
               32'shd172124d, 32'shd170fe61, 32'shd16fea7c, 32'shd16ed69e, 32'shd16dc2c7, 32'shd16caef7, 32'shd16b9b2f, 32'shd16a876d, 
               32'shd16973b3, 32'shd1686000, 32'shd1674c54, 32'shd16638b0, 32'shd1652512, 32'shd164117c, 32'shd162fded, 32'shd161ea65, 
               32'shd160d6e5, 32'shd15fc36b, 32'shd15eaff9, 32'shd15d9c8e, 32'shd15c892a, 32'shd15b75cd, 32'shd15a6278, 32'shd1594f29, 
               32'shd1583be2, 32'shd15728a2, 32'shd156156a, 32'shd1550238, 32'shd153ef0e, 32'shd152dbeb, 32'shd151c8cf, 32'shd150b5ba, 
               32'shd14fa2ad, 32'shd14e8fa6, 32'shd14d7ca7, 32'shd14c69af, 32'shd14b56be, 32'shd14a43d5, 32'shd14930f3, 32'shd1481e17, 
               32'shd1470b44, 32'shd145f877, 32'shd144e5b1, 32'shd143d2f3, 32'shd142c03c, 32'shd141ad8c, 32'shd1409ae3, 32'shd13f8842, 
               32'shd13e75a8, 32'shd13d6315, 32'shd13c5089, 32'shd13b3e04, 32'shd13a2b87, 32'shd1391911, 32'shd13806a2, 32'shd136f43a, 
               32'shd135e1d9, 32'shd134cf80, 32'shd133bd2e, 32'shd132aae3, 32'shd131989f, 32'shd1308663, 32'shd12f742d, 32'shd12e61ff, 
               32'shd12d4fd9, 32'shd12c3db9, 32'shd12b2ba1, 32'shd12a198f, 32'shd1290786, 32'shd127f583, 32'shd126e387, 32'shd125d193, 
               32'shd124bfa6, 32'shd123adc0, 32'shd1229be2, 32'shd1218a0a, 32'shd120783a, 32'shd11f6671, 32'shd11e54b0, 32'shd11d42f5, 
               32'shd11c3142, 32'shd11b1f96, 32'shd11a0df1, 32'shd118fc54, 32'shd117eabd, 32'shd116d92e, 32'shd115c7a7, 32'shd114b626, 
               32'shd113a4ad, 32'shd112933b, 32'shd11181d0, 32'shd110706c, 32'shd10f5f10, 32'shd10e4dbb, 32'shd10d3c6d, 32'shd10c2b26, 
               32'shd10b19e7, 32'shd10a08ae, 32'shd108f77d, 32'shd107e654, 32'shd106d531, 32'shd105c416, 32'shd104b302, 32'shd103a1f5, 
               32'shd10290f0, 32'shd1017ff2, 32'shd1006efb, 32'shd0ff5e0b, 32'shd0fe4d22, 32'shd0fd3c41, 32'shd0fc2b67, 32'shd0fb1a94, 
               32'shd0fa09c9, 32'shd0f8f905, 32'shd0f7e848, 32'shd0f6d792, 32'shd0f5c6e3, 32'shd0f4b63c, 32'shd0f3a59c, 32'shd0f29503, 
               32'shd0f18472, 32'shd0f073e8, 32'shd0ef6365, 32'shd0ee52e9, 32'shd0ed4275, 32'shd0ec3208, 32'shd0eb21a2, 32'shd0ea1143, 
               32'shd0e900ec, 32'shd0e7f09b, 32'shd0e6e053, 32'shd0e5d011, 32'shd0e4bfd7, 32'shd0e3afa4, 32'shd0e29f78, 32'shd0e18f53, 
               32'shd0e07f36, 32'shd0df6f20, 32'shd0de5f11, 32'shd0dd4f0a, 32'shd0dc3f0a, 32'shd0db2f11, 32'shd0da1f1f, 32'shd0d90f35, 
               32'shd0d7ff51, 32'shd0d6ef76, 32'shd0d5dfa1, 32'shd0d4cfd4, 32'shd0d3c00e, 32'shd0d2b04f, 32'shd0d1a097, 32'shd0d090e7, 
               32'shd0cf813e, 32'shd0ce719d, 32'shd0cd6202, 32'shd0cc526f, 32'shd0cb42e3, 32'shd0ca335f, 32'shd0c923e1, 32'shd0c8146c, 
               32'shd0c704fd, 32'shd0c5f595, 32'shd0c4e635, 32'shd0c3d6dc, 32'shd0c2c78b, 32'shd0c1b841, 32'shd0c0a8fe, 32'shd0bf99c2, 
               32'shd0be8a8d, 32'shd0bd7b60, 32'shd0bc6c3a, 32'shd0bb5d1c, 32'shd0ba4e05, 32'shd0b93ef5, 32'shd0b82fec, 32'shd0b720eb, 
               32'shd0b611f1, 32'shd0b502fe, 32'shd0b3f412, 32'shd0b2e52e, 32'shd0b1d651, 32'shd0b0c77b, 32'shd0afb8ad, 32'shd0aea9e6, 
               32'shd0ad9b26, 32'shd0ac8c6e, 32'shd0ab7dbd, 32'shd0aa6f13, 32'shd0a96070, 32'shd0a851d5, 32'shd0a74341, 32'shd0a634b4, 
               32'shd0a5262f, 32'shd0a417b1, 32'shd0a3093a, 32'shd0a1facb, 32'shd0a0ec63, 32'shd09fde02, 32'shd09ecfa8, 32'shd09dc156, 
               32'shd09cb30b, 32'shd09ba4c8, 32'shd09a968b, 32'shd0998856, 32'shd0987a29, 32'shd0976c02, 32'shd0965de3, 32'shd0954fcc, 
               32'shd09441bb, 32'shd09333b2, 32'shd09225b0, 32'shd09117b6, 32'shd09009c3, 32'shd08efbd7, 32'shd08dedf2, 32'shd08ce015, 
               32'shd08bd23f, 32'shd08ac470, 32'shd089b6a9, 32'shd088a8e9, 32'shd0879b31, 32'shd0868d7f, 32'shd0857fd5, 32'shd0847233, 
               32'shd0836497, 32'shd0825703, 32'shd0814977, 32'shd0803bf1, 32'shd07f2e73, 32'shd07e20fc, 32'shd07d138d, 32'shd07c0625, 
               32'shd07af8c4, 32'shd079eb6b, 32'shd078de19, 32'shd077d0ce, 32'shd076c38b, 32'shd075b64f, 32'shd074a91a, 32'shd0739bec, 
               32'shd0728ec6, 32'shd07181a7, 32'shd0707490, 32'shd06f6780, 32'shd06e5a77, 32'shd06d4d76, 32'shd06c407c, 32'shd06b3389, 
               32'shd06a269d, 32'shd06919b9, 32'shd0680cdd, 32'shd0670007, 32'shd065f339, 32'shd064e673, 32'shd063d9b3, 32'shd062ccfb, 
               32'shd061c04a, 32'shd060b3a1, 32'shd05fa6ff, 32'shd05e9a64, 32'shd05d8dd1, 32'shd05c8145, 32'shd05b74c0, 32'shd05a6843, 
               32'shd0595bcd, 32'shd0584f5f, 32'shd05742f7, 32'shd0563698, 32'shd0552a3f, 32'shd0541dee, 32'shd05311a4, 32'shd0520562, 
               32'shd050f926, 32'shd04fecf3, 32'shd04ee0c6, 32'shd04dd4a1, 32'shd04cc884, 32'shd04bbc6d, 32'shd04ab05e, 32'shd049a457, 
               32'shd0489856, 32'shd0478c5d, 32'shd046806c, 32'shd0457482, 32'shd044689f, 32'shd0435cc3, 32'shd04250ef, 32'shd0414522, 
               32'shd040395d, 32'shd03f2d9f, 32'shd03e21e8, 32'shd03d1639, 32'shd03c0a91, 32'shd03afef1, 32'shd039f357, 32'shd038e7c5, 
               32'shd037dc3b, 32'shd036d0b8, 32'shd035c53c, 32'shd034b9c8, 32'shd033ae5b, 32'shd032a2f5, 32'shd0319797, 32'shd0308c40, 
               32'shd02f80f1, 32'shd02e75a8, 32'shd02d6a68, 32'shd02c5f2e, 32'shd02b53fc, 32'shd02a48d2, 32'shd0293dae, 32'shd0283293, 
               32'shd027277e, 32'shd0261c71, 32'shd025116b, 32'shd024066d, 32'shd022fb76, 32'shd021f086, 32'shd020e59e, 32'shd01fdabd, 
               32'shd01ecfe4, 32'shd01dc512, 32'shd01cba47, 32'shd01baf84, 32'shd01aa4c8, 32'shd0199a13, 32'shd0188f66, 32'shd01784c1, 
               32'shd0167a22, 32'shd0156f8b, 32'shd01464fc, 32'shd0135a73, 32'shd0124ff3, 32'shd0114579, 32'shd0103b07, 32'shd00f309d, 
               32'shd00e2639, 32'shd00d1bdd, 32'shd00c1189, 32'shd00b073c, 32'shd009fcf6, 32'shd008f2b8, 32'shd007e881, 32'shd006de52, 
               32'shd005d42a, 32'shd004ca09, 32'shd003bff0, 32'shd002b5de, 32'shd001abd3, 32'shd000a1d0, 32'shcfff97d5, 32'shcffe8de0, 
               32'shcffd83f4, 32'shcffc7a0e, 32'shcffb7030, 32'shcffa6659, 32'shcff95c8a, 32'shcff852c2, 32'shcff74902, 32'shcff63f49, 
               32'shcff53597, 32'shcff42bed, 32'shcff3224a, 32'shcff218af, 32'shcff10f1b, 32'shcff0058e, 32'shcfeefc09, 32'shcfedf28b, 
               32'shcfece915, 32'shcfebdfa6, 32'shcfead63f, 32'shcfe9ccdf, 32'shcfe8c386, 32'shcfe7ba35, 32'shcfe6b0eb, 32'shcfe5a7a8, 
               32'shcfe49e6d, 32'shcfe3953a, 32'shcfe28c0e, 32'shcfe182e9, 32'shcfe079cc, 32'shcfdf70b6, 32'shcfde67a7, 32'shcfdd5ea0, 
               32'shcfdc55a1, 32'shcfdb4ca8, 32'shcfda43b8, 32'shcfd93ace, 32'shcfd831ec, 32'shcfd72912, 32'shcfd6203f, 32'shcfd51773, 
               32'shcfd40eaf, 32'shcfd305f2, 32'shcfd1fd3d, 32'shcfd0f48f, 32'shcfcfebe8, 32'shcfcee349, 32'shcfcddab2, 32'shcfccd221, 
               32'shcfcbc999, 32'shcfcac117, 32'shcfc9b89d, 32'shcfc8b02b, 32'shcfc7a7c0, 32'shcfc69f5c, 32'shcfc59700, 32'shcfc48eab, 
               32'shcfc3865e, 32'shcfc27e18, 32'shcfc175da, 32'shcfc06da3, 32'shcfbf6573, 32'shcfbe5d4b, 32'shcfbd552b, 32'shcfbc4d11, 
               32'shcfbb4500, 32'shcfba3cf5, 32'shcfb934f2, 32'shcfb82cf7, 32'shcfb72503, 32'shcfb61d16, 32'shcfb51531, 32'shcfb40d54, 
               32'shcfb3057d, 32'shcfb1fdaf, 32'shcfb0f5e7, 32'shcfafee28, 32'shcfaee66f, 32'shcfaddebe, 32'shcfacd715, 32'shcfabcf73, 
               32'shcfaac7d8, 32'shcfa9c045, 32'shcfa8b8b9, 32'shcfa7b135, 32'shcfa6a9b8, 32'shcfa5a243, 32'shcfa49ad5, 32'shcfa3936f, 
               32'shcfa28c10, 32'shcfa184b8, 32'shcfa07d68, 32'shcf9f7620, 32'shcf9e6edf, 32'shcf9d67a5, 32'shcf9c6073, 32'shcf9b5948, 
               32'shcf9a5225, 32'shcf994b09, 32'shcf9843f5, 32'shcf973ce8, 32'shcf9635e2, 32'shcf952ee4, 32'shcf9427ee, 32'shcf9320ff, 
               32'shcf921a17, 32'shcf911337, 32'shcf900c5f, 32'shcf8f058e, 32'shcf8dfec4, 32'shcf8cf802, 32'shcf8bf147, 32'shcf8aea94, 
               32'shcf89e3e8, 32'shcf88dd44, 32'shcf87d6a7, 32'shcf86d012, 32'shcf85c984, 32'shcf84c2fd, 32'shcf83bc7e, 32'shcf82b607, 
               32'shcf81af97, 32'shcf80a92e, 32'shcf7fa2cd, 32'shcf7e9c74, 32'shcf7d9622, 32'shcf7c8fd7, 32'shcf7b8994, 32'shcf7a8359, 
               32'shcf797d24, 32'shcf7876f8, 32'shcf7770d3, 32'shcf766ab5, 32'shcf75649f, 32'shcf745e90, 32'shcf735889, 32'shcf725289, 
               32'shcf714c91, 32'shcf7046a0, 32'shcf6f40b7, 32'shcf6e3ad5, 32'shcf6d34fb, 32'shcf6c2f28, 32'shcf6b295d, 32'shcf6a2399, 
               32'shcf691ddd, 32'shcf681828, 32'shcf67127a, 32'shcf660cd5, 32'shcf650736, 32'shcf64019f, 32'shcf62fc10, 32'shcf61f688, 
               32'shcf60f108, 32'shcf5feb8f, 32'shcf5ee61e, 32'shcf5de0b4, 32'shcf5cdb51, 32'shcf5bd5f7, 32'shcf5ad0a3, 32'shcf59cb57, 
               32'shcf58c613, 32'shcf57c0d6, 32'shcf56bba1, 32'shcf55b673, 32'shcf54b14d, 32'shcf53ac2e, 32'shcf52a716, 32'shcf51a207, 
               32'shcf509cfe, 32'shcf4f97fe, 32'shcf4e9304, 32'shcf4d8e12, 32'shcf4c8928, 32'shcf4b8445, 32'shcf4a7f6a, 32'shcf497a96, 
               32'shcf4875ca, 32'shcf477105, 32'shcf466c48, 32'shcf456793, 32'shcf4462e4, 32'shcf435e3e, 32'shcf42599f, 32'shcf415507, 
               32'shcf405077, 32'shcf3f4bee, 32'shcf3e476d, 32'shcf3d42f4, 32'shcf3c3e82, 32'shcf3b3a17, 32'shcf3a35b4, 32'shcf393159, 
               32'shcf382d05, 32'shcf3728b8, 32'shcf362473, 32'shcf352036, 32'shcf341c00, 32'shcf3317d2, 32'shcf3213ab, 32'shcf310f8c, 
               32'shcf300b74, 32'shcf2f0764, 32'shcf2e035b, 32'shcf2cff5a, 32'shcf2bfb60, 32'shcf2af76e, 32'shcf29f383, 32'shcf28efa0, 
               32'shcf27ebc5, 32'shcf26e7f1, 32'shcf25e424, 32'shcf24e05f, 32'shcf23dca2, 32'shcf22d8ec, 32'shcf21d53e, 32'shcf20d197, 
               32'shcf1fcdf8, 32'shcf1eca60, 32'shcf1dc6d0, 32'shcf1cc347, 32'shcf1bbfc6, 32'shcf1abc4d, 32'shcf19b8db, 32'shcf18b570, 
               32'shcf17b20d, 32'shcf16aeb2, 32'shcf15ab5e, 32'shcf14a812, 32'shcf13a4cd, 32'shcf12a190, 32'shcf119e5a, 32'shcf109b2c, 
               32'shcf0f9805, 32'shcf0e94e6, 32'shcf0d91cf, 32'shcf0c8ebf, 32'shcf0b8bb7, 32'shcf0a88b6, 32'shcf0985bc, 32'shcf0882cb, 
               32'shcf077fe1, 32'shcf067cfe, 32'shcf057a23, 32'shcf04774f, 32'shcf037483, 32'shcf0271bf, 32'shcf016f02, 32'shcf006c4d, 
               32'shceff699f, 32'shcefe66f9, 32'shcefd645a, 32'shcefc61c3, 32'shcefb5f34, 32'shcefa5cac, 32'shcef95a2b, 32'shcef857b2, 
               32'shcef75541, 32'shcef652d7, 32'shcef55075, 32'shcef44e1b, 32'shcef34bc8, 32'shcef2497c, 32'shcef14738, 32'shcef044fc, 
               32'shceef42c7, 32'shceee409a, 32'shceed3e74, 32'shceec3c56, 32'shceeb3a40, 32'shceea3831, 32'shcee93629, 32'shcee8342a, 
               32'shcee73231, 32'shcee63041, 32'shcee52e58, 32'shcee42c76, 32'shcee32a9c, 32'shcee228ca, 32'shcee126ff, 32'shcee0253c, 
               32'shcedf2380, 32'shcede21cc, 32'shcedd2020, 32'shcedc1e7b, 32'shcedb1cde, 32'shceda1b48, 32'shced919ba, 32'shced81833, 
               32'shced716b4, 32'shced6153d, 32'shced513cd, 32'shced41265, 32'shced31104, 32'shced20fab, 32'shced10e59, 32'shced00d0f, 
               32'shcecf0bcd, 32'shcece0a92, 32'shcecd095f, 32'shcecc0833, 32'shcecb070f, 32'shceca05f3, 32'shcec904de, 32'shcec803d1, 
               32'shcec702cb, 32'shcec601cd, 32'shcec500d7, 32'shcec3ffe8, 32'shcec2ff01, 32'shcec1fe21, 32'shcec0fd49, 32'shcebffc79, 
               32'shcebefbb0, 32'shcebdfaee, 32'shcebcfa35, 32'shcebbf983, 32'shcebaf8d8, 32'shceb9f835, 32'shceb8f79a, 32'shceb7f706, 
               32'shceb6f67a, 32'shceb5f5f5, 32'shceb4f579, 32'shceb3f503, 32'shceb2f496, 32'shceb1f42f, 32'shceb0f3d1, 32'shceaff37a, 
               32'shceaef32b, 32'shceadf2e3, 32'shceacf2a3, 32'shceabf26b, 32'shceaaf23a, 32'shcea9f210, 32'shcea8f1ef, 32'shcea7f1d5, 
               32'shcea6f1c2, 32'shcea5f1b7, 32'shcea4f1b4, 32'shcea3f1b9, 32'shcea2f1c5, 32'shcea1f1d8, 32'shcea0f1f4, 32'shce9ff216, 
               32'shce9ef241, 32'shce9df273, 32'shce9cf2ad, 32'shce9bf2ee, 32'shce9af337, 32'shce99f387, 32'shce98f3e0, 32'shce97f43f, 
               32'shce96f4a7, 32'shce95f516, 32'shce94f58c, 32'shce93f60b, 32'shce92f691, 32'shce91f71e, 32'shce90f7b3, 32'shce8ff850, 
               32'shce8ef8f4, 32'shce8df9a0, 32'shce8cfa54, 32'shce8bfb0f, 32'shce8afbd2, 32'shce89fc9d, 32'shce88fd6f, 32'shce87fe48, 
               32'shce86ff2a, 32'shce860013, 32'shce850104, 32'shce8401fc, 32'shce8302fc, 32'shce820403, 32'shce810512, 32'shce800629, 
               32'shce7f0748, 32'shce7e086e, 32'shce7d099b, 32'shce7c0ad1, 32'shce7b0c0e, 32'shce7a0d52, 32'shce790e9f, 32'shce780ff3, 
               32'shce77114e, 32'shce7612b1, 32'shce75141c, 32'shce74158e, 32'shce731709, 32'shce72188a, 32'shce711a14, 32'shce701ba5, 
               32'shce6f1d3d, 32'shce6e1ede, 32'shce6d2086, 32'shce6c2235, 32'shce6b23ec, 32'shce6a25ab, 32'shce692772, 32'shce682940, 
               32'shce672b16, 32'shce662cf3, 32'shce652ed8, 32'shce6430c5, 32'shce6332ba, 32'shce6234b6, 32'shce6136b9, 32'shce6038c5, 
               32'shce5f3ad8, 32'shce5e3cf2, 32'shce5d3f15, 32'shce5c413f, 32'shce5b4370, 32'shce5a45aa, 32'shce5947eb, 32'shce584a33, 
               32'shce574c84, 32'shce564edc, 32'shce55513b, 32'shce5453a2, 32'shce535611, 32'shce525888, 32'shce515b06, 32'shce505d8c, 
               32'shce4f6019, 32'shce4e62af, 32'shce4d654c, 32'shce4c67f0, 32'shce4b6a9c, 32'shce4a6d50, 32'shce49700c, 32'shce4872cf, 
               32'shce47759a, 32'shce46786c, 32'shce457b47, 32'shce447e28, 32'shce438112, 32'shce428403, 32'shce4186fc, 32'shce4089fd, 
               32'shce3f8d05, 32'shce3e9015, 32'shce3d932c, 32'shce3c964c, 32'shce3b9973, 32'shce3a9ca1, 32'shce399fd7, 32'shce38a315, 
               32'shce37a65b, 32'shce36a9a8, 32'shce35acfd, 32'shce34b05a, 32'shce33b3be, 32'shce32b72a, 32'shce31ba9e, 32'shce30be19, 
               32'shce2fc19c, 32'shce2ec527, 32'shce2dc8ba, 32'shce2ccc54, 32'shce2bcff5, 32'shce2ad39f, 32'shce29d750, 32'shce28db09, 
               32'shce27dec9, 32'shce26e292, 32'shce25e662, 32'shce24ea39, 32'shce23ee18, 32'shce22f1ff, 32'shce21f5ee, 32'shce20f9e4, 
               32'shce1ffde2, 32'shce1f01e8, 32'shce1e05f6, 32'shce1d0a0b, 32'shce1c0e28, 32'shce1b124c, 32'shce1a1678, 32'shce191aac, 
               32'shce181ee8, 32'shce17232b, 32'shce162776, 32'shce152bc9, 32'shce143023, 32'shce133485, 32'shce1238ef, 32'shce113d60, 
               32'shce1041d9, 32'shce0f465a, 32'shce0e4ae3, 32'shce0d4f73, 32'shce0c540b, 32'shce0b58ab, 32'shce0a5d52, 32'shce096201, 
               32'shce0866b8, 32'shce076b77, 32'shce06703d, 32'shce05750b, 32'shce0479e0, 32'shce037ebe, 32'shce0283a3, 32'shce01888f, 
               32'shce008d84, 32'shcdff9280, 32'shcdfe9784, 32'shcdfd9c90, 32'shcdfca1a3, 32'shcdfba6be, 32'shcdfaabe1, 32'shcdf9b10b, 
               32'shcdf8b63d, 32'shcdf7bb77, 32'shcdf6c0b9, 32'shcdf5c602, 32'shcdf4cb53, 32'shcdf3d0ac, 32'shcdf2d60c, 32'shcdf1db74, 
               32'shcdf0e0e4, 32'shcdefe65c, 32'shcdeeebdb, 32'shcdedf162, 32'shcdecf6f1, 32'shcdebfc87, 32'shcdeb0226, 32'shcdea07cc, 
               32'shcde90d79, 32'shcde8132f, 32'shcde718ec, 32'shcde61eb1, 32'shcde5247d, 32'shcde42a52, 32'shcde3302e, 32'shcde23611, 
               32'shcde13bfd, 32'shcde041f0, 32'shcddf47eb, 32'shcdde4dee, 32'shcddd53f8, 32'shcddc5a0a, 32'shcddb6024, 32'shcdda6646, 
               32'shcdd96c6f, 32'shcdd872a0, 32'shcdd778d9, 32'shcdd67f19, 32'shcdd58562, 32'shcdd48bb2, 32'shcdd39209, 32'shcdd29869, 
               32'shcdd19ed0, 32'shcdd0a53f, 32'shcdcfabb6, 32'shcdceb234, 32'shcdcdb8ba, 32'shcdccbf48, 32'shcdcbc5de, 32'shcdcacc7b, 
               32'shcdc9d320, 32'shcdc8d9cd, 32'shcdc7e082, 32'shcdc6e73e, 32'shcdc5ee02, 32'shcdc4f4ce, 32'shcdc3fba2, 32'shcdc3027d, 
               32'shcdc20960, 32'shcdc1104b, 32'shcdc0173e, 32'shcdbf1e38, 32'shcdbe253a, 32'shcdbd2c44, 32'shcdbc3356, 32'shcdbb3a6f, 
               32'shcdba4190, 32'shcdb948b9, 32'shcdb84fea, 32'shcdb75722, 32'shcdb65e62, 32'shcdb565aa, 32'shcdb46cfa, 32'shcdb37451, 
               32'shcdb27bb0, 32'shcdb18317, 32'shcdb08a86, 32'shcdaf91fc, 32'shcdae997a, 32'shcdada100, 32'shcdaca88e, 32'shcdabb023, 
               32'shcdaab7c0, 32'shcda9bf65, 32'shcda8c712, 32'shcda7cec7, 32'shcda6d683, 32'shcda5de47, 32'shcda4e613, 32'shcda3ede6, 
               32'shcda2f5c2, 32'shcda1fda5, 32'shcda10590, 32'shcda00d82, 32'shcd9f157d, 32'shcd9e1d7f, 32'shcd9d2589, 32'shcd9c2d9a, 
               32'shcd9b35b4, 32'shcd9a3dd5, 32'shcd9945fe, 32'shcd984e2f, 32'shcd975668, 32'shcd965ea8, 32'shcd9566f0, 32'shcd946f40, 
               32'shcd937798, 32'shcd927ff7, 32'shcd91885e, 32'shcd9090cd, 32'shcd8f9944, 32'shcd8ea1c3, 32'shcd8daa49, 32'shcd8cb2d7, 
               32'shcd8bbb6d, 32'shcd8ac40b, 32'shcd89ccb0, 32'shcd88d55d, 32'shcd87de12, 32'shcd86e6cf, 32'shcd85ef94, 32'shcd84f860, 
               32'shcd840134, 32'shcd830a10, 32'shcd8212f4, 32'shcd811bdf, 32'shcd8024d3, 32'shcd7f2dce, 32'shcd7e36d1, 32'shcd7d3fdb, 
               32'shcd7c48ee, 32'shcd7b5208, 32'shcd7a5b2a, 32'shcd796454, 32'shcd786d85, 32'shcd7776bf, 32'shcd768000, 32'shcd758949, 
               32'shcd74929a, 32'shcd739bf2, 32'shcd72a553, 32'shcd71aebb, 32'shcd70b82b, 32'shcd6fc1a3, 32'shcd6ecb22, 32'shcd6dd4a9, 
               32'shcd6cde39, 32'shcd6be7d0, 32'shcd6af16e, 32'shcd69fb15, 32'shcd6904c3, 32'shcd680e79, 32'shcd671837, 32'shcd6621fd, 
               32'shcd652bcb, 32'shcd6435a0, 32'shcd633f7d, 32'shcd624962, 32'shcd61534f, 32'shcd605d44, 32'shcd5f6740, 32'shcd5e7144, 
               32'shcd5d7b50, 32'shcd5c8564, 32'shcd5b8f80, 32'shcd5a99a3, 32'shcd59a3ce, 32'shcd58ae01, 32'shcd57b83c, 32'shcd56c27f, 
               32'shcd55ccca, 32'shcd54d71c, 32'shcd53e176, 32'shcd52ebd8, 32'shcd51f642, 32'shcd5100b3, 32'shcd500b2d, 32'shcd4f15ae, 
               32'shcd4e2037, 32'shcd4d2ac8, 32'shcd4c3560, 32'shcd4b4001, 32'shcd4a4aa9, 32'shcd495559, 32'shcd486011, 32'shcd476ad1, 
               32'shcd467599, 32'shcd458068, 32'shcd448b3f, 32'shcd43961e, 32'shcd42a105, 32'shcd41abf4, 32'shcd40b6ea, 32'shcd3fc1e9, 
               32'shcd3eccef, 32'shcd3dd7fd, 32'shcd3ce313, 32'shcd3bee30, 32'shcd3af956, 32'shcd3a0483, 32'shcd390fb8, 32'shcd381af5, 
               32'shcd37263a, 32'shcd363187, 32'shcd353cdb, 32'shcd344837, 32'shcd33539c, 32'shcd325f08, 32'shcd316a7b, 32'shcd3075f7, 
               32'shcd2f817b, 32'shcd2e8d06, 32'shcd2d9899, 32'shcd2ca434, 32'shcd2bafd7, 32'shcd2abb81, 32'shcd29c734, 32'shcd28d2ee, 
               32'shcd27deb0, 32'shcd26ea7b, 32'shcd25f64c, 32'shcd250226, 32'shcd240e08, 32'shcd2319f1, 32'shcd2225e2, 32'shcd2131db, 
               32'shcd203ddc, 32'shcd1f49e5, 32'shcd1e55f6, 32'shcd1d620e, 32'shcd1c6e2e, 32'shcd1b7a57, 32'shcd1a8687, 32'shcd1992be, 
               32'shcd189efe, 32'shcd17ab46, 32'shcd16b795, 32'shcd15c3ec, 32'shcd14d04b, 32'shcd13dcb2, 32'shcd12e921, 32'shcd11f598, 
               32'shcd110216, 32'shcd100e9d, 32'shcd0f1b2b, 32'shcd0e27c1, 32'shcd0d345f, 32'shcd0c4105, 32'shcd0b4db3, 32'shcd0a5a68, 
               32'shcd096725, 32'shcd0873eb, 32'shcd0780b8, 32'shcd068d8d, 32'shcd059a6a, 32'shcd04a74e, 32'shcd03b43b, 32'shcd02c12f, 
               32'shcd01ce2b, 32'shcd00db30, 32'shccffe83c, 32'shccfef54f, 32'shccfe026b, 32'shccfd0f8f, 32'shccfc1cba, 32'shccfb29ed, 
               32'shccfa3729, 32'shccf9446c, 32'shccf851b7, 32'shccf75f09, 32'shccf66c64, 32'shccf579c7, 32'shccf48731, 32'shccf394a3, 
               32'shccf2a21d, 32'shccf1af9f, 32'shccf0bd29, 32'shccefcabb, 32'shcceed855, 32'shccede5f6, 32'shccecf3a0, 32'shccec0151, 
               32'shcceb0f0a, 32'shccea1ccb, 32'shcce92a94, 32'shcce83865, 32'shcce7463e, 32'shcce6541e, 32'shcce56206, 32'shcce46ff7, 
               32'shcce37def, 32'shcce28bef, 32'shcce199f7, 32'shcce0a807, 32'shccdfb61f, 32'shccdec43e, 32'shccddd266, 32'shccdce095, 
               32'shccdbeecc, 32'shccdafd0b, 32'shccda0b52, 32'shccd919a1, 32'shccd827f8, 32'shccd73657, 32'shccd644bd, 32'shccd5532c, 
               32'shccd461a2, 32'shccd37021, 32'shccd27ea7, 32'shccd18d35, 32'shccd09bcb, 32'shcccfaa69, 32'shccceb90e, 32'shcccdc7bc, 
               32'shccccd671, 32'shcccbe52f, 32'shcccaf3f4, 32'shccca02c1, 32'shccc91196, 32'shccc82073, 32'shccc72f58, 32'shccc63e45, 
               32'shccc54d3a, 32'shccc45c36, 32'shccc36b3b, 32'shccc27a47, 32'shccc1895c, 32'shccc09878, 32'shccbfa79c, 32'shccbeb6c8, 
               32'shccbdc5fc, 32'shccbcd538, 32'shccbbe47b, 32'shccbaf3c7, 32'shccba031a, 32'shccb91276, 32'shccb821d9, 32'shccb73144, 
               32'shccb640b8, 32'shccb55033, 32'shccb45fb6, 32'shccb36f41, 32'shccb27ed3, 32'shccb18e6e, 32'shccb09e11, 32'shccafadbb, 
               32'shccaebd6e, 32'shccadcd28, 32'shccacdcea, 32'shccabecb5, 32'shccaafc87, 32'shccaa0c61, 32'shcca91c43, 32'shcca82c2d, 
               32'shcca73c1e, 32'shcca64c18, 32'shcca55c1a, 32'shcca46c23, 32'shcca37c35, 32'shcca28c4e, 32'shcca19c6f, 32'shcca0ac99, 
               32'shcc9fbcca, 32'shcc9ecd03, 32'shcc9ddd44, 32'shcc9ced8d, 32'shcc9bfddd, 32'shcc9b0e36, 32'shcc9a1e97, 32'shcc992f00, 
               32'shcc983f70, 32'shcc974fe9, 32'shcc966069, 32'shcc9570f1, 32'shcc948182, 32'shcc93921a, 32'shcc92a2ba, 32'shcc91b362, 
               32'shcc90c412, 32'shcc8fd4ca, 32'shcc8ee58a, 32'shcc8df651, 32'shcc8d0721, 32'shcc8c17f9, 32'shcc8b28d8, 32'shcc8a39c0, 
               32'shcc894aaf, 32'shcc885ba7, 32'shcc876ca6, 32'shcc867dad, 32'shcc858ebc, 32'shcc849fd4, 32'shcc83b0f3, 32'shcc82c21a, 
               32'shcc81d349, 32'shcc80e47f, 32'shcc7ff5be, 32'shcc7f0705, 32'shcc7e1854, 32'shcc7d29aa, 32'shcc7c3b09, 32'shcc7b4c70, 
               32'shcc7a5dde, 32'shcc796f55, 32'shcc7880d3, 32'shcc779259, 32'shcc76a3e8, 32'shcc75b57e, 32'shcc74c71c, 32'shcc73d8c2, 
               32'shcc72ea70, 32'shcc71fc26, 32'shcc710de4, 32'shcc701faa, 32'shcc6f3178, 32'shcc6e434e, 32'shcc6d552c, 32'shcc6c6711, 
               32'shcc6b78ff, 32'shcc6a8af5, 32'shcc699cf2, 32'shcc68aef8, 32'shcc67c105, 32'shcc66d31b, 32'shcc65e538, 32'shcc64f75e, 
               32'shcc64098b, 32'shcc631bc0, 32'shcc622dfd, 32'shcc614043, 32'shcc605290, 32'shcc5f64e5, 32'shcc5e7742, 32'shcc5d89a7, 
               32'shcc5c9c14, 32'shcc5bae89, 32'shcc5ac106, 32'shcc59d38b, 32'shcc58e618, 32'shcc57f8ad, 32'shcc570b4a, 32'shcc561dee, 
               32'shcc55309b, 32'shcc544350, 32'shcc53560c, 32'shcc5268d1, 32'shcc517b9e, 32'shcc508e72, 32'shcc4fa14f, 32'shcc4eb433, 
               32'shcc4dc720, 32'shcc4cda14, 32'shcc4bed11, 32'shcc4b0015, 32'shcc4a1322, 32'shcc492636, 32'shcc483952, 32'shcc474c77, 
               32'shcc465fa3, 32'shcc4572d7, 32'shcc448614, 32'shcc439958, 32'shcc42aca4, 32'shcc41bff8, 32'shcc40d354, 32'shcc3fe6b8, 
               32'shcc3efa25, 32'shcc3e0d99, 32'shcc3d2115, 32'shcc3c3499, 32'shcc3b4825, 32'shcc3a5bb9, 32'shcc396f55, 32'shcc3882f9, 
               32'shcc3796a5, 32'shcc36aa59, 32'shcc35be15, 32'shcc34d1d9, 32'shcc33e5a5, 32'shcc32f979, 32'shcc320d55, 32'shcc312139, 
               32'shcc303524, 32'shcc2f4918, 32'shcc2e5d14, 32'shcc2d7118, 32'shcc2c8524, 32'shcc2b9938, 32'shcc2aad54, 32'shcc29c177, 
               32'shcc28d5a3, 32'shcc27e9d7, 32'shcc26fe13, 32'shcc261257, 32'shcc2526a2, 32'shcc243af6, 32'shcc234f52, 32'shcc2263b6, 
               32'shcc217822, 32'shcc208c95, 32'shcc1fa111, 32'shcc1eb595, 32'shcc1dca21, 32'shcc1cdeb5, 32'shcc1bf350, 32'shcc1b07f4, 
               32'shcc1a1ca0, 32'shcc193154, 32'shcc184610, 32'shcc175ad3, 32'shcc166f9f, 32'shcc158473, 32'shcc14994f, 32'shcc13ae33, 
               32'shcc12c31f, 32'shcc11d813, 32'shcc10ed0e, 32'shcc100212, 32'shcc0f171e, 32'shcc0e2c32, 32'shcc0d414e, 32'shcc0c5672, 
               32'shcc0b6b9e, 32'shcc0a80d2, 32'shcc09960e, 32'shcc08ab52, 32'shcc07c09e, 32'shcc06d5f2, 32'shcc05eb4e, 32'shcc0500b2, 
               32'shcc04161e, 32'shcc032b92, 32'shcc02410e, 32'shcc015692, 32'shcc006c1e, 32'shcbff81b2, 32'shcbfe974e, 32'shcbfdacf2, 
               32'shcbfcc29f, 32'shcbfbd853, 32'shcbfaee0f, 32'shcbfa03d3, 32'shcbf919a0, 32'shcbf82f74, 32'shcbf74550, 32'shcbf65b34, 
               32'shcbf57121, 32'shcbf48715, 32'shcbf39d12, 32'shcbf2b316, 32'shcbf1c923, 32'shcbf0df37, 32'shcbeff554, 32'shcbef0b78, 
               32'shcbee21a5, 32'shcbed37d9, 32'shcbec4e16, 32'shcbeb645b, 32'shcbea7aa7, 32'shcbe990fc, 32'shcbe8a759, 32'shcbe7bdbe, 
               32'shcbe6d42b, 32'shcbe5ea9f, 32'shcbe5011c, 32'shcbe417a1, 32'shcbe32e2e, 32'shcbe244c3, 32'shcbe15b60, 32'shcbe07205, 
               32'shcbdf88b3, 32'shcbde9f68, 32'shcbddb625, 32'shcbdcccea, 32'shcbdbe3b7, 32'shcbdafa8d, 32'shcbda116a, 32'shcbd92850, 
               32'shcbd83f3d, 32'shcbd75633, 32'shcbd66d30, 32'shcbd58436, 32'shcbd49b43, 32'shcbd3b259, 32'shcbd2c977, 32'shcbd1e09c, 
               32'shcbd0f7ca, 32'shcbd00f00, 32'shcbcf263e, 32'shcbce3d84, 32'shcbcd54d2, 32'shcbcc6c28, 32'shcbcb8386, 32'shcbca9aec, 
               32'shcbc9b25a, 32'shcbc8c9d1, 32'shcbc7e14f, 32'shcbc6f8d5, 32'shcbc61064, 32'shcbc527fa, 32'shcbc43f99, 32'shcbc3573f, 
               32'shcbc26eee, 32'shcbc186a5, 32'shcbc09e64, 32'shcbbfb62a, 32'shcbbecdf9, 32'shcbbde5d0, 32'shcbbcfdaf, 32'shcbbc1596, 
               32'shcbbb2d85, 32'shcbba457c, 32'shcbb95d7c, 32'shcbb87583, 32'shcbb78d92, 32'shcbb6a5aa, 32'shcbb5bdc9, 32'shcbb4d5f1, 
               32'shcbb3ee20, 32'shcbb30658, 32'shcbb21e98, 32'shcbb136df, 32'shcbb04f2f, 32'shcbaf6787, 32'shcbae7fe7, 32'shcbad984f, 
               32'shcbacb0bf, 32'shcbabc938, 32'shcbaae1b8, 32'shcba9fa40, 32'shcba912d1, 32'shcba82b69, 32'shcba7440a, 32'shcba65cb2, 
               32'shcba57563, 32'shcba48e1c, 32'shcba3a6dd, 32'shcba2bfa6, 32'shcba1d877, 32'shcba0f150, 32'shcba00a31, 32'shcb9f231a, 
               32'shcb9e3c0b, 32'shcb9d5505, 32'shcb9c6e06, 32'shcb9b8710, 32'shcb9aa021, 32'shcb99b93b, 32'shcb98d25d, 32'shcb97eb87, 
               32'shcb9704b9, 32'shcb961df3, 32'shcb953735, 32'shcb94507f, 32'shcb9369d1, 32'shcb92832c, 32'shcb919c8e, 32'shcb90b5f9, 
               32'shcb8fcf6b, 32'shcb8ee8e6, 32'shcb8e0269, 32'shcb8d1bf4, 32'shcb8c3587, 32'shcb8b4f22, 32'shcb8a68c5, 32'shcb898270, 
               32'shcb889c23, 32'shcb87b5df, 32'shcb86cfa2, 32'shcb85e96e, 32'shcb850342, 32'shcb841d1d, 32'shcb833701, 32'shcb8250ed, 
               32'shcb816ae1, 32'shcb8084de, 32'shcb7f9ee2, 32'shcb7eb8ee, 32'shcb7dd303, 32'shcb7ced1f, 32'shcb7c0744, 32'shcb7b2171, 
               32'shcb7a3ba5, 32'shcb7955e2, 32'shcb787027, 32'shcb778a75, 32'shcb76a4ca, 32'shcb75bf27, 32'shcb74d98d, 32'shcb73f3fa, 
               32'shcb730e70, 32'shcb7228ee, 32'shcb714373, 32'shcb705e01, 32'shcb6f7898, 32'shcb6e9336, 32'shcb6daddc, 32'shcb6cc88a, 
               32'shcb6be341, 32'shcb6afe00, 32'shcb6a18c6, 32'shcb693395, 32'shcb684e6c, 32'shcb67694b, 32'shcb668432, 32'shcb659f22, 
               32'shcb64ba19, 32'shcb63d518, 32'shcb62f020, 32'shcb620b30, 32'shcb612648, 32'shcb604168, 32'shcb5f5c90, 32'shcb5e77c0, 
               32'shcb5d92f8, 32'shcb5cae39, 32'shcb5bc981, 32'shcb5ae4d2, 32'shcb5a002b, 32'shcb591b8b, 32'shcb5836f4, 32'shcb575266, 
               32'shcb566ddf, 32'shcb558960, 32'shcb54a4ea, 32'shcb53c07b, 32'shcb52dc15, 32'shcb51f7b7, 32'shcb511361, 32'shcb502f13, 
               32'shcb4f4acd, 32'shcb4e6690, 32'shcb4d825a, 32'shcb4c9e2d, 32'shcb4bba08, 32'shcb4ad5ea, 32'shcb49f1d5, 32'shcb490dc9, 
               32'shcb4829c4, 32'shcb4745c7, 32'shcb4661d3, 32'shcb457de6, 32'shcb449a02, 32'shcb43b626, 32'shcb42d252, 32'shcb41ee86, 
               32'shcb410ac3, 32'shcb402707, 32'shcb3f4354, 32'shcb3e5fa8, 32'shcb3d7c05, 32'shcb3c986a, 32'shcb3bb4d7, 32'shcb3ad14d, 
               32'shcb39edca, 32'shcb390a50, 32'shcb3826dd, 32'shcb374373, 32'shcb366011, 32'shcb357cb7, 32'shcb349965, 32'shcb33b61c, 
               32'shcb32d2da, 32'shcb31efa1, 32'shcb310c70, 32'shcb302947, 32'shcb2f4626, 32'shcb2e630d, 32'shcb2d7ffc, 32'shcb2c9cf4, 
               32'shcb2bb9f4, 32'shcb2ad6fb, 32'shcb29f40b, 32'shcb291123, 32'shcb282e44, 32'shcb274b6c, 32'shcb26689d, 32'shcb2585d5, 
               32'shcb24a316, 32'shcb23c05f, 32'shcb22ddb1, 32'shcb21fb0a, 32'shcb21186b, 32'shcb2035d5, 32'shcb1f5347, 32'shcb1e70c1, 
               32'shcb1d8e43, 32'shcb1cabcd, 32'shcb1bc95f, 32'shcb1ae6fa, 32'shcb1a049d, 32'shcb192248, 32'shcb183ffb, 32'shcb175db6, 
               32'shcb167b79, 32'shcb159945, 32'shcb14b718, 32'shcb13d4f4, 32'shcb12f2d8, 32'shcb1210c4, 32'shcb112eb9, 32'shcb104cb5, 
               32'shcb0f6aba, 32'shcb0e88c7, 32'shcb0da6dc, 32'shcb0cc4f9, 32'shcb0be31e, 32'shcb0b014b, 32'shcb0a1f81, 32'shcb093dbf, 
               32'shcb085c05, 32'shcb077a53, 32'shcb0698a9, 32'shcb05b708, 32'shcb04d56e, 32'shcb03f3dd, 32'shcb031254, 32'shcb0230d3, 
               32'shcb014f5b, 32'shcb006dea, 32'shcaff8c82, 32'shcafeab22, 32'shcafdc9ca, 32'shcafce87a, 32'shcafc0732, 32'shcafb25f3, 
               32'shcafa44bc, 32'shcaf9638d, 32'shcaf88266, 32'shcaf7a147, 32'shcaf6c030, 32'shcaf5df22, 32'shcaf4fe1c, 32'shcaf41d1e, 
               32'shcaf33c28, 32'shcaf25b3a, 32'shcaf17a55, 32'shcaf09977, 32'shcaefb8a2, 32'shcaeed7d5, 32'shcaedf711, 32'shcaed1654, 
               32'shcaec35a0, 32'shcaeb54f3, 32'shcaea744f, 32'shcae993b4, 32'shcae8b320, 32'shcae7d295, 32'shcae6f211, 32'shcae61196, 
               32'shcae53123, 32'shcae450b9, 32'shcae37056, 32'shcae28ffc, 32'shcae1afaa, 32'shcae0cf60, 32'shcadfef1e, 32'shcadf0ee4, 
               32'shcade2eb3, 32'shcadd4e8a, 32'shcadc6e69, 32'shcadb8e50, 32'shcadaae40, 32'shcad9ce37, 32'shcad8ee37, 32'shcad80e3f, 
               32'shcad72e4f, 32'shcad64e68, 32'shcad56e88, 32'shcad48eb1, 32'shcad3aee2, 32'shcad2cf1b, 32'shcad1ef5d, 32'shcad10fa6, 
               32'shcad02ff8, 32'shcacf5052, 32'shcace70b4, 32'shcacd911f, 32'shcaccb191, 32'shcacbd20c, 32'shcacaf28f, 32'shcaca131a, 
               32'shcac933ae, 32'shcac8544a, 32'shcac774ed, 32'shcac69599, 32'shcac5b64e, 32'shcac4d70a, 32'shcac3f7cf, 32'shcac3189c, 
               32'shcac23971, 32'shcac15a4e, 32'shcac07b34, 32'shcabf9c21, 32'shcabebd17, 32'shcabdde16, 32'shcabcff1c, 32'shcabc202a, 
               32'shcabb4141, 32'shcaba6260, 32'shcab98388, 32'shcab8a4b7, 32'shcab7c5ef, 32'shcab6e72f, 32'shcab60877, 32'shcab529c7, 
               32'shcab44b1f, 32'shcab36c80, 32'shcab28de9, 32'shcab1af5a, 32'shcab0d0d4, 32'shcaaff255, 32'shcaaf13df, 32'shcaae3571, 
               32'shcaad570c, 32'shcaac78ae, 32'shcaab9a59, 32'shcaaabc0c, 32'shcaa9ddc7, 32'shcaa8ff8a, 32'shcaa82156, 32'shcaa7432a, 
               32'shcaa66506, 32'shcaa586ea, 32'shcaa4a8d7, 32'shcaa3cacc, 32'shcaa2ecc9, 32'shcaa20ece, 32'shcaa130db, 32'shcaa052f1, 
               32'shca9f750f, 32'shca9e9735, 32'shca9db964, 32'shca9cdb9a, 32'shca9bfdd9, 32'shca9b2020, 32'shca9a4270, 32'shca9964c7, 
               32'shca988727, 32'shca97a98f, 32'shca96cbff, 32'shca95ee78, 32'shca9510f8, 32'shca943381, 32'shca935613, 32'shca9278ac, 
               32'shca919b4e, 32'shca90bdf8, 32'shca8fe0aa, 32'shca8f0364, 32'shca8e2627, 32'shca8d48f2, 32'shca8c6bc5, 32'shca8b8ea0, 
               32'shca8ab184, 32'shca89d470, 32'shca88f764, 32'shca881a60, 32'shca873d65, 32'shca866072, 32'shca858387, 32'shca84a6a4, 
               32'shca83c9ca, 32'shca82ecf8, 32'shca82102e, 32'shca81336c, 32'shca8056b3, 32'shca7f7a02, 32'shca7e9d59, 32'shca7dc0b8, 
               32'shca7ce420, 32'shca7c078f, 32'shca7b2b08, 32'shca7a4e88, 32'shca797211, 32'shca7895a1, 32'shca77b93b, 32'shca76dcdc, 
               32'shca760086, 32'shca752437, 32'shca7447f2, 32'shca736bb4, 32'shca728f7f, 32'shca71b351, 32'shca70d72d, 32'shca6ffb10, 
               32'shca6f1efc, 32'shca6e42f0, 32'shca6d66ec, 32'shca6c8af0, 32'shca6baefd, 32'shca6ad312, 32'shca69f72f, 32'shca691b55, 
               32'shca683f83, 32'shca6763b9, 32'shca6687f7, 32'shca65ac3e, 32'shca64d08d, 32'shca63f4e4, 32'shca631943, 32'shca623dab, 
               32'shca61621b, 32'shca608693, 32'shca5fab13, 32'shca5ecf9c, 32'shca5df42d, 32'shca5d18c6, 32'shca5c3d68, 32'shca5b6212, 
               32'shca5a86c4, 32'shca59ab7e, 32'shca58d041, 32'shca57f50c, 32'shca5719df, 32'shca563eba, 32'shca55639e, 32'shca54888a, 
               32'shca53ad7e, 32'shca52d27b, 32'shca51f780, 32'shca511c8d, 32'shca5041a2, 32'shca4f66c0, 32'shca4e8be6, 32'shca4db114, 
               32'shca4cd64b, 32'shca4bfb89, 32'shca4b20d0, 32'shca4a4620, 32'shca496b77, 32'shca4890d7, 32'shca47b640, 32'shca46dbb0, 
               32'shca460129, 32'shca4526aa, 32'shca444c33, 32'shca4371c5, 32'shca42975f, 32'shca41bd01, 32'shca40e2ac, 32'shca40085e, 
               32'shca3f2e19, 32'shca3e53dd, 32'shca3d79a8, 32'shca3c9f7c, 32'shca3bc559, 32'shca3aeb3d, 32'shca3a112a, 32'shca39371f, 
               32'shca385d1d, 32'shca378322, 32'shca36a930, 32'shca35cf47, 32'shca34f565, 32'shca341b8c, 32'shca3341bb, 32'shca3267f3, 
               32'shca318e32, 32'shca30b47a, 32'shca2fdacb, 32'shca2f0123, 32'shca2e2784, 32'shca2d4dee, 32'shca2c745f, 32'shca2b9ad9, 
               32'shca2ac15b, 32'shca29e7e6, 32'shca290e79, 32'shca283514, 32'shca275bb7, 32'shca268263, 32'shca25a917, 32'shca24cfd3, 
               32'shca23f698, 32'shca231d64, 32'shca22443a, 32'shca216b17, 32'shca2091fd, 32'shca1fb8eb, 32'shca1edfe2, 32'shca1e06e0, 
               32'shca1d2de7, 32'shca1c54f7, 32'shca1b7c0e, 32'shca1aa32e, 32'shca19ca57, 32'shca18f187, 32'shca1818c0, 32'shca174001, 
               32'shca16674b, 32'shca158e9d, 32'shca14b5f7, 32'shca13dd59, 32'shca1304c4, 32'shca122c37, 32'shca1153b3, 32'shca107b37, 
               32'shca0fa2c3, 32'shca0eca57, 32'shca0df1f4, 32'shca0d1999, 32'shca0c4146, 32'shca0b68fc, 32'shca0a90ba, 32'shca09b880, 
               32'shca08e04f, 32'shca080826, 32'shca073005, 32'shca0657ed, 32'shca057fdd, 32'shca04a7d5, 32'shca03cfd5, 32'shca02f7de, 
               32'shca021fef, 32'shca014809, 32'shca00702b, 32'shc9ff9855, 32'shc9fec088, 32'shc9fde8c2, 32'shc9fd1106, 32'shc9fc3951, 
               32'shc9fb61a5, 32'shc9fa8a01, 32'shc9f9b266, 32'shc9f8dad3, 32'shc9f80348, 32'shc9f72bc5, 32'shc9f6544b, 32'shc9f57cd9, 
               32'shc9f4a570, 32'shc9f3ce0f, 32'shc9f2f6b6, 32'shc9f21f65, 32'shc9f1481d, 32'shc9f070dd, 32'shc9ef99a6, 32'shc9eec277, 
               32'shc9edeb50, 32'shc9ed1431, 32'shc9ec3d1b, 32'shc9eb660d, 32'shc9ea8f08, 32'shc9e9b80b, 32'shc9e8e116, 32'shc9e80a2a, 
               32'shc9e73346, 32'shc9e65c6a, 32'shc9e58596, 32'shc9e4aecb, 32'shc9e3d809, 32'shc9e3014e, 32'shc9e22a9c, 32'shc9e153f3, 
               32'shc9e07d51, 32'shc9dfa6b8, 32'shc9ded028, 32'shc9ddf99f, 32'shc9dd231f, 32'shc9dc4ca8, 32'shc9db7639, 32'shc9da9fd2, 
               32'shc9d9c973, 32'shc9d8f31d, 32'shc9d81ccf, 32'shc9d7468a, 32'shc9d6704c, 32'shc9d59a18, 32'shc9d4c3eb, 32'shc9d3edc7, 
               32'shc9d317ab, 32'shc9d24198, 32'shc9d16b8d, 32'shc9d0958a, 32'shc9cfbf90, 32'shc9cee99e, 32'shc9ce13b4, 32'shc9cd3dd3, 
               32'shc9cc67fa, 32'shc9cb922a, 32'shc9cabc62, 32'shc9c9e6a2, 32'shc9c910ea, 32'shc9c83b3b, 32'shc9c76595, 32'shc9c68ff6, 
               32'shc9c5ba60, 32'shc9c4e4d3, 32'shc9c40f4d, 32'shc9c339d0, 32'shc9c2645c, 32'shc9c18ef0, 32'shc9c0b98c, 32'shc9bfe430, 
               32'shc9bf0edd, 32'shc9be3993, 32'shc9bd6450, 32'shc9bc8f16, 32'shc9bbb9e5, 32'shc9bae4bc, 32'shc9ba0f9b, 32'shc9b93a82, 
               32'shc9b86572, 32'shc9b7906a, 32'shc9b6bb6b, 32'shc9b5e674, 32'shc9b51185, 32'shc9b43c9f, 32'shc9b367c1, 32'shc9b292eb, 
               32'shc9b1be1e, 32'shc9b0e95a, 32'shc9b0149d, 32'shc9af3fe9, 32'shc9ae6b3d, 32'shc9ad969a, 32'shc9acc1ff, 32'shc9abed6d, 
               32'shc9ab18e3, 32'shc9aa4461, 32'shc9a96fe7, 32'shc9a89b76, 32'shc9a7c70e, 32'shc9a6f2ae, 32'shc9a61e56, 32'shc9a54a06, 
               32'shc9a475bf, 32'shc9a3a180, 32'shc9a2cd4a, 32'shc9a1f91c, 32'shc9a124f7, 32'shc9a050d9, 32'shc99f7cc5, 32'shc99ea8b8, 
               32'shc99dd4b4, 32'shc99d00b8, 32'shc99c2cc5, 32'shc99b58da, 32'shc99a84f8, 32'shc999b11e, 32'shc998dd4c, 32'shc9980983, 
               32'shc99735c2, 32'shc9966209, 32'shc9958e59, 32'shc994bab1, 32'shc993e712, 32'shc993137b, 32'shc9923fed, 32'shc9916c66, 
               32'shc99098e9, 32'shc98fc573, 32'shc98ef206, 32'shc98e1ea2, 32'shc98d4b45, 32'shc98c77f2, 32'shc98ba4a6, 32'shc98ad163, 
               32'shc989fe29, 32'shc9892af6, 32'shc98857cd, 32'shc98784ab, 32'shc986b192, 32'shc985de82, 32'shc9850b79, 32'shc9843879, 
               32'shc9836582, 32'shc9829293, 32'shc981bfac, 32'shc980ecce, 32'shc98019f8, 32'shc97f472b, 32'shc97e7466, 32'shc97da1aa, 
               32'shc97ccef5, 32'shc97bfc4a, 32'shc97b29a6, 32'shc97a570b, 32'shc9798479, 32'shc978b1ef, 32'shc977df6d, 32'shc9770cf4, 
               32'shc9763a83, 32'shc975681a, 32'shc97495ba, 32'shc973c362, 32'shc972f113, 32'shc9721ecc, 32'shc9714c8e, 32'shc9707a58, 
               32'shc96fa82a, 32'shc96ed605, 32'shc96e03e8, 32'shc96d31d4, 32'shc96c5fc8, 32'shc96b8dc4, 32'shc96abbc9, 32'shc969e9d7, 
               32'shc96917ec, 32'shc968460a, 32'shc9677431, 32'shc966a260, 32'shc965d097, 32'shc964fed7, 32'shc9642d1f, 32'shc9635b70, 
               32'shc96289c9, 32'shc961b82b, 32'shc960e695, 32'shc9601507, 32'shc95f4382, 32'shc95e7205, 32'shc95da090, 32'shc95ccf25, 
               32'shc95bfdc1, 32'shc95b2c66, 32'shc95a5b13, 32'shc95989c9, 32'shc958b887, 32'shc957e74e, 32'shc957161d, 32'shc95644f4, 
               32'shc95573d4, 32'shc954a2bc, 32'shc953d1ad, 32'shc95300a6, 32'shc9522fa8, 32'shc9515eb2, 32'shc9508dc5, 32'shc94fbce0, 
               32'shc94eec03, 32'shc94e1b2f, 32'shc94d4a63, 32'shc94c79a0, 32'shc94ba8e5, 32'shc94ad832, 32'shc94a0788, 32'shc94936e7, 
               32'shc948664d, 32'shc94795bd, 32'shc946c534, 32'shc945f4b4, 32'shc945243d, 32'shc94453ce, 32'shc9438368, 32'shc942b30a, 
               32'shc941e2b4, 32'shc9411267, 32'shc9404222, 32'shc93f71e6, 32'shc93ea1b2, 32'shc93dd186, 32'shc93d0163, 32'shc93c3149, 
               32'shc93b6137, 32'shc93a912d, 32'shc939c12c, 32'shc938f133, 32'shc9382143, 32'shc937515b, 32'shc936817b, 32'shc935b1a5, 
               32'shc934e1d6, 32'shc9341210, 32'shc9334252, 32'shc932729d, 32'shc931a2f0, 32'shc930d34c, 32'shc93003b0, 32'shc92f341d, 
               32'shc92e6492, 32'shc92d9510, 32'shc92cc596, 32'shc92bf624, 32'shc92b26bb, 32'shc92a575a, 32'shc9298802, 32'shc928b8b3, 
               32'shc927e96b, 32'shc9271a2d, 32'shc9264af6, 32'shc9257bc8, 32'shc924aca3, 32'shc923dd86, 32'shc9230e71, 32'shc9223f65, 
               32'shc9217062, 32'shc920a167, 32'shc91fd274, 32'shc91f038a, 32'shc91e34a8, 32'shc91d65cf, 32'shc91c96fe, 32'shc91bc836, 
               32'shc91af976, 32'shc91a2abe, 32'shc9195c0f, 32'shc9188d69, 32'shc917becb, 32'shc916f035, 32'shc91621a8, 32'shc9155324, 
               32'shc91484a8, 32'shc913b634, 32'shc912e7c9, 32'shc9121966, 32'shc9114b0c, 32'shc9107cba, 32'shc90fae71, 32'shc90ee030, 
               32'shc90e11f7, 32'shc90d43c8, 32'shc90c75a0, 32'shc90ba781, 32'shc90ad96b, 32'shc90a0b5d, 32'shc9093d57, 32'shc9086f5a, 
               32'shc907a166, 32'shc906d379, 32'shc9060596, 32'shc90537bb, 32'shc90469e8, 32'shc9039c1e, 32'shc902ce5c, 32'shc90200a3, 
               32'shc90132f2, 32'shc900654a, 32'shc8ff97aa, 32'shc8feca13, 32'shc8fdfc84, 32'shc8fd2efe, 32'shc8fc6180, 32'shc8fb940b, 
               32'shc8fac69e, 32'shc8f9f939, 32'shc8f92bdd, 32'shc8f85e8a, 32'shc8f7913f, 32'shc8f6c3fd, 32'shc8f5f6c3, 32'shc8f52991, 
               32'shc8f45c68, 32'shc8f38f48, 32'shc8f2c230, 32'shc8f1f520, 32'shc8f12819, 32'shc8f05b1a, 32'shc8ef8e24, 32'shc8eec137, 
               32'shc8edf452, 32'shc8ed2775, 32'shc8ec5aa1, 32'shc8eb8dd6, 32'shc8eac112, 32'shc8e9f458, 32'shc8e927a6, 32'shc8e85afc, 
               32'shc8e78e5b, 32'shc8e6c1c2, 32'shc8e5f532, 32'shc8e528ab, 32'shc8e45c2c, 32'shc8e38fb5, 32'shc8e2c347, 32'shc8e1f6e1, 
               32'shc8e12a84, 32'shc8e05e2f, 32'shc8df91e3, 32'shc8dec5a0, 32'shc8ddf965, 32'shc8dd2d32, 32'shc8dc6108, 32'shc8db94e6, 
               32'shc8dac8cd, 32'shc8d9fcbd, 32'shc8d930b4, 32'shc8d864b5, 32'shc8d798be, 32'shc8d6cccf, 32'shc8d600e9, 32'shc8d5350c, 
               32'shc8d46936, 32'shc8d39d6a, 32'shc8d2d1a6, 32'shc8d205ea, 32'shc8d13a37, 32'shc8d06e8d, 32'shc8cfa2eb, 32'shc8ced751, 
               32'shc8ce0bc0, 32'shc8cd4038, 32'shc8cc74b8, 32'shc8cba940, 32'shc8caddd1, 32'shc8ca126b, 32'shc8c9470d, 32'shc8c87bb8, 
               32'shc8c7b06b, 32'shc8c6e527, 32'shc8c619eb, 32'shc8c54eb7, 32'shc8c4838d, 32'shc8c3b86a, 32'shc8c2ed50, 32'shc8c2223f, 
               32'shc8c15736, 32'shc8c08c36, 32'shc8bfc13f, 32'shc8bef64f, 32'shc8be2b69, 32'shc8bd608b, 32'shc8bc95b5, 32'shc8bbcae8, 
               32'shc8bb0023, 32'shc8ba3567, 32'shc8b96ab4, 32'shc8b8a009, 32'shc8b7d566, 32'shc8b70acc, 32'shc8b6403b, 32'shc8b575b2, 
               32'shc8b4ab32, 32'shc8b3e0ba, 32'shc8b3164a, 32'shc8b24be4, 32'shc8b18185, 32'shc8b0b730, 32'shc8afece2, 32'shc8af229e, 
               32'shc8ae5862, 32'shc8ad8e2e, 32'shc8acc403, 32'shc8abf9e0, 32'shc8ab2fc6, 32'shc8aa65b5, 32'shc8a99bac, 32'shc8a8d1ac, 
               32'shc8a807b4, 32'shc8a73dc4, 32'shc8a673dd, 32'shc8a5a9ff, 32'shc8a4e029, 32'shc8a4165c, 32'shc8a34c98, 32'shc8a282db, 
               32'shc8a1b928, 32'shc8a0ef7d, 32'shc8a025da, 32'shc89f5c40, 32'shc89e92af, 32'shc89dc926, 32'shc89cffa6, 32'shc89c362e, 
               32'shc89b6cbf, 32'shc89aa358, 32'shc899d9fa, 32'shc89910a4, 32'shc8984757, 32'shc8977e12, 32'shc896b4d6, 32'shc895eba3, 
               32'shc8952278, 32'shc8945956, 32'shc893903c, 32'shc892c72b, 32'shc891fe22, 32'shc8913522, 32'shc8906c2a, 32'shc88fa33b, 
               32'shc88eda54, 32'shc88e1176, 32'shc88d48a1, 32'shc88c7fd4, 32'shc88bb710, 32'shc88aee54, 32'shc88a25a1, 32'shc8895cf6, 
               32'shc8889454, 32'shc887cbba, 32'shc8870329, 32'shc8863aa1, 32'shc8857221, 32'shc884a9aa, 32'shc883e13b, 32'shc88318d5, 
               32'shc8825077, 32'shc8818822, 32'shc880bfd5, 32'shc87ff791, 32'shc87f2f56, 32'shc87e6723, 32'shc87d9ef8, 32'shc87cd6d7, 
               32'shc87c0ebd, 32'shc87b46ad, 32'shc87a7ea5, 32'shc879b6a5, 32'shc878eeae, 32'shc87826c0, 32'shc8775eda, 32'shc87696fd, 
               32'shc875cf28, 32'shc875075c, 32'shc8743f98, 32'shc87377dd, 32'shc872b02b, 32'shc871e881, 32'shc87120e0, 32'shc8705947, 
               32'shc86f91b7, 32'shc86eca2f, 32'shc86e02b0, 32'shc86d3b3a, 32'shc86c73cc, 32'shc86bac66, 32'shc86ae50a, 32'shc86a1db6, 
               32'shc869566a, 32'shc8688f27, 32'shc867c7ec, 32'shc86700ba, 32'shc8663991, 32'shc8657270, 32'shc864ab58, 32'shc863e449, 
               32'shc8631d42, 32'shc8625643, 32'shc8618f4d, 32'shc860c860, 32'shc860017b, 32'shc85f3a9f, 32'shc85e73cc, 32'shc85dad01, 
               32'shc85ce63e, 32'shc85c1f84, 32'shc85b58d3, 32'shc85a922b, 32'shc859cb8a, 32'shc85904f3, 32'shc8583e64, 32'shc85777de, 
               32'shc856b160, 32'shc855eaeb, 32'shc855247e, 32'shc8545e1a, 32'shc85397bf, 32'shc852d16c, 32'shc8520b22, 32'shc85144e0, 
               32'shc8507ea7, 32'shc84fb877, 32'shc84ef24f, 32'shc84e2c2f, 32'shc84d6619, 32'shc84ca00b, 32'shc84bda05, 32'shc84b1408, 
               32'shc84a4e14, 32'shc8498828, 32'shc848c245, 32'shc847fc6a, 32'shc8473698, 32'shc84670cf, 32'shc845ab0e, 32'shc844e556, 
               32'shc8441fa6, 32'shc84359ff, 32'shc8429461, 32'shc841cecb, 32'shc841093e, 32'shc84043b9, 32'shc83f7e3d, 32'shc83eb8ca, 
               32'shc83df35f, 32'shc83d2dfd, 32'shc83c68a3, 32'shc83ba352, 32'shc83ade0a, 32'shc83a18ca, 32'shc8395393, 32'shc8388e64, 
               32'shc837c93e, 32'shc8370420, 32'shc8363f0c, 32'shc83579ff, 32'shc834b4fc, 32'shc833f001, 32'shc8332b0e, 32'shc8326625, 
               32'shc831a143, 32'shc830dc6b, 32'shc830179b, 32'shc82f52d3, 32'shc82e8e15, 32'shc82dc95e, 32'shc82d04b1, 32'shc82c400c, 
               32'shc82b7b70, 32'shc82ab6dc, 32'shc829f251, 32'shc8292dce, 32'shc8286954, 32'shc827a4e3, 32'shc826e07a, 32'shc8261c1a, 
               32'shc82557c3, 32'shc8249374, 32'shc823cf2e, 32'shc8230af0, 32'shc82246bb, 32'shc821828f, 32'shc820be6b, 32'shc81ffa50, 
               32'shc81f363d, 32'shc81e7233, 32'shc81dae32, 32'shc81cea39, 32'shc81c2649, 32'shc81b6262, 32'shc81a9e83, 32'shc819daad, 
               32'shc81916df, 32'shc818531a, 32'shc8178f5e, 32'shc816cbaa, 32'shc81607ff, 32'shc815445d, 32'shc81480c3, 32'shc813bd32, 
               32'shc812f9a9, 32'shc8123629, 32'shc81172b2, 32'shc810af43, 32'shc80febdd, 32'shc80f287f, 32'shc80e652b, 32'shc80da1de, 
               32'shc80cde9b, 32'shc80c1b60, 32'shc80b582e, 32'shc80a9504, 32'shc809d1e3, 32'shc8090eca, 32'shc8084bba, 32'shc80788b3, 
               32'shc806c5b5, 32'shc80602bf, 32'shc8053fd2, 32'shc8047ced, 32'shc803ba11, 32'shc802f73d, 32'shc8023473, 32'shc80171b1, 
               32'shc800aef7, 32'shc7ffec46, 32'shc7ff299e, 32'shc7fe66fe, 32'shc7fda468, 32'shc7fce1d9, 32'shc7fc1f54, 32'shc7fb5cd7, 
               32'shc7fa9a62, 32'shc7f9d7f6, 32'shc7f91593, 32'shc7f85339, 32'shc7f790e7, 32'shc7f6ce9e, 32'shc7f60c5d, 32'shc7f54a25, 
               32'shc7f487f6, 32'shc7f3c5cf, 32'shc7f303b1, 32'shc7f2419c, 32'shc7f17f8f, 32'shc7f0bd8b, 32'shc7effb90, 32'shc7ef399d, 
               32'shc7ee77b3, 32'shc7edb5d2, 32'shc7ecf3f9, 32'shc7ec3229, 32'shc7eb7061, 32'shc7eaaea2, 32'shc7e9ecec, 32'shc7e92b3e, 
               32'shc7e8699a, 32'shc7e7a7fd, 32'shc7e6e66a, 32'shc7e624df, 32'shc7e5635c, 32'shc7e4a1e3, 32'shc7e3e072, 32'shc7e31f09, 
               32'shc7e25daa, 32'shc7e19c53, 32'shc7e0db04, 32'shc7e019be, 32'shc7df5881, 32'shc7de974d, 32'shc7ddd621, 32'shc7dd14fe, 
               32'shc7dc53e3, 32'shc7db92d2, 32'shc7dad1c9, 32'shc7da10c8, 32'shc7d94fd0, 32'shc7d88ee1, 32'shc7d7cdfb, 32'shc7d70d1d, 
               32'shc7d64c47, 32'shc7d58b7b, 32'shc7d4cab7, 32'shc7d409fc, 32'shc7d34949, 32'shc7d2889f, 32'shc7d1c7fe, 32'shc7d10766, 
               32'shc7d046d6, 32'shc7cf864e, 32'shc7cec5d0, 32'shc7ce055a, 32'shc7cd44ed, 32'shc7cc8488, 32'shc7cbc42c, 32'shc7cb03d9, 
               32'shc7ca438f, 32'shc7c9834d, 32'shc7c8c313, 32'shc7c802e3, 32'shc7c742bb, 32'shc7c6829c, 32'shc7c5c285, 32'shc7c50277, 
               32'shc7c44272, 32'shc7c38276, 32'shc7c2c282, 32'shc7c20297, 32'shc7c142b4, 32'shc7c082da, 32'shc7bfc309, 32'shc7bf0340, 
               32'shc7be4381, 32'shc7bd83ca, 32'shc7bcc41b, 32'shc7bc0475, 32'shc7bb44d8, 32'shc7ba8544, 32'shc7b9c5b8, 32'shc7b90635, 
               32'shc7b846ba, 32'shc7b78749, 32'shc7b6c7e0, 32'shc7b6087f, 32'shc7b54928, 32'shc7b489d9, 32'shc7b3ca92, 32'shc7b30b55, 
               32'shc7b24c20, 32'shc7b18cf3, 32'shc7b0cdd0, 32'shc7b00eb5, 32'shc7af4fa3, 32'shc7ae9099, 32'shc7add198, 32'shc7ad12a0, 
               32'shc7ac53b1, 32'shc7ab94ca, 32'shc7aad5ec, 32'shc7aa1716, 32'shc7a9584a, 32'shc7a89986, 32'shc7a7daca, 32'shc7a71c18, 
               32'shc7a65d6e, 32'shc7a59ecc, 32'shc7a4e034, 32'shc7a421a4, 32'shc7a3631d, 32'shc7a2a49e, 32'shc7a1e628, 32'shc7a127bb, 
               32'shc7a06957, 32'shc79faafb, 32'shc79eeca8, 32'shc79e2e5d, 32'shc79d701c, 32'shc79cb1e3, 32'shc79bf3b3, 32'shc79b358b, 
               32'shc79a776c, 32'shc799b956, 32'shc798fb48, 32'shc7983d44, 32'shc7977f48, 32'shc796c154, 32'shc7960369, 32'shc7954587, 
               32'shc79487ae, 32'shc793c9de, 32'shc7930c16, 32'shc7924e56, 32'shc79190a0, 32'shc790d2f2, 32'shc790154d, 32'shc78f57b1, 
               32'shc78e9a1d, 32'shc78ddc92, 32'shc78d1f10, 32'shc78c6196, 32'shc78ba425, 32'shc78ae6bd, 32'shc78a295e, 32'shc7896c07, 
               32'shc788aeb9, 32'shc787f174, 32'shc7873437, 32'shc7867703, 32'shc785b9d8, 32'shc784fcb5, 32'shc7843f9c, 32'shc783828b, 
               32'shc782c582, 32'shc7820883, 32'shc7814b8c, 32'shc7808e9d, 32'shc77fd1b8, 32'shc77f14db, 32'shc77e5807, 32'shc77d9b3c, 
               32'shc77cde79, 32'shc77c21bf, 32'shc77b650e, 32'shc77aa865, 32'shc779ebc5, 32'shc7792f2e, 32'shc77872a0, 32'shc777b61a, 
               32'shc776f99d, 32'shc7763d29, 32'shc77580be, 32'shc774c45b, 32'shc7740801, 32'shc7734bb0, 32'shc7728f67, 32'shc771d327, 
               32'shc77116f0, 32'shc7705ac2, 32'shc76f9e9c, 32'shc76ee27f, 32'shc76e266b, 32'shc76d6a5f, 32'shc76cae5c, 32'shc76bf262, 
               32'shc76b3671, 32'shc76a7a88, 32'shc769bea8, 32'shc76902d1, 32'shc7684702, 32'shc7678b3d, 32'shc766cf80, 32'shc76613cb, 
               32'shc7655820, 32'shc7649c7d, 32'shc763e0e3, 32'shc7632552, 32'shc76269c9, 32'shc761ae49, 32'shc760f2d2, 32'shc7603763, 
               32'shc75f7bfe, 32'shc75ec0a1, 32'shc75e054c, 32'shc75d4a01, 32'shc75c8ebe, 32'shc75bd384, 32'shc75b1853, 32'shc75a5d2a, 
               32'shc759a20a, 32'shc758e6f3, 32'shc7582be5, 32'shc75770df, 32'shc756b5e2, 32'shc755faee, 32'shc7554003, 32'shc7548520, 
               32'shc753ca46, 32'shc7530f75, 32'shc75254ac, 32'shc75199ed, 32'shc750df36, 32'shc7502488, 32'shc74f69e2, 32'shc74eaf45, 
               32'shc74df4b1, 32'shc74d3a26, 32'shc74c7fa4, 32'shc74bc52a, 32'shc74b0ab9, 32'shc74a5050, 32'shc74995f1, 32'shc748db9a, 
               32'shc748214c, 32'shc7476707, 32'shc746acca, 32'shc745f296, 32'shc745386b, 32'shc7447e49, 32'shc743c42f, 32'shc7430a1f, 
               32'shc7425016, 32'shc7419617, 32'shc740dc21, 32'shc7402233, 32'shc73f684e, 32'shc73eae71, 32'shc73df49e, 32'shc73d3ad3, 
               32'shc73c8111, 32'shc73bc758, 32'shc73b0da7, 32'shc73a53ff, 32'shc7399a60, 32'shc738e0ca, 32'shc738273d, 32'shc7376db8, 
               32'shc736b43c, 32'shc735fac8, 32'shc735415e, 32'shc73487fc, 32'shc733cea3, 32'shc7331553, 32'shc7325c0c, 32'shc731a2cd, 
               32'shc730e997, 32'shc730306a, 32'shc72f7745, 32'shc72ebe2a, 32'shc72e0517, 32'shc72d4c0d, 32'shc72c930b, 32'shc72bda13, 
               32'shc72b2123, 32'shc72a683c, 32'shc729af5d, 32'shc728f688, 32'shc7283dbb, 32'shc72784f7, 32'shc726cc3c, 32'shc7261389, 
               32'shc7255ae0, 32'shc724a23f, 32'shc723e9a6, 32'shc7233117, 32'shc7227890, 32'shc721c013, 32'shc721079d, 32'shc7204f31, 
               32'shc71f96ce, 32'shc71ede73, 32'shc71e2621, 32'shc71d6dd7, 32'shc71cb597, 32'shc71bfd5f, 32'shc71b4530, 32'shc71a8d0a, 
               32'shc719d4ed, 32'shc7191cd8, 32'shc71864cc, 32'shc717acc9, 32'shc716f4cf, 32'shc7163cdd, 32'shc71584f5, 32'shc714cd15, 
               32'shc714153e, 32'shc7135d6f, 32'shc712a5aa, 32'shc711eded, 32'shc7113639, 32'shc7107e8d, 32'shc70fc6eb, 32'shc70f0f51, 
               32'shc70e57c0, 32'shc70da038, 32'shc70ce8b9, 32'shc70c3142, 32'shc70b79d4, 32'shc70ac26f, 32'shc70a0b13, 32'shc70953c0, 
               32'shc7089c75, 32'shc707e533, 32'shc7072dfa, 32'shc70676ca, 32'shc705bfa2, 32'shc7050883, 32'shc704516d, 32'shc7039a60, 
               32'shc702e35c, 32'shc7022c60, 32'shc701756d, 32'shc700be83, 32'shc70007a2, 32'shc6ff50ca, 32'shc6fe99fa, 32'shc6fde333, 
               32'shc6fd2c75, 32'shc6fc75c0, 32'shc6fbbf13, 32'shc6fb0870, 32'shc6fa51d5, 32'shc6f99b43, 32'shc6f8e4b9, 32'shc6f82e39, 
               32'shc6f777c1, 32'shc6f6c152, 32'shc6f60aec, 32'shc6f5548f, 32'shc6f49e3a, 32'shc6f3e7ee, 32'shc6f331ab, 32'shc6f27b71, 
               32'shc6f1c540, 32'shc6f10f17, 32'shc6f058f8, 32'shc6efa2e1, 32'shc6eeecd3, 32'shc6ee36cd, 32'shc6ed80d1, 32'shc6eccadd, 
               32'shc6ec14f2, 32'shc6eb5f10, 32'shc6eaa936, 32'shc6e9f366, 32'shc6e93d9e, 32'shc6e887df, 32'shc6e7d229, 32'shc6e71c7c, 
               32'shc6e666d7, 32'shc6e5b13c, 32'shc6e4fba9, 32'shc6e4461f, 32'shc6e3909d, 32'shc6e2db25, 32'shc6e225b5, 32'shc6e1704e, 
               32'shc6e0baf0, 32'shc6e0059b, 32'shc6df504f, 32'shc6de9b0b, 32'shc6dde5d0, 32'shc6dd309e, 32'shc6dc7b75, 32'shc6dbc654, 
               32'shc6db113d, 32'shc6da5c2e, 32'shc6d9a728, 32'shc6d8f22b, 32'shc6d83d37, 32'shc6d7884b, 32'shc6d6d369, 32'shc6d61e8f, 
               32'shc6d569be, 32'shc6d4b4f5, 32'shc6d40036, 32'shc6d34b7f, 32'shc6d296d1, 32'shc6d1e22d, 32'shc6d12d90, 32'shc6d078fd, 
               32'shc6cfc472, 32'shc6cf0ff1, 32'shc6ce5b78, 32'shc6cda708, 32'shc6ccf2a1, 32'shc6cc3e42, 32'shc6cb89ed, 32'shc6cad5a0, 
               32'shc6ca215c, 32'shc6c96d21, 32'shc6c8b8ee, 32'shc6c804c5, 32'shc6c750a4, 32'shc6c69c8c, 32'shc6c5e87d, 32'shc6c53477, 
               32'shc6c4807a, 32'shc6c3cc85, 32'shc6c31899, 32'shc6c264b7, 32'shc6c1b0dd, 32'shc6c0fd0b, 32'shc6c04943, 32'shc6bf9583, 
               32'shc6bee1cd, 32'shc6be2e1f, 32'shc6bd7a7a, 32'shc6bcc6dd, 32'shc6bc134a, 32'shc6bb5fbf, 32'shc6baac3d, 32'shc6b9f8c5, 
               32'shc6b94554, 32'shc6b891ed, 32'shc6b7de8f, 32'shc6b72b39, 32'shc6b677ec, 32'shc6b5c4a8, 32'shc6b5116d, 32'shc6b45e3b, 
               32'shc6b3ab12, 32'shc6b2f7f1, 32'shc6b244d9, 32'shc6b191ca, 32'shc6b0dec4, 32'shc6b02bc7, 32'shc6af78d3, 32'shc6aec5e7, 
               32'shc6ae1304, 32'shc6ad602a, 32'shc6acad59, 32'shc6abfa91, 32'shc6ab47d2, 32'shc6aa951b, 32'shc6a9e26e, 32'shc6a92fc9, 
               32'shc6a87d2d, 32'shc6a7ca9a, 32'shc6a7180f, 32'shc6a6658e, 32'shc6a5b315, 32'shc6a500a5, 32'shc6a44e3e, 32'shc6a39be0, 
               32'shc6a2e98b, 32'shc6a2373f, 32'shc6a184fb, 32'shc6a0d2c0, 32'shc6a0208f, 32'shc69f6e66, 32'shc69ebc45, 32'shc69e0a2e, 
               32'shc69d5820, 32'shc69ca61a, 32'shc69bf41d, 32'shc69b4229, 32'shc69a903e, 32'shc699de5c, 32'shc6992c83, 32'shc6987ab2, 
               32'shc697c8eb, 32'shc697172c, 32'shc6966576, 32'shc695b3c9, 32'shc6950224, 32'shc6945089, 32'shc6939ef6, 32'shc692ed6d, 
               32'shc6923bec, 32'shc6918a74, 32'shc690d905, 32'shc690279f, 32'shc68f7641, 32'shc68ec4ed, 32'shc68e13a1, 32'shc68d625e, 
               32'shc68cb124, 32'shc68bfff3, 32'shc68b4ecb, 32'shc68a9dac, 32'shc689ec95, 32'shc6893b87, 32'shc6888a83, 32'shc687d987, 
               32'shc6872894, 32'shc68677a9, 32'shc685c6c8, 32'shc68515f0, 32'shc6846520, 32'shc683b459, 32'shc683039b, 32'shc68252e6, 
               32'shc681a23a, 32'shc680f197, 32'shc68040fc, 32'shc67f906b, 32'shc67edfe2, 32'shc67e2f62, 32'shc67d7eeb, 32'shc67cce7d, 
               32'shc67c1e18, 32'shc67b6dbc, 32'shc67abd68, 32'shc67a0d1e, 32'shc6795cdc, 32'shc678aca3, 32'shc677fc73, 32'shc6774c4c, 
               32'shc6769c2e, 32'shc675ec18, 32'shc6753c0c, 32'shc6748c08, 32'shc673dc0d, 32'shc6732c1b, 32'shc6727c32, 32'shc671cc52, 
               32'shc6711c7b, 32'shc6706cad, 32'shc66fbce7, 32'shc66f0d2b, 32'shc66e5d77, 32'shc66dadcc, 32'shc66cfe2a, 32'shc66c4e91, 
               32'shc66b9f01, 32'shc66aef79, 32'shc66a3ffb, 32'shc6699085, 32'shc668e119, 32'shc66831b5, 32'shc667825a, 32'shc666d308, 
               32'shc66623be, 32'shc665747e, 32'shc664c547, 32'shc6641618, 32'shc66366f3, 32'shc662b7d6, 32'shc66208c2, 32'shc66159b7, 
               32'shc660aab5, 32'shc65ffbbc, 32'shc65f4ccb, 32'shc65e9de4, 32'shc65def05, 32'shc65d4030, 32'shc65c9163, 32'shc65be29f, 
               32'shc65b33e4, 32'shc65a8532, 32'shc659d688, 32'shc65927e8, 32'shc6587951, 32'shc657cac2, 32'shc6571c3c, 32'shc6566dc0, 
               32'shc655bf4c, 32'shc65510e1, 32'shc654627f, 32'shc653b426, 32'shc65305d5, 32'shc652578e, 32'shc651a94f, 32'shc650fb1a, 
               32'shc6504ced, 32'shc64f9ec9, 32'shc64ef0ae, 32'shc64e429c, 32'shc64d9493, 32'shc64ce693, 32'shc64c389b, 32'shc64b8aad, 
               32'shc64adcc7, 32'shc64a2eeb, 32'shc6498117, 32'shc648d34c, 32'shc648258a, 32'shc64777d1, 32'shc646ca21, 32'shc6461c7a, 
               32'shc6456edb, 32'shc644c146, 32'shc64413b9, 32'shc6436636, 32'shc642b8bb, 32'shc6420b49, 32'shc6415de0, 32'shc640b080, 
               32'shc6400329, 32'shc63f55db, 32'shc63ea896, 32'shc63dfb59, 32'shc63d4e26, 32'shc63ca0fb, 32'shc63bf3d9, 32'shc63b46c1, 
               32'shc63a99b1, 32'shc639ecaa, 32'shc6393fac, 32'shc63892b7, 32'shc637e5ca, 32'shc63738e7, 32'shc6368c0d, 32'shc635df3b, 
               32'shc6353273, 32'shc63485b3, 32'shc633d8fc, 32'shc6332c4e, 32'shc6327faa, 32'shc631d30e, 32'shc631267a, 32'shc63079f0, 
               32'shc62fcd6f, 32'shc62f20f7, 32'shc62e7487, 32'shc62dc821, 32'shc62d1bc3, 32'shc62c6f6e, 32'shc62bc323, 32'shc62b16e0, 
               32'shc62a6aa6, 32'shc629be75, 32'shc629124d, 32'shc628662e, 32'shc627ba17, 32'shc6270e0a, 32'shc6266206, 32'shc625b60a, 
               32'shc6250a18, 32'shc6245e2e, 32'shc623b24d, 32'shc6230675, 32'shc6225aa6, 32'shc621aee1, 32'shc6210323, 32'shc620576f, 
               32'shc61fabc4, 32'shc61f0022, 32'shc61e5489, 32'shc61da8f8, 32'shc61cfd71, 32'shc61c51f2, 32'shc61ba67d, 32'shc61afb10, 
               32'shc61a4fac, 32'shc619a451, 32'shc618f8ff, 32'shc6184db6, 32'shc617a276, 32'shc616f73f, 32'shc6164c11, 32'shc615a0ec, 
               32'shc614f5cf, 32'shc6144abc, 32'shc6139fb2, 32'shc612f4b0, 32'shc61249b7, 32'shc6119ec8, 32'shc610f3e1, 32'shc6104903, 
               32'shc60f9e2e, 32'shc60ef362, 32'shc60e489f, 32'shc60d9de5, 32'shc60cf334, 32'shc60c488c, 32'shc60b9ded, 32'shc60af357, 
               32'shc60a48c9, 32'shc6099e45, 32'shc608f3c9, 32'shc6084957, 32'shc6079eed, 32'shc606f48c, 32'shc6064a35, 32'shc6059fe6, 
               32'shc604f5a0, 32'shc6044b63, 32'shc603a12f, 32'shc602f704, 32'shc6024ce2, 32'shc601a2c9, 32'shc600f8b9, 32'shc6004eb1, 
               32'shc5ffa4b3, 32'shc5fefabe, 32'shc5fe50d1, 32'shc5fda6ee, 32'shc5fcfd13, 32'shc5fc5342, 32'shc5fba979, 32'shc5faffb9, 
               32'shc5fa5603, 32'shc5f9ac55, 32'shc5f902b0, 32'shc5f85914, 32'shc5f7af81, 32'shc5f705f7, 32'shc5f65c76, 32'shc5f5b2fe, 
               32'shc5f5098f, 32'shc5f46029, 32'shc5f3b6cb, 32'shc5f30d77, 32'shc5f2642c, 32'shc5f1bae9, 32'shc5f111b0, 32'shc5f0687f, 
               32'shc5efbf58, 32'shc5ef1639, 32'shc5ee6d24, 32'shc5edc417, 32'shc5ed1b13, 32'shc5ec7218, 32'shc5ebc927, 32'shc5eb203e, 
               32'shc5ea775e, 32'shc5e9ce87, 32'shc5e925b9, 32'shc5e87cf4, 32'shc5e7d438, 32'shc5e72b85, 32'shc5e682db, 32'shc5e5da3a, 
               32'shc5e531a1, 32'shc5e48912, 32'shc5e3e08c, 32'shc5e3380e, 32'shc5e28f9a, 32'shc5e1e72f, 32'shc5e13ecc, 32'shc5e09673, 
               32'shc5dfee22, 32'shc5df45db, 32'shc5de9d9c, 32'shc5ddf566, 32'shc5dd4d3a, 32'shc5dca516, 32'shc5dbfcfb, 32'shc5db54e9, 
               32'shc5daace1, 32'shc5da04e1, 32'shc5d95cea, 32'shc5d8b4fc, 32'shc5d80d17, 32'shc5d7653b, 32'shc5d6bd68, 32'shc5d6159e, 
               32'shc5d56ddd, 32'shc5d4c625, 32'shc5d41e76, 32'shc5d376d0, 32'shc5d2cf33, 32'shc5d2279e, 32'shc5d18013, 32'shc5d0d891, 
               32'shc5d03118, 32'shc5cf89a7, 32'shc5cee240, 32'shc5ce3ae1, 32'shc5cd938c, 32'shc5ccec40, 32'shc5cc44fc, 32'shc5cb9dc2, 
               32'shc5caf690, 32'shc5ca4f68, 32'shc5c9a848, 32'shc5c90132, 32'shc5c85a24, 32'shc5c7b31f, 32'shc5c70c24, 32'shc5c66531, 
               32'shc5c5be47, 32'shc5c51767, 32'shc5c4708f, 32'shc5c3c9c0, 32'shc5c322fb, 32'shc5c27c3e, 32'shc5c1d58a, 32'shc5c12edf, 
               32'shc5c0883d, 32'shc5bfe1a5, 32'shc5bf3b15, 32'shc5be948e, 32'shc5bdee10, 32'shc5bd479b, 32'shc5bca12f, 32'shc5bbfacc, 
               32'shc5bb5472, 32'shc5baae21, 32'shc5ba07d9, 32'shc5b9619a, 32'shc5b8bb64, 32'shc5b81537, 32'shc5b76f13, 32'shc5b6c8f8, 
               32'shc5b622e6, 32'shc5b57cdd, 32'shc5b4d6dd, 32'shc5b430e6, 32'shc5b38af8, 32'shc5b2e513, 32'shc5b23f37, 32'shc5b19963, 
               32'shc5b0f399, 32'shc5b04dd8, 32'shc5afa820, 32'shc5af0271, 32'shc5ae5ccb, 32'shc5adb72d, 32'shc5ad1199, 32'shc5ac6c0e, 
               32'shc5abc68c, 32'shc5ab2113, 32'shc5aa7ba3, 32'shc5a9d63b, 32'shc5a930dd, 32'shc5a88b88, 32'shc5a7e63c, 32'shc5a740f8, 
               32'shc5a69bbe, 32'shc5a5f68d, 32'shc5a55165, 32'shc5a4ac46, 32'shc5a4072f, 32'shc5a36222, 32'shc5a2bd1e, 32'shc5a21823, 
               32'shc5a17330, 32'shc5a0ce47, 32'shc5a02967, 32'shc59f8490, 32'shc59edfc2, 32'shc59e3afc, 32'shc59d9640, 32'shc59cf18d, 
               32'shc59c4ce3, 32'shc59ba842, 32'shc59b03a9, 32'shc59a5f1a, 32'shc599ba94, 32'shc5991617, 32'shc59871a3, 32'shc597cd38, 
               32'shc59728d5, 32'shc596847c, 32'shc595e02c, 32'shc5953be5, 32'shc59497a7, 32'shc593f372, 32'shc5934f46, 32'shc592ab22, 
               32'shc5920708, 32'shc59162f7, 32'shc590beef, 32'shc5901af0, 32'shc58f76fa, 32'shc58ed30d, 32'shc58e2f29, 32'shc58d8b4e, 
               32'shc58ce77c, 32'shc58c43b3, 32'shc58b9ff3, 32'shc58afc3c, 32'shc58a588e, 32'shc589b4e9, 32'shc589114e, 32'shc5886dbb, 
               32'shc587ca31, 32'shc58726b0, 32'shc5868338, 32'shc585dfc9, 32'shc5853c63, 32'shc5849907, 32'shc583f5b3, 32'shc5835268, 
               32'shc582af26, 32'shc5820bee, 32'shc58168be, 32'shc580c597, 32'shc580227a, 32'shc57f7f65, 32'shc57edc5a, 32'shc57e3957, 
               32'shc57d965d, 32'shc57cf36d, 32'shc57c5085, 32'shc57bada7, 32'shc57b0ad1, 32'shc57a6805, 32'shc579c542, 32'shc5792287, 
               32'shc5787fd6, 32'shc577dd2d, 32'shc5773a8e, 32'shc57697f8, 32'shc575f56b, 32'shc57552e6, 32'shc574b06b, 32'shc5740df9, 
               32'shc5736b90, 32'shc572c930, 32'shc57226d9, 32'shc571848b, 32'shc570e246, 32'shc570400a, 32'shc56f9dd7, 32'shc56efbad, 
               32'shc56e598c, 32'shc56db774, 32'shc56d1565, 32'shc56c735f, 32'shc56bd163, 32'shc56b2f6f, 32'shc56a8d84, 32'shc569eba2, 
               32'shc56949ca, 32'shc568a7fa, 32'shc5680634, 32'shc5676476, 32'shc566c2c2, 32'shc5662116, 32'shc5657f74, 32'shc564ddda, 
               32'shc5643c4a, 32'shc5639ac3, 32'shc562f944, 32'shc56257cf, 32'shc561b663, 32'shc5611500, 32'shc56073a6, 32'shc55fd255, 
               32'shc55f310d, 32'shc55e8fce, 32'shc55dee98, 32'shc55d4d6b, 32'shc55cac47, 32'shc55c0b2c, 32'shc55b6a1a, 32'shc55ac912, 
               32'shc55a2812, 32'shc559871b, 32'shc558e62e, 32'shc5584549, 32'shc557a46e, 32'shc557039b, 32'shc55662d2, 32'shc555c211, 
               32'shc555215a, 32'shc55480ac, 32'shc553e007, 32'shc5533f6b, 32'shc5529ed7, 32'shc551fe4d, 32'shc5515dcc, 32'shc550bd54, 
               32'shc5501ce5, 32'shc54f7c7f, 32'shc54edc23, 32'shc54e3bcf, 32'shc54d9b84, 32'shc54cfb42, 32'shc54c5b0a, 32'shc54bbada, 
               32'shc54b1ab4, 32'shc54a7a96, 32'shc549da82, 32'shc5493a76, 32'shc5489a74, 32'shc547fa7b, 32'shc5475a8b, 32'shc546baa4, 
               32'shc5461ac6, 32'shc5457af1, 32'shc544db25, 32'shc5443b62, 32'shc5439ba8, 32'shc542fbf7, 32'shc5425c4f, 32'shc541bcb1, 
               32'shc5411d1b, 32'shc5407d8e, 32'shc53fde0b, 32'shc53f3e90, 32'shc53e9f1f, 32'shc53dffb7, 32'shc53d6057, 32'shc53cc101, 
               32'shc53c21b4, 32'shc53b8270, 32'shc53ae335, 32'shc53a4403, 32'shc539a4da, 32'shc53905ba, 32'shc53866a4, 32'shc537c796, 
               32'shc5372891, 32'shc5368996, 32'shc535eaa3, 32'shc5354bba, 32'shc534acd9, 32'shc5340e02, 32'shc5336f34, 32'shc532d06f, 
               32'shc53231b3, 32'shc5319300, 32'shc530f456, 32'shc53055b5, 32'shc52fb71d, 32'shc52f188e, 32'shc52e7a09, 32'shc52ddb8c, 
               32'shc52d3d18, 32'shc52c9eae, 32'shc52c004d, 32'shc52b61f4, 32'shc52ac3a5, 32'shc52a255f, 32'shc5298722, 32'shc528e8ee, 
               32'shc5284ac3, 32'shc527aca1, 32'shc5270e88, 32'shc5267078, 32'shc525d272, 32'shc5253474, 32'shc5249680, 32'shc523f894, 
               32'shc5235ab2, 32'shc522bcd9, 32'shc5221f08, 32'shc5218141, 32'shc520e383, 32'shc52045ce, 32'shc51fa822, 32'shc51f0a7f, 
               32'shc51e6ce6, 32'shc51dcf55, 32'shc51d31ce, 32'shc51c944f, 32'shc51bf6da, 32'shc51b596d, 32'shc51abc0a, 32'shc51a1eb0, 
               32'shc519815f, 32'shc518e417, 32'shc51846d8, 32'shc517a9a2, 32'shc5170c75, 32'shc5166f52, 32'shc515d237, 32'shc5153526, 
               32'shc514981d, 32'shc513fb1e, 32'shc5135e28, 32'shc512c13b, 32'shc5122457, 32'shc511877c, 32'shc510eaaa, 32'shc5104de1, 
               32'shc50fb121, 32'shc50f146b, 32'shc50e77bd, 32'shc50ddb19, 32'shc50d3e7d, 32'shc50ca1eb, 32'shc50c0562, 32'shc50b68e2, 
               32'shc50acc6b, 32'shc50a2ffd, 32'shc5099398, 32'shc508f73d, 32'shc5085aea, 32'shc507bea1, 32'shc5072260, 32'shc5068629, 
               32'shc505e9fb, 32'shc5054dd5, 32'shc504b1b9, 32'shc50415a6, 32'shc503799d, 32'shc502dd9c, 32'shc50241a4, 32'shc501a5b6, 
               32'shc50109d0, 32'shc5006df4, 32'shc4ffd221, 32'shc4ff3656, 32'shc4fe9a95, 32'shc4fdfedd, 32'shc4fd632f, 32'shc4fcc789, 
               32'shc4fc2bec, 32'shc4fb9059, 32'shc4faf4ce, 32'shc4fa594d, 32'shc4f9bdd4, 32'shc4f92265, 32'shc4f886ff, 32'shc4f7eba2, 
               32'shc4f7504e, 32'shc4f6b504, 32'shc4f619c2, 32'shc4f57e8a, 32'shc4f4e35a, 32'shc4f44834, 32'shc4f3ad17, 32'shc4f31202, 
               32'shc4f276f7, 32'shc4f1dbf6, 32'shc4f140fd, 32'shc4f0a60d, 32'shc4f00b27, 32'shc4ef7049, 32'shc4eed575, 32'shc4ee3aa9, 
               32'shc4ed9fe7, 32'shc4ed052e, 32'shc4ec6a7e, 32'shc4ebcfd8, 32'shc4eb353a, 32'shc4ea9aa5, 32'shc4ea001a, 32'shc4e96597, 
               32'shc4e8cb1e, 32'shc4e830ae, 32'shc4e79647, 32'shc4e6fbe9, 32'shc4e66194, 32'shc4e5c749, 32'shc4e52d06, 32'shc4e492cd, 
               32'shc4e3f89c, 32'shc4e35e75, 32'shc4e2c457, 32'shc4e22a42, 32'shc4e19036, 32'shc4e0f633, 32'shc4e05c3a, 32'shc4dfc249, 
               32'shc4df2862, 32'shc4de8e83, 32'shc4ddf4ae, 32'shc4dd5ae2, 32'shc4dcc11f, 32'shc4dc2765, 32'shc4db8db5, 32'shc4daf40d, 
               32'shc4da5a6f, 32'shc4d9c0d9, 32'shc4d9274d, 32'shc4d88dca, 32'shc4d7f450, 32'shc4d75adf, 32'shc4d6c177, 32'shc4d62819, 
               32'shc4d58ec3, 32'shc4d4f577, 32'shc4d45c34, 32'shc4d3c2fa, 32'shc4d329c9, 32'shc4d290a1, 32'shc4d1f782, 32'shc4d15e6d, 
               32'shc4d0c560, 32'shc4d02c5d, 32'shc4cf9363, 32'shc4cefa71, 32'shc4ce6189, 32'shc4cdc8ab, 32'shc4cd2fd5, 32'shc4cc9708, 
               32'shc4cbfe45, 32'shc4cb658b, 32'shc4caccd9, 32'shc4ca3431, 32'shc4c99b92, 32'shc4c902fd, 32'shc4c86a70, 32'shc4c7d1ec, 
               32'shc4c73972, 32'shc4c6a101, 32'shc4c60899, 32'shc4c5703a, 32'shc4c4d7e4, 32'shc4c43f97, 32'shc4c3a753, 32'shc4c30f19, 
               32'shc4c276e8, 32'shc4c1dec0, 32'shc4c146a0, 32'shc4c0ae8b, 32'shc4c0167e, 32'shc4bf7e7a, 32'shc4bee680, 32'shc4be4e8e, 
               32'shc4bdb6a6, 32'shc4bd1ec7, 32'shc4bc86f1, 32'shc4bbef24, 32'shc4bb5760, 32'shc4babfa6, 32'shc4ba27f5, 32'shc4b9904c, 
               32'shc4b8f8ad, 32'shc4b86117, 32'shc4b7c98a, 32'shc4b73207, 32'shc4b69a8c, 32'shc4b6031b, 32'shc4b56bb3, 32'shc4b4d453, 
               32'shc4b43cfd, 32'shc4b3a5b1, 32'shc4b30e6d, 32'shc4b27732, 32'shc4b1e001, 32'shc4b148d9, 32'shc4b0b1ba, 32'shc4b01aa4, 
               32'shc4af8397, 32'shc4aeec93, 32'shc4ae5599, 32'shc4adbea7, 32'shc4ad27bf, 32'shc4ac90e0, 32'shc4abfa0a, 32'shc4ab633d, 
               32'shc4aacc7a, 32'shc4aa35bf, 32'shc4a99f0e, 32'shc4a90866, 32'shc4a871c7, 32'shc4a7db31, 32'shc4a744a4, 32'shc4a6ae21, 
               32'shc4a617a6, 32'shc4a58135, 32'shc4a4eacd, 32'shc4a4546e, 32'shc4a3be18, 32'shc4a327cb, 32'shc4a29188, 32'shc4a1fb4e, 
               32'shc4a1651c, 32'shc4a0cef4, 32'shc4a038d6, 32'shc49fa2c0, 32'shc49f0cb3, 32'shc49e76b0, 32'shc49de0b6, 32'shc49d4ac5, 
               32'shc49cb4dd, 32'shc49c1efe, 32'shc49b8928, 32'shc49af35c, 32'shc49a5d98, 32'shc499c7de, 32'shc499322d, 32'shc4989c86, 
               32'shc49806e7, 32'shc4977151, 32'shc496dbc5, 32'shc4964642, 32'shc495b0c8, 32'shc4951b57, 32'shc49485ef, 32'shc493f091, 
               32'shc4935b3c, 32'shc492c5ef, 32'shc49230ac, 32'shc4919b72, 32'shc4910642, 32'shc490711a, 32'shc48fdbfc, 32'shc48f46e7, 
               32'shc48eb1db, 32'shc48e1cd8, 32'shc48d87de, 32'shc48cf2ee, 32'shc48c5e06, 32'shc48bc928, 32'shc48b3453, 32'shc48a9f87, 
               32'shc48a0ac4, 32'shc489760b, 32'shc488e15b, 32'shc4884cb3, 32'shc487b815, 32'shc4872381, 32'shc4868ef5, 32'shc485fa72, 
               32'shc48565f9, 32'shc484d189, 32'shc4843d22, 32'shc483a8c4, 32'shc4831470, 32'shc4828024, 32'shc481ebe2, 32'shc48157a9, 
               32'shc480c379, 32'shc4802f52, 32'shc47f9b34, 32'shc47f0720, 32'shc47e7315, 32'shc47ddf13, 32'shc47d4b1a, 32'shc47cb72a, 
               32'shc47c2344, 32'shc47b8f66, 32'shc47afb92, 32'shc47a67c7, 32'shc479d405, 32'shc479404d, 32'shc478ac9d, 32'shc47818f7, 
               32'shc477855a, 32'shc476f1c6, 32'shc4765e3b, 32'shc475caba, 32'shc4753741, 32'shc474a3d2, 32'shc474106c, 32'shc4737d10, 
               32'shc472e9bc, 32'shc4725671, 32'shc471c330, 32'shc4712ff8, 32'shc4709cc9, 32'shc47009a4, 32'shc46f7687, 32'shc46ee374, 
               32'shc46e5069, 32'shc46dbd69, 32'shc46d2a71, 32'shc46c9782, 32'shc46c049d, 32'shc46b71c1, 32'shc46adeee, 32'shc46a4c24, 
               32'shc469b963, 32'shc46926ac, 32'shc46893fd, 32'shc4680158, 32'shc4676ebc, 32'shc466dc2a, 32'shc46649a0, 32'shc465b720, 
               32'shc46524a9, 32'shc464923b, 32'shc463ffd6, 32'shc4636d7a, 32'shc462db28, 32'shc46248df, 32'shc461b69f, 32'shc4612468, 
               32'shc460923b, 32'shc4600016, 32'shc45f6dfb, 32'shc45edbe9, 32'shc45e49e0, 32'shc45db7e1, 32'shc45d25ea, 32'shc45c93fd, 
               32'shc45c0219, 32'shc45b703e, 32'shc45ade6c, 32'shc45a4ca4, 32'shc459bae5, 32'shc459292f, 32'shc4589782, 32'shc45805de, 
               32'shc4577444, 32'shc456e2b3, 32'shc456512b, 32'shc455bfac, 32'shc4552e36, 32'shc4549cca, 32'shc4540b67, 32'shc4537a0d, 
               32'shc452e8bc, 32'shc4525774, 32'shc451c636, 32'shc4513500, 32'shc450a3d4, 32'shc45012b2, 32'shc44f8198, 32'shc44ef088, 
               32'shc44e5f80, 32'shc44dce82, 32'shc44d3d8e, 32'shc44caca2, 32'shc44c1bc0, 32'shc44b8ae7, 32'shc44afa17, 32'shc44a6950, 
               32'shc449d892, 32'shc44947de, 32'shc448b733, 32'shc4482691, 32'shc44795f8, 32'shc4470569, 32'shc44674e3, 32'shc445e466, 
               32'shc44553f2, 32'shc444c387, 32'shc4443326, 32'shc443a2cd, 32'shc443127e, 32'shc4428239, 32'shc441f1fc, 32'shc44161c9, 
               32'shc440d19e, 32'shc440417d, 32'shc43fb166, 32'shc43f2157, 32'shc43e9152, 32'shc43e0156, 32'shc43d7163, 32'shc43ce179, 
               32'shc43c5199, 32'shc43bc1c2, 32'shc43b31f4, 32'shc43aa22f, 32'shc43a1273, 32'shc43982c1, 32'shc438f318, 32'shc4386378, 
               32'shc437d3e1, 32'shc4374454, 32'shc436b4cf, 32'shc4362554, 32'shc43595e3, 32'shc435067a, 32'shc434771b, 32'shc433e7c4, 
               32'shc4335877, 32'shc432c934, 32'shc43239f9, 32'shc431aac8, 32'shc4311ba0, 32'shc4308c81, 32'shc42ffd6b, 32'shc42f6e5f, 
               32'shc42edf5c, 32'shc42e5062, 32'shc42dc171, 32'shc42d328a, 32'shc42ca3ac, 32'shc42c14d7, 32'shc42b860b, 32'shc42af748, 
               32'shc42a688f, 32'shc429d9df, 32'shc4294b38, 32'shc428bc9a, 32'shc4282e06, 32'shc4279f7b, 32'shc42710f9, 32'shc4268280, 
               32'shc425f410, 32'shc42565aa, 32'shc424d74d, 32'shc42448f9, 32'shc423baae, 32'shc4232c6d, 32'shc4229e35, 32'shc4221006, 
               32'shc42181e0, 32'shc420f3c4, 32'shc42065b1, 32'shc41fd7a7, 32'shc41f49a6, 32'shc41ebbaf, 32'shc41e2dc0, 32'shc41d9fdb, 
               32'shc41d11ff, 32'shc41c842d, 32'shc41bf664, 32'shc41b68a3, 32'shc41adaed, 32'shc41a4d3f, 32'shc419bf9b, 32'shc41931ff, 
               32'shc418a46d, 32'shc41816e5, 32'shc4178965, 32'shc416fbef, 32'shc4166e82, 32'shc415e11f, 32'shc41553c4, 32'shc414c673, 
               32'shc414392b, 32'shc413abec, 32'shc4131eb7, 32'shc412918a, 32'shc4120467, 32'shc411774d, 32'shc410ea3d, 32'shc4105d36, 
               32'shc40fd037, 32'shc40f4343, 32'shc40eb657, 32'shc40e2975, 32'shc40d9c9c, 32'shc40d0fcc, 32'shc40c8305, 32'shc40bf648, 
               32'shc40b6994, 32'shc40adce9, 32'shc40a5047, 32'shc409c3af, 32'shc4093720, 32'shc408aa9a, 32'shc4081e1d, 32'shc40791aa, 
               32'shc4070540, 32'shc40678df, 32'shc405ec87, 32'shc4056039, 32'shc404d3f4, 32'shc40447b8, 32'shc403bb85, 32'shc4032f5c, 
               32'shc402a33c, 32'shc4021725, 32'shc4018b17, 32'shc400ff13, 32'shc4007318, 32'shc3ffe726, 32'shc3ff5b3d, 32'shc3fecf5e, 
               32'shc3fe4388, 32'shc3fdb7bb, 32'shc3fd2bf7, 32'shc3fca03d, 32'shc3fc148c, 32'shc3fb88e4, 32'shc3fafd45, 32'shc3fa71b0, 
               32'shc3f9e624, 32'shc3f95aa1, 32'shc3f8cf27, 32'shc3f843b7, 32'shc3f7b850, 32'shc3f72cf2, 32'shc3f6a19e, 32'shc3f61652, 
               32'shc3f58b10, 32'shc3f4ffd8, 32'shc3f474a8, 32'shc3f3e982, 32'shc3f35e65, 32'shc3f2d351, 32'shc3f24847, 32'shc3f1bd46, 
               32'shc3f1324e, 32'shc3f0a75f, 32'shc3f01c7a, 32'shc3ef919d, 32'shc3ef06cb, 32'shc3ee7c01, 32'shc3edf141, 32'shc3ed6689, 
               32'shc3ecdbdc, 32'shc3ec5137, 32'shc3ebc69c, 32'shc3eb3c0a, 32'shc3eab181, 32'shc3ea2701, 32'shc3e99c8b, 32'shc3e9121e, 
               32'shc3e887bb, 32'shc3e7fd60, 32'shc3e7730f, 32'shc3e6e8c7, 32'shc3e65e88, 32'shc3e5d453, 32'shc3e54a27, 32'shc3e4c004, 
               32'shc3e435ea, 32'shc3e3abda, 32'shc3e321d3, 32'shc3e297d5, 32'shc3e20de1, 32'shc3e183f6, 32'shc3e0fa14, 32'shc3e0703b, 
               32'shc3dfe66c, 32'shc3df5ca6, 32'shc3ded2e9, 32'shc3de4935, 32'shc3ddbf8b, 32'shc3dd35ea, 32'shc3dcac52, 32'shc3dc22c4, 
               32'shc3db993e, 32'shc3db0fc2, 32'shc3da8650, 32'shc3d9fce6, 32'shc3d97386, 32'shc3d8ea2f, 32'shc3d860e2, 32'shc3d7d79d, 
               32'shc3d74e62, 32'shc3d6c531, 32'shc3d63c08, 32'shc3d5b2e9, 32'shc3d529d3, 32'shc3d4a0c7, 32'shc3d417c3, 32'shc3d38ec9, 
               32'shc3d305d8, 32'shc3d27cf1, 32'shc3d1f413, 32'shc3d16b3e, 32'shc3d0e272, 32'shc3d059b0, 32'shc3cfd0f7, 32'shc3cf4847, 
               32'shc3cebfa0, 32'shc3ce3703, 32'shc3cdae6f, 32'shc3cd25e4, 32'shc3cc9d63, 32'shc3cc14eb, 32'shc3cb8c7c, 32'shc3cb0416, 
               32'shc3ca7bba, 32'shc3c9f367, 32'shc3c96b1e, 32'shc3c8e2dd, 32'shc3c85aa6, 32'shc3c7d278, 32'shc3c74a54, 32'shc3c6c238, 
               32'shc3c63a26, 32'shc3c5b21e, 32'shc3c52a1e, 32'shc3c4a228, 32'shc3c41a3b, 32'shc3c39258, 32'shc3c30a7e, 32'shc3c282ad, 
               32'shc3c1fae5, 32'shc3c17327, 32'shc3c0eb71, 32'shc3c063c6, 32'shc3bfdc23, 32'shc3bf548a, 32'shc3beccfa, 32'shc3be4573, 
               32'shc3bdbdf6, 32'shc3bd3682, 32'shc3bcaf17, 32'shc3bc27b6, 32'shc3bba05e, 32'shc3bb190f, 32'shc3ba91c9, 32'shc3ba0a8d, 
               32'shc3b9835a, 32'shc3b8fc30, 32'shc3b87510, 32'shc3b7edf9, 32'shc3b766eb, 32'shc3b6dfe6, 32'shc3b658eb, 32'shc3b5d1f9, 
               32'shc3b54b11, 32'shc3b4c431, 32'shc3b43d5b, 32'shc3b3b68f, 32'shc3b32fcb, 32'shc3b2a911, 32'shc3b22260, 32'shc3b19bb9, 
               32'shc3b1151b, 32'shc3b08e86, 32'shc3b007fa, 32'shc3af8178, 32'shc3aefaff, 32'shc3ae748f, 32'shc3adee28, 32'shc3ad67cb, 
               32'shc3ace178, 32'shc3ac5b2d, 32'shc3abd4ec, 32'shc3ab4eb4, 32'shc3aac885, 32'shc3aa4260, 32'shc3a9bc44, 32'shc3a93631, 
               32'shc3a8b028, 32'shc3a82a28, 32'shc3a7a431, 32'shc3a71e44, 32'shc3a6985f, 32'shc3a61285, 32'shc3a58cb3, 32'shc3a506eb, 
               32'shc3a4812c, 32'shc3a3fb76, 32'shc3a375ca, 32'shc3a2f027, 32'shc3a26a8d, 32'shc3a1e4fd, 32'shc3a15f76, 32'shc3a0d9f8, 
               32'shc3a05484, 32'shc39fcf18, 32'shc39f49b7, 32'shc39ec45e, 32'shc39e3f0f, 32'shc39db9c9, 32'shc39d348c, 32'shc39caf59, 
               32'shc39c2a2f, 32'shc39ba50e, 32'shc39b1ff7, 32'shc39a9ae9, 32'shc39a15e4, 32'shc39990e9, 32'shc3990bf7, 32'shc398870e, 
               32'shc398022f, 32'shc3977d59, 32'shc396f88c, 32'shc39673c8, 32'shc395ef0e, 32'shc3956a5d, 32'shc394e5b6, 32'shc3946117, 
               32'shc393dc82, 32'shc39357f7, 32'shc392d375, 32'shc3924efc, 32'shc391ca8c, 32'shc3914626, 32'shc390c1c9, 32'shc3903d75, 
               32'shc38fb92a, 32'shc38f34e9, 32'shc38eb0b2, 32'shc38e2c83, 32'shc38da85e, 32'shc38d2442, 32'shc38ca030, 32'shc38c1c27, 
               32'shc38b9827, 32'shc38b1431, 32'shc38a9043, 32'shc38a0c60, 32'shc3898885, 32'shc38904b4, 32'shc38880ec, 32'shc387fd2e, 
               32'shc3877978, 32'shc386f5cc, 32'shc386722a, 32'shc385ee91, 32'shc3856b01, 32'shc384e77a, 32'shc38463fd, 32'shc383e089, 
               32'shc3835d1e, 32'shc382d9bd, 32'shc3825665, 32'shc381d317, 32'shc3814fd1, 32'shc380cc95, 32'shc3804963, 32'shc37fc639, 
               32'shc37f4319, 32'shc37ec003, 32'shc37e3cf6, 32'shc37db9f2, 32'shc37d36f7, 32'shc37cb406, 32'shc37c311e, 32'shc37bae3f, 
               32'shc37b2b6a, 32'shc37aa89e, 32'shc37a25db, 32'shc379a322, 32'shc3792072, 32'shc3789dcb, 32'shc3781b2e, 32'shc377989a, 
               32'shc377160f, 32'shc376938e, 32'shc3761116, 32'shc3758ea7, 32'shc3750c42, 32'shc37489e6, 32'shc3740793, 32'shc373854a, 
               32'shc373030a, 32'shc37280d3, 32'shc371fea6, 32'shc3717c82, 32'shc370fa68, 32'shc3707856, 32'shc36ff64e, 32'shc36f7450, 
               32'shc36ef25b, 32'shc36e706f, 32'shc36dee8c, 32'shc36d6cb3, 32'shc36ceae3, 32'shc36c691d, 32'shc36be75f, 32'shc36b65ab, 
               32'shc36ae401, 32'shc36a6260, 32'shc369e0c8, 32'shc3695f3a, 32'shc368ddb4, 32'shc3685c39, 32'shc367dac6, 32'shc367595d, 
               32'shc366d7fd, 32'shc36656a7, 32'shc365d55a, 32'shc3655416, 32'shc364d2dc, 32'shc36451ab, 32'shc363d083, 32'shc3634f65, 
               32'shc362ce50, 32'shc3624d44, 32'shc361cc42, 32'shc3614b49, 32'shc360ca59, 32'shc3604973, 32'shc35fc896, 32'shc35f47c2, 
               32'shc35ec6f8, 32'shc35e4637, 32'shc35dc580, 32'shc35d44d2, 32'shc35cc42d, 32'shc35c4391, 32'shc35bc2ff, 32'shc35b4277, 
               32'shc35ac1f7, 32'shc35a4181, 32'shc359c114, 32'shc35940b1, 32'shc358c057, 32'shc3584006, 32'shc357bfbf, 32'shc3573f81, 
               32'shc356bf4d, 32'shc3563f21, 32'shc355bf00, 32'shc3553ee7, 32'shc354bed8, 32'shc3543ed2, 32'shc353bed6, 32'shc3533ee3, 
               32'shc352bef9, 32'shc3523f18, 32'shc351bf41, 32'shc3513f74, 32'shc350bfaf, 32'shc3503ff5, 32'shc34fc043, 32'shc34f409b, 
               32'shc34ec0fc, 32'shc34e4166, 32'shc34dc1da, 32'shc34d4257, 32'shc34cc2de, 32'shc34c436e, 32'shc34bc407, 32'shc34b44aa, 
               32'shc34ac556, 32'shc34a460b, 32'shc349c6ca, 32'shc3494792, 32'shc348c864, 32'shc348493f, 32'shc347ca23, 32'shc3474b10, 
               32'shc346cc07, 32'shc3464d07, 32'shc345ce11, 32'shc3454f24, 32'shc344d041, 32'shc3445166, 32'shc343d295, 32'shc34353ce, 
               32'shc342d510, 32'shc342565b, 32'shc341d7b0, 32'shc341590e, 32'shc340da75, 32'shc3405be6, 32'shc33fdd60, 32'shc33f5ee3, 
               32'shc33ee070, 32'shc33e6206, 32'shc33de3a5, 32'shc33d654e, 32'shc33ce701, 32'shc33c68bc, 32'shc33bea81, 32'shc33b6c50, 
               32'shc33aee27, 32'shc33a7009, 32'shc339f1f3, 32'shc33973e7, 32'shc338f5e4, 32'shc33877eb, 32'shc337f9fb, 32'shc3377c14, 
               32'shc336fe37, 32'shc3368063, 32'shc3360298, 32'shc33584d7, 32'shc3350720, 32'shc3348971, 32'shc3340bcc, 32'shc3338e30, 
               32'shc333109e, 32'shc3329315, 32'shc3321596, 32'shc3319820, 32'shc3311ab3, 32'shc3309d50, 32'shc3301ff5, 32'shc32fa2a5, 
               32'shc32f255e, 32'shc32ea820, 32'shc32e2aeb, 32'shc32dadc0, 32'shc32d309e, 32'shc32cb386, 32'shc32c3677, 32'shc32bb971, 
               32'shc32b3c75, 32'shc32abf82, 32'shc32a4299, 32'shc329c5b9, 32'shc32948e2, 32'shc328cc15, 32'shc3284f51, 32'shc327d296, 
               32'shc32755e5, 32'shc326d93e, 32'shc3265c9f, 32'shc325e00a, 32'shc325637f, 32'shc324e6fc, 32'shc3246a83, 32'shc323ee14, 
               32'shc32371ae, 32'shc322f551, 32'shc32278fe, 32'shc321fcb4, 32'shc3218073, 32'shc321043c, 32'shc320880e, 32'shc3200bea, 
               32'shc31f8fcf, 32'shc31f13bd, 32'shc31e97b5, 32'shc31e1bb6, 32'shc31d9fc1, 32'shc31d23d5, 32'shc31ca7f2, 32'shc31c2c19, 
               32'shc31bb049, 32'shc31b3483, 32'shc31ab8c6, 32'shc31a3d12, 32'shc319c168, 32'shc31945c7, 32'shc318ca2f, 32'shc3184ea1, 
               32'shc317d31c, 32'shc31757a1, 32'shc316dc2f, 32'shc31660c6, 32'shc315e567, 32'shc3156a11, 32'shc314eec5, 32'shc3147382, 
               32'shc313f848, 32'shc3137d18, 32'shc31301f1, 32'shc31286d4, 32'shc3120bc0, 32'shc31190b5, 32'shc31115b4, 32'shc3109abc, 
               32'shc3101fce, 32'shc30fa4e9, 32'shc30f2a0d, 32'shc30eaf3b, 32'shc30e3472, 32'shc30db9b3, 32'shc30d3efd, 32'shc30cc450, 
               32'shc30c49ad, 32'shc30bcf13, 32'shc30b5482, 32'shc30ad9fb, 32'shc30a5f7e, 32'shc309e509, 32'shc3096a9f, 32'shc308f03d, 
               32'shc30875e5, 32'shc307fb97, 32'shc3078151, 32'shc3070715, 32'shc3068ce3, 32'shc30612ba, 32'shc305989a, 32'shc3051e84, 
               32'shc304a477, 32'shc3042a74, 32'shc303b07a, 32'shc3033689, 32'shc302bca2, 32'shc30242c4, 32'shc301c8f0, 32'shc3014f25, 
               32'shc300d563, 32'shc3005bab, 32'shc2ffe1fc, 32'shc2ff6857, 32'shc2feeebb, 32'shc2fe7529, 32'shc2fdfb9f, 32'shc2fd8220, 
               32'shc2fd08a9, 32'shc2fc8f3c, 32'shc2fc15d9, 32'shc2fb9c7f, 32'shc2fb232e, 32'shc2faa9e7, 32'shc2fa30a9, 32'shc2f9b775, 
               32'shc2f93e4a, 32'shc2f8c528, 32'shc2f84c10, 32'shc2f7d301, 32'shc2f759fc, 32'shc2f6e100, 32'shc2f6680d, 32'shc2f5ef24, 
               32'shc2f57644, 32'shc2f4fd6e, 32'shc2f484a1, 32'shc2f40bdd, 32'shc2f39323, 32'shc2f31a73, 32'shc2f2a1cb, 32'shc2f2292e, 
               32'shc2f1b099, 32'shc2f1380e, 32'shc2f0bf8c, 32'shc2f04714, 32'shc2efcea6, 32'shc2ef5640, 32'shc2eedde4, 32'shc2ee6592, 
               32'shc2eded49, 32'shc2ed7509, 32'shc2ecfcd3, 32'shc2ec84a6, 32'shc2ec0c82, 32'shc2eb9468, 32'shc2eb1c58, 32'shc2eaa451, 
               32'shc2ea2c53, 32'shc2e9b45f, 32'shc2e93c74, 32'shc2e8c492, 32'shc2e84cba, 32'shc2e7d4ec, 32'shc2e75d26, 32'shc2e6e56b, 
               32'shc2e66db8, 32'shc2e5f60f, 32'shc2e57e70, 32'shc2e506da, 32'shc2e48f4d, 32'shc2e417ca, 32'shc2e3a050, 32'shc2e328df, 
               32'shc2e2b178, 32'shc2e23a1b, 32'shc2e1c2c7, 32'shc2e14b7c, 32'shc2e0d43b, 32'shc2e05d03, 32'shc2dfe5d4, 32'shc2df6eaf, 
               32'shc2def794, 32'shc2de8082, 32'shc2de0979, 32'shc2dd927a, 32'shc2dd1b84, 32'shc2dca497, 32'shc2dc2db4, 32'shc2dbb6db, 
               32'shc2db400a, 32'shc2dac944, 32'shc2da5286, 32'shc2d9dbd3, 32'shc2d96528, 32'shc2d8ee87, 32'shc2d877f0, 32'shc2d80161, 
               32'shc2d78add, 32'shc2d71461, 32'shc2d69df0, 32'shc2d62787, 32'shc2d5b128, 32'shc2d53ad3, 32'shc2d4c486, 32'shc2d44e44, 
               32'shc2d3d80a, 32'shc2d361db, 32'shc2d2ebb4, 32'shc2d27597, 32'shc2d1ff84, 32'shc2d1897a, 32'shc2d11379, 32'shc2d09d82, 
               32'shc2d02794, 32'shc2cfb1b0, 32'shc2cf3bd5, 32'shc2cec603, 32'shc2ce503b, 32'shc2cdda7d, 32'shc2cd64c7, 32'shc2ccef1c, 
               32'shc2cc7979, 32'shc2cc03e1, 32'shc2cb8e51, 32'shc2cb18cb, 32'shc2caa34f, 32'shc2ca2ddc, 32'shc2c9b872, 32'shc2c94312, 
               32'shc2c8cdbb, 32'shc2c8586e, 32'shc2c7e32a, 32'shc2c76def, 32'shc2c6f8be, 32'shc2c68397, 32'shc2c60e78, 32'shc2c59964, 
               32'shc2c52459, 32'shc2c4af57, 32'shc2c43a5e, 32'shc2c3c56f, 32'shc2c3508a, 32'shc2c2dbae, 32'shc2c266db, 32'shc2c1f212, 
               32'shc2c17d52, 32'shc2c1089c, 32'shc2c093ef, 32'shc2c01f4c, 32'shc2bfaab2, 32'shc2bf3622, 32'shc2bec19b, 32'shc2be4d1d, 
               32'shc2bdd8a9, 32'shc2bd643e, 32'shc2bcefdd, 32'shc2bc7b85, 32'shc2bc0737, 32'shc2bb92f2, 32'shc2bb1eb6, 32'shc2baaa84, 
               32'shc2ba365c, 32'shc2b9c23d, 32'shc2b94e27, 32'shc2b8da1b, 32'shc2b86618, 32'shc2b7f21f, 32'shc2b77e2f, 32'shc2b70a49, 
               32'shc2b6966c, 32'shc2b62298, 32'shc2b5aece, 32'shc2b53b0d, 32'shc2b4c756, 32'shc2b453a9, 32'shc2b3e004, 32'shc2b36c6a, 
               32'shc2b2f8d8, 32'shc2b28550, 32'shc2b211d2, 32'shc2b19e5d, 32'shc2b12af1, 32'shc2b0b78f, 32'shc2b04437, 32'shc2afd0e8, 
               32'shc2af5da2, 32'shc2aeea66, 32'shc2ae7733, 32'shc2ae0409, 32'shc2ad90ea, 32'shc2ad1dd3, 32'shc2acaac6, 32'shc2ac37c3, 
               32'shc2abc4c9, 32'shc2ab51d8, 32'shc2aadef1, 32'shc2aa6c13, 32'shc2a9f93f, 32'shc2a98674, 32'shc2a913b3, 32'shc2a8a0fb, 
               32'shc2a82e4d, 32'shc2a7bba8, 32'shc2a7490c, 32'shc2a6d67a, 32'shc2a663f2, 32'shc2a5f173, 32'shc2a57efd, 32'shc2a50c91, 
               32'shc2a49a2e, 32'shc2a427d5, 32'shc2a3b585, 32'shc2a3433f, 32'shc2a2d102, 32'shc2a25ecf, 32'shc2a1eca5, 32'shc2a17a84, 
               32'shc2a1086d, 32'shc2a09660, 32'shc2a0245c, 32'shc29fb261, 32'shc29f4070, 32'shc29ece88, 32'shc29e5caa, 32'shc29dead5, 
               32'shc29d790a, 32'shc29d0748, 32'shc29c9590, 32'shc29c23e1, 32'shc29bb23c, 32'shc29b40a0, 32'shc29acf0d, 32'shc29a5d84, 
               32'shc299ec05, 32'shc2997a8f, 32'shc2990922, 32'shc29897bf, 32'shc2982665, 32'shc297b515, 32'shc29743ce, 32'shc296d291, 
               32'shc296615d, 32'shc295f033, 32'shc2957f12, 32'shc2950dfb, 32'shc2949ced, 32'shc2942be8, 32'shc293baed, 32'shc29349fc, 
               32'shc292d914, 32'shc2926835, 32'shc291f760, 32'shc2918695, 32'shc29115d3, 32'shc290a51a, 32'shc290346b, 32'shc28fc3c5, 
               32'shc28f5329, 32'shc28ee296, 32'shc28e720d, 32'shc28e018d, 32'shc28d9117, 32'shc28d20aa, 32'shc28cb047, 32'shc28c3fed, 
               32'shc28bcf9c, 32'shc28b5f55, 32'shc28aef18, 32'shc28a7ee4, 32'shc28a0eb9, 32'shc2899e98, 32'shc2892e81, 32'shc288be73, 
               32'shc2884e6e, 32'shc287de73, 32'shc2876e82, 32'shc286fe99, 32'shc2868ebb, 32'shc2861ee6, 32'shc285af1a, 32'shc2853f58, 
               32'shc284cf9f, 32'shc2845ff0, 32'shc283f04a, 32'shc28380ad, 32'shc283111b, 32'shc282a191, 32'shc2823211, 32'shc281c29b, 
               32'shc281532e, 32'shc280e3cb, 32'shc2807471, 32'shc2800520, 32'shc27f95d9, 32'shc27f269c, 32'shc27eb768, 32'shc27e483d, 
               32'shc27dd91c, 32'shc27d6a05, 32'shc27cfaf7, 32'shc27c8bf2, 32'shc27c1cf7, 32'shc27bae06, 32'shc27b3f1e, 32'shc27ad03f, 
               32'shc27a616a, 32'shc279f29e, 32'shc27983dc, 32'shc2791523, 32'shc278a674, 32'shc27837ce, 32'shc277c932, 32'shc2775aa0, 
               32'shc276ec16, 32'shc2767d97, 32'shc2760f20, 32'shc275a0b4, 32'shc2753250, 32'shc274c3f7, 32'shc27455a6, 32'shc273e760, 
               32'shc2737922, 32'shc2730aee, 32'shc2729cc4, 32'shc2722ea3, 32'shc271c08c, 32'shc271527e, 32'shc270e47a, 32'shc270767f, 
               32'shc270088e, 32'shc26f9aa6, 32'shc26f2cc7, 32'shc26ebef2, 32'shc26e5127, 32'shc26de365, 32'shc26d75ad, 32'shc26d07fe, 
               32'shc26c9a58, 32'shc26c2cbd, 32'shc26bbf2a, 32'shc26b51a1, 32'shc26ae422, 32'shc26a76ac, 32'shc26a093f, 32'shc2699bdd, 
               32'shc2692e83, 32'shc268c133, 32'shc26853ed, 32'shc267e6b0, 32'shc267797c, 32'shc2670c52, 32'shc2669f32, 32'shc266321b, 
               32'shc265c50e, 32'shc265580a, 32'shc264eb0f, 32'shc2647e1e, 32'shc2641137, 32'shc263a459, 32'shc2633785, 32'shc262caba, 
               32'shc2625df8, 32'shc261f140, 32'shc2618492, 32'shc26117ed, 32'shc260ab51, 32'shc2603ec0, 32'shc25fd237, 32'shc25f65b8, 
               32'shc25ef943, 32'shc25e8cd7, 32'shc25e2074, 32'shc25db41c, 32'shc25d47cc, 32'shc25cdb86, 32'shc25c6f4a, 32'shc25c0317, 
               32'shc25b96ee, 32'shc25b2ace, 32'shc25abeb7, 32'shc25a52ab, 32'shc259e6a7, 32'shc2597aad, 32'shc2590ebd, 32'shc258a2d6, 
               32'shc25836f9, 32'shc257cb25, 32'shc2575f5b, 32'shc256f39a, 32'shc25687e3, 32'shc2561c35, 32'shc255b091, 32'shc25544f6, 
               32'shc254d965, 32'shc2546ddd, 32'shc254025f, 32'shc25396ea, 32'shc2532b7f, 32'shc252c01d, 32'shc25254c5, 32'shc251e976, 
               32'shc2517e31, 32'shc25112f6, 32'shc250a7c3, 32'shc2503c9b, 32'shc24fd17c, 32'shc24f6666, 32'shc24efb5a, 32'shc24e9057, 
               32'shc24e255e, 32'shc24dba6f, 32'shc24d4f89, 32'shc24ce4ac, 32'shc24c79d9, 32'shc24c0f10, 32'shc24ba450, 32'shc24b3999, 
               32'shc24aceed, 32'shc24a6449, 32'shc249f9af, 32'shc2498f1f, 32'shc2492498, 32'shc248ba1b, 32'shc2484fa7, 32'shc247e53c, 
               32'shc2477adc, 32'shc2471084, 32'shc246a637, 32'shc2463bf2, 32'shc245d1b8, 32'shc2456786, 32'shc244fd5f, 32'shc2449341, 
               32'shc244292c, 32'shc243bf21, 32'shc243551f, 32'shc242eb27, 32'shc2428139, 32'shc2421754, 32'shc241ad78, 32'shc24143a6, 
               32'shc240d9de, 32'shc240701f, 32'shc2400669, 32'shc23f9cbd, 32'shc23f331b, 32'shc23ec982, 32'shc23e5ff3, 32'shc23df66d, 
               32'shc23d8cf1, 32'shc23d237e, 32'shc23cba15, 32'shc23c50b5, 32'shc23be75f, 32'shc23b7e12, 32'shc23b14cf, 32'shc23aab95, 
               32'shc23a4265, 32'shc239d93f, 32'shc2397021, 32'shc239070e, 32'shc2389e04, 32'shc2383504, 32'shc237cc0d, 32'shc237631f, 
               32'shc236fa3b, 32'shc2369161, 32'shc2362890, 32'shc235bfc9, 32'shc235570b, 32'shc234ee57, 32'shc23485ac, 32'shc2341d0b, 
               32'shc233b473, 32'shc2334be5, 32'shc232e361, 32'shc2327ae6, 32'shc2321274, 32'shc231aa0c, 32'shc23141ae, 32'shc230d959, 
               32'shc230710d, 32'shc23008cb, 32'shc22fa093, 32'shc22f3864, 32'shc22ed03f, 32'shc22e6823, 32'shc22e0011, 32'shc22d9808, 
               32'shc22d3009, 32'shc22cc814, 32'shc22c6028, 32'shc22bf845, 32'shc22b906c, 32'shc22b289d, 32'shc22ac0d7, 32'shc22a591a, 
               32'shc229f167, 32'shc22989be, 32'shc229221e, 32'shc228ba88, 32'shc22852fb, 32'shc227eb78, 32'shc22783fe, 32'shc2271c8e, 
               32'shc226b528, 32'shc2264dcb, 32'shc225e677, 32'shc2257f2d, 32'shc22517ed, 32'shc224b0b6, 32'shc2244989, 32'shc223e265, 
               32'shc2237b4b, 32'shc223143a, 32'shc222ad33, 32'shc2224635, 32'shc221df41, 32'shc2217857, 32'shc2211176, 32'shc220aa9e, 
               32'shc22043d0, 32'shc21fdd0c, 32'shc21f7651, 32'shc21f0fa0, 32'shc21ea8f8, 32'shc21e425a, 32'shc21ddbc5, 32'shc21d753a, 
               32'shc21d0eb8, 32'shc21ca840, 32'shc21c41d2, 32'shc21bdb6d, 32'shc21b7511, 32'shc21b0ebf, 32'shc21aa877, 32'shc21a4238, 
               32'shc219dc03, 32'shc21975d7, 32'shc2190fb5, 32'shc218a99d, 32'shc218438e, 32'shc217dd88, 32'shc217778c, 32'shc217119a, 
               32'shc216abb1, 32'shc21645d2, 32'shc215dffc, 32'shc2157a30, 32'shc215146d, 32'shc214aeb4, 32'shc2144904, 32'shc213e35e, 
               32'shc2137dc2, 32'shc213182f, 32'shc212b2a5, 32'shc2124d26, 32'shc211e7af, 32'shc2118243, 32'shc2111cdf, 32'shc210b786, 
               32'shc2105236, 32'shc20fecef, 32'shc20f87b2, 32'shc20f227f, 32'shc20ebd55, 32'shc20e5835, 32'shc20df31e, 32'shc20d8e11, 
               32'shc20d290d, 32'shc20cc413, 32'shc20c5f22, 32'shc20bfa3b, 32'shc20b955e, 32'shc20b308a, 32'shc20acbc0, 32'shc20a66ff, 
               32'shc20a0248, 32'shc2099d9a, 32'shc20938f6, 32'shc208d45b, 32'shc2086fca, 32'shc2080b43, 32'shc207a6c5, 32'shc2074251, 
               32'shc206dde6, 32'shc2067985, 32'shc206152d, 32'shc205b0df, 32'shc2054c9b, 32'shc204e860, 32'shc204842e, 32'shc2042006, 
               32'shc203bbe8, 32'shc20357d3, 32'shc202f3c8, 32'shc2028fc6, 32'shc2022bce, 32'shc201c7e0, 32'shc20163fb, 32'shc201001f, 
               32'shc2009c4e, 32'shc2003885, 32'shc1ffd4c7, 32'shc1ff7111, 32'shc1ff0d66, 32'shc1fea9c4, 32'shc1fe462b, 32'shc1fde29c, 
               32'shc1fd7f17, 32'shc1fd1b9b, 32'shc1fcb829, 32'shc1fc54c0, 32'shc1fbf161, 32'shc1fb8e0c, 32'shc1fb2ac0, 32'shc1fac77e, 
               32'shc1fa6445, 32'shc1fa0115, 32'shc1f99df0, 32'shc1f93ad4, 32'shc1f8d7c1, 32'shc1f874b8, 32'shc1f811b9, 32'shc1f7aec3, 
               32'shc1f74bd6, 32'shc1f6e8f4, 32'shc1f6861a, 32'shc1f6234b, 32'shc1f5c085, 32'shc1f55dc8, 32'shc1f4fb15, 32'shc1f4986c, 
               32'shc1f435cc, 32'shc1f3d336, 32'shc1f370a9, 32'shc1f30e26, 32'shc1f2abad, 32'shc1f2493d, 32'shc1f1e6d7, 32'shc1f1847a, 
               32'shc1f12227, 32'shc1f0bfdd, 32'shc1f05d9d, 32'shc1effb66, 32'shc1ef9939, 32'shc1ef3716, 32'shc1eed4fc, 32'shc1ee72ec, 
               32'shc1ee10e5, 32'shc1edaee8, 32'shc1ed4cf5, 32'shc1eceb0b, 32'shc1ec892b, 32'shc1ec2754, 32'shc1ebc587, 32'shc1eb63c3, 
               32'shc1eb0209, 32'shc1eaa058, 32'shc1ea3eb1, 32'shc1e9dd14, 32'shc1e97b80, 32'shc1e919f6, 32'shc1e8b876, 32'shc1e856fe, 
               32'shc1e7f591, 32'shc1e7942d, 32'shc1e732d3, 32'shc1e6d182, 32'shc1e6703b, 32'shc1e60efd, 32'shc1e5adc9, 32'shc1e54c9f, 
               32'shc1e4eb7e, 32'shc1e48a67, 32'shc1e42959, 32'shc1e3c855, 32'shc1e3675a, 32'shc1e30669, 32'shc1e2a582, 32'shc1e244a4, 
               32'shc1e1e3d0, 32'shc1e18305, 32'shc1e12244, 32'shc1e0c18d, 32'shc1e060df, 32'shc1e0003a, 32'shc1df9fa0, 32'shc1df3f0f, 
               32'shc1dede87, 32'shc1de7e09, 32'shc1de1d94, 32'shc1ddbd2a, 32'shc1dd5cc8, 32'shc1dcfc71, 32'shc1dc9c23, 32'shc1dc3bde, 
               32'shc1dbdba3, 32'shc1db7b72, 32'shc1db1b4a, 32'shc1dabb2c, 32'shc1da5b17, 32'shc1d9fb0c, 32'shc1d99b0b, 32'shc1d93b13, 
               32'shc1d8db25, 32'shc1d87b40, 32'shc1d81b65, 32'shc1d7bb93, 32'shc1d75bcb, 32'shc1d6fc0d, 32'shc1d69c58, 32'shc1d63cad, 
               32'shc1d5dd0c, 32'shc1d57d74, 32'shc1d51de5, 32'shc1d4be60, 32'shc1d45ee5, 32'shc1d3ff73, 32'shc1d3a00b, 32'shc1d340ad, 
               32'shc1d2e158, 32'shc1d2820d, 32'shc1d222cb, 32'shc1d1c393, 32'shc1d16464, 32'shc1d1053f, 32'shc1d0a624, 32'shc1d04712, 
               32'shc1cfe80a, 32'shc1cf890c, 32'shc1cf2a17, 32'shc1cecb2b, 32'shc1ce6c49, 32'shc1ce0d71, 32'shc1cdaea3, 32'shc1cd4fde, 
               32'shc1ccf122, 32'shc1cc9270, 32'shc1cc33c8, 32'shc1cbd529, 32'shc1cb7694, 32'shc1cb1809, 32'shc1cab987, 32'shc1ca5b0f, 
               32'shc1c9fca0, 32'shc1c99e3b, 32'shc1c93fdf, 32'shc1c8e18d, 32'shc1c88345, 32'shc1c82506, 32'shc1c7c6d1, 32'shc1c768a6, 
               32'shc1c70a84, 32'shc1c6ac6b, 32'shc1c64e5d, 32'shc1c5f057, 32'shc1c5925c, 32'shc1c5346a, 32'shc1c4d682, 32'shc1c478a3, 
               32'shc1c41ace, 32'shc1c3bd02, 32'shc1c35f40, 32'shc1c30188, 32'shc1c2a3d9, 32'shc1c24634, 32'shc1c1e898, 32'shc1c18b06, 
               32'shc1c12d7e, 32'shc1c0cfff, 32'shc1c0728a, 32'shc1c0151e, 32'shc1bfb7bc, 32'shc1bf5a64, 32'shc1befd15, 32'shc1be9fd0, 
               32'shc1be4294, 32'shc1bde562, 32'shc1bd883a, 32'shc1bd2b1b, 32'shc1bcce06, 32'shc1bc70fa, 32'shc1bc13f8, 32'shc1bbb700, 
               32'shc1bb5a11, 32'shc1bafd2c, 32'shc1baa050, 32'shc1ba437e, 32'shc1b9e6b6, 32'shc1b989f7, 32'shc1b92d42, 32'shc1b8d097, 
               32'shc1b873f5, 32'shc1b8175c, 32'shc1b7bacd, 32'shc1b75e48, 32'shc1b701cd, 32'shc1b6a55b, 32'shc1b648f3, 32'shc1b5ec94, 
               32'shc1b5903f, 32'shc1b533f3, 32'shc1b4d7b1, 32'shc1b47b79, 32'shc1b41f4a, 32'shc1b3c325, 32'shc1b3670a, 32'shc1b30af8, 
               32'shc1b2aef0, 32'shc1b252f1, 32'shc1b1f6fc, 32'shc1b19b10, 32'shc1b13f2f, 32'shc1b0e356, 32'shc1b08788, 32'shc1b02bc3, 
               32'shc1afd007, 32'shc1af7456, 32'shc1af18ae, 32'shc1aebd0f, 32'shc1ae617a, 32'shc1ae05ef, 32'shc1adaa6d, 32'shc1ad4ef5, 
               32'shc1acf386, 32'shc1ac9821, 32'shc1ac3cc6, 32'shc1abe174, 32'shc1ab862c, 32'shc1ab2aee, 32'shc1aacfb9, 32'shc1aa748e, 
               32'shc1aa196c, 32'shc1a9be54, 32'shc1a96346, 32'shc1a90841, 32'shc1a8ad46, 32'shc1a85254, 32'shc1a7f76c, 32'shc1a79c8e, 
               32'shc1a741b9, 32'shc1a6e6ee, 32'shc1a68c2d, 32'shc1a63175, 32'shc1a5d6c7, 32'shc1a57c22, 32'shc1a52187, 32'shc1a4c6f6, 
               32'shc1a46c6e, 32'shc1a411f0, 32'shc1a3b77b, 32'shc1a35d10, 32'shc1a302af, 32'shc1a2a857, 32'shc1a24e09, 32'shc1a1f3c5, 
               32'shc1a1998a, 32'shc1a13f59, 32'shc1a0e531, 32'shc1a08b13, 32'shc1a030ff, 32'shc19fd6f4, 32'shc19f7cf3, 32'shc19f22fb, 
               32'shc19ec90d, 32'shc19e6f29, 32'shc19e154e, 32'shc19dbb7d, 32'shc19d61b6, 32'shc19d07f8, 32'shc19cae44, 32'shc19c549a, 
               32'shc19bfaf9, 32'shc19ba161, 32'shc19b47d4, 32'shc19aee50, 32'shc19a94d5, 32'shc19a3b64, 32'shc199e1fd, 32'shc199889f, 
               32'shc1992f4c, 32'shc198d601, 32'shc1987cc1, 32'shc1982389, 32'shc197ca5c, 32'shc1977138, 32'shc197181e, 32'shc196bf0d, 
               32'shc1966606, 32'shc1960d09, 32'shc195b415, 32'shc1955b2b, 32'shc195024b, 32'shc194a974, 32'shc19450a7, 32'shc193f7e3, 
               32'shc1939f29, 32'shc1934679, 32'shc192edd2, 32'shc1929535, 32'shc1923ca2, 32'shc191e418, 32'shc1918b98, 32'shc1913321, 
               32'shc190dab4, 32'shc1908251, 32'shc19029f7, 32'shc18fd1a7, 32'shc18f7961, 32'shc18f2124, 32'shc18ec8f1, 32'shc18e70c7, 
               32'shc18e18a7, 32'shc18dc091, 32'shc18d6884, 32'shc18d1081, 32'shc18cb888, 32'shc18c6098, 32'shc18c08b2, 32'shc18bb0d5, 
               32'shc18b5903, 32'shc18b0139, 32'shc18aa97a, 32'shc18a51c4, 32'shc189fa17, 32'shc189a275, 32'shc1894adc, 32'shc188f34c, 
               32'shc1889bc6, 32'shc188444a, 32'shc187ecd8, 32'shc187956f, 32'shc1873e10, 32'shc186e6ba, 32'shc1868f6e, 32'shc186382c, 
               32'shc185e0f3, 32'shc18589c4, 32'shc185329e, 32'shc184db82, 32'shc1848470, 32'shc1842d68, 32'shc183d669, 32'shc1837f73, 
               32'shc1832888, 32'shc182d1a6, 32'shc1827acd, 32'shc18223ff, 32'shc181cd3a, 32'shc181767e, 32'shc1811fcc, 32'shc180c924, 
               32'shc1807285, 32'shc1801bf1, 32'shc17fc565, 32'shc17f6ee4, 32'shc17f186c, 32'shc17ec1fd, 32'shc17e6b99, 32'shc17e153d, 
               32'shc17dbeec, 32'shc17d68a4, 32'shc17d1266, 32'shc17cbc32, 32'shc17c6607, 32'shc17c0fe5, 32'shc17bb9ce, 32'shc17b63c0, 
               32'shc17b0dbb, 32'shc17ab7c1, 32'shc17a61d0, 32'shc17a0be8, 32'shc179b60b, 32'shc1796036, 32'shc1790a6c, 32'shc178b4ab, 
               32'shc1785ef4, 32'shc1780946, 32'shc177b3a3, 32'shc1775e08, 32'shc1770878, 32'shc176b2f1, 32'shc1765d73, 32'shc1760800, 
               32'shc175b296, 32'shc1755d35, 32'shc17507df, 32'shc174b291, 32'shc1745d4e, 32'shc1740814, 32'shc173b2e4, 32'shc1735dbd, 
               32'shc17308a1, 32'shc172b38d, 32'shc1725e84, 32'shc1720984, 32'shc171b48e, 32'shc1715fa1, 32'shc1710abe, 32'shc170b5e5, 
               32'shc1706115, 32'shc1700c4f, 32'shc16fb792, 32'shc16f62e0, 32'shc16f0e36, 32'shc16eb997, 32'shc16e6501, 32'shc16e1075, 
               32'shc16dbbf3, 32'shc16d677a, 32'shc16d130a, 32'shc16cbea5, 32'shc16c6a49, 32'shc16c15f7, 32'shc16bc1ae, 32'shc16b6d6f, 
               32'shc16b193a, 32'shc16ac50e, 32'shc16a70ec, 32'shc16a1cd4, 32'shc169c8c5, 32'shc16974c0, 32'shc16920c5, 32'shc168ccd3, 
               32'shc16878eb, 32'shc168250c, 32'shc167d137, 32'shc1677d6c, 32'shc16729ab, 32'shc166d5f3, 32'shc1668245, 32'shc1662ea0, 
               32'shc165db05, 32'shc1658774, 32'shc16533ed, 32'shc164e06f, 32'shc1648cfa, 32'shc1643990, 32'shc163e62f, 32'shc16392d8, 
               32'shc1633f8a, 32'shc162ec46, 32'shc162990c, 32'shc16245db, 32'shc161f2b4, 32'shc1619f97, 32'shc1614c83, 32'shc160f979, 
               32'shc160a678, 32'shc1605382, 32'shc1600095, 32'shc15fadb1, 32'shc15f5ad7, 32'shc15f0807, 32'shc15eb541, 32'shc15e6284, 
               32'shc15e0fd1, 32'shc15dbd27, 32'shc15d6a88, 32'shc15d17f2, 32'shc15cc565, 32'shc15c72e2, 32'shc15c2069, 32'shc15bcdfa, 
               32'shc15b7b94, 32'shc15b2937, 32'shc15ad6e5, 32'shc15a849c, 32'shc15a325d, 32'shc159e027, 32'shc1598dfb, 32'shc1593bd9, 
               32'shc158e9c1, 32'shc15897b2, 32'shc15845ac, 32'shc157f3b1, 32'shc157a1bf, 32'shc1574fd7, 32'shc156fdf8, 32'shc156ac23, 
               32'shc1565a58, 32'shc1560896, 32'shc155b6de, 32'shc1556530, 32'shc155138c, 32'shc154c1f1, 32'shc154705f, 32'shc1541ed8, 
               32'shc153cd5a, 32'shc1537be5, 32'shc1532a7b, 32'shc152d91a, 32'shc15287c3, 32'shc1523675, 32'shc151e531, 32'shc15193f7, 
               32'shc15142c6, 32'shc150f19f, 32'shc150a082, 32'shc1504f6e, 32'shc14ffe64, 32'shc14fad64, 32'shc14f5c6d, 32'shc14f0b80, 
               32'shc14eba9d, 32'shc14e69c3, 32'shc14e18f3, 32'shc14dc82d, 32'shc14d7771, 32'shc14d26be, 32'shc14cd614, 32'shc14c8575, 
               32'shc14c34df, 32'shc14be453, 32'shc14b93d0, 32'shc14b4357, 32'shc14af2e8, 32'shc14aa282, 32'shc14a5226, 32'shc14a01d4, 
               32'shc149b18b, 32'shc149614c, 32'shc1491117, 32'shc148c0ec, 32'shc14870ca, 32'shc14820b2, 32'shc147d0a3, 32'shc147809e, 
               32'shc14730a3, 32'shc146e0b1, 32'shc14690ca, 32'shc14640eb, 32'shc145f117, 32'shc145a14c, 32'shc145518b, 32'shc14501d3, 
               32'shc144b225, 32'shc1446281, 32'shc14412e7, 32'shc143c356, 32'shc14373cf, 32'shc1432451, 32'shc142d4de, 32'shc1428574, 
               32'shc1423613, 32'shc141e6bc, 32'shc141976f, 32'shc141482c, 32'shc140f8f2, 32'shc140a9c2, 32'shc1405a9c, 32'shc1400b7f, 
               32'shc13fbc6c, 32'shc13f6d63, 32'shc13f1e63, 32'shc13ecf6d, 32'shc13e8081, 32'shc13e319e, 32'shc13de2c5, 32'shc13d93f6, 
               32'shc13d4530, 32'shc13cf674, 32'shc13ca7c2, 32'shc13c591a, 32'shc13c0a7b, 32'shc13bbbe6, 32'shc13b6d5a, 32'shc13b1ed8, 
               32'shc13ad060, 32'shc13a81f2, 32'shc13a338d, 32'shc139e532, 32'shc13996e0, 32'shc1394898, 32'shc138fa5a, 32'shc138ac26, 
               32'shc1385dfb, 32'shc1380fda, 32'shc137c1c3, 32'shc13773b5, 32'shc13725b1, 32'shc136d7b7, 32'shc13689c6, 32'shc1363bdf, 
               32'shc135ee02, 32'shc135a02f, 32'shc1355265, 32'shc13504a4, 32'shc134b6ee, 32'shc1346941, 32'shc1341b9e, 32'shc133ce04, 
               32'shc1338075, 32'shc13332ef, 32'shc132e572, 32'shc13297ff, 32'shc1324a96, 32'shc131fd37, 32'shc131afe1, 32'shc1316295, 
               32'shc1311553, 32'shc130c81a, 32'shc1307aeb, 32'shc1302dc6, 32'shc12fe0ab, 32'shc12f9399, 32'shc12f4690, 32'shc12ef992, 
               32'shc12eac9d, 32'shc12e5fb2, 32'shc12e12d1, 32'shc12dc5f9, 32'shc12d792b, 32'shc12d2c66, 32'shc12cdfac, 32'shc12c92fb, 
               32'shc12c4653, 32'shc12bf9b6, 32'shc12bad22, 32'shc12b6098, 32'shc12b1417, 32'shc12ac7a0, 32'shc12a7b33, 32'shc12a2ecf, 
               32'shc129e276, 32'shc1299626, 32'shc12949df, 32'shc128fda2, 32'shc128b16f, 32'shc1286546, 32'shc1281926, 32'shc127cd10, 
               32'shc1278104, 32'shc1273501, 32'shc126e909, 32'shc1269d19, 32'shc1265134, 32'shc1260558, 32'shc125b986, 32'shc1256dbe, 
               32'shc12521ff, 32'shc124d64a, 32'shc1248a9e, 32'shc1243efd, 32'shc123f365, 32'shc123a7d7, 32'shc1235c52, 32'shc12310d7, 
               32'shc122c566, 32'shc12279fe, 32'shc1222ea1, 32'shc121e34c, 32'shc1219802, 32'shc1214cc1, 32'shc121018a, 32'shc120b65d, 
               32'shc1206b39, 32'shc120201f, 32'shc11fd50f, 32'shc11f8a09, 32'shc11f3f0c, 32'shc11ef419, 32'shc11ea92f, 32'shc11e5e4f, 
               32'shc11e1379, 32'shc11dc8ad, 32'shc11d7dea, 32'shc11d3331, 32'shc11ce882, 32'shc11c9ddd, 32'shc11c5341, 32'shc11c08af, 
               32'shc11bbe26, 32'shc11b73a7, 32'shc11b2932, 32'shc11adec7, 32'shc11a9465, 32'shc11a4a0d, 32'shc119ffbf, 32'shc119b57a, 
               32'shc1196b3f, 32'shc119210e, 32'shc118d6e7, 32'shc1188cc9, 32'shc11842b5, 32'shc117f8ab, 32'shc117aeaa, 32'shc11764b3, 
               32'shc1171ac6, 32'shc116d0e2, 32'shc1168708, 32'shc1163d38, 32'shc115f372, 32'shc115a9b5, 32'shc1156002, 32'shc1151658, 
               32'shc114ccb9, 32'shc1148323, 32'shc1143997, 32'shc113f014, 32'shc113a69b, 32'shc1135d2c, 32'shc11313c7, 32'shc112ca6b, 
               32'shc1128119, 32'shc11237d0, 32'shc111ee92, 32'shc111a55d, 32'shc1115c32, 32'shc1111310, 32'shc110c9f8, 32'shc11080ea, 
               32'shc11037e6, 32'shc10feeeb, 32'shc10fa5fa, 32'shc10f5d13, 32'shc10f1435, 32'shc10ecb62, 32'shc10e8297, 32'shc10e39d7, 
               32'shc10df120, 32'shc10da873, 32'shc10d5fd0, 32'shc10d1736, 32'shc10ccea6, 32'shc10c8620, 32'shc10c3da4, 32'shc10bf531, 
               32'shc10bacc8, 32'shc10b6468, 32'shc10b1c13, 32'shc10ad3c7, 32'shc10a8b85, 32'shc10a434c, 32'shc109fb1d, 32'shc109b2f8, 
               32'shc1096add, 32'shc10922cb, 32'shc108dac3, 32'shc10892c5, 32'shc1084ad0, 32'shc10802e5, 32'shc107bb04, 32'shc107732d, 
               32'shc1072b5f, 32'shc106e39b, 32'shc1069be1, 32'shc1065430, 32'shc1060c89, 32'shc105c4ec, 32'shc1057d59, 32'shc10535cf, 
               32'shc104ee4f, 32'shc104a6d8, 32'shc1045f6c, 32'shc1041809, 32'shc103d0b0, 32'shc1038960, 32'shc103421b, 32'shc102fadf, 
               32'shc102b3ac, 32'shc1026c84, 32'shc1022565, 32'shc101de50, 32'shc1019744, 32'shc1015042, 32'shc101094a, 32'shc100c25c, 
               32'shc1007b77, 32'shc100349c, 32'shc0ffedcb, 32'shc0ffa704, 32'shc0ff6046, 32'shc0ff1992, 32'shc0fed2e8, 32'shc0fe8c47, 
               32'shc0fe45b0, 32'shc0fdff23, 32'shc0fdb8a0, 32'shc0fd7226, 32'shc0fd2bb6, 32'shc0fce54f, 32'shc0fc9ef3, 32'shc0fc58a0, 
               32'shc0fc1257, 32'shc0fbcc17, 32'shc0fb85e2, 32'shc0fb3fb6, 32'shc0faf993, 32'shc0fab37b, 32'shc0fa6d6c, 32'shc0fa2767, 
               32'shc0f9e16b, 32'shc0f99b7a, 32'shc0f95592, 32'shc0f90fb4, 32'shc0f8c9df, 32'shc0f88414, 32'shc0f83e53, 32'shc0f7f89c, 
               32'shc0f7b2ee, 32'shc0f76d4a, 32'shc0f727b0, 32'shc0f6e220, 32'shc0f69c99, 32'shc0f6571c, 32'shc0f611a8, 32'shc0f5cc3f, 
               32'shc0f586df, 32'shc0f54189, 32'shc0f4fc3c, 32'shc0f4b6fa, 32'shc0f471c1, 32'shc0f42c91, 32'shc0f3e76c, 32'shc0f3a250, 
               32'shc0f35d3e, 32'shc0f31836, 32'shc0f2d337, 32'shc0f28e42, 32'shc0f24957, 32'shc0f20475, 32'shc0f1bf9d, 32'shc0f17acf, 
               32'shc0f1360b, 32'shc0f0f151, 32'shc0f0aca0, 32'shc0f067f9, 32'shc0f0235b, 32'shc0efdec7, 32'shc0ef9a3d, 32'shc0ef55bd, 
               32'shc0ef1147, 32'shc0eeccda, 32'shc0ee8877, 32'shc0ee441e, 32'shc0edffce, 32'shc0edbb88, 32'shc0ed774c, 32'shc0ed3319, 
               32'shc0eceef1, 32'shc0ecaad2, 32'shc0ec66bc, 32'shc0ec22b1, 32'shc0ebdeaf, 32'shc0eb9ab7, 32'shc0eb56c9, 32'shc0eb12e4, 
               32'shc0eacf09, 32'shc0ea8b38, 32'shc0ea4771, 32'shc0ea03b3, 32'shc0e9bfff, 32'shc0e97c55, 32'shc0e938b4, 32'shc0e8f51d, 
               32'shc0e8b190, 32'shc0e86e0d, 32'shc0e82a93, 32'shc0e7e724, 32'shc0e7a3bd, 32'shc0e76061, 32'shc0e71d0e, 32'shc0e6d9c5, 
               32'shc0e69686, 32'shc0e65351, 32'shc0e61025, 32'shc0e5cd03, 32'shc0e589eb, 32'shc0e546dc, 32'shc0e503d7, 32'shc0e4c0dc, 
               32'shc0e47deb, 32'shc0e43b03, 32'shc0e3f825, 32'shc0e3b551, 32'shc0e37287, 32'shc0e32fc6, 32'shc0e2ed0f, 32'shc0e2aa62, 
               32'shc0e267be, 32'shc0e22525, 32'shc0e1e294, 32'shc0e1a00e, 32'shc0e15d92, 32'shc0e11b1f, 32'shc0e0d8b6, 32'shc0e09656, 
               32'shc0e05401, 32'shc0e011b5, 32'shc0dfcf73, 32'shc0df8d3a, 32'shc0df4b0b, 32'shc0df08e6, 32'shc0dec6cb, 32'shc0de84ba, 
               32'shc0de42b2, 32'shc0de00b4, 32'shc0ddbec0, 32'shc0dd7cd5, 32'shc0dd3af4, 32'shc0dcf91d, 32'shc0dcb750, 32'shc0dc758c, 
               32'shc0dc33d2, 32'shc0dbf222, 32'shc0dbb07c, 32'shc0db6edf, 32'shc0db2d4c, 32'shc0daebc3, 32'shc0daaa44, 32'shc0da68ce, 
               32'shc0da2762, 32'shc0d9e600, 32'shc0d9a4a7, 32'shc0d96359, 32'shc0d92214, 32'shc0d8e0d8, 32'shc0d89fa7, 32'shc0d85e7f, 
               32'shc0d81d61, 32'shc0d7dc4d, 32'shc0d79b42, 32'shc0d75a41, 32'shc0d7194a, 32'shc0d6d85d, 32'shc0d69779, 32'shc0d6569f, 
               32'shc0d615cf, 32'shc0d5d509, 32'shc0d5944c, 32'shc0d55399, 32'shc0d512f0, 32'shc0d4d251, 32'shc0d491bb, 32'shc0d4512f, 
               32'shc0d410ad, 32'shc0d3d034, 32'shc0d38fc6, 32'shc0d34f61, 32'shc0d30f05, 32'shc0d2ceb4, 32'shc0d28e6c, 32'shc0d24e2e, 
               32'shc0d20dfa, 32'shc0d1cdcf, 32'shc0d18dae, 32'shc0d14d97, 32'shc0d10d8a, 32'shc0d0cd87, 32'shc0d08d8d, 32'shc0d04d9d, 
               32'shc0d00db6, 32'shc0cfcdda, 32'shc0cf8e07, 32'shc0cf4e3e, 32'shc0cf0e7f, 32'shc0cecec9, 32'shc0ce8f1d, 32'shc0ce4f7b, 
               32'shc0ce0fe3, 32'shc0cdd054, 32'shc0cd90cf, 32'shc0cd5154, 32'shc0cd11e3, 32'shc0ccd27b, 32'shc0cc931d, 32'shc0cc53c9, 
               32'shc0cc147f, 32'shc0cbd53e, 32'shc0cb9607, 32'shc0cb56da, 32'shc0cb17b7, 32'shc0cad89d, 32'shc0ca998d, 32'shc0ca5a87, 
               32'shc0ca1b8a, 32'shc0c9dc98, 32'shc0c99daf, 32'shc0c95ed0, 32'shc0c91ffa, 32'shc0c8e12f, 32'shc0c8a26d, 32'shc0c863b4, 
               32'shc0c82506, 32'shc0c7e661, 32'shc0c7a7c6, 32'shc0c76935, 32'shc0c72aae, 32'shc0c6ec30, 32'shc0c6adbc, 32'shc0c66f52, 
               32'shc0c630f2, 32'shc0c5f29b, 32'shc0c5b44e, 32'shc0c5760b, 32'shc0c537d1, 32'shc0c4f9a2, 32'shc0c4bb7c, 32'shc0c47d60, 
               32'shc0c43f4d, 32'shc0c40144, 32'shc0c3c346, 32'shc0c38550, 32'shc0c34765, 32'shc0c30983, 32'shc0c2cbab, 32'shc0c28ddd, 
               32'shc0c25019, 32'shc0c2125e, 32'shc0c1d4ad, 32'shc0c19706, 32'shc0c15969, 32'shc0c11bd5, 32'shc0c0de4b, 32'shc0c0a0cb, 
               32'shc0c06355, 32'shc0c025e8, 32'shc0bfe885, 32'shc0bfab2c, 32'shc0bf6ddd, 32'shc0bf3097, 32'shc0bef35b, 32'shc0beb629, 
               32'shc0be7901, 32'shc0be3be2, 32'shc0bdfecd, 32'shc0bdc1c2, 32'shc0bd84c1, 32'shc0bd47c9, 32'shc0bd0adb, 32'shc0bccdf7, 
               32'shc0bc911d, 32'shc0bc544d, 32'shc0bc1786, 32'shc0bbdac9, 32'shc0bb9e15, 32'shc0bb616c, 32'shc0bb24cc, 32'shc0bae836, 
               32'shc0baabaa, 32'shc0ba6f27, 32'shc0ba32af, 32'shc0b9f640, 32'shc0b9b9da, 32'shc0b97d7f, 32'shc0b9412d, 32'shc0b904e5, 
               32'shc0b8c8a7, 32'shc0b88c73, 32'shc0b85048, 32'shc0b81427, 32'shc0b7d810, 32'shc0b79c02, 32'shc0b75fff, 32'shc0b72405, 
               32'shc0b6e815, 32'shc0b6ac2e, 32'shc0b67052, 32'shc0b6347f, 32'shc0b5f8b6, 32'shc0b5bcf7, 32'shc0b58141, 32'shc0b54595, 
               32'shc0b509f3, 32'shc0b4ce5b, 32'shc0b492cc, 32'shc0b45748, 32'shc0b41bcd, 32'shc0b3e05b, 32'shc0b3a4f4, 32'shc0b36996, 
               32'shc0b32e42, 32'shc0b2f2f8, 32'shc0b2b7b8, 32'shc0b27c81, 32'shc0b24154, 32'shc0b20631, 32'shc0b1cb17, 32'shc0b19008, 
               32'shc0b15502, 32'shc0b11a06, 32'shc0b0df13, 32'shc0b0a42b, 32'shc0b0694c, 32'shc0b02e77, 32'shc0aff3ac, 32'shc0afb8ea, 
               32'shc0af7e33, 32'shc0af4385, 32'shc0af08e0, 32'shc0aece46, 32'shc0ae93b5, 32'shc0ae592e, 32'shc0ae1eb1, 32'shc0ade43e, 
               32'shc0ada9d4, 32'shc0ad6f74, 32'shc0ad351e, 32'shc0acfad2, 32'shc0acc08f, 32'shc0ac8656, 32'shc0ac4c27, 32'shc0ac1202, 
               32'shc0abd7e6, 32'shc0ab9dd5, 32'shc0ab63cd, 32'shc0ab29ce, 32'shc0aaefda, 32'shc0aab5ef, 32'shc0aa7c0e, 32'shc0aa4237, 
               32'shc0aa086a, 32'shc0a9cea6, 32'shc0a994ec, 32'shc0a95b3c, 32'shc0a92196, 32'shc0a8e7f9, 32'shc0a8ae67, 32'shc0a874de, 
               32'shc0a83b5e, 32'shc0a801e9, 32'shc0a7c87d, 32'shc0a78f1b, 32'shc0a755c3, 32'shc0a71c75, 32'shc0a6e330, 32'shc0a6a9f5, 
               32'shc0a670c4, 32'shc0a6379d, 32'shc0a5fe7f, 32'shc0a5c56c, 32'shc0a58c62, 32'shc0a55361, 32'shc0a51a6b, 32'shc0a4e17e, 
               32'shc0a4a89b, 32'shc0a46fc2, 32'shc0a436f3, 32'shc0a3fe2d, 32'shc0a3c571, 32'shc0a38cbf, 32'shc0a35417, 32'shc0a31b78, 
               32'shc0a2e2e3, 32'shc0a2aa58, 32'shc0a271d7, 32'shc0a23960, 32'shc0a200f2, 32'shc0a1c88e, 32'shc0a19034, 32'shc0a157e4, 
               32'shc0a11f9d, 32'shc0a0e760, 32'shc0a0af2d, 32'shc0a07704, 32'shc0a03ee4, 32'shc0a006cf, 32'shc09fcec3, 32'shc09f96c1, 
               32'shc09f5ec8, 32'shc09f26da, 32'shc09eeef5, 32'shc09eb71a, 32'shc09e7f48, 32'shc09e4781, 32'shc09e0fc3, 32'shc09dd80f, 
               32'shc09da065, 32'shc09d68c4, 32'shc09d312e, 32'shc09cf9a1, 32'shc09cc21e, 32'shc09c8aa4, 32'shc09c5335, 32'shc09c1bcf, 
               32'shc09be473, 32'shc09bad21, 32'shc09b75d8, 32'shc09b3e9a, 32'shc09b0765, 32'shc09ad03a, 32'shc09a9918, 32'shc09a6201, 
               32'shc09a2af3, 32'shc099f3ef, 32'shc099bcf5, 32'shc0998604, 32'shc0994f1d, 32'shc0991840, 32'shc098e16d, 32'shc098aaa4, 
               32'shc09873e4, 32'shc0983d2f, 32'shc0980683, 32'shc097cfe0, 32'shc0979948, 32'shc09762b9, 32'shc0972c34, 32'shc096f5b9, 
               32'shc096bf48, 32'shc09688e0, 32'shc0965282, 32'shc0961c2e, 32'shc095e5e4, 32'shc095afa4, 32'shc095796d, 32'shc0954340, 
               32'shc0950d1d, 32'shc094d703, 32'shc094a0f4, 32'shc0946aee, 32'shc09434f2, 32'shc093ff00, 32'shc093c917, 32'shc0939339, 
               32'shc0935d64, 32'shc0932799, 32'shc092f1d7, 32'shc092bc20, 32'shc0928672, 32'shc09250ce, 32'shc0921b34, 32'shc091e5a4, 
               32'shc091b01d, 32'shc0917aa0, 32'shc091452d, 32'shc0910fc4, 32'shc090da64, 32'shc090a50e, 32'shc0906fc3, 32'shc0903a80, 
               32'shc0900548, 32'shc08fd019, 32'shc08f9af5, 32'shc08f65da, 32'shc08f30c8, 32'shc08efbc1, 32'shc08ec6c3, 32'shc08e91cf, 
               32'shc08e5ce5, 32'shc08e2805, 32'shc08df32e, 32'shc08dbe62, 32'shc08d899f, 32'shc08d54e5, 32'shc08d2036, 32'shc08ceb90, 
               32'shc08cb6f5, 32'shc08c8262, 32'shc08c4dda, 32'shc08c195c, 32'shc08be4e7, 32'shc08bb07c, 32'shc08b7c1b, 32'shc08b47c4, 
               32'shc08b1376, 32'shc08adf32, 32'shc08aaaf8, 32'shc08a76c8, 32'shc08a42a2, 32'shc08a0e85, 32'shc089da72, 32'shc089a669, 
               32'shc089726a, 32'shc0893e75, 32'shc0890a89, 32'shc088d6a7, 32'shc088a2cf, 32'shc0886f00, 32'shc0883b3c, 32'shc0880781, 
               32'shc087d3d0, 32'shc087a029, 32'shc0876c8c, 32'shc08738f8, 32'shc087056e, 32'shc086d1ee, 32'shc0869e78, 32'shc0866b0c, 
               32'shc08637a9, 32'shc0860450, 32'shc085d101, 32'shc0859dbc, 32'shc0856a80, 32'shc085374e, 32'shc0850426, 32'shc084d108, 
               32'shc0849df4, 32'shc0846ae9, 32'shc08437e9, 32'shc08404f2, 32'shc083d204, 32'shc0839f21, 32'shc0836c47, 32'shc0833978, 
               32'shc08306b2, 32'shc082d3f5, 32'shc082a143, 32'shc0826e9a, 32'shc0823bfb, 32'shc0820966, 32'shc081d6db, 32'shc081a45a, 
               32'shc08171e2, 32'shc0813f74, 32'shc0810d10, 32'shc080dab6, 32'shc080a865, 32'shc080761e, 32'shc08043e1, 32'shc08011ae, 
               32'shc07fdf85, 32'shc07fad65, 32'shc07f7b50, 32'shc07f4944, 32'shc07f1741, 32'shc07ee549, 32'shc07eb35a, 32'shc07e8176, 
               32'shc07e4f9b, 32'shc07e1dc9, 32'shc07dec02, 32'shc07dba44, 32'shc07d8890, 32'shc07d56e6, 32'shc07d2546, 32'shc07cf3b0, 
               32'shc07cc223, 32'shc07c90a0, 32'shc07c5f27, 32'shc07c2db8, 32'shc07bfc52, 32'shc07bcaf7, 32'shc07b99a5, 32'shc07b685d, 
               32'shc07b371e, 32'shc07b05ea, 32'shc07ad4bf, 32'shc07aa39e, 32'shc07a7287, 32'shc07a417a, 32'shc07a1076, 32'shc079df7c, 
               32'shc079ae8c, 32'shc0797da6, 32'shc0794cca, 32'shc0791bf7, 32'shc078eb2f, 32'shc078ba70, 32'shc07889bb, 32'shc078590f, 
               32'shc078286e, 32'shc077f7d6, 32'shc077c748, 32'shc07796c4, 32'shc0776649, 32'shc07735d9, 32'shc0770572, 32'shc076d515, 
               32'shc076a4c2, 32'shc0767478, 32'shc0764439, 32'shc0761403, 32'shc075e3d7, 32'shc075b3b5, 32'shc075839c, 32'shc075538e, 
               32'shc0752389, 32'shc074f38e, 32'shc074c39d, 32'shc07493b5, 32'shc07463d8, 32'shc0743404, 32'shc074043a, 32'shc073d47a, 
               32'shc073a4c3, 32'shc0737517, 32'shc0734574, 32'shc07315db, 32'shc072e64c, 32'shc072b6c6, 32'shc072874b, 32'shc07257d9, 
               32'shc0722871, 32'shc071f913, 32'shc071c9be, 32'shc0719a74, 32'shc0716b33, 32'shc0713bfc, 32'shc0710ccf, 32'shc070ddab, 
               32'shc070ae92, 32'shc0707f82, 32'shc070507c, 32'shc0702180, 32'shc06ff28e, 32'shc06fc3a5, 32'shc06f94c6, 32'shc06f65f1, 
               32'shc06f3726, 32'shc06f0865, 32'shc06ed9ad, 32'shc06eaaff, 32'shc06e7c5b, 32'shc06e4dc1, 32'shc06e1f31, 32'shc06df0aa, 
               32'shc06dc22e, 32'shc06d93bb, 32'shc06d6551, 32'shc06d36f2, 32'shc06d089d, 32'shc06cda51, 32'shc06cac0f, 32'shc06c7dd7, 
               32'shc06c4fa8, 32'shc06c2184, 32'shc06bf369, 32'shc06bc558, 32'shc06b9751, 32'shc06b6954, 32'shc06b3b60, 32'shc06b0d77, 
               32'shc06adf97, 32'shc06ab1c1, 32'shc06a83f5, 32'shc06a5632, 32'shc06a2879, 32'shc069facb, 32'shc069cd26, 32'shc0699f8a, 
               32'shc06971f9, 32'shc0694471, 32'shc06916f3, 32'shc068e97f, 32'shc068bc15, 32'shc0688eb5, 32'shc068615e, 32'shc0683411, 
               32'shc06806ce, 32'shc067d995, 32'shc067ac66, 32'shc0677f40, 32'shc0675225, 32'shc0672513, 32'shc066f80a, 32'shc066cb0c, 
               32'shc0669e18, 32'shc066712d, 32'shc066444c, 32'shc0661775, 32'shc065eaa8, 32'shc065bde4, 32'shc065912a, 32'shc065647b, 
               32'shc06537d4, 32'shc0650b38, 32'shc064dea6, 32'shc064b21d, 32'shc064859e, 32'shc0645929, 32'shc0642cbe, 32'shc064005d, 
               32'shc063d405, 32'shc063a7b7, 32'shc0637b73, 32'shc0634f39, 32'shc0632309, 32'shc062f6e2, 32'shc062cac6, 32'shc0629eb3, 
               32'shc06272aa, 32'shc06246aa, 32'shc0621ab5, 32'shc061eec9, 32'shc061c2e7, 32'shc061970f, 32'shc0616b41, 32'shc0613f7d, 
               32'shc06113c2, 32'shc060e811, 32'shc060bc6a, 32'shc06090cd, 32'shc060653a, 32'shc06039b0, 32'shc0600e30, 32'shc05fe2ba, 
               32'shc05fb74e, 32'shc05f8bec, 32'shc05f6093, 32'shc05f3545, 32'shc05f0a00, 32'shc05edec5, 32'shc05eb393, 32'shc05e886c, 
               32'shc05e5d4e, 32'shc05e323a, 32'shc05e0730, 32'shc05ddc30, 32'shc05db13a, 32'shc05d864d, 32'shc05d5b6b, 32'shc05d3092, 
               32'shc05d05c3, 32'shc05cdafd, 32'shc05cb042, 32'shc05c8590, 32'shc05c5ae8, 32'shc05c304a, 32'shc05c05b6, 32'shc05bdb2b, 
               32'shc05bb0ab, 32'shc05b8634, 32'shc05b5bc7, 32'shc05b3164, 32'shc05b070a, 32'shc05adcbb, 32'shc05ab275, 32'shc05a8839, 
               32'shc05a5e07, 32'shc05a33df, 32'shc05a09c0, 32'shc059dfac, 32'shc059b5a1, 32'shc0598ba0, 32'shc05961a9, 32'shc05937bb, 
               32'shc0590dd8, 32'shc058e3fe, 32'shc058ba2e, 32'shc0589068, 32'shc05866ac, 32'shc0583cf9, 32'shc0581350, 32'shc057e9b2, 
               32'shc057c01d, 32'shc0579691, 32'shc0576d10, 32'shc0574398, 32'shc0571a2b, 32'shc056f0c7, 32'shc056c76c, 32'shc0569e1c, 
               32'shc05674d6, 32'shc0564b99, 32'shc0562266, 32'shc055f93d, 32'shc055d01e, 32'shc055a708, 32'shc0557dfd, 32'shc05554fb, 
               32'shc0552c03, 32'shc0550315, 32'shc054da30, 32'shc054b156, 32'shc0548885, 32'shc0545fbe, 32'shc0543701, 32'shc0540e4e, 
               32'shc053e5a5, 32'shc053bd05, 32'shc053946f, 32'shc0536be3, 32'shc0534361, 32'shc0531ae9, 32'shc052f27a, 32'shc052ca16, 
               32'shc052a1bb, 32'shc052796a, 32'shc0525123, 32'shc05228e5, 32'shc05200b2, 32'shc051d888, 32'shc051b068, 32'shc0518852, 
               32'shc0516045, 32'shc0513843, 32'shc051104a, 32'shc050e85c, 32'shc050c077, 32'shc050989b, 32'shc05070ca, 32'shc0504902, 
               32'shc0502145, 32'shc04ff991, 32'shc04fd1e7, 32'shc04faa46, 32'shc04f82b0, 32'shc04f5b23, 32'shc04f33a1, 32'shc04f0c28, 
               32'shc04ee4b8, 32'shc04ebd53, 32'shc04e95f8, 32'shc04e6ea6, 32'shc04e475e, 32'shc04e2020, 32'shc04df8ec, 32'shc04dd1c1, 
               32'shc04daaa1, 32'shc04d838a, 32'shc04d5c7d, 32'shc04d357a, 32'shc04d0e81, 32'shc04ce791, 32'shc04cc0ac, 32'shc04c99d0, 
               32'shc04c72fe, 32'shc04c4c36, 32'shc04c2577, 32'shc04bfec3, 32'shc04bd818, 32'shc04bb177, 32'shc04b8ae0, 32'shc04b6453, 
               32'shc04b3dcf, 32'shc04b1756, 32'shc04af0e6, 32'shc04aca80, 32'shc04aa424, 32'shc04a7dd2, 32'shc04a5789, 32'shc04a314b, 
               32'shc04a0b16, 32'shc049e4eb, 32'shc049beca, 32'shc04998b2, 32'shc04972a5, 32'shc0494ca1, 32'shc04926a7, 32'shc04900b7, 
               32'shc048dad1, 32'shc048b4f5, 32'shc0488f22, 32'shc0486959, 32'shc048439b, 32'shc0481de5, 32'shc047f83a, 32'shc047d299, 
               32'shc047ad01, 32'shc0478773, 32'shc04761ef, 32'shc0473c75, 32'shc0471705, 32'shc046f19f, 32'shc046cc42, 32'shc046a6ef, 
               32'shc04681a6, 32'shc0465c67, 32'shc0463732, 32'shc0461206, 32'shc045ece5, 32'shc045c7cd, 32'shc045a2bf, 32'shc0457dba, 
               32'shc04558c0, 32'shc04533d0, 32'shc0450ee9, 32'shc044ea0c, 32'shc044c539, 32'shc044a070, 32'shc0447bb0, 32'shc04456fb, 
               32'shc044324f, 32'shc0440dad, 32'shc043e915, 32'shc043c487, 32'shc043a002, 32'shc0437b88, 32'shc0435717, 32'shc04332b0, 
               32'shc0430e53, 32'shc042ea00, 32'shc042c5b6, 32'shc042a177, 32'shc0427d41, 32'shc0425915, 32'shc04234f3, 32'shc04210da, 
               32'shc041eccc, 32'shc041c8c7, 32'shc041a4cd, 32'shc04180dc, 32'shc0415cf4, 32'shc0413917, 32'shc0411544, 32'shc040f17a, 
               32'shc040cdba, 32'shc040aa04, 32'shc0408658, 32'shc04062b6, 32'shc0403f1d, 32'shc0401b8e, 32'shc03ff80a, 32'shc03fd48f, 
               32'shc03fb11d, 32'shc03f8db6, 32'shc03f6a58, 32'shc03f4705, 32'shc03f23bb, 32'shc03f007b, 32'shc03edd45, 32'shc03eba18, 
               32'shc03e96f6, 32'shc03e73dd, 32'shc03e50ce, 32'shc03e2dc9, 32'shc03e0ace, 32'shc03de7dd, 32'shc03dc4f5, 32'shc03da217, 
               32'shc03d7f44, 32'shc03d5c79, 32'shc03d39b9, 32'shc03d1703, 32'shc03cf456, 32'shc03cd1b4, 32'shc03caf1b, 32'shc03c8c8c, 
               32'shc03c6a07, 32'shc03c478b, 32'shc03c251a, 32'shc03c02b2, 32'shc03be054, 32'shc03bbe00, 32'shc03b9bb6, 32'shc03b7975, 
               32'shc03b573f, 32'shc03b3512, 32'shc03b12ef, 32'shc03af0d6, 32'shc03acec7, 32'shc03aacc2, 32'shc03a8ac6, 32'shc03a68d4, 
               32'shc03a46ed, 32'shc03a250e, 32'shc03a033a, 32'shc039e170, 32'shc039bfaf, 32'shc0399df9, 32'shc0397c4c, 32'shc0395aa9, 
               32'shc0393910, 32'shc0391780, 32'shc038f5fb, 32'shc038d47f, 32'shc038b30d, 32'shc03891a5, 32'shc0387047, 32'shc0384ef3, 
               32'shc0382da8, 32'shc0380c68, 32'shc037eb31, 32'shc037ca04, 32'shc037a8e1, 32'shc03787c7, 32'shc03766b8, 32'shc03745b2, 
               32'shc03724b6, 32'shc03703c4, 32'shc036e2dc, 32'shc036c1fe, 32'shc036a129, 32'shc036805f, 32'shc0365f9e, 32'shc0363ee7, 
               32'shc0361e3a, 32'shc035fd96, 32'shc035dcfd, 32'shc035bc6d, 32'shc0359be8, 32'shc0357b6c, 32'shc0355afa, 32'shc0353a91, 
               32'shc0351a33, 32'shc034f9de, 32'shc034d994, 32'shc034b953, 32'shc034991c, 32'shc03478ee, 32'shc03458cb, 32'shc03438b1, 
               32'shc03418a2, 32'shc033f89c, 32'shc033d8a0, 32'shc033b8ad, 32'shc03398c5, 32'shc03378e7, 32'shc0335912, 32'shc0333947, 
               32'shc0331986, 32'shc032f9cf, 32'shc032da22, 32'shc032ba7e, 32'shc0329ae4, 32'shc0327b55, 32'shc0325bcf, 32'shc0323c52, 
               32'shc0321ce0, 32'shc031fd78, 32'shc031de19, 32'shc031bec4, 32'shc0319f79, 32'shc0318038, 32'shc0316101, 32'shc03141d3, 
               32'shc03122b0, 32'shc0310396, 32'shc030e486, 32'shc030c580, 32'shc030a684, 32'shc0308792, 32'shc03068a9, 32'shc03049ca, 
               32'shc0302af5, 32'shc0300c2a, 32'shc02fed69, 32'shc02fceb2, 32'shc02fb004, 32'shc02f9161, 32'shc02f72c7, 32'shc02f5437, 
               32'shc02f35b1, 32'shc02f1734, 32'shc02ef8c2, 32'shc02eda59, 32'shc02ebbfb, 32'shc02e9da6, 32'shc02e7f5b, 32'shc02e6119, 
               32'shc02e42e2, 32'shc02e24b4, 32'shc02e0691, 32'shc02de877, 32'shc02dca67, 32'shc02dac61, 32'shc02d8e64, 32'shc02d7072, 
               32'shc02d5289, 32'shc02d34aa, 32'shc02d16d5, 32'shc02cf90a, 32'shc02cdb49, 32'shc02cbd91, 32'shc02c9fe4, 32'shc02c8240, 
               32'shc02c64a6, 32'shc02c4716, 32'shc02c2990, 32'shc02c0c13, 32'shc02beea1, 32'shc02bd138, 32'shc02bb3d9, 32'shc02b9684, 
               32'shc02b7939, 32'shc02b5bf8, 32'shc02b3ec0, 32'shc02b2192, 32'shc02b046f, 32'shc02ae755, 32'shc02aca44, 32'shc02aad3e, 
               32'shc02a9042, 32'shc02a734f, 32'shc02a5666, 32'shc02a3988, 32'shc02a1cb2, 32'shc029ffe7, 32'shc029e326, 32'shc029c66e, 
               32'shc029a9c1, 32'shc0298d1d, 32'shc0297083, 32'shc02953f3, 32'shc029376c, 32'shc0291af0, 32'shc028fe7d, 32'shc028e215, 
               32'shc028c5b6, 32'shc028a961, 32'shc0288d15, 32'shc02870d4, 32'shc028549c, 32'shc028386f, 32'shc0281c4b, 32'shc0280031, 
               32'shc027e421, 32'shc027c81a, 32'shc027ac1e, 32'shc027902b, 32'shc0277442, 32'shc0275864, 32'shc0273c8e, 32'shc02720c3, 
               32'shc0270502, 32'shc026e94a, 32'shc026cd9d, 32'shc026b1f9, 32'shc026965f, 32'shc0267acf, 32'shc0265f48, 32'shc02643cc, 
               32'shc0262859, 32'shc0260cf0, 32'shc025f191, 32'shc025d63c, 32'shc025baf1, 32'shc0259fb0, 32'shc0258478, 32'shc025694a, 
               32'shc0254e27, 32'shc025330d, 32'shc02517fc, 32'shc024fcf6, 32'shc024e1fa, 32'shc024c707, 32'shc024ac1e, 32'shc024913f, 
               32'shc024766a, 32'shc0245b9f, 32'shc02440de, 32'shc0242626, 32'shc0240b78, 32'shc023f0d5, 32'shc023d63b, 32'shc023bbab, 
               32'shc023a124, 32'shc02386a8, 32'shc0236c35, 32'shc02351cc, 32'shc023376e, 32'shc0231d18, 32'shc02302cd, 32'shc022e88c, 
               32'shc022ce54, 32'shc022b427, 32'shc0229a03, 32'shc0227fe9, 32'shc02265d9, 32'shc0224bd3, 32'shc02231d6, 32'shc02217e4, 
               32'shc021fdfb, 32'shc021e41c, 32'shc021ca47, 32'shc021b07c, 32'shc02196bb, 32'shc0217d03, 32'shc0216356, 32'shc02149b2, 
               32'shc0213018, 32'shc0211688, 32'shc020fd02, 32'shc020e385, 32'shc020ca13, 32'shc020b0aa, 32'shc020974b, 32'shc0207df6, 
               32'shc02064ab, 32'shc0204b6a, 32'shc0203232, 32'shc0201905, 32'shc01fffe1, 32'shc01fe6c7, 32'shc01fcdb7, 32'shc01fb4b1, 
               32'shc01f9bb5, 32'shc01f82c2, 32'shc01f69da, 32'shc01f50fb, 32'shc01f3826, 32'shc01f1f5b, 32'shc01f069a, 32'shc01eede2, 
               32'shc01ed535, 32'shc01ebc91, 32'shc01ea3f7, 32'shc01e8b67, 32'shc01e72e1, 32'shc01e5a65, 32'shc01e41f3, 32'shc01e298a, 
               32'shc01e112b, 32'shc01df8d7, 32'shc01de08c, 32'shc01dc84a, 32'shc01db013, 32'shc01d97e6, 32'shc01d7fc2, 32'shc01d67a8, 
               32'shc01d4f99, 32'shc01d3792, 32'shc01d1f96, 32'shc01d07a4, 32'shc01cefbb, 32'shc01cd7dd, 32'shc01cc008, 32'shc01ca83d, 
               32'shc01c907c, 32'shc01c78c5, 32'shc01c6118, 32'shc01c4974, 32'shc01c31da, 32'shc01c1a4b, 32'shc01c02c5, 32'shc01beb48, 
               32'shc01bd3d6, 32'shc01bbc6e, 32'shc01ba50f, 32'shc01b8dbb, 32'shc01b7670, 32'shc01b5f2f, 32'shc01b47f8, 32'shc01b30ca, 
               32'shc01b19a7, 32'shc01b028d, 32'shc01aeb7e, 32'shc01ad478, 32'shc01abd7c, 32'shc01aa68a, 32'shc01a8fa1, 32'shc01a78c3, 
               32'shc01a61ee, 32'shc01a4b24, 32'shc01a3463, 32'shc01a1dac, 32'shc01a06fe, 32'shc019f05b, 32'shc019d9c2, 32'shc019c332, 
               32'shc019acac, 32'shc0199630, 32'shc0197fbe, 32'shc0196956, 32'shc01952f8, 32'shc0193ca3, 32'shc0192659, 32'shc0191018, 
               32'shc018f9e1, 32'shc018e3b4, 32'shc018cd91, 32'shc018b777, 32'shc018a168, 32'shc0188b62, 32'shc0187566, 32'shc0185f74, 
               32'shc018498c, 32'shc01833ae, 32'shc0181dda, 32'shc018080f, 32'shc017f24e, 32'shc017dc98, 32'shc017c6eb, 32'shc017b148, 
               32'shc0179bae, 32'shc017861f, 32'shc0177099, 32'shc0175b1e, 32'shc01745ac, 32'shc0173044, 32'shc0171ae6, 32'shc0170591, 
               32'shc016f047, 32'shc016db07, 32'shc016c5d0, 32'shc016b0a3, 32'shc0169b80, 32'shc0168667, 32'shc0167158, 32'shc0165c52, 
               32'shc0164757, 32'shc0163265, 32'shc0161d7d, 32'shc016089f, 32'shc015f3cb, 32'shc015df01, 32'shc015ca40, 32'shc015b58a, 
               32'shc015a0dd, 32'shc0158c3a, 32'shc01577a1, 32'shc0156312, 32'shc0154e8d, 32'shc0153a11, 32'shc01525a0, 32'shc0151138, 
               32'shc014fcda, 32'shc014e886, 32'shc014d43c, 32'shc014bffc, 32'shc014abc5, 32'shc0149799, 32'shc0148376, 32'shc0146f5d, 
               32'shc0145b4e, 32'shc0144749, 32'shc014334e, 32'shc0141f5c, 32'shc0140b75, 32'shc013f797, 32'shc013e3c3, 32'shc013cff9, 
               32'shc013bc39, 32'shc013a883, 32'shc01394d6, 32'shc0138134, 32'shc0136d9b, 32'shc0135a0c, 32'shc0134687, 32'shc013330c, 
               32'shc0131f9b, 32'shc0130c33, 32'shc012f8d6, 32'shc012e582, 32'shc012d238, 32'shc012bef8, 32'shc012abc2, 32'shc0129896, 
               32'shc0128574, 32'shc012725b, 32'shc0125f4c, 32'shc0124c47, 32'shc012394c, 32'shc012265b, 32'shc0121374, 32'shc0120097, 
               32'shc011edc3, 32'shc011daf9, 32'shc011c83a, 32'shc011b584, 32'shc011a2d8, 32'shc0119035, 32'shc0117d9d, 32'shc0116b0e, 
               32'shc011588a, 32'shc011460f, 32'shc011339e, 32'shc0112137, 32'shc0110eda, 32'shc010fc86, 32'shc010ea3d, 32'shc010d7fd, 
               32'shc010c5c7, 32'shc010b39b, 32'shc010a179, 32'shc0108f61, 32'shc0107d53, 32'shc0106b4e, 32'shc0105954, 32'shc0104763, 
               32'shc010357c, 32'shc010239f, 32'shc01011cc, 32'shc0100002, 32'shc00fee43, 32'shc00fdc8d, 32'shc00fcae2, 32'shc00fb940, 
               32'shc00fa7a8, 32'shc00f9619, 32'shc00f8495, 32'shc00f731b, 32'shc00f61aa, 32'shc00f5043, 32'shc00f3ee6, 32'shc00f2d93, 
               32'shc00f1c4a, 32'shc00f0b0b, 32'shc00ef9d6, 32'shc00ee8aa, 32'shc00ed788, 32'shc00ec670, 32'shc00eb562, 32'shc00ea45e, 
               32'shc00e9364, 32'shc00e8274, 32'shc00e718d, 32'shc00e60b0, 32'shc00e4fde, 32'shc00e3f15, 32'shc00e2e56, 32'shc00e1da0, 
               32'shc00e0cf5, 32'shc00dfc53, 32'shc00debbc, 32'shc00ddb2e, 32'shc00dcaaa, 32'shc00dba30, 32'shc00da9c0, 32'shc00d9959, 
               32'shc00d88fd, 32'shc00d78aa, 32'shc00d6861, 32'shc00d5823, 32'shc00d47ed, 32'shc00d37c2, 32'shc00d27a1, 32'shc00d178a, 
               32'shc00d077c, 32'shc00cf778, 32'shc00ce77e, 32'shc00cd78e, 32'shc00cc7a8, 32'shc00cb7cc, 32'shc00ca7f9, 32'shc00c9831, 
               32'shc00c8872, 32'shc00c78bd, 32'shc00c6912, 32'shc00c5971, 32'shc00c49da, 32'shc00c3a4d, 32'shc00c2ac9, 32'shc00c1b4f, 
               32'shc00c0be0, 32'shc00bfc7a, 32'shc00bed1e, 32'shc00bddcb, 32'shc00bce83, 32'shc00bbf44, 32'shc00bb010, 32'shc00ba0e5, 
               32'shc00b91c4, 32'shc00b82ad, 32'shc00b73a0, 32'shc00b649d, 32'shc00b55a3, 32'shc00b46b4, 32'shc00b37ce, 32'shc00b28f2, 
               32'shc00b1a20, 32'shc00b0b58, 32'shc00afc9a, 32'shc00aede5, 32'shc00adf3b, 32'shc00ad09a, 32'shc00ac203, 32'shc00ab376, 
               32'shc00aa4f3, 32'shc00a967a, 32'shc00a880a, 32'shc00a79a5, 32'shc00a6b49, 32'shc00a5cf8, 32'shc00a4eb0, 32'shc00a4072, 
               32'shc00a323d, 32'shc00a2413, 32'shc00a15f3, 32'shc00a07dc, 32'shc009f9cf, 32'shc009ebcc, 32'shc009ddd3, 32'shc009cfe4, 
               32'shc009c1ff, 32'shc009b423, 32'shc009a652, 32'shc009988a, 32'shc0098acc, 32'shc0097d18, 32'shc0096f6e, 32'shc00961ce, 
               32'shc0095438, 32'shc00946ab, 32'shc0093929, 32'shc0092bb0, 32'shc0091e41, 32'shc00910dc, 32'shc0090381, 32'shc008f62f, 
               32'shc008e8e8, 32'shc008dbaa, 32'shc008ce76, 32'shc008c14d, 32'shc008b42d, 32'shc008a716, 32'shc0089a0a, 32'shc0088d08, 
               32'shc008800f, 32'shc0087321, 32'shc008663c, 32'shc0085961, 32'shc0084c90, 32'shc0083fc8, 32'shc008330b, 32'shc0082658, 
               32'shc00819ae, 32'shc0080d0e, 32'shc0080078, 32'shc007f3ec, 32'shc007e76a, 32'shc007daf2, 32'shc007ce83, 32'shc007c21f, 
               32'shc007b5c4, 32'shc007a973, 32'shc0079d2c, 32'shc00790ef, 32'shc00784bc, 32'shc0077893, 32'shc0076c73, 32'shc007605d, 
               32'shc0075452, 32'shc0074850, 32'shc0073c58, 32'shc0073069, 32'shc0072485, 32'shc00718ab, 32'shc0070cda, 32'shc0070113, 
               32'shc006f556, 32'shc006e9a3, 32'shc006ddfa, 32'shc006d25b, 32'shc006c6c6, 32'shc006bb3a, 32'shc006afb8, 32'shc006a441, 
               32'shc00698d3, 32'shc0068d6f, 32'shc0068214, 32'shc00676c4, 32'shc0066b7d, 32'shc0066041, 32'shc006550e, 32'shc00649e5, 
               32'shc0063ec6, 32'shc00633b1, 32'shc00628a6, 32'shc0061da4, 32'shc00612ad, 32'shc00607bf, 32'shc005fcdb, 32'shc005f201, 
               32'shc005e731, 32'shc005dc6b, 32'shc005d1af, 32'shc005c6fc, 32'shc005bc54, 32'shc005b1b5, 32'shc005a720, 32'shc0059c95, 
               32'shc0059214, 32'shc005879c, 32'shc0057d2f, 32'shc00572cb, 32'shc0056872, 32'shc0055e22, 32'shc00553dc, 32'shc00549a0, 
               32'shc0053f6e, 32'shc0053545, 32'shc0052b27, 32'shc0052112, 32'shc0051707, 32'shc0050d06, 32'shc005030f, 32'shc004f922, 
               32'shc004ef3f, 32'shc004e566, 32'shc004db96, 32'shc004d1d0, 32'shc004c814, 32'shc004be62, 32'shc004b4ba, 32'shc004ab1c, 
               32'shc004a188, 32'shc00497fd, 32'shc0048e7d, 32'shc0048506, 32'shc0047b99, 32'shc0047236, 32'shc00468dd, 32'shc0045f8d, 
               32'shc0045648, 32'shc0044d0d, 32'shc00443db, 32'shc0043ab3, 32'shc0043195, 32'shc0042881, 32'shc0041f77, 32'shc0041676, 
               32'shc0040d80, 32'shc0040493, 32'shc003fbb0, 32'shc003f2d8, 32'shc003ea09, 32'shc003e143, 32'shc003d888, 32'shc003cfd7, 
               32'shc003c72f, 32'shc003be91, 32'shc003b5fe, 32'shc003ad74, 32'shc003a4f4, 32'shc0039c7d, 32'shc0039411, 32'shc0038baf, 
               32'shc0038356, 32'shc0037b07, 32'shc00372c2, 32'shc0036a87, 32'shc0036256, 32'shc0035a2f, 32'shc0035211, 32'shc00349fe, 
               32'shc00341f4, 32'shc00339f4, 32'shc00331fe, 32'shc0032a12, 32'shc0032230, 32'shc0031a58, 32'shc0031289, 32'shc0030ac5, 
               32'shc003030a, 32'shc002fb59, 32'shc002f3b2, 32'shc002ec15, 32'shc002e482, 32'shc002dcf8, 32'shc002d579, 32'shc002ce03, 
               32'shc002c697, 32'shc002bf35, 32'shc002b7dd, 32'shc002b08f, 32'shc002a94b, 32'shc002a210, 32'shc0029ae0, 32'shc00293b9, 
               32'shc0028c9c, 32'shc0028589, 32'shc0027e80, 32'shc0027781, 32'shc002708c, 32'shc00269a0, 32'shc00262be, 32'shc0025be7, 
               32'shc0025519, 32'shc0024e55, 32'shc002479b, 32'shc00240ea, 32'shc0023a44, 32'shc00233a7, 32'shc0022d15, 32'shc002268c, 
               32'shc002200d, 32'shc0021998, 32'shc002132d, 32'shc0020ccb, 32'shc0020674, 32'shc0020026, 32'shc001f9e2, 32'shc001f3a8, 
               32'shc001ed78, 32'shc001e752, 32'shc001e136, 32'shc001db24, 32'shc001d51b, 32'shc001cf1c, 32'shc001c928, 32'shc001c33d, 
               32'shc001bd5c, 32'shc001b784, 32'shc001b1b7, 32'shc001abf4, 32'shc001a63a, 32'shc001a08a, 32'shc0019ae5, 32'shc0019549, 
               32'shc0018fb6, 32'shc0018a2e, 32'shc00184b0, 32'shc0017f3b, 32'shc00179d1, 32'shc0017470, 32'shc0016f19, 32'shc00169cc, 
               32'shc0016489, 32'shc0015f50, 32'shc0015a20, 32'shc00154fb, 32'shc0014fdf, 32'shc0014acd, 32'shc00145c5, 32'shc00140c7, 
               32'shc0013bd3, 32'shc00136e8, 32'shc0013208, 32'shc0012d31, 32'shc0012865, 32'shc00123a2, 32'shc0011ee9, 32'shc0011a3a, 
               32'shc0011594, 32'shc00110f9, 32'shc0010c67, 32'shc00107e0, 32'shc0010362, 32'shc000feee, 32'shc000fa84, 32'shc000f624, 
               32'shc000f1ce, 32'shc000ed81, 32'shc000e93f, 32'shc000e506, 32'shc000e0d7, 32'shc000dcb2, 32'shc000d897, 32'shc000d486, 
               32'shc000d07e, 32'shc000cc81, 32'shc000c88d, 32'shc000c4a4, 32'shc000c0c4, 32'shc000bcee, 32'shc000b921, 32'shc000b55f, 
               32'shc000b1a7, 32'shc000adf8, 32'shc000aa54, 32'shc000a6b9, 32'shc000a328, 32'shc0009fa1, 32'shc0009c24, 32'shc00098b0, 
               32'shc0009547, 32'shc00091e7, 32'shc0008e92, 32'shc0008b46, 32'shc0008804, 32'shc00084cc, 32'shc000819d, 32'shc0007e79, 
               32'shc0007b5f, 32'shc000784e, 32'shc0007547, 32'shc000724a, 32'shc0006f57, 32'shc0006c6e, 32'shc000698f, 32'shc00066b9, 
               32'shc00063ee, 32'shc000612c, 32'shc0005e74, 32'shc0005bc7, 32'shc0005922, 32'shc0005688, 32'shc00053f8, 32'shc0005171, 
               32'shc0004ef5, 32'shc0004c82, 32'shc0004a19, 32'shc00047ba, 32'shc0004565, 32'shc000431a, 32'shc00040d9, 32'shc0003ea1, 
               32'shc0003c74, 32'shc0003a50, 32'shc0003836, 32'shc0003626, 32'shc0003420, 32'shc0003223, 32'shc0003031, 32'shc0002e48, 
               32'shc0002c6a, 32'shc0002a95, 32'shc00028ca, 32'shc0002709, 32'shc0002552, 32'shc00023a4, 32'shc0002201, 32'shc0002067, 
               32'shc0001ed8, 32'shc0001d52, 32'shc0001bd6, 32'shc0001a64, 32'shc00018fb, 32'shc000179d, 32'shc0001649, 32'shc00014fe, 
               32'shc00013bd, 32'shc0001286, 32'shc0001159, 32'shc0001036, 32'shc0000f1d, 32'shc0000e0d, 32'shc0000d08, 32'shc0000c0c, 
               32'shc0000b1a, 32'shc0000a33, 32'shc0000954, 32'shc0000880, 32'shc00007b6, 32'shc00006f5, 32'shc000063f, 32'shc0000592, 
               32'shc00004ef, 32'shc0000456, 32'shc00003c7, 32'shc0000342, 32'shc00002c7, 32'shc0000255, 32'shc00001ed, 32'shc0000190, 
               32'shc000013c, 32'shc00000f2, 32'shc00000b2, 32'shc000007b, 32'shc000004f, 32'shc000002c, 32'shc0000014, 32'shc0000005
            };

            reg signed [31:0] W_Im_table[32768] = '{
               32'sh00000000, 32'shfffe6de0, 32'shfffcdbc1, 32'shfffb49a1, 32'shfff9b781, 32'shfff82561, 32'shfff69342, 32'shfff50122, 
               32'shfff36f02, 32'shfff1dce3, 32'shfff04ac3, 32'shffeeb8a3, 32'shffed2684, 32'shffeb9464, 32'shffea0245, 32'shffe87025, 
               32'shffe6de05, 32'shffe54be6, 32'shffe3b9c6, 32'shffe227a7, 32'shffe09587, 32'shffdf0368, 32'shffdd7148, 32'shffdbdf29, 
               32'shffda4d09, 32'shffd8baea, 32'shffd728ca, 32'shffd596ab, 32'shffd4048c, 32'shffd2726c, 32'shffd0e04d, 32'shffcf4e2e, 
               32'shffcdbc0f, 32'shffcc29ef, 32'shffca97d0, 32'shffc905b1, 32'shffc77392, 32'shffc5e173, 32'shffc44f54, 32'shffc2bd35, 
               32'shffc12b16, 32'shffbf98f7, 32'shffbe06d8, 32'shffbc74b9, 32'shffbae29a, 32'shffb9507c, 32'shffb7be5d, 32'shffb62c3e, 
               32'shffb49a1f, 32'shffb30801, 32'shffb175e2, 32'shffafe3c4, 32'shffae51a5, 32'shffacbf87, 32'shffab2d69, 32'shffa99b4a, 
               32'shffa8092c, 32'shffa6770e, 32'shffa4e4f0, 32'shffa352d2, 32'shffa1c0b4, 32'shffa02e96, 32'shff9e9c78, 32'shff9d0a5a, 
               32'shff9b783c, 32'shff99e61e, 32'shff985401, 32'shff96c1e3, 32'shff952fc5, 32'shff939da8, 32'shff920b8b, 32'shff90796d, 
               32'shff8ee750, 32'shff8d5533, 32'shff8bc316, 32'shff8a30f8, 32'shff889edb, 32'shff870cbe, 32'shff857aa2, 32'shff83e885, 
               32'shff825668, 32'shff80c44b, 32'shff7f322f, 32'shff7da012, 32'shff7c0df6, 32'shff7a7bda, 32'shff78e9bd, 32'shff7757a1, 
               32'shff75c585, 32'shff743369, 32'shff72a14d, 32'shff710f31, 32'shff6f7d16, 32'shff6deafa, 32'shff6c58de, 32'shff6ac6c3, 
               32'shff6934a8, 32'shff67a28c, 32'shff661071, 32'shff647e56, 32'shff62ec3b, 32'shff615a20, 32'shff5fc805, 32'shff5e35ea, 
               32'shff5ca3d0, 32'shff5b11b5, 32'shff597f9b, 32'shff57ed80, 32'shff565b66, 32'shff54c94c, 32'shff533732, 32'shff51a518, 
               32'shff5012fe, 32'shff4e80e5, 32'shff4ceecb, 32'shff4b5cb1, 32'shff49ca98, 32'shff48387f, 32'shff46a666, 32'shff45144c, 
               32'shff438234, 32'shff41f01b, 32'shff405e02, 32'shff3ecbe9, 32'shff3d39d1, 32'shff3ba7b9, 32'shff3a15a0, 32'shff388388, 
               32'shff36f170, 32'shff355f58, 32'shff33cd40, 32'shff323b29, 32'shff30a911, 32'shff2f16fa, 32'shff2d84e3, 32'shff2bf2cb, 
               32'shff2a60b4, 32'shff28ce9e, 32'shff273c87, 32'shff25aa70, 32'shff24185a, 32'shff228643, 32'shff20f42d, 32'shff1f6217, 
               32'shff1dd001, 32'shff1c3deb, 32'shff1aabd5, 32'shff1919c0, 32'shff1787aa, 32'shff15f595, 32'shff146380, 32'shff12d16b, 
               32'shff113f56, 32'shff0fad41, 32'shff0e1b2d, 32'shff0c8919, 32'shff0af704, 32'shff0964f0, 32'shff07d2dc, 32'shff0640c8, 
               32'shff04aeb5, 32'shff031ca1, 32'shff018a8e, 32'shfefff87b, 32'shfefe6668, 32'shfefcd455, 32'shfefb4242, 32'shfef9b02f, 
               32'shfef81e1d, 32'shfef68c0b, 32'shfef4f9f8, 32'shfef367e6, 32'shfef1d5d5, 32'shfef043c3, 32'shfeeeb1b2, 32'shfeed1fa0, 
               32'shfeeb8d8f, 32'shfee9fb7e, 32'shfee8696d, 32'shfee6d75d, 32'shfee5454c, 32'shfee3b33c, 32'shfee2212c, 32'shfee08f1c, 
               32'shfedefd0c, 32'shfedd6afd, 32'shfedbd8ed, 32'shfeda46de, 32'shfed8b4cf, 32'shfed722c0, 32'shfed590b1, 32'shfed3fea3, 
               32'shfed26c94, 32'shfed0da86, 32'shfecf4878, 32'shfecdb66a, 32'shfecc245d, 32'shfeca924f, 32'shfec90042, 32'shfec76e35, 
               32'shfec5dc28, 32'shfec44a1b, 32'shfec2b80f, 32'shfec12603, 32'shfebf93f6, 32'shfebe01ea, 32'shfebc6fdf, 32'shfebaddd3, 
               32'shfeb94bc8, 32'shfeb7b9bd, 32'shfeb627b2, 32'shfeb495a7, 32'shfeb3039d, 32'shfeb17192, 32'shfeafdf88, 32'shfeae4d7e, 
               32'shfeacbb74, 32'shfeab296b, 32'shfea99761, 32'shfea80558, 32'shfea6734f, 32'shfea4e147, 32'shfea34f3e, 32'shfea1bd36, 
               32'shfea02b2e, 32'shfe9e9926, 32'shfe9d071e, 32'shfe9b7517, 32'shfe99e310, 32'shfe985109, 32'shfe96bf02, 32'shfe952cfb, 
               32'shfe939af5, 32'shfe9208ef, 32'shfe9076e9, 32'shfe8ee4e3, 32'shfe8d52de, 32'shfe8bc0d9, 32'shfe8a2ed4, 32'shfe889ccf, 
               32'shfe870aca, 32'shfe8578c6, 32'shfe83e6c2, 32'shfe8254be, 32'shfe80c2ba, 32'shfe7f30b7, 32'shfe7d9eb4, 32'shfe7c0cb1, 
               32'shfe7a7aae, 32'shfe78e8ab, 32'shfe7756a9, 32'shfe75c4a7, 32'shfe7432a5, 32'shfe72a0a4, 32'shfe710ea2, 32'shfe6f7ca1, 
               32'shfe6deaa1, 32'shfe6c58a0, 32'shfe6ac6a0, 32'shfe6934a0, 32'shfe67a2a0, 32'shfe6610a0, 32'shfe647ea1, 32'shfe62eca2, 
               32'shfe615aa3, 32'shfe5fc8a4, 32'shfe5e36a6, 32'shfe5ca4a8, 32'shfe5b12aa, 32'shfe5980ac, 32'shfe57eeaf, 32'shfe565cb2, 
               32'shfe54cab5, 32'shfe5338b8, 32'shfe51a6bc, 32'shfe5014c0, 32'shfe4e82c4, 32'shfe4cf0c9, 32'shfe4b5ecd, 32'shfe49ccd2, 
               32'shfe483ad8, 32'shfe46a8dd, 32'shfe4516e3, 32'shfe4384e9, 32'shfe41f2ef, 32'shfe4060f6, 32'shfe3ecefd, 32'shfe3d3d04, 
               32'shfe3bab0b, 32'shfe3a1913, 32'shfe38871b, 32'shfe36f523, 32'shfe35632c, 32'shfe33d134, 32'shfe323f3d, 32'shfe30ad47, 
               32'shfe2f1b50, 32'shfe2d895a, 32'shfe2bf764, 32'shfe2a656f, 32'shfe28d379, 32'shfe274184, 32'shfe25af90, 32'shfe241d9b, 
               32'shfe228ba7, 32'shfe20f9b3, 32'shfe1f67c0, 32'shfe1dd5cd, 32'shfe1c43da, 32'shfe1ab1e7, 32'shfe191ff5, 32'shfe178e02, 
               32'shfe15fc11, 32'shfe146a1f, 32'shfe12d82e, 32'shfe11463d, 32'shfe0fb44c, 32'shfe0e225c, 32'shfe0c906c, 32'shfe0afe7c, 
               32'shfe096c8d, 32'shfe07da9e, 32'shfe0648af, 32'shfe04b6c0, 32'shfe0324d2, 32'shfe0192e4, 32'shfe0000f7, 32'shfdfe6f0a, 
               32'shfdfcdd1d, 32'shfdfb4b30, 32'shfdf9b944, 32'shfdf82758, 32'shfdf6956c, 32'shfdf50380, 32'shfdf37195, 32'shfdf1dfab, 
               32'shfdf04dc0, 32'shfdeebbd6, 32'shfded29ec, 32'shfdeb9803, 32'shfdea0619, 32'shfde87431, 32'shfde6e248, 32'shfde55060, 
               32'shfde3be78, 32'shfde22c90, 32'shfde09aa9, 32'shfddf08c2, 32'shfddd76dc, 32'shfddbe4f5, 32'shfdda530f, 32'shfdd8c12a, 
               32'shfdd72f45, 32'shfdd59d60, 32'shfdd40b7b, 32'shfdd27997, 32'shfdd0e7b3, 32'shfdcf55cf, 32'shfdcdc3ec, 32'shfdcc3209, 
               32'shfdcaa027, 32'shfdc90e44, 32'shfdc77c62, 32'shfdc5ea81, 32'shfdc458a0, 32'shfdc2c6bf, 32'shfdc134de, 32'shfdbfa2fe, 
               32'shfdbe111e, 32'shfdbc7f3f, 32'shfdbaed60, 32'shfdb95b81, 32'shfdb7c9a3, 32'shfdb637c5, 32'shfdb4a5e7, 32'shfdb31409, 
               32'shfdb1822c, 32'shfdaff050, 32'shfdae5e74, 32'shfdaccc98, 32'shfdab3abc, 32'shfda9a8e1, 32'shfda81706, 32'shfda6852b, 
               32'shfda4f351, 32'shfda36178, 32'shfda1cf9e, 32'shfda03dc5, 32'shfd9eabec, 32'shfd9d1a14, 32'shfd9b883c, 32'shfd99f665, 
               32'shfd98648d, 32'shfd96d2b7, 32'shfd9540e0, 32'shfd93af0a, 32'shfd921d34, 32'shfd908b5f, 32'shfd8ef98a, 32'shfd8d67b5, 
               32'shfd8bd5e1, 32'shfd8a440d, 32'shfd88b23a, 32'shfd872067, 32'shfd858e94, 32'shfd83fcc2, 32'shfd826af0, 32'shfd80d91e, 
               32'shfd7f474d, 32'shfd7db57c, 32'shfd7c23ac, 32'shfd7a91dc, 32'shfd79000d, 32'shfd776e3d, 32'shfd75dc6e, 32'shfd744aa0, 
               32'shfd72b8d2, 32'shfd712704, 32'shfd6f9537, 32'shfd6e036a, 32'shfd6c719e, 32'shfd6adfd2, 32'shfd694e06, 32'shfd67bc3b, 
               32'shfd662a70, 32'shfd6498a5, 32'shfd6306db, 32'shfd617512, 32'shfd5fe348, 32'shfd5e5180, 32'shfd5cbfb7, 32'shfd5b2def, 
               32'shfd599c28, 32'shfd580a60, 32'shfd56789a, 32'shfd54e6d3, 32'shfd53550d, 32'shfd51c348, 32'shfd503182, 32'shfd4e9fbe, 
               32'shfd4d0df9, 32'shfd4b7c35, 32'shfd49ea72, 32'shfd4858af, 32'shfd46c6ec, 32'shfd45352a, 32'shfd43a368, 32'shfd4211a7, 
               32'shfd407fe6, 32'shfd3eee25, 32'shfd3d5c65, 32'shfd3bcaa5, 32'shfd3a38e6, 32'shfd38a727, 32'shfd371569, 32'shfd3583ab, 
               32'shfd33f1ed, 32'shfd326030, 32'shfd30ce73, 32'shfd2f3cb7, 32'shfd2daafb, 32'shfd2c1940, 32'shfd2a8785, 32'shfd28f5ca, 
               32'shfd276410, 32'shfd25d257, 32'shfd24409d, 32'shfd22aee5, 32'shfd211d2c, 32'shfd1f8b74, 32'shfd1df9bd, 32'shfd1c6806, 
               32'shfd1ad650, 32'shfd194499, 32'shfd17b2e4, 32'shfd16212f, 32'shfd148f7a, 32'shfd12fdc6, 32'shfd116c12, 32'shfd0fda5e, 
               32'shfd0e48ab, 32'shfd0cb6f9, 32'shfd0b2547, 32'shfd099395, 32'shfd0801e4, 32'shfd067033, 32'shfd04de83, 32'shfd034cd3, 
               32'shfd01bb24, 32'shfd002975, 32'shfcfe97c7, 32'shfcfd0619, 32'shfcfb746c, 32'shfcf9e2bf, 32'shfcf85112, 32'shfcf6bf66, 
               32'shfcf52dbb, 32'shfcf39c0f, 32'shfcf20a65, 32'shfcf078bb, 32'shfceee711, 32'shfced5568, 32'shfcebc3bf, 32'shfcea3217, 
               32'shfce8a06f, 32'shfce70ec8, 32'shfce57d21, 32'shfce3eb7a, 32'shfce259d5, 32'shfce0c82f, 32'shfcdf368a, 32'shfcdda4e6, 
               32'shfcdc1342, 32'shfcda819e, 32'shfcd8effb, 32'shfcd75e59, 32'shfcd5ccb7, 32'shfcd43b15, 32'shfcd2a974, 32'shfcd117d4, 
               32'shfccf8634, 32'shfccdf494, 32'shfccc62f5, 32'shfccad157, 32'shfcc93fb9, 32'shfcc7ae1b, 32'shfcc61c7e, 32'shfcc48ae1, 
               32'shfcc2f945, 32'shfcc167aa, 32'shfcbfd60e, 32'shfcbe4474, 32'shfcbcb2da, 32'shfcbb2140, 32'shfcb98fa7, 32'shfcb7fe0f, 
               32'shfcb66c77, 32'shfcb4dadf, 32'shfcb34948, 32'shfcb1b7b1, 32'shfcb0261b, 32'shfcae9486, 32'shfcad02f1, 32'shfcab715c, 
               32'shfca9dfc8, 32'shfca84e35, 32'shfca6bca2, 32'shfca52b0f, 32'shfca3997e, 32'shfca207ec, 32'shfca0765b, 32'shfc9ee4cb, 
               32'shfc9d533b, 32'shfc9bc1ac, 32'shfc9a301d, 32'shfc989e8f, 32'shfc970d01, 32'shfc957b74, 32'shfc93e9e7, 32'shfc92585b, 
               32'shfc90c6cf, 32'shfc8f3544, 32'shfc8da3ba, 32'shfc8c122f, 32'shfc8a80a6, 32'shfc88ef1d, 32'shfc875d95, 32'shfc85cc0d, 
               32'shfc843a85, 32'shfc82a8fe, 32'shfc811778, 32'shfc7f85f2, 32'shfc7df46d, 32'shfc7c62e8, 32'shfc7ad164, 32'shfc793fe1, 
               32'shfc77ae5e, 32'shfc761cdb, 32'shfc748b59, 32'shfc72f9d8, 32'shfc716857, 32'shfc6fd6d7, 32'shfc6e4557, 32'shfc6cb3d8, 
               32'shfc6b2259, 32'shfc6990db, 32'shfc67ff5d, 32'shfc666de0, 32'shfc64dc64, 32'shfc634ae8, 32'shfc61b96d, 32'shfc6027f2, 
               32'shfc5e9678, 32'shfc5d04fe, 32'shfc5b7385, 32'shfc59e20c, 32'shfc585094, 32'shfc56bf1d, 32'shfc552da6, 32'shfc539c30, 
               32'shfc520aba, 32'shfc507945, 32'shfc4ee7d0, 32'shfc4d565c, 32'shfc4bc4e9, 32'shfc4a3376, 32'shfc48a204, 32'shfc471092, 
               32'shfc457f21, 32'shfc43edb0, 32'shfc425c40, 32'shfc40cad1, 32'shfc3f3962, 32'shfc3da7f4, 32'shfc3c1686, 32'shfc3a8519, 
               32'shfc38f3ac, 32'shfc376240, 32'shfc35d0d5, 32'shfc343f6a, 32'shfc32ae00, 32'shfc311c97, 32'shfc2f8b2e, 32'shfc2df9c5, 
               32'shfc2c685d, 32'shfc2ad6f6, 32'shfc29458f, 32'shfc27b429, 32'shfc2622c4, 32'shfc24915f, 32'shfc22fffb, 32'shfc216e97, 
               32'shfc1fdd34, 32'shfc1e4bd1, 32'shfc1cba6f, 32'shfc1b290e, 32'shfc1997ae, 32'shfc18064d, 32'shfc1674ee, 32'shfc14e38f, 
               32'shfc135231, 32'shfc11c0d3, 32'shfc102f76, 32'shfc0e9e1a, 32'shfc0d0cbe, 32'shfc0b7b62, 32'shfc09ea08, 32'shfc0858ae, 
               32'shfc06c754, 32'shfc0535fc, 32'shfc03a4a3, 32'shfc02134c, 32'shfc0081f5, 32'shfbfef09f, 32'shfbfd5f49, 32'shfbfbcdf4, 
               32'shfbfa3c9f, 32'shfbf8ab4b, 32'shfbf719f8, 32'shfbf588a5, 32'shfbf3f753, 32'shfbf26602, 32'shfbf0d4b1, 32'shfbef4361, 
               32'shfbedb212, 32'shfbec20c3, 32'shfbea8f75, 32'shfbe8fe27, 32'shfbe76cda, 32'shfbe5db8e, 32'shfbe44a42, 32'shfbe2b8f7, 
               32'shfbe127ac, 32'shfbdf9663, 32'shfbde0519, 32'shfbdc73d1, 32'shfbdae289, 32'shfbd95142, 32'shfbd7bffb, 32'shfbd62eb5, 
               32'shfbd49d70, 32'shfbd30c2b, 32'shfbd17ae7, 32'shfbcfe9a4, 32'shfbce5861, 32'shfbccc71f, 32'shfbcb35dd, 32'shfbc9a49d, 
               32'shfbc8135c, 32'shfbc6821d, 32'shfbc4f0de, 32'shfbc35fa0, 32'shfbc1ce62, 32'shfbc03d25, 32'shfbbeabe9, 32'shfbbd1aad, 
               32'shfbbb8973, 32'shfbb9f838, 32'shfbb866ff, 32'shfbb6d5c6, 32'shfbb5448d, 32'shfbb3b356, 32'shfbb2221f, 32'shfbb090e8, 
               32'shfbaeffb3, 32'shfbad6e7e, 32'shfbabdd49, 32'shfbaa4c16, 32'shfba8bae3, 32'shfba729b1, 32'shfba5987f, 32'shfba4074e, 
               32'shfba2761e, 32'shfba0e4ee, 32'shfb9f53bf, 32'shfb9dc291, 32'shfb9c3163, 32'shfb9aa036, 32'shfb990f0a, 32'shfb977ddf, 
               32'shfb95ecb4, 32'shfb945b89, 32'shfb92ca60, 32'shfb913937, 32'shfb8fa80f, 32'shfb8e16e7, 32'shfb8c85c1, 32'shfb8af49b, 
               32'shfb896375, 32'shfb87d250, 32'shfb86412c, 32'shfb84b009, 32'shfb831ee6, 32'shfb818dc4, 32'shfb7ffca3, 32'shfb7e6b83, 
               32'shfb7cda63, 32'shfb7b4944, 32'shfb79b825, 32'shfb782707, 32'shfb7695ea, 32'shfb7504ce, 32'shfb7373b2, 32'shfb71e297, 
               32'shfb70517d, 32'shfb6ec063, 32'shfb6d2f4a, 32'shfb6b9e32, 32'shfb6a0d1b, 32'shfb687c04, 32'shfb66eaee, 32'shfb6559d9, 
               32'shfb63c8c4, 32'shfb6237b0, 32'shfb60a69d, 32'shfb5f158a, 32'shfb5d8479, 32'shfb5bf368, 32'shfb5a6257, 32'shfb58d148, 
               32'shfb574039, 32'shfb55af2a, 32'shfb541e1d, 32'shfb528d10, 32'shfb50fc04, 32'shfb4f6af9, 32'shfb4dd9ee, 32'shfb4c48e4, 
               32'shfb4ab7db, 32'shfb4926d3, 32'shfb4795cb, 32'shfb4604c4, 32'shfb4473be, 32'shfb42e2b9, 32'shfb4151b4, 32'shfb3fc0b0, 
               32'shfb3e2fac, 32'shfb3c9eaa, 32'shfb3b0da8, 32'shfb397ca7, 32'shfb37eba7, 32'shfb365aa7, 32'shfb34c9a8, 32'shfb3338aa, 
               32'shfb31a7ac, 32'shfb3016b0, 32'shfb2e85b4, 32'shfb2cf4b9, 32'shfb2b63be, 32'shfb29d2c5, 32'shfb2841cc, 32'shfb26b0d3, 
               32'shfb251fdc, 32'shfb238ee5, 32'shfb21fdef, 32'shfb206cfa, 32'shfb1edc06, 32'shfb1d4b12, 32'shfb1bba1f, 32'shfb1a292d, 
               32'shfb18983b, 32'shfb17074b, 32'shfb15765b, 32'shfb13e56c, 32'shfb12547d, 32'shfb10c38f, 32'shfb0f32a3, 32'shfb0da1b6, 
               32'shfb0c10cb, 32'shfb0a7fe1, 32'shfb08eef7, 32'shfb075e0e, 32'shfb05cd25, 32'shfb043c3e, 32'shfb02ab57, 32'shfb011a71, 
               32'shfaff898c, 32'shfafdf8a7, 32'shfafc67c4, 32'shfafad6e1, 32'shfaf945ff, 32'shfaf7b51d, 32'shfaf6243d, 32'shfaf4935d, 
               32'shfaf3027e, 32'shfaf171a0, 32'shfaefe0c2, 32'shfaee4fe5, 32'shfaecbf0a, 32'shfaeb2e2e, 32'shfae99d54, 32'shfae80c7a, 
               32'shfae67ba2, 32'shfae4eaca, 32'shfae359f3, 32'shfae1c91c, 32'shfae03847, 32'shfadea772, 32'shfadd169e, 32'shfadb85ca, 
               32'shfad9f4f8, 32'shfad86426, 32'shfad6d355, 32'shfad54285, 32'shfad3b1b6, 32'shfad220e8, 32'shfad0901a, 32'shfaceff4d, 
               32'shfacd6e81, 32'shfacbddb6, 32'shfaca4ceb, 32'shfac8bc22, 32'shfac72b59, 32'shfac59a91, 32'shfac409c9, 32'shfac27903, 
               32'shfac0e83d, 32'shfabf5778, 32'shfabdc6b4, 32'shfabc35f1, 32'shfabaa52f, 32'shfab9146d, 32'shfab783ad, 32'shfab5f2ed, 
               32'shfab4622d, 32'shfab2d16f, 32'shfab140b2, 32'shfaafaff5, 32'shfaae1f39, 32'shfaac8e7e, 32'shfaaafdc4, 32'shfaa96d0a, 
               32'shfaa7dc52, 32'shfaa64b9a, 32'shfaa4bae3, 32'shfaa32a2d, 32'shfaa19978, 32'shfaa008c3, 32'shfa9e7810, 32'shfa9ce75d, 
               32'shfa9b56ab, 32'shfa99c5fa, 32'shfa98354a, 32'shfa96a49a, 32'shfa9513eb, 32'shfa93833e, 32'shfa91f291, 32'shfa9061e5, 
               32'shfa8ed139, 32'shfa8d408f, 32'shfa8bafe5, 32'shfa8a1f3c, 32'shfa888e95, 32'shfa86fded, 32'shfa856d47, 32'shfa83dca2, 
               32'shfa824bfd, 32'shfa80bb5a, 32'shfa7f2ab7, 32'shfa7d9a15, 32'shfa7c0974, 32'shfa7a78d3, 32'shfa78e834, 32'shfa775795, 
               32'shfa75c6f8, 32'shfa74365b, 32'shfa72a5bf, 32'shfa711524, 32'shfa6f8489, 32'shfa6df3f0, 32'shfa6c6357, 32'shfa6ad2bf, 
               32'shfa694229, 32'shfa67b193, 32'shfa6620fd, 32'shfa649069, 32'shfa62ffd6, 32'shfa616f43, 32'shfa5fdeb1, 32'shfa5e4e21, 
               32'shfa5cbd91, 32'shfa5b2d02, 32'shfa599c73, 32'shfa580be6, 32'shfa567b5a, 32'shfa54eace, 32'shfa535a43, 32'shfa51c9b9, 
               32'shfa503930, 32'shfa4ea8a8, 32'shfa4d1821, 32'shfa4b879b, 32'shfa49f715, 32'shfa486691, 32'shfa46d60d, 32'shfa45458a, 
               32'shfa43b508, 32'shfa422487, 32'shfa409407, 32'shfa3f0388, 32'shfa3d7309, 32'shfa3be28c, 32'shfa3a520f, 32'shfa38c194, 
               32'shfa373119, 32'shfa35a09f, 32'shfa341026, 32'shfa327fae, 32'shfa30ef36, 32'shfa2f5ec0, 32'shfa2dce4b, 32'shfa2c3dd6, 
               32'shfa2aad62, 32'shfa291cf0, 32'shfa278c7e, 32'shfa25fc0d, 32'shfa246b9d, 32'shfa22db2d, 32'shfa214abf, 32'shfa1fba52, 
               32'shfa1e29e5, 32'shfa1c997a, 32'shfa1b090f, 32'shfa1978a6, 32'shfa17e83d, 32'shfa1657d5, 32'shfa14c76e, 32'shfa133708, 
               32'shfa11a6a3, 32'shfa10163e, 32'shfa0e85db, 32'shfa0cf579, 32'shfa0b6517, 32'shfa09d4b7, 32'shfa084457, 32'shfa06b3f8, 
               32'shfa05239a, 32'shfa03933d, 32'shfa0202e1, 32'shfa007286, 32'shf9fee22c, 32'shf9fd51d3, 32'shf9fbc17b, 32'shf9fa3123, 
               32'shf9f8a0cd, 32'shf9f71078, 32'shf9f58023, 32'shf9f3efcf, 32'shf9f25f7d, 32'shf9f0cf2b, 32'shf9ef3eda, 32'shf9edae8a, 
               32'shf9ec1e3b, 32'shf9ea8ded, 32'shf9e8fda0, 32'shf9e76d54, 32'shf9e5dd09, 32'shf9e44cbf, 32'shf9e2bc75, 32'shf9e12c2d, 
               32'shf9df9be6, 32'shf9de0b9f, 32'shf9dc7b5a, 32'shf9daeb15, 32'shf9d95ad1, 32'shf9d7ca8f, 32'shf9d63a4d, 32'shf9d4aa0c, 
               32'shf9d319cc, 32'shf9d1898d, 32'shf9cff94f, 32'shf9ce6912, 32'shf9ccd8d6, 32'shf9cb489b, 32'shf9c9b861, 32'shf9c82828, 
               32'shf9c697f0, 32'shf9c507b9, 32'shf9c37782, 32'shf9c1e74d, 32'shf9c05719, 32'shf9bec6e5, 32'shf9bd36b3, 32'shf9bba681, 
               32'shf9ba1651, 32'shf9b88621, 32'shf9b6f5f3, 32'shf9b565c5, 32'shf9b3d599, 32'shf9b2456d, 32'shf9b0b542, 32'shf9af2519, 
               32'shf9ad94f0, 32'shf9ac04c8, 32'shf9aa74a1, 32'shf9a8e47c, 32'shf9a75457, 32'shf9a5c433, 32'shf9a43410, 32'shf9a2a3ee, 
               32'shf9a113cd, 32'shf99f83ad, 32'shf99df38e, 32'shf99c6371, 32'shf99ad354, 32'shf9994338, 32'shf997b31d, 32'shf9962303, 
               32'shf99492ea, 32'shf99302d2, 32'shf99172bb, 32'shf98fe2a5, 32'shf98e528f, 32'shf98cc27b, 32'shf98b3268, 32'shf989a256, 
               32'shf9881245, 32'shf9868235, 32'shf984f226, 32'shf9836218, 32'shf981d20b, 32'shf98041ff, 32'shf97eb1f4, 32'shf97d21ea, 
               32'shf97b91e1, 32'shf97a01d9, 32'shf97871d2, 32'shf976e1cc, 32'shf97551c6, 32'shf973c1c2, 32'shf97231bf, 32'shf970a1bd, 
               32'shf96f11bc, 32'shf96d81bc, 32'shf96bf1be, 32'shf96a61c0, 32'shf968d1c3, 32'shf96741c7, 32'shf965b1cc, 32'shf96421d2, 
               32'shf96291d9, 32'shf96101e1, 32'shf95f71ea, 32'shf95de1f5, 32'shf95c5200, 32'shf95ac20c, 32'shf9593219, 32'shf957a228, 
               32'shf9561237, 32'shf9548247, 32'shf952f259, 32'shf951626b, 32'shf94fd27f, 32'shf94e4293, 32'shf94cb2a8, 32'shf94b22bf, 
               32'shf94992d7, 32'shf94802ef, 32'shf9467309, 32'shf944e323, 32'shf943533f, 32'shf941c35c, 32'shf940337a, 32'shf93ea399, 
               32'shf93d13b8, 32'shf93b83d9, 32'shf939f3fb, 32'shf938641e, 32'shf936d442, 32'shf9354468, 32'shf933b48e, 32'shf93224b5, 
               32'shf93094dd, 32'shf92f0506, 32'shf92d7531, 32'shf92be55c, 32'shf92a5589, 32'shf928c5b6, 32'shf92735e5, 32'shf925a614, 
               32'shf9241645, 32'shf9228677, 32'shf920f6a9, 32'shf91f66dd, 32'shf91dd712, 32'shf91c4748, 32'shf91ab77f, 32'shf91927b7, 
               32'shf91797f0, 32'shf916082b, 32'shf9147866, 32'shf912e8a2, 32'shf91158e0, 32'shf90fc91e, 32'shf90e395e, 32'shf90ca99e, 
               32'shf90b19e0, 32'shf9098a23, 32'shf907fa67, 32'shf9066aac, 32'shf904daf2, 32'shf9034b39, 32'shf901bb81, 32'shf9002bca, 
               32'shf8fe9c15, 32'shf8fd0c60, 32'shf8fb7cac, 32'shf8f9ecfa, 32'shf8f85d49, 32'shf8f6cd98, 32'shf8f53de9, 32'shf8f3ae3b, 
               32'shf8f21e8e, 32'shf8f08ee2, 32'shf8eeff37, 32'shf8ed6f8e, 32'shf8ebdfe5, 32'shf8ea503d, 32'shf8e8c097, 32'shf8e730f2, 
               32'shf8e5a14d, 32'shf8e411aa, 32'shf8e28208, 32'shf8e0f267, 32'shf8df62c7, 32'shf8ddd328, 32'shf8dc438b, 32'shf8dab3ee, 
               32'shf8d92452, 32'shf8d794b8, 32'shf8d6051f, 32'shf8d47587, 32'shf8d2e5f0, 32'shf8d1565a, 32'shf8cfc6c5, 32'shf8ce3731, 
               32'shf8cca79e, 32'shf8cb180d, 32'shf8c9887c, 32'shf8c7f8ed, 32'shf8c6695f, 32'shf8c4d9d2, 32'shf8c34a46, 32'shf8c1babb, 
               32'shf8c02b31, 32'shf8be9ba9, 32'shf8bd0c21, 32'shf8bb7c9b, 32'shf8b9ed15, 32'shf8b85d91, 32'shf8b6ce0e, 32'shf8b53e8c, 
               32'shf8b3af0c, 32'shf8b21f8c, 32'shf8b0900d, 32'shf8af0090, 32'shf8ad7114, 32'shf8abe199, 32'shf8aa521f, 32'shf8a8c2a6, 
               32'shf8a7332e, 32'shf8a5a3b8, 32'shf8a41442, 32'shf8a284ce, 32'shf8a0f55b, 32'shf89f65e8, 32'shf89dd678, 32'shf89c4708, 
               32'shf89ab799, 32'shf899282c, 32'shf89798bf, 32'shf8960954, 32'shf89479ea, 32'shf892ea81, 32'shf8915b19, 32'shf88fcbb3, 
               32'shf88e3c4d, 32'shf88cace9, 32'shf88b1d86, 32'shf8898e23, 32'shf887fec3, 32'shf8866f63, 32'shf884e004, 32'shf88350a7, 
               32'shf881c14b, 32'shf88031ef, 32'shf87ea295, 32'shf87d133d, 32'shf87b83e5, 32'shf879f48e, 32'shf8786539, 32'shf876d5e5, 
               32'shf8754692, 32'shf873b740, 32'shf87227ef, 32'shf87098a0, 32'shf86f0952, 32'shf86d7a04, 32'shf86beab8, 32'shf86a5b6d, 
               32'shf868cc24, 32'shf8673cdb, 32'shf865ad94, 32'shf8641e4e, 32'shf8628f09, 32'shf860ffc5, 32'shf85f7082, 32'shf85de141, 
               32'shf85c5201, 32'shf85ac2c1, 32'shf8593383, 32'shf857a447, 32'shf856150b, 32'shf85485d1, 32'shf852f698, 32'shf8516760, 
               32'shf84fd829, 32'shf84e48f3, 32'shf84cb9bf, 32'shf84b2a8b, 32'shf8499b59, 32'shf8480c28, 32'shf8467cf9, 32'shf844edca, 
               32'shf8435e9d, 32'shf841cf71, 32'shf8404046, 32'shf83eb11c, 32'shf83d21f3, 32'shf83b92cc, 32'shf83a03a6, 32'shf8387481, 
               32'shf836e55d, 32'shf835563b, 32'shf833c719, 32'shf83237f9, 32'shf830a8da, 32'shf82f19bc, 32'shf82d8aa0, 32'shf82bfb84, 
               32'shf82a6c6a, 32'shf828dd51, 32'shf8274e3a, 32'shf825bf23, 32'shf824300e, 32'shf822a0fa, 32'shf82111e7, 32'shf81f82d5, 
               32'shf81df3c5, 32'shf81c64b6, 32'shf81ad5a8, 32'shf819469b, 32'shf817b78f, 32'shf8162885, 32'shf814997c, 32'shf8130a74, 
               32'shf8117b6d, 32'shf80fec68, 32'shf80e5d64, 32'shf80cce61, 32'shf80b3f5f, 32'shf809b05e, 32'shf808215f, 32'shf8069261, 
               32'shf8050364, 32'shf8037468, 32'shf801e56e, 32'shf8005675, 32'shf7fec77d, 32'shf7fd3886, 32'shf7fba991, 32'shf7fa1a9c, 
               32'shf7f88ba9, 32'shf7f6fcb8, 32'shf7f56dc7, 32'shf7f3ded8, 32'shf7f24fea, 32'shf7f0c0fd, 32'shf7ef3211, 32'shf7eda327, 
               32'shf7ec143e, 32'shf7ea8556, 32'shf7e8f670, 32'shf7e7678a, 32'shf7e5d8a6, 32'shf7e449c3, 32'shf7e2bae2, 32'shf7e12c01, 
               32'shf7df9d22, 32'shf7de0e44, 32'shf7dc7f68, 32'shf7daf08d, 32'shf7d961b3, 32'shf7d7d2da, 32'shf7d64402, 32'shf7d4b52c, 
               32'shf7d32657, 32'shf7d19783, 32'shf7d008b1, 32'shf7ce79df, 32'shf7cceb0f, 32'shf7cb5c41, 32'shf7c9cd73, 32'shf7c83ea7, 
               32'shf7c6afdc, 32'shf7c52112, 32'shf7c3924a, 32'shf7c20383, 32'shf7c074bd, 32'shf7bee5f9, 32'shf7bd5735, 32'shf7bbc873, 
               32'shf7ba39b3, 32'shf7b8aaf3, 32'shf7b71c35, 32'shf7b58d78, 32'shf7b3febc, 32'shf7b27002, 32'shf7b0e149, 32'shf7af5291, 
               32'shf7adc3db, 32'shf7ac3525, 32'shf7aaa671, 32'shf7a917bf, 32'shf7a7890d, 32'shf7a5fa5d, 32'shf7a46baf, 32'shf7a2dd01, 
               32'shf7a14e55, 32'shf79fbfaa, 32'shf79e3100, 32'shf79ca258, 32'shf79b13b1, 32'shf799850b, 32'shf797f667, 32'shf79667c4, 
               32'shf794d922, 32'shf7934a81, 32'shf791bbe2, 32'shf7902d44, 32'shf78e9ea7, 32'shf78d100c, 32'shf78b8172, 32'shf789f2d9, 
               32'shf7886442, 32'shf786d5ab, 32'shf7854717, 32'shf783b883, 32'shf78229f1, 32'shf7809b60, 32'shf77f0cd0, 32'shf77d7e42, 
               32'shf77befb5, 32'shf77a6129, 32'shf778d29f, 32'shf7774416, 32'shf775b58e, 32'shf7742708, 32'shf7729883, 32'shf77109ff, 
               32'shf76f7b7d, 32'shf76decfb, 32'shf76c5e7c, 32'shf76acffd, 32'shf7694180, 32'shf767b304, 32'shf766248a, 32'shf7649610, 
               32'shf7630799, 32'shf7617922, 32'shf75feaad, 32'shf75e5c39, 32'shf75ccdc6, 32'shf75b3f55, 32'shf759b0e5, 32'shf7582277, 
               32'shf756940a, 32'shf755059e, 32'shf7537733, 32'shf751e8ca, 32'shf7505a62, 32'shf74ecbfc, 32'shf74d3d96, 32'shf74baf33, 
               32'shf74a20d0, 32'shf748926f, 32'shf747040f, 32'shf74575b1, 32'shf743e754, 32'shf74258f8, 32'shf740ca9d, 32'shf73f3c44, 
               32'shf73daded, 32'shf73c1f96, 32'shf73a9141, 32'shf73902ee, 32'shf737749b, 32'shf735e64a, 32'shf73457fb, 32'shf732c9ad, 
               32'shf7313b60, 32'shf72fad14, 32'shf72e1eca, 32'shf72c9081, 32'shf72b023a, 32'shf72973f4, 32'shf727e5af, 32'shf726576c, 
               32'shf724c92a, 32'shf7233ae9, 32'shf721acaa, 32'shf7201e6c, 32'shf71e902f, 32'shf71d01f4, 32'shf71b73ba, 32'shf719e582, 
               32'shf718574b, 32'shf716c915, 32'shf7153ae1, 32'shf713acae, 32'shf7121e7c, 32'shf710904c, 32'shf70f021d, 32'shf70d73f0, 
               32'shf70be5c4, 32'shf70a5799, 32'shf708c970, 32'shf7073b48, 32'shf705ad22, 32'shf7041efd, 32'shf70290d9, 32'shf70102b6, 
               32'shf6ff7496, 32'shf6fde676, 32'shf6fc5858, 32'shf6faca3b, 32'shf6f93c20, 32'shf6f7ae06, 32'shf6f61fed, 32'shf6f491d6, 
               32'shf6f303c0, 32'shf6f175ac, 32'shf6efe798, 32'shf6ee5987, 32'shf6eccb77, 32'shf6eb3d68, 32'shf6e9af5a, 32'shf6e8214e, 
               32'shf6e69344, 32'shf6e5053a, 32'shf6e37733, 32'shf6e1e92c, 32'shf6e05b27, 32'shf6decd24, 32'shf6dd3f21, 32'shf6dbb121, 
               32'shf6da2321, 32'shf6d89523, 32'shf6d70727, 32'shf6d5792c, 32'shf6d3eb32, 32'shf6d25d39, 32'shf6d0cf43, 32'shf6cf414d, 
               32'shf6cdb359, 32'shf6cc2566, 32'shf6ca9775, 32'shf6c90985, 32'shf6c77b97, 32'shf6c5edaa, 32'shf6c45fbe, 32'shf6c2d1d4, 
               32'shf6c143ec, 32'shf6bfb604, 32'shf6be281e, 32'shf6bc9a3a, 32'shf6bb0c57, 32'shf6b97e76, 32'shf6b7f095, 32'shf6b662b7, 
               32'shf6b4d4d9, 32'shf6b346fe, 32'shf6b1b923, 32'shf6b02b4a, 32'shf6ae9d73, 32'shf6ad0f9d, 32'shf6ab81c8, 32'shf6a9f3f5, 
               32'shf6a86623, 32'shf6a6d853, 32'shf6a54a84, 32'shf6a3bcb6, 32'shf6a22eea, 32'shf6a0a120, 32'shf69f1357, 32'shf69d858f, 
               32'shf69bf7c9, 32'shf69a6a04, 32'shf698dc41, 32'shf6974e7f, 32'shf695c0be, 32'shf69432ff, 32'shf692a542, 32'shf6911786, 
               32'shf68f89cb, 32'shf68dfc12, 32'shf68c6e5a, 32'shf68ae0a4, 32'shf68952ef, 32'shf687c53c, 32'shf686378a, 32'shf684a9da, 
               32'shf6831c2b, 32'shf6818e7d, 32'shf68000d1, 32'shf67e7327, 32'shf67ce57e, 32'shf67b57d6, 32'shf679ca30, 32'shf6783c8b, 
               32'shf676aee8, 32'shf6752146, 32'shf67393a6, 32'shf6720607, 32'shf670786a, 32'shf66eeace, 32'shf66d5d34, 32'shf66bcf9b, 
               32'shf66a4203, 32'shf668b46d, 32'shf66726d9, 32'shf6659946, 32'shf6640bb4, 32'shf6627e24, 32'shf660f096, 32'shf65f6309, 
               32'shf65dd57d, 32'shf65c47f3, 32'shf65aba6b, 32'shf6592ce4, 32'shf6579f5e, 32'shf65611da, 32'shf6548457, 32'shf652f6d6, 
               32'shf6516956, 32'shf64fdbd8, 32'shf64e4e5c, 32'shf64cc0e0, 32'shf64b3367, 32'shf649a5ef, 32'shf6481878, 32'shf6468b03, 
               32'shf644fd8f, 32'shf643701d, 32'shf641e2ac, 32'shf640553d, 32'shf63ec7cf, 32'shf63d3a63, 32'shf63bacf8, 32'shf63a1f8f, 
               32'shf6389228, 32'shf63704c1, 32'shf635775d, 32'shf633e9fa, 32'shf6325c98, 32'shf630cf38, 32'shf62f41d9, 32'shf62db47c, 
               32'shf62c2721, 32'shf62a99c7, 32'shf6290c6e, 32'shf6277f17, 32'shf625f1c2, 32'shf624646e, 32'shf622d71b, 32'shf62149ca, 
               32'shf61fbc7b, 32'shf61e2f2d, 32'shf61ca1e1, 32'shf61b1496, 32'shf619874c, 32'shf617fa05, 32'shf6166cbe, 32'shf614df7a, 
               32'shf6135237, 32'shf611c4f5, 32'shf61037b5, 32'shf60eaa76, 32'shf60d1d39, 32'shf60b8ffd, 32'shf60a02c3, 32'shf608758b, 
               32'shf606e854, 32'shf6055b1f, 32'shf603cdeb, 32'shf60240b9, 32'shf600b388, 32'shf5ff2659, 32'shf5fd992b, 32'shf5fc0bff, 
               32'shf5fa7ed4, 32'shf5f8f1ab, 32'shf5f76484, 32'shf5f5d75e, 32'shf5f44a39, 32'shf5f2bd16, 32'shf5f12ff5, 32'shf5efa2d5, 
               32'shf5ee15b7, 32'shf5ec889a, 32'shf5eafb7f, 32'shf5e96e66, 32'shf5e7e14e, 32'shf5e65437, 32'shf5e4c722, 32'shf5e33a0f, 
               32'shf5e1acfd, 32'shf5e01fed, 32'shf5de92de, 32'shf5dd05d1, 32'shf5db78c6, 32'shf5d9ebbc, 32'shf5d85eb3, 32'shf5d6d1ad, 
               32'shf5d544a7, 32'shf5d3b7a4, 32'shf5d22aa2, 32'shf5d09da1, 32'shf5cf10a2, 32'shf5cd83a5, 32'shf5cbf6a9, 32'shf5ca69af, 
               32'shf5c8dcb6, 32'shf5c74fbf, 32'shf5c5c2c9, 32'shf5c435d5, 32'shf5c2a8e3, 32'shf5c11bf2, 32'shf5bf8f03, 32'shf5be0215, 
               32'shf5bc7529, 32'shf5bae83f, 32'shf5b95b56, 32'shf5b7ce6f, 32'shf5b64189, 32'shf5b4b4a5, 32'shf5b327c2, 32'shf5b19ae1, 
               32'shf5b00e02, 32'shf5ae8124, 32'shf5acf448, 32'shf5ab676d, 32'shf5a9da94, 32'shf5a84dbd, 32'shf5a6c0e7, 32'shf5a53413, 
               32'shf5a3a740, 32'shf5a21a6f, 32'shf5a08da0, 32'shf59f00d2, 32'shf59d7406, 32'shf59be73b, 32'shf59a5a72, 32'shf598cdab, 
               32'shf59740e5, 32'shf595b421, 32'shf594275e, 32'shf5929a9d, 32'shf5910dde, 32'shf58f8120, 32'shf58df464, 32'shf58c67a9, 
               32'shf58adaf0, 32'shf5894e39, 32'shf587c183, 32'shf58634cf, 32'shf584a81d, 32'shf5831b6c, 32'shf5818ebd, 32'shf580020f, 
               32'shf57e7563, 32'shf57ce8b9, 32'shf57b5c10, 32'shf579cf69, 32'shf57842c3, 32'shf576b61f, 32'shf575297d, 32'shf5739cdc, 
               32'shf572103d, 32'shf57083a0, 32'shf56ef704, 32'shf56d6a6a, 32'shf56bddd1, 32'shf56a513b, 32'shf568c4a5, 32'shf5673812, 
               32'shf565ab80, 32'shf5641eef, 32'shf5629261, 32'shf56105d4, 32'shf55f7948, 32'shf55decbe, 32'shf55c6036, 32'shf55ad3b0, 
               32'shf559472b, 32'shf557baa8, 32'shf5562e26, 32'shf554a1a6, 32'shf5531528, 32'shf55188ab, 32'shf54ffc30, 32'shf54e6fb7, 
               32'shf54ce33f, 32'shf54b56c9, 32'shf549ca55, 32'shf5483de2, 32'shf546b171, 32'shf5452501, 32'shf5439893, 32'shf5420c27, 
               32'shf5407fbd, 32'shf53ef354, 32'shf53d66ed, 32'shf53bda87, 32'shf53a4e24, 32'shf538c1c1, 32'shf5373561, 32'shf535a902, 
               32'shf5341ca5, 32'shf5329049, 32'shf53103ef, 32'shf52f7797, 32'shf52deb41, 32'shf52c5eec, 32'shf52ad299, 32'shf5294647, 
               32'shf527b9f7, 32'shf5262da9, 32'shf524a15d, 32'shf5231512, 32'shf52188c9, 32'shf51ffc81, 32'shf51e703b, 32'shf51ce3f7, 
               32'shf51b57b5, 32'shf519cb74, 32'shf5183f35, 32'shf516b2f7, 32'shf51526bc, 32'shf5139a82, 32'shf5120e49, 32'shf5108213, 
               32'shf50ef5de, 32'shf50d69aa, 32'shf50bdd79, 32'shf50a5149, 32'shf508c51b, 32'shf50738ee, 32'shf505acc3, 32'shf504209a, 
               32'shf5029473, 32'shf501084d, 32'shf4ff7c29, 32'shf4fdf007, 32'shf4fc63e6, 32'shf4fad7c7, 32'shf4f94baa, 32'shf4f7bf8e, 
               32'shf4f63374, 32'shf4f4a75c, 32'shf4f31b46, 32'shf4f18f31, 32'shf4f0031e, 32'shf4ee770c, 32'shf4eceafd, 32'shf4eb5eef, 
               32'shf4e9d2e3, 32'shf4e846d8, 32'shf4e6bacf, 32'shf4e52ec8, 32'shf4e3a2c3, 32'shf4e216bf, 32'shf4e08abd, 32'shf4defebd, 
               32'shf4dd72be, 32'shf4dbe6c2, 32'shf4da5ac7, 32'shf4d8cecd, 32'shf4d742d6, 32'shf4d5b6e0, 32'shf4d42aeb, 32'shf4d29ef9, 
               32'shf4d11308, 32'shf4cf8719, 32'shf4cdfb2c, 32'shf4cc6f40, 32'shf4cae356, 32'shf4c9576e, 32'shf4c7cb88, 32'shf4c63fa3, 
               32'shf4c4b3c0, 32'shf4c327df, 32'shf4c19c00, 32'shf4c01022, 32'shf4be8446, 32'shf4bcf86c, 32'shf4bb6c93, 32'shf4b9e0bc, 
               32'shf4b854e7, 32'shf4b6c914, 32'shf4b53d42, 32'shf4b3b173, 32'shf4b225a4, 32'shf4b099d8, 32'shf4af0e0d, 32'shf4ad8245, 
               32'shf4abf67e, 32'shf4aa6ab8, 32'shf4a8def5, 32'shf4a75333, 32'shf4a5c773, 32'shf4a43bb4, 32'shf4a2aff8, 32'shf4a1243d, 
               32'shf49f9884, 32'shf49e0ccc, 32'shf49c8117, 32'shf49af563, 32'shf49969b1, 32'shf497de00, 32'shf4965252, 32'shf494c6a5, 
               32'shf4933afa, 32'shf491af51, 32'shf49023a9, 32'shf48e9803, 32'shf48d0c5f, 32'shf48b80bd, 32'shf489f51d, 32'shf488697e, 
               32'shf486dde1, 32'shf4855246, 32'shf483c6ad, 32'shf4823b15, 32'shf480af7f, 32'shf47f23eb, 32'shf47d9859, 32'shf47c0cc8, 
               32'shf47a8139, 32'shf478f5ad, 32'shf4776a21, 32'shf475de98, 32'shf4745310, 32'shf472c78a, 32'shf4713c06, 32'shf46fb084, 
               32'shf46e2504, 32'shf46c9985, 32'shf46b0e08, 32'shf469828d, 32'shf467f713, 32'shf4666b9c, 32'shf464e026, 32'shf46354b2, 
               32'shf461c940, 32'shf4603dcf, 32'shf45eb261, 32'shf45d26f4, 32'shf45b9b89, 32'shf45a1020, 32'shf45884b8, 32'shf456f953, 
               32'shf4556def, 32'shf453e28d, 32'shf452572c, 32'shf450cbce, 32'shf44f4071, 32'shf44db517, 32'shf44c29be, 32'shf44a9e66, 
               32'shf4491311, 32'shf44787bd, 32'shf445fc6b, 32'shf444711b, 32'shf442e5cd, 32'shf4415a81, 32'shf43fcf36, 32'shf43e43ed, 
               32'shf43cb8a7, 32'shf43b2d61, 32'shf439a21e, 32'shf43816dd, 32'shf4368b9d, 32'shf435005f, 32'shf4337523, 32'shf431e9e9, 
               32'shf4305eb0, 32'shf42ed37a, 32'shf42d4845, 32'shf42bbd12, 32'shf42a31e1, 32'shf428a6b2, 32'shf4271b84, 32'shf4259058, 
               32'shf424052f, 32'shf4227a07, 32'shf420eee1, 32'shf41f63bc, 32'shf41dd89a, 32'shf41c4d79, 32'shf41ac25a, 32'shf419373d, 
               32'shf417ac22, 32'shf4162109, 32'shf41495f1, 32'shf4130adc, 32'shf4117fc8, 32'shf40ff4b6, 32'shf40e69a6, 32'shf40cde97, 
               32'shf40b538b, 32'shf409c880, 32'shf4083d78, 32'shf406b271, 32'shf405276c, 32'shf4039c68, 32'shf4021167, 32'shf4008668, 
               32'shf3fefb6a, 32'shf3fd706e, 32'shf3fbe574, 32'shf3fa5a7c, 32'shf3f8cf86, 32'shf3f74491, 32'shf3f5b99f, 32'shf3f42eae, 
               32'shf3f2a3bf, 32'shf3f118d2, 32'shf3ef8de7, 32'shf3ee02fe, 32'shf3ec7817, 32'shf3eaed31, 32'shf3e9624d, 32'shf3e7d76c, 
               32'shf3e64c8c, 32'shf3e4c1ae, 32'shf3e336d1, 32'shf3e1abf7, 32'shf3e0211f, 32'shf3de9648, 32'shf3dd0b73, 32'shf3db80a0, 
               32'shf3d9f5cf, 32'shf3d86b00, 32'shf3d6e033, 32'shf3d55568, 32'shf3d3ca9e, 32'shf3d23fd7, 32'shf3d0b511, 32'shf3cf2a4d, 
               32'shf3cd9f8b, 32'shf3cc14cb, 32'shf3ca8a0d, 32'shf3c8ff51, 32'shf3c77496, 32'shf3c5e9de, 32'shf3c45f27, 32'shf3c2d472, 
               32'shf3c149bf, 32'shf3bfbf0e, 32'shf3be345f, 32'shf3bca9b2, 32'shf3bb1f07, 32'shf3b9945d, 32'shf3b809b6, 32'shf3b67f10, 
               32'shf3b4f46c, 32'shf3b369ca, 32'shf3b1df2a, 32'shf3b0548c, 32'shf3aec9f0, 32'shf3ad3f56, 32'shf3abb4bd, 32'shf3aa2a27, 
               32'shf3a89f92, 32'shf3a71500, 32'shf3a58a6f, 32'shf3a3ffe0, 32'shf3a27553, 32'shf3a0eac8, 32'shf39f603f, 32'shf39dd5b8, 
               32'shf39c4b32, 32'shf39ac0af, 32'shf399362d, 32'shf397abae, 32'shf3962130, 32'shf39496b4, 32'shf3930c3b, 32'shf39181c3, 
               32'shf38ff74d, 32'shf38e6cd9, 32'shf38ce266, 32'shf38b57f6, 32'shf389cd88, 32'shf388431b, 32'shf386b8b1, 32'shf3852e48, 
               32'shf383a3e2, 32'shf382197d, 32'shf3808f1a, 32'shf37f04b9, 32'shf37d7a5b, 32'shf37beffe, 32'shf37a65a2, 32'shf378db49, 
               32'shf37750f2, 32'shf375c69d, 32'shf3743c49, 32'shf372b1f8, 32'shf37127a9, 32'shf36f9d5b, 32'shf36e130f, 32'shf36c88c6, 
               32'shf36afe7e, 32'shf3697438, 32'shf367e9f4, 32'shf3665fb3, 32'shf364d573, 32'shf3634b35, 32'shf361c0f9, 32'shf36036be, 
               32'shf35eac86, 32'shf35d2250, 32'shf35b981c, 32'shf35a0de9, 32'shf35883b9, 32'shf356f98b, 32'shf3556f5e, 32'shf353e534, 
               32'shf3525b0b, 32'shf350d0e5, 32'shf34f46c0, 32'shf34dbc9d, 32'shf34c327c, 32'shf34aa85e, 32'shf3491e41, 32'shf3479426, 
               32'shf3460a0d, 32'shf3447ff6, 32'shf342f5e1, 32'shf3416bce, 32'shf33fe1bd, 32'shf33e57ae, 32'shf33ccda1, 32'shf33b4396, 
               32'shf339b98d, 32'shf3382f86, 32'shf336a580, 32'shf3351b7d, 32'shf333917c, 32'shf332077c, 32'shf3307d7f, 32'shf32ef384, 
               32'shf32d698a, 32'shf32bdf93, 32'shf32a559e, 32'shf328cbaa, 32'shf32741b9, 32'shf325b7c9, 32'shf3242ddc, 32'shf322a3f0, 
               32'shf3211a07, 32'shf31f901f, 32'shf31e0639, 32'shf31c7c56, 32'shf31af274, 32'shf3196895, 32'shf317deb7, 32'shf31654db, 
               32'shf314cb02, 32'shf313412a, 32'shf311b755, 32'shf3102d81, 32'shf30ea3af, 32'shf30d19e0, 32'shf30b9012, 32'shf30a0646, 
               32'shf3087c7d, 32'shf306f2b5, 32'shf30568ef, 32'shf303df2c, 32'shf302556a, 32'shf300cbaa, 32'shf2ff41ed, 32'shf2fdb831, 
               32'shf2fc2e77, 32'shf2faa4c0, 32'shf2f91b0a, 32'shf2f79156, 32'shf2f607a5, 32'shf2f47df5, 32'shf2f2f448, 32'shf2f16a9c, 
               32'shf2efe0f2, 32'shf2ee574b, 32'shf2eccda5, 32'shf2eb4402, 32'shf2e9ba60, 32'shf2e830c1, 32'shf2e6a723, 32'shf2e51d88, 
               32'shf2e393ef, 32'shf2e20a57, 32'shf2e080c2, 32'shf2def72e, 32'shf2dd6d9d, 32'shf2dbe40e, 32'shf2da5a81, 32'shf2d8d0f5, 
               32'shf2d7476c, 32'shf2d5bde5, 32'shf2d43460, 32'shf2d2aadd, 32'shf2d1215b, 32'shf2cf97dc, 32'shf2ce0e5f, 32'shf2cc84e4, 
               32'shf2cafb6b, 32'shf2c971f5, 32'shf2c7e880, 32'shf2c65f0d, 32'shf2c4d59c, 32'shf2c34c2d, 32'shf2c1c2c0, 32'shf2c03956, 
               32'shf2beafed, 32'shf2bd2687, 32'shf2bb9d22, 32'shf2ba13c0, 32'shf2b88a5f, 32'shf2b70101, 32'shf2b577a4, 32'shf2b3ee4a, 
               32'shf2b264f2, 32'shf2b0db9b, 32'shf2af5247, 32'shf2adc8f5, 32'shf2ac3fa5, 32'shf2aab657, 32'shf2a92d0b, 32'shf2a7a3c1, 
               32'shf2a61a7a, 32'shf2a49134, 32'shf2a307f0, 32'shf2a17eae, 32'shf29ff56f, 32'shf29e6c31, 32'shf29ce2f6, 32'shf29b59bc, 
               32'shf299d085, 32'shf2984750, 32'shf296be1d, 32'shf29534ec, 32'shf293abbd, 32'shf2922290, 32'shf2909965, 32'shf28f103c, 
               32'shf28d8715, 32'shf28bfdf0, 32'shf28a74ce, 32'shf288ebad, 32'shf287628f, 32'shf285d972, 32'shf2845058, 32'shf282c740, 
               32'shf2813e2a, 32'shf27fb516, 32'shf27e2c04, 32'shf27ca2f4, 32'shf27b19e6, 32'shf27990da, 32'shf27807d0, 32'shf2767ec9, 
               32'shf274f5c3, 32'shf2736cc0, 32'shf271e3bf, 32'shf2705abf, 32'shf26ed1c2, 32'shf26d48c7, 32'shf26bbfce, 32'shf26a36d8, 
               32'shf268ade3, 32'shf26724f0, 32'shf2659c00, 32'shf2641311, 32'shf2628a25, 32'shf261013b, 32'shf25f7852, 32'shf25def6c, 
               32'shf25c6688, 32'shf25adda7, 32'shf25954c7, 32'shf257cbe9, 32'shf256430e, 32'shf254ba34, 32'shf253315d, 32'shf251a888, 
               32'shf2501fb5, 32'shf24e96e4, 32'shf24d0e15, 32'shf24b8548, 32'shf249fc7d, 32'shf24873b5, 32'shf246eaee, 32'shf245622a, 
               32'shf243d968, 32'shf24250a8, 32'shf240c7ea, 32'shf23f3f2e, 32'shf23db674, 32'shf23c2dbd, 32'shf23aa507, 32'shf2391c54, 
               32'shf23793a3, 32'shf2360af4, 32'shf2348247, 32'shf232f99c, 32'shf23170f3, 32'shf22fe84c, 32'shf22e5fa8, 32'shf22cd706, 
               32'shf22b4e66, 32'shf229c5c7, 32'shf2283d2c, 32'shf226b492, 32'shf2252bfa, 32'shf223a365, 32'shf2221ad1, 32'shf2209240, 
               32'shf21f09b1, 32'shf21d8124, 32'shf21bf899, 32'shf21a7010, 32'shf218e78a, 32'shf2175f06, 32'shf215d683, 32'shf2144e03, 
               32'shf212c585, 32'shf2113d09, 32'shf20fb490, 32'shf20e2c18, 32'shf20ca3a3, 32'shf20b1b30, 32'shf20992bf, 32'shf2080a50, 
               32'shf20681e3, 32'shf204f978, 32'shf2037110, 32'shf201e8aa, 32'shf2006046, 32'shf1fed7e4, 32'shf1fd4f84, 32'shf1fbc726, 
               32'shf1fa3ecb, 32'shf1f8b671, 32'shf1f72e1a, 32'shf1f5a5c5, 32'shf1f41d72, 32'shf1f29522, 32'shf1f10cd3, 32'shf1ef8487, 
               32'shf1edfc3d, 32'shf1ec73f5, 32'shf1eaebaf, 32'shf1e9636b, 32'shf1e7db2a, 32'shf1e652eb, 32'shf1e4caae, 32'shf1e34273, 
               32'shf1e1ba3a, 32'shf1e03203, 32'shf1dea9cf, 32'shf1dd219d, 32'shf1db996d, 32'shf1da113f, 32'shf1d88913, 32'shf1d700ea, 
               32'shf1d578c2, 32'shf1d3f09d, 32'shf1d2687a, 32'shf1d0e059, 32'shf1cf583b, 32'shf1cdd01e, 32'shf1cc4804, 32'shf1cabfec, 
               32'shf1c937d6, 32'shf1c7afc3, 32'shf1c627b1, 32'shf1c49fa2, 32'shf1c31795, 32'shf1c18f8a, 32'shf1c00781, 32'shf1be7f7b, 
               32'shf1bcf777, 32'shf1bb6f75, 32'shf1b9e775, 32'shf1b85f77, 32'shf1b6d77c, 32'shf1b54f82, 32'shf1b3c78b, 32'shf1b23f97, 
               32'shf1b0b7a4, 32'shf1af2fb3, 32'shf1ada7c5, 32'shf1ac1fd9, 32'shf1aa97ef, 32'shf1a91008, 32'shf1a78822, 32'shf1a6003f, 
               32'shf1a4785e, 32'shf1a2f080, 32'shf1a168a3, 32'shf19fe0c9, 32'shf19e58f1, 32'shf19cd11b, 32'shf19b4947, 32'shf199c176, 
               32'shf19839a6, 32'shf196b1d9, 32'shf1952a0f, 32'shf193a246, 32'shf1921a80, 32'shf19092bc, 32'shf18f0afa, 32'shf18d833a, 
               32'shf18bfb7d, 32'shf18a73c2, 32'shf188ec09, 32'shf1876452, 32'shf185dc9d, 32'shf18454eb, 32'shf182cd3b, 32'shf181458d, 
               32'shf17fbde2, 32'shf17e3638, 32'shf17cae91, 32'shf17b26ec, 32'shf1799f4a, 32'shf17817a9, 32'shf176900b, 32'shf175086f, 
               32'shf17380d6, 32'shf171f93e, 32'shf17071a9, 32'shf16eea16, 32'shf16d6286, 32'shf16bdaf7, 32'shf16a536b, 32'shf168cbe1, 
               32'shf1674459, 32'shf165bcd4, 32'shf1643551, 32'shf162add0, 32'shf1612651, 32'shf15f9ed5, 32'shf15e175b, 32'shf15c8fe3, 
               32'shf15b086d, 32'shf15980fa, 32'shf157f989, 32'shf156721a, 32'shf154eaad, 32'shf1536343, 32'shf151dbdb, 32'shf1505475, 
               32'shf14ecd11, 32'shf14d45b0, 32'shf14bbe51, 32'shf14a36f4, 32'shf148af9a, 32'shf1472842, 32'shf145a0ec, 32'shf1441998, 
               32'shf1429247, 32'shf1410af8, 32'shf13f83ab, 32'shf13dfc60, 32'shf13c7518, 32'shf13aedd2, 32'shf139668e, 32'shf137df4d, 
               32'shf136580d, 32'shf134d0d0, 32'shf1334996, 32'shf131c25d, 32'shf1303b27, 32'shf12eb3f4, 32'shf12d2cc2, 32'shf12ba593, 
               32'shf12a1e66, 32'shf128973b, 32'shf1271013, 32'shf12588ed, 32'shf12401c9, 32'shf1227aa8, 32'shf120f389, 32'shf11f6c6c, 
               32'shf11de551, 32'shf11c5e39, 32'shf11ad723, 32'shf119500f, 32'shf117c8fe, 32'shf11641ef, 32'shf114bae2, 32'shf11333d7, 
               32'shf111accf, 32'shf11025c9, 32'shf10e9ec6, 32'shf10d17c4, 32'shf10b90c5, 32'shf10a09c9, 32'shf10882ce, 32'shf106fbd6, 
               32'shf10574e0, 32'shf103eded, 32'shf10266fc, 32'shf100e00d, 32'shf0ff5921, 32'shf0fdd236, 32'shf0fc4b4f, 32'shf0fac469, 
               32'shf0f93d86, 32'shf0f7b6a5, 32'shf0f62fc6, 32'shf0f4a8ea, 32'shf0f32210, 32'shf0f19b38, 32'shf0f01463, 32'shf0ee8d90, 
               32'shf0ed06bf, 32'shf0eb7ff1, 32'shf0e9f925, 32'shf0e8725b, 32'shf0e6eb94, 32'shf0e564cf, 32'shf0e3de0c, 32'shf0e2574c, 
               32'shf0e0d08d, 32'shf0df49d2, 32'shf0ddc318, 32'shf0dc3c61, 32'shf0dab5ad, 32'shf0d92efa, 32'shf0d7a84a, 32'shf0d6219c, 
               32'shf0d49af1, 32'shf0d31448, 32'shf0d18da1, 32'shf0d006fd, 32'shf0ce805b, 32'shf0ccf9bb, 32'shf0cb731e, 32'shf0c9ec83, 
               32'shf0c865ea, 32'shf0c6df54, 32'shf0c558c0, 32'shf0c3d22e, 32'shf0c24b9f, 32'shf0c0c512, 32'shf0bf3e88, 32'shf0bdb7ff, 
               32'shf0bc317a, 32'shf0baaaf6, 32'shf0b92475, 32'shf0b79df6, 32'shf0b6177a, 32'shf0b49100, 32'shf0b30a88, 32'shf0b18413, 
               32'shf0affda0, 32'shf0ae772f, 32'shf0acf0c1, 32'shf0ab6a55, 32'shf0a9e3eb, 32'shf0a85d84, 32'shf0a6d71f, 32'shf0a550bd, 
               32'shf0a3ca5d, 32'shf0a243ff, 32'shf0a0bda4, 32'shf09f374b, 32'shf09db0f4, 32'shf09c2aa0, 32'shf09aa44e, 32'shf0991dff, 
               32'shf09797b2, 32'shf0961167, 32'shf0948b1f, 32'shf09304d9, 32'shf0917e95, 32'shf08ff854, 32'shf08e7215, 32'shf08cebd9, 
               32'shf08b659f, 32'shf089df67, 32'shf0885932, 32'shf086d2ff, 32'shf0854cce, 32'shf083c6a0, 32'shf0824074, 32'shf080ba4b, 
               32'shf07f3424, 32'shf07dadff, 32'shf07c27dd, 32'shf07aa1bd, 32'shf0791ba0, 32'shf0779585, 32'shf0760f6c, 32'shf0748956, 
               32'shf0730342, 32'shf0717d31, 32'shf06ff722, 32'shf06e7115, 32'shf06ceb0b, 32'shf06b6503, 32'shf069defe, 32'shf06858fb, 
               32'shf066d2fa, 32'shf0654cfc, 32'shf063c700, 32'shf0624107, 32'shf060bb10, 32'shf05f351b, 32'shf05daf29, 32'shf05c293a, 
               32'shf05aa34c, 32'shf0591d61, 32'shf0579779, 32'shf0561193, 32'shf0548baf, 32'shf05305ce, 32'shf0517fef, 32'shf04ffa12, 
               32'shf04e7438, 32'shf04cee61, 32'shf04b688c, 32'shf049e2b9, 32'shf0485ce9, 32'shf046d71b, 32'shf045514f, 32'shf043cb86, 
               32'shf04245c0, 32'shf040bffb, 32'shf03f3a3a, 32'shf03db47a, 32'shf03c2ebd, 32'shf03aa903, 32'shf039234b, 32'shf0379d95, 
               32'shf03617e2, 32'shf0349231, 32'shf0330c83, 32'shf03186d7, 32'shf030012e, 32'shf02e7b87, 32'shf02cf5e2, 32'shf02b7040, 
               32'shf029eaa1, 32'shf0286503, 32'shf026df68, 32'shf02559d0, 32'shf023d43a, 32'shf0224ea7, 32'shf020c916, 32'shf01f4387, 
               32'shf01dbdfb, 32'shf01c3871, 32'shf01ab2ea, 32'shf0192d66, 32'shf017a7e3, 32'shf0162263, 32'shf0149ce6, 32'shf013176b, 
               32'shf01191f3, 32'shf0100c7d, 32'shf00e8709, 32'shf00d0198, 32'shf00b7c29, 32'shf009f6bd, 32'shf0087153, 32'shf006ebec, 
               32'shf0056687, 32'shf003e125, 32'shf0025bc5, 32'shf000d668, 32'shefff510d, 32'sheffdcbb4, 32'sheffc465e, 32'sheffac10b, 
               32'sheff93bba, 32'sheff7b66b, 32'sheff6311f, 32'sheff4abd5, 32'sheff3268e, 32'sheff1a149, 32'sheff01c07, 32'shefee96c7, 
               32'shefed118a, 32'shefeb8c4f, 32'shefea0717, 32'shefe881e1, 32'shefe6fcae, 32'shefe5777d, 32'shefe3f24f, 32'shefe26d23, 
               32'shefe0e7f9, 32'shefdf62d2, 32'shefddddae, 32'shefdc588c, 32'shefdad36c, 32'shefd94e50, 32'shefd7c935, 32'shefd6441d, 
               32'shefd4bf08, 32'shefd339f5, 32'shefd1b4e4, 32'shefd02fd6, 32'shefceaacb, 32'shefcd25c1, 32'shefcba0bb, 32'shefca1bb7, 
               32'shefc896b5, 32'shefc711b6, 32'shefc58cba, 32'shefc407c0, 32'shefc282c8, 32'shefc0fdd3, 32'shefbf78e1, 32'shefbdf3f1, 
               32'shefbc6f03, 32'shefbaea18, 32'shefb96530, 32'shefb7e04a, 32'shefb65b66, 32'shefb4d686, 32'shefb351a7, 32'shefb1cccb, 
               32'shefb047f2, 32'shefaec31b, 32'shefad3e47, 32'shefabb975, 32'shefaa34a5, 32'shefa8afd9, 32'shefa72b0e, 32'shefa5a646, 
               32'shefa42181, 32'shefa29cbe, 32'shefa117fe, 32'shef9f9341, 32'shef9e0e85, 32'shef9c89cd, 32'shef9b0517, 32'shef998063, 
               32'shef97fbb2, 32'shef967704, 32'shef94f258, 32'shef936dae, 32'shef91e907, 32'shef906463, 32'shef8edfc1, 32'shef8d5b22, 
               32'shef8bd685, 32'shef8a51eb, 32'shef88cd53, 32'shef8748be, 32'shef85c42b, 32'shef843f9b, 32'shef82bb0e, 32'shef813683, 
               32'shef7fb1fa, 32'shef7e2d74, 32'shef7ca8f1, 32'shef7b2470, 32'shef799ff2, 32'shef781b76, 32'shef7696fd, 32'shef751286, 
               32'shef738e12, 32'shef7209a1, 32'shef708532, 32'shef6f00c5, 32'shef6d7c5b, 32'shef6bf7f4, 32'shef6a738f, 32'shef68ef2d, 
               32'shef676ace, 32'shef65e670, 32'shef646216, 32'shef62ddbe, 32'shef615969, 32'shef5fd516, 32'shef5e50c6, 32'shef5ccc78, 
               32'shef5b482d, 32'shef59c3e4, 32'shef583f9e, 32'shef56bb5b, 32'shef55371a, 32'shef53b2dc, 32'shef522ea0, 32'shef50aa67, 
               32'shef4f2630, 32'shef4da1fc, 32'shef4c1dcb, 32'shef4a999c, 32'shef491570, 32'shef479146, 32'shef460d1f, 32'shef4488fa, 
               32'shef4304d8, 32'shef4180b9, 32'shef3ffc9c, 32'shef3e7882, 32'shef3cf46a, 32'shef3b7055, 32'shef39ec43, 32'shef386833, 
               32'shef36e426, 32'shef35601b, 32'shef33dc13, 32'shef32580d, 32'shef30d40a, 32'shef2f500a, 32'shef2dcc0c, 32'shef2c4811, 
               32'shef2ac419, 32'shef294023, 32'shef27bc2f, 32'shef26383f, 32'shef24b451, 32'shef233065, 32'shef21ac7c, 32'shef202896, 
               32'shef1ea4b2, 32'shef1d20d1, 32'shef1b9cf2, 32'shef1a1916, 32'shef18953d, 32'shef171166, 32'shef158d92, 32'shef1409c1, 
               32'shef1285f2, 32'shef110225, 32'shef0f7e5c, 32'shef0dfa95, 32'shef0c76d0, 32'shef0af30e, 32'shef096f4f, 32'shef07eb93, 
               32'shef0667d9, 32'shef04e421, 32'shef03606c, 32'shef01dcba, 32'shef00590b, 32'sheefed55e, 32'sheefd51b4, 32'sheefbce0c, 
               32'sheefa4a67, 32'sheef8c6c5, 32'sheef74325, 32'sheef5bf88, 32'sheef43bed, 32'sheef2b855, 32'sheef134c0, 32'sheeefb12d, 
               32'sheeee2d9d, 32'sheeecaa10, 32'sheeeb2685, 32'sheee9a2fd, 32'sheee81f78, 32'sheee69bf5, 32'sheee51875, 32'sheee394f7, 
               32'sheee2117c, 32'sheee08e04, 32'sheedf0a8e, 32'sheedd871b, 32'sheedc03ab, 32'sheeda803d, 32'sheed8fcd2, 32'sheed7796a, 
               32'sheed5f604, 32'sheed472a1, 32'sheed2ef40, 32'sheed16be3, 32'sheecfe887, 32'sheece652f, 32'sheecce1d9, 32'sheecb5e86, 
               32'sheec9db35, 32'sheec857e7, 32'sheec6d49c, 32'sheec55153, 32'sheec3ce0d, 32'sheec24aca, 32'sheec0c78a, 32'sheebf444c, 
               32'sheebdc110, 32'sheebc3dd8, 32'sheebabaa2, 32'sheeb9376e, 32'sheeb7b43e, 32'sheeb63110, 32'sheeb4ade4, 32'sheeb32abc, 
               32'sheeb1a796, 32'sheeb02472, 32'sheeaea152, 32'sheead1e34, 32'sheeab9b18, 32'sheeaa1800, 32'sheea894ea, 32'sheea711d6, 
               32'sheea58ec6, 32'sheea40bb8, 32'sheea288ad, 32'sheea105a4, 32'shee9f829e, 32'shee9dff9b, 32'shee9c7c9a, 32'shee9af99d, 
               32'shee9976a1, 32'shee97f3a9, 32'shee9670b3, 32'shee94edc0, 32'shee936acf, 32'shee91e7e2, 32'shee9064f7, 32'shee8ee20e, 
               32'shee8d5f29, 32'shee8bdc46, 32'shee8a5965, 32'shee88d688, 32'shee8753ad, 32'shee85d0d4, 32'shee844dff, 32'shee82cb2c, 
               32'shee81485c, 32'shee7fc58f, 32'shee7e42c4, 32'shee7cbffc, 32'shee7b3d36, 32'shee79ba74, 32'shee7837b4, 32'shee76b4f7, 
               32'shee75323c, 32'shee73af84, 32'shee722ccf, 32'shee70aa1d, 32'shee6f276d, 32'shee6da4c0, 32'shee6c2216, 32'shee6a9f6e, 
               32'shee691cc9, 32'shee679a27, 32'shee661788, 32'shee6494eb, 32'shee631251, 32'shee618fba, 32'shee600d25, 32'shee5e8a93, 
               32'shee5d0804, 32'shee5b8578, 32'shee5a02ee, 32'shee588067, 32'shee56fde3, 32'shee557b61, 32'shee53f8e2, 32'shee527666, 
               32'shee50f3ed, 32'shee4f7176, 32'shee4def02, 32'shee4c6c91, 32'shee4aea23, 32'shee4967b7, 32'shee47e54e, 32'shee4662e8, 
               32'shee44e084, 32'shee435e24, 32'shee41dbc6, 32'shee40596a, 32'shee3ed712, 32'shee3d54bc, 32'shee3bd269, 32'shee3a5018, 
               32'shee38cdcb, 32'shee374b80, 32'shee35c938, 32'shee3446f2, 32'shee32c4b0, 32'shee314270, 32'shee2fc033, 32'shee2e3df8, 
               32'shee2cbbc1, 32'shee2b398c, 32'shee29b75a, 32'shee28352a, 32'shee26b2fe, 32'shee2530d4, 32'shee23aead, 32'shee222c88, 
               32'shee20aa67, 32'shee1f2848, 32'shee1da62c, 32'shee1c2412, 32'shee1aa1fc, 32'shee191fe8, 32'shee179dd7, 32'shee161bc8, 
               32'shee1499bd, 32'shee1317b4, 32'shee1195ae, 32'shee1013ab, 32'shee0e91aa, 32'shee0d0fac, 32'shee0b8db1, 32'shee0a0bb9, 
               32'shee0889c4, 32'shee0707d1, 32'shee0585e1, 32'shee0403f4, 32'shee02820a, 32'shee010022, 32'shedff7e3d, 32'shedfdfc5b, 
               32'shedfc7a7c, 32'shedfaf8a0, 32'shedf976c6, 32'shedf7f4ef, 32'shedf6731b, 32'shedf4f14a, 32'shedf36f7b, 32'shedf1edaf, 
               32'shedf06be6, 32'shedeeea20, 32'sheded685d, 32'shedebe69c, 32'shedea64de, 32'shede8e323, 32'shede7616b, 32'shede5dfb5, 
               32'shede45e03, 32'shede2dc53, 32'shede15aa6, 32'sheddfd8fb, 32'shedde5754, 32'sheddcd5af, 32'sheddb540d, 32'shedd9d26e, 
               32'shedd850d2, 32'shedd6cf38, 32'shedd54da2, 32'shedd3cc0e, 32'shedd24a7d, 32'shedd0c8ee, 32'shedcf4763, 32'shedcdc5da, 
               32'shedcc4454, 32'shedcac2d1, 32'shedc94151, 32'shedc7bfd3, 32'shedc63e59, 32'shedc4bce1, 32'shedc33b6c, 32'shedc1b9fa, 
               32'shedc0388a, 32'shedbeb71e, 32'shedbd35b4, 32'shedbbb44d, 32'shedba32e9, 32'shedb8b187, 32'shedb73029, 32'shedb5aecd, 
               32'shedb42d74, 32'shedb2ac1e, 32'shedb12acb, 32'shedafa97b, 32'shedae282d, 32'shedaca6e2, 32'shedab259a, 32'sheda9a455, 
               32'sheda82313, 32'sheda6a1d4, 32'sheda52097, 32'sheda39f5d, 32'sheda21e26, 32'sheda09cf2, 32'shed9f1bc1, 32'shed9d9a92, 
               32'shed9c1967, 32'shed9a983e, 32'shed991718, 32'shed9795f5, 32'shed9614d5, 32'shed9493b7, 32'shed93129d, 32'shed919185, 
               32'shed901070, 32'shed8e8f5e, 32'shed8d0e4f, 32'shed8b8d42, 32'shed8a0c39, 32'shed888b32, 32'shed870a2e, 32'shed85892d, 
               32'shed84082f, 32'shed828734, 32'shed81063b, 32'shed7f8546, 32'shed7e0453, 32'shed7c8363, 32'shed7b0276, 32'shed79818c, 
               32'shed7800a5, 32'shed767fc0, 32'shed74fedf, 32'shed737e00, 32'shed71fd24, 32'shed707c4b, 32'shed6efb75, 32'shed6d7aa2, 
               32'shed6bf9d1, 32'shed6a7904, 32'shed68f839, 32'shed677771, 32'shed65f6ac, 32'shed6475ea, 32'shed62f52b, 32'shed61746f, 
               32'shed5ff3b5, 32'shed5e72fe, 32'shed5cf24b, 32'shed5b719a, 32'shed59f0ec, 32'shed587041, 32'shed56ef99, 32'shed556ef3, 
               32'shed53ee51, 32'shed526db1, 32'shed50ed14, 32'shed4f6c7b, 32'shed4debe4, 32'shed4c6b50, 32'shed4aeabe, 32'shed496a30, 
               32'shed47e9a5, 32'shed46691c, 32'shed44e897, 32'shed436814, 32'shed41e794, 32'shed406717, 32'shed3ee69d, 32'shed3d6626, 
               32'shed3be5b1, 32'shed3a6540, 32'shed38e4d2, 32'shed376466, 32'shed35e3fd, 32'shed346397, 32'shed32e334, 32'shed3162d4, 
               32'shed2fe277, 32'shed2e621d, 32'shed2ce1c6, 32'shed2b6171, 32'shed29e120, 32'shed2860d1, 32'shed26e086, 32'shed25603d, 
               32'shed23dff7, 32'shed225fb4, 32'shed20df74, 32'shed1f5f37, 32'shed1ddefd, 32'shed1c5ec5, 32'shed1ade91, 32'shed195e5f, 
               32'shed17de31, 32'shed165e05, 32'shed14dddc, 32'shed135db6, 32'shed11dd94, 32'shed105d74, 32'shed0edd56, 32'shed0d5d3c, 
               32'shed0bdd25, 32'shed0a5d11, 32'shed08dcff, 32'shed075cf1, 32'shed05dce5, 32'shed045cdd, 32'shed02dcd7, 32'shed015cd4, 
               32'shecffdcd4, 32'shecfe5cd8, 32'shecfcdcde, 32'shecfb5ce7, 32'shecf9dcf3, 32'shecf85d01, 32'shecf6dd13, 32'shecf55d28, 
               32'shecf3dd3f, 32'shecf25d5a, 32'shecf0dd78, 32'shecef5d98, 32'shecedddbb, 32'shecec5de2, 32'sheceade0b, 32'shece95e37, 
               32'shece7de66, 32'shece65e98, 32'shece4dece, 32'shece35f06, 32'shece1df40, 32'shece05f7e, 32'shecdedfbf, 32'shecdd6003, 
               32'shecdbe04a, 32'shecda6093, 32'shecd8e0e0, 32'shecd76130, 32'shecd5e182, 32'shecd461d8, 32'shecd2e230, 32'shecd1628c, 
               32'sheccfe2ea, 32'shecce634b, 32'sheccce3b0, 32'sheccb6417, 32'shecc9e481, 32'shecc864ee, 32'shecc6e55f, 32'shecc565d2, 
               32'shecc3e648, 32'shecc266c1, 32'shecc0e73d, 32'shecbf67bc, 32'shecbde83e, 32'shecbc68c3, 32'shecbae94b, 32'shecb969d5, 
               32'shecb7ea63, 32'shecb66af4, 32'shecb4eb88, 32'shecb36c1f, 32'shecb1ecb8, 32'shecb06d55, 32'shecaeedf5, 32'shecad6e97, 
               32'shecabef3d, 32'shecaa6fe6, 32'sheca8f091, 32'sheca77140, 32'sheca5f1f2, 32'sheca472a6, 32'sheca2f35e, 32'sheca17418, 
               32'shec9ff4d6, 32'shec9e7596, 32'shec9cf65a, 32'shec9b7720, 32'shec99f7ea, 32'shec9878b6, 32'shec96f986, 32'shec957a58, 
               32'shec93fb2e, 32'shec927c06, 32'shec90fce1, 32'shec8f7dc0, 32'shec8dfea1, 32'shec8c7f86, 32'shec8b006d, 32'shec898158, 
               32'shec880245, 32'shec868335, 32'shec850429, 32'shec83851f, 32'shec820619, 32'shec808715, 32'shec7f0815, 32'shec7d8917, 
               32'shec7c0a1d, 32'shec7a8b25, 32'shec790c31, 32'shec778d3f, 32'shec760e51, 32'shec748f65, 32'shec73107d, 32'shec719197, 
               32'shec7012b5, 32'shec6e93d6, 32'shec6d14f9, 32'shec6b9620, 32'shec6a1749, 32'shec689876, 32'shec6719a6, 32'shec659ad9, 
               32'shec641c0e, 32'shec629d47, 32'shec611e83, 32'shec5f9fc2, 32'shec5e2103, 32'shec5ca248, 32'shec5b2390, 32'shec59a4db, 
               32'shec582629, 32'shec56a77a, 32'shec5528ce, 32'shec53aa25, 32'shec522b7f, 32'shec50acdc, 32'shec4f2e3d, 32'shec4dafa0, 
               32'shec4c3106, 32'shec4ab26f, 32'shec4933dc, 32'shec47b54b, 32'shec4636bd, 32'shec44b833, 32'shec4339ab, 32'shec41bb27, 
               32'shec403ca5, 32'shec3ebe27, 32'shec3d3fac, 32'shec3bc133, 32'shec3a42be, 32'shec38c44c, 32'shec3745dd, 32'shec35c771, 
               32'shec344908, 32'shec32caa2, 32'shec314c3f, 32'shec2fcddf, 32'shec2e4f82, 32'shec2cd128, 32'shec2b52d1, 32'shec29d47e, 
               32'shec28562d, 32'shec26d7e0, 32'shec255995, 32'shec23db4e, 32'shec225d09, 32'shec20dec8, 32'shec1f608a, 32'shec1de24f, 
               32'shec1c6417, 32'shec1ae5e2, 32'shec1967b0, 32'shec17e981, 32'shec166b55, 32'shec14ed2c, 32'shec136f06, 32'shec11f0e4, 
               32'shec1072c4, 32'shec0ef4a8, 32'shec0d768e, 32'shec0bf878, 32'shec0a7a65, 32'shec08fc55, 32'shec077e48, 32'shec06003e, 
               32'shec048237, 32'shec030433, 32'shec018632, 32'shec000835, 32'shebfe8a3a, 32'shebfd0c42, 32'shebfb8e4e, 32'shebfa105d, 
               32'shebf8926f, 32'shebf71483, 32'shebf5969b, 32'shebf418b6, 32'shebf29ad4, 32'shebf11cf6, 32'shebef9f1a, 32'shebee2141, 
               32'shebeca36c, 32'shebeb259a, 32'shebe9a7ca, 32'shebe829fe, 32'shebe6ac35, 32'shebe52e6f, 32'shebe3b0ac, 32'shebe232ec, 
               32'shebe0b52f, 32'shebdf3776, 32'shebddb9bf, 32'shebdc3c0c, 32'shebdabe5c, 32'shebd940ae, 32'shebd7c304, 32'shebd6455d, 
               32'shebd4c7ba, 32'shebd34a19, 32'shebd1cc7b, 32'shebd04ee1, 32'shebced149, 32'shebcd53b5, 32'shebcbd624, 32'shebca5896, 
               32'shebc8db0b, 32'shebc75d83, 32'shebc5dffe, 32'shebc4627d, 32'shebc2e4fe, 32'shebc16783, 32'shebbfea0b, 32'shebbe6c95, 
               32'shebbcef23, 32'shebbb71b5, 32'shebb9f449, 32'shebb876e0, 32'shebb6f97b, 32'shebb57c18, 32'shebb3feb9, 32'shebb2815d, 
               32'shebb10404, 32'shebaf86ae, 32'shebae095c, 32'shebac8c0c, 32'shebab0ec0, 32'sheba99176, 32'sheba81430, 32'sheba696ed, 
               32'sheba519ad, 32'sheba39c71, 32'sheba21f37, 32'sheba0a200, 32'sheb9f24cd, 32'sheb9da79d, 32'sheb9c2a70, 32'sheb9aad46, 
               32'sheb99301f, 32'sheb97b2fc, 32'sheb9635db, 32'sheb94b8be, 32'sheb933ba4, 32'sheb91be8d, 32'sheb904179, 32'sheb8ec468, 
               32'sheb8d475b, 32'sheb8bca50, 32'sheb8a4d49, 32'sheb88d045, 32'sheb875344, 32'sheb85d646, 32'sheb84594c, 32'sheb82dc54, 
               32'sheb815f60, 32'sheb7fe26f, 32'sheb7e6581, 32'sheb7ce896, 32'sheb7b6bae, 32'sheb79eeca, 32'sheb7871e8, 32'sheb76f50a, 
               32'sheb75782f, 32'sheb73fb57, 32'sheb727e83, 32'sheb7101b1, 32'sheb6f84e3, 32'sheb6e0818, 32'sheb6c8b50, 32'sheb6b0e8b, 
               32'sheb6991ca, 32'sheb68150b, 32'sheb669850, 32'sheb651b98, 32'sheb639ee3, 32'sheb622231, 32'sheb60a582, 32'sheb5f28d7, 
               32'sheb5dac2f, 32'sheb5c2f8a, 32'sheb5ab2e8, 32'sheb593649, 32'sheb57b9ae, 32'sheb563d16, 32'sheb54c081, 32'sheb5343ef, 
               32'sheb51c760, 32'sheb504ad4, 32'sheb4ece4c, 32'sheb4d51c7, 32'sheb4bd545, 32'sheb4a58c6, 32'sheb48dc4b, 32'sheb475fd2, 
               32'sheb45e35d, 32'sheb4466eb, 32'sheb42ea7c, 32'sheb416e11, 32'sheb3ff1a8, 32'sheb3e7543, 32'sheb3cf8e1, 32'sheb3b7c82, 
               32'sheb3a0027, 32'sheb3883ce, 32'sheb370779, 32'sheb358b27, 32'sheb340ed9, 32'sheb32928d, 32'sheb311645, 32'sheb2f99ff, 
               32'sheb2e1dbe, 32'sheb2ca17f, 32'sheb2b2543, 32'sheb29a90b, 32'sheb282cd6, 32'sheb26b0a4, 32'sheb253475, 32'sheb23b84a, 
               32'sheb223c22, 32'sheb20bffd, 32'sheb1f43db, 32'sheb1dc7bc, 32'sheb1c4ba1, 32'sheb1acf89, 32'sheb195374, 32'sheb17d762, 
               32'sheb165b54, 32'sheb14df49, 32'sheb136341, 32'sheb11e73c, 32'sheb106b3a, 32'sheb0eef3c, 32'sheb0d7341, 32'sheb0bf749, 
               32'sheb0a7b54, 32'sheb08ff63, 32'sheb078375, 32'sheb06078a, 32'sheb048ba2, 32'sheb030fbe, 32'sheb0193dd, 32'sheb0017ff, 
               32'sheafe9c24, 32'sheafd204c, 32'sheafba478, 32'sheafa28a7, 32'sheaf8acd9, 32'sheaf7310f, 32'sheaf5b547, 32'sheaf43983, 
               32'sheaf2bdc3, 32'sheaf14205, 32'sheaefc64b, 32'sheaee4a94, 32'sheaeccee0, 32'sheaeb532f, 32'sheae9d782, 32'sheae85bd8, 
               32'sheae6e031, 32'sheae5648e, 32'sheae3e8ed, 32'sheae26d50, 32'sheae0f1b6, 32'sheadf7620, 32'sheaddfa8d, 32'sheadc7efd, 
               32'sheadb0370, 32'shead987e6, 32'shead80c60, 32'shead690dd, 32'shead5155d, 32'shead399e1, 32'shead21e68, 32'shead0a2f2, 
               32'sheacf277f, 32'sheacdac10, 32'sheacc30a4, 32'sheacab53b, 32'sheac939d5, 32'sheac7be73, 32'sheac64314, 32'sheac4c7b8, 
               32'sheac34c60, 32'sheac1d10b, 32'sheac055b9, 32'sheabeda6a, 32'sheabd5f1f, 32'sheabbe3d7, 32'sheaba6892, 32'sheab8ed50, 
               32'sheab77212, 32'sheab5f6d7, 32'sheab47b9f, 32'sheab3006b, 32'sheab1853a, 32'sheab00a0c, 32'sheaae8ee2, 32'sheaad13ba, 
               32'sheaab9896, 32'sheaaa1d76, 32'sheaa8a258, 32'sheaa7273e, 32'sheaa5ac27, 32'sheaa43114, 32'sheaa2b604, 32'sheaa13af7, 
               32'shea9fbfed, 32'shea9e44e7, 32'shea9cc9e4, 32'shea9b4ee4, 32'shea99d3e8, 32'shea9858ee, 32'shea96ddf9, 32'shea956306, 
               32'shea93e817, 32'shea926d2b, 32'shea90f242, 32'shea8f775d, 32'shea8dfc7b, 32'shea8c819c, 32'shea8b06c1, 32'shea898be9, 
               32'shea881114, 32'shea869642, 32'shea851b74, 32'shea83a0a9, 32'shea8225e2, 32'shea80ab1e, 32'shea7f305d, 32'shea7db59f, 
               32'shea7c3ae5, 32'shea7ac02e, 32'shea79457a, 32'shea77caca, 32'shea76501d, 32'shea74d573, 32'shea735acd, 32'shea71e02a, 
               32'shea70658a, 32'shea6eeaee, 32'shea6d7055, 32'shea6bf5bf, 32'shea6a7b2d, 32'shea69009e, 32'shea678612, 32'shea660b8a, 
               32'shea649105, 32'shea631683, 32'shea619c04, 32'shea602189, 32'shea5ea712, 32'shea5d2c9d, 32'shea5bb22c, 32'shea5a37be, 
               32'shea58bd54, 32'shea5742ed, 32'shea55c889, 32'shea544e29, 32'shea52d3cc, 32'shea515972, 32'shea4fdf1c, 32'shea4e64c9, 
               32'shea4cea79, 32'shea4b702d, 32'shea49f5e4, 32'shea487b9e, 32'shea47015c, 32'shea45871d, 32'shea440ce1, 32'shea4292a9, 
               32'shea411874, 32'shea3f9e43, 32'shea3e2415, 32'shea3ca9ea, 32'shea3b2fc2, 32'shea39b59e, 32'shea383b7e, 32'shea36c160, 
               32'shea354746, 32'shea33cd30, 32'shea32531c, 32'shea30d90c, 32'shea2f5f00, 32'shea2de4f7, 32'shea2c6af1, 32'shea2af0ee, 
               32'shea2976ef, 32'shea27fcf4, 32'shea2682fb, 32'shea250906, 32'shea238f15, 32'shea221526, 32'shea209b3b, 32'shea1f2154, 
               32'shea1da770, 32'shea1c2d8f, 32'shea1ab3b2, 32'shea1939d8, 32'shea17c001, 32'shea16462e, 32'shea14cc5e, 32'shea135291, 
               32'shea11d8c8, 32'shea105f03, 32'shea0ee540, 32'shea0d6b81, 32'shea0bf1c6, 32'shea0a780e, 32'shea08fe59, 32'shea0784a7, 
               32'shea060af9, 32'shea04914f, 32'shea0317a7, 32'shea019e04, 32'shea002463, 32'she9feaac6, 32'she9fd312c, 32'she9fbb796, 
               32'she9fa3e03, 32'she9f8c474, 32'she9f74ae8, 32'she9f5d15f, 32'she9f457da, 32'she9f2de58, 32'she9f164d9, 32'she9efeb5e, 
               32'she9ee71e6, 32'she9ecf872, 32'she9eb7f01, 32'she9ea0594, 32'she9e88c2a, 32'she9e712c3, 32'she9e59960, 32'she9e42000, 
               32'she9e2a6a3, 32'she9e12d4a, 32'she9dfb3f5, 32'she9de3aa3, 32'she9dcc154, 32'she9db4808, 32'she9d9cec0, 32'she9d8557c, 
               32'she9d6dc3b, 32'she9d562fd, 32'she9d3e9c3, 32'she9d2708c, 32'she9d0f758, 32'she9cf7e28, 32'she9ce04fc, 32'she9cc8bd3, 
               32'she9cb12ad, 32'she9c9998a, 32'she9c8206b, 32'she9c6a750, 32'she9c52e38, 32'she9c3b523, 32'she9c23c12, 32'she9c0c304, 
               32'she9bf49fa, 32'she9bdd0f3, 32'she9bc57f0, 32'she9badeef, 32'she9b965f3, 32'she9b7ecfa, 32'she9b67404, 32'she9b4fb12, 
               32'she9b38223, 32'she9b20937, 32'she9b0904f, 32'she9af176b, 32'she9ad9e8a, 32'she9ac25ac, 32'she9aaacd2, 32'she9a933fb, 
               32'she9a7bb28, 32'she9a64258, 32'she9a4c98b, 32'she9a350c2, 32'she9a1d7fd, 32'she9a05f3b, 32'she99ee67c, 32'she99d6dc1, 
               32'she99bf509, 32'she99a7c55, 32'she99903a4, 32'she9978af7, 32'she996124d, 32'she99499a6, 32'she9932103, 32'she991a864, 
               32'she9902fc7, 32'she98eb72f, 32'she98d3e9a, 32'she98bc608, 32'she98a4d7a, 32'she988d4ef, 32'she9875c68, 32'she985e3e4, 
               32'she9846b63, 32'she982f2e6, 32'she9817a6d, 32'she98001f7, 32'she97e8984, 32'she97d1115, 32'she97b98aa, 32'she97a2042, 
               32'she978a7dd, 32'she9772f7c, 32'she975b71e, 32'she9743ec4, 32'she972c66d, 32'she9714e1a, 32'she96fd5ca, 32'she96e5d7e, 
               32'she96ce535, 32'she96b6cf0, 32'she969f4ae, 32'she9687c70, 32'she9670435, 32'she9658bfd, 32'she96413c9, 32'she9629b99, 
               32'she961236c, 32'she95fab43, 32'she95e331d, 32'she95cbafa, 32'she95b42db, 32'she959cac0, 32'she95852a8, 32'she956da93, 
               32'she9556282, 32'she953ea75, 32'she952726b, 32'she950fa64, 32'she94f8261, 32'she94e0a62, 32'she94c9266, 32'she94b1a6d, 
               32'she949a278, 32'she9482a87, 32'she946b299, 32'she9453aae, 32'she943c2c7, 32'she9424ae4, 32'she940d304, 32'she93f5b27, 
               32'she93de34e, 32'she93c6b79, 32'she93af3a7, 32'she9397bd8, 32'she938040d, 32'she9368c46, 32'she9351482, 32'she9339cc2, 
               32'she9322505, 32'she930ad4b, 32'she92f3596, 32'she92dbde3, 32'she92c4634, 32'she92ace89, 32'she92956e1, 32'she927df3d, 
               32'she926679c, 32'she924efff, 32'she9237866, 32'she92200cf, 32'she920893d, 32'she91f11ae, 32'she91d9a22, 32'she91c229a, 
               32'she91aab16, 32'she9193395, 32'she917bc17, 32'she916449d, 32'she914cd27, 32'she91355b4, 32'she911de45, 32'she91066d9, 
               32'she90eef71, 32'she90d780c, 32'she90c00ab, 32'she90a894d, 32'she90911f3, 32'she9079a9d, 32'she906234a, 32'she904abfa, 
               32'she90334af, 32'she901bd66, 32'she9004621, 32'she8fecee0, 32'she8fd57a2, 32'she8fbe068, 32'she8fa6932, 32'she8f8f1ff, 
               32'she8f77acf, 32'she8f603a3, 32'she8f48c7b, 32'she8f31556, 32'she8f19e34, 32'she8f02717, 32'she8eeaffd, 32'she8ed38e6, 
               32'she8ebc1d3, 32'she8ea4ac3, 32'she8e8d3b7, 32'she8e75caf, 32'she8e5e5aa, 32'she8e46ea9, 32'she8e2f7ab, 32'she8e180b1, 
               32'she8e009ba, 32'she8de92c7, 32'she8dd1bd8, 32'she8dba4ec, 32'she8da2e04, 32'she8d8b71f, 32'she8d7403e, 32'she8d5c960, 
               32'she8d45286, 32'she8d2dbb0, 32'she8d164dd, 32'she8cfee0e, 32'she8ce7742, 32'she8cd007a, 32'she8cb89b5, 32'she8ca12f4, 
               32'she8c89c37, 32'she8c7257d, 32'she8c5aec7, 32'she8c43814, 32'she8c2c165, 32'she8c14aba, 32'she8bfd412, 32'she8be5d6d, 
               32'she8bce6cd, 32'she8bb702f, 32'she8b9f996, 32'she8b88300, 32'she8b70c6d, 32'she8b595df, 32'she8b41f53, 32'she8b2a8cc, 
               32'she8b13248, 32'she8afbbc7, 32'she8ae454b, 32'she8acced1, 32'she8ab585c, 32'she8a9e1ea, 32'she8a86b7b, 32'she8a6f510, 
               32'she8a57ea9, 32'she8a40845, 32'she8a291e5, 32'she8a11b89, 32'she89fa530, 32'she89e2edb, 32'she89cb889, 32'she89b423b, 
               32'she899cbf1, 32'she89855aa, 32'she896df67, 32'she8956927, 32'she893f2eb, 32'she8927cb3, 32'she891067e, 32'she88f904d, 
               32'she88e1a20, 32'she88ca3f6, 32'she88b2dcf, 32'she889b7ad, 32'she888418e, 32'she886cb72, 32'she885555a, 32'she883df46, 
               32'she8826936, 32'she880f329, 32'she87f7d1f, 32'she87e071a, 32'she87c9118, 32'she87b1b19, 32'she879a51e, 32'she8782f27, 
               32'she876b934, 32'she8754344, 32'she873cd57, 32'she872576f, 32'she870e18a, 32'she86f6ba8, 32'she86df5cb, 32'she86c7ff0, 
               32'she86b0a1a, 32'she8699447, 32'she8681e78, 32'she866a8ac, 32'she86532e4, 32'she863bd20, 32'she862475f, 32'she860d1a2, 
               32'she85f5be9, 32'she85de633, 32'she85c7081, 32'she85afad3, 32'she8598528, 32'she8580f81, 32'she85699dd, 32'she855243d, 
               32'she853aea1, 32'she8523909, 32'she850c374, 32'she84f4de2, 32'she84dd855, 32'she84c62cb, 32'she84aed45, 32'she84977c2, 
               32'she8480243, 32'she8468cc8, 32'she8451750, 32'she843a1dc, 32'she8422c6c, 32'she840b6ff, 32'she83f4196, 32'she83dcc31, 
               32'she83c56cf, 32'she83ae171, 32'she8396c16, 32'she837f6c0, 32'she836816d, 32'she8350c1d, 32'she83396d2, 32'she832218a, 
               32'she830ac45, 32'she82f3705, 32'she82dc1c8, 32'she82c4c8e, 32'she82ad759, 32'she8296227, 32'she827ecf8, 32'she82677ce, 
               32'she82502a7, 32'she8238d84, 32'she8221864, 32'she820a348, 32'she81f2e30, 32'she81db91b, 32'she81c440a, 32'she81acefd, 
               32'she81959f4, 32'she817e4ee, 32'she8166fec, 32'she814faed, 32'she81385f3, 32'she81210fc, 32'she8109c08, 32'she80f2719, 
               32'she80db22d, 32'she80c3d44, 32'she80ac860, 32'she809537f, 32'she807dea2, 32'she80669c8, 32'she804f4f2, 32'she8038020, 
               32'she8020b52, 32'she8009687, 32'she7ff21c0, 32'she7fdacfd, 32'she7fc383d, 32'she7fac381, 32'she7f94ec9, 32'she7f7da14, 
               32'she7f66564, 32'she7f4f0b7, 32'she7f37c0d, 32'she7f20768, 32'she7f092c6, 32'she7ef1e27, 32'she7eda98d, 32'she7ec34f6, 
               32'she7eac063, 32'she7e94bd3, 32'she7e7d748, 32'she7e662c0, 32'she7e4ee3c, 32'she7e379bb, 32'she7e2053e, 32'she7e090c5, 
               32'she7df1c50, 32'she7dda7de, 32'she7dc3370, 32'she7dabf06, 32'she7d94a9f, 32'she7d7d63d, 32'she7d661de, 32'she7d4ed82, 
               32'she7d3792b, 32'she7d204d7, 32'she7d09087, 32'she7cf1c3a, 32'she7cda7f2, 32'she7cc33ad, 32'she7cabf6c, 32'she7c94b2e, 
               32'she7c7d6f4, 32'she7c662be, 32'she7c4ee8c, 32'she7c37a5e, 32'she7c20633, 32'she7c0920c, 32'she7bf1de8, 32'she7bda9c9, 
               32'she7bc35ad, 32'she7bac195, 32'she7b94d80, 32'she7b7d970, 32'she7b66563, 32'she7b4f15a, 32'she7b37d55, 32'she7b20953, 
               32'she7b09555, 32'she7af215b, 32'she7adad65, 32'she7ac3972, 32'she7aac583, 32'she7a95198, 32'she7a7ddb1, 32'she7a669cd, 
               32'she7a4f5ed, 32'she7a38211, 32'she7a20e39, 32'she7a09a64, 32'she79f2693, 32'she79db2c6, 32'she79c3efd, 32'she79acb37, 
               32'she7995776, 32'she797e3b8, 32'she7966ffd, 32'she794fc47, 32'she7938894, 32'she79214e5, 32'she790a13a, 32'she78f2d92, 
               32'she78db9ef, 32'she78c464f, 32'she78ad2b3, 32'she7895f1a, 32'she787eb86, 32'she78677f5, 32'she7850468, 32'she78390df, 
               32'she7821d59, 32'she780a9d8, 32'she77f365a, 32'she77dc2e0, 32'she77c4f69, 32'she77adbf7, 32'she7796888, 32'she777f51d, 
               32'she77681b6, 32'she7750e52, 32'she7739af2, 32'she7722797, 32'she770b43e, 32'she76f40ea, 32'she76dcd9a, 32'she76c5a4d, 
               32'she76ae704, 32'she76973bf, 32'she768007e, 32'she7668d40, 32'she7651a06, 32'she763a6d0, 32'she762339e, 32'she760c070, 
               32'she75f4d45, 32'she75dda1e, 32'she75c66fb, 32'she75af3dc, 32'she75980c1, 32'she7580da9, 32'she7569a95, 32'she7552785, 
               32'she753b479, 32'she7524171, 32'she750ce6c, 32'she74f5b6b, 32'she74de86f, 32'she74c7575, 32'she74b0280, 32'she7498f8f, 
               32'she7481ca1, 32'she746a9b7, 32'she74536d1, 32'she743c3ef, 32'she7425110, 32'she740de35, 32'she73f6b5f, 32'she73df88c, 
               32'she73c85bc, 32'she73b12f1, 32'she739a029, 32'she7382d66, 32'she736baa6, 32'she73547ea, 32'she733d531, 32'she732627d, 
               32'she730efcc, 32'she72f7d20, 32'she72e0a77, 32'she72c97d1, 32'she72b2530, 32'she729b293, 32'she7283ff9, 32'she726cd63, 
               32'she7255ad1, 32'she723e843, 32'she72275b9, 32'she7210332, 32'she71f90b0, 32'she71e1e31, 32'she71cabb6, 32'she71b393f, 
               32'she719c6cb, 32'she718545c, 32'she716e1f0, 32'she7156f89, 32'she713fd25, 32'she7128ac4, 32'she7111868, 32'she70fa610, 
               32'she70e33bb, 32'she70cc16b, 32'she70b4f1e, 32'she709dcd5, 32'she7086a8f, 32'she706f84e, 32'she7058611, 32'she70413d7, 
               32'she702a1a1, 32'she7012f6f, 32'she6ffbd41, 32'she6fe4b17, 32'she6fcd8f1, 32'she6fb66ce, 32'she6f9f4b0, 32'she6f88295, 
               32'she6f7107e, 32'she6f59e6b, 32'she6f42c5c, 32'she6f2ba51, 32'she6f14849, 32'she6efd645, 32'she6ee6446, 32'she6ecf24a, 
               32'she6eb8052, 32'she6ea0e5e, 32'she6e89c6d, 32'she6e72a81, 32'she6e5b899, 32'she6e446b4, 32'she6e2d4d3, 32'she6e162f6, 
               32'she6dff11d, 32'she6de7f48, 32'she6dd0d77, 32'she6db9ba9, 32'she6da29e0, 32'she6d8b81a, 32'she6d74658, 32'she6d5d49b, 
               32'she6d462e1, 32'she6d2f12a, 32'she6d17f78, 32'she6d00dca, 32'she6ce9c1f, 32'she6cd2a79, 32'she6cbb8d6, 32'she6ca4737, 
               32'she6c8d59c, 32'she6c76405, 32'she6c5f272, 32'she6c480e3, 32'she6c30f57, 32'she6c19dd0, 32'she6c02c4c, 32'she6bebacd, 
               32'she6bd4951, 32'she6bbd7d9, 32'she6ba6665, 32'she6b8f4f5, 32'she6b78389, 32'she6b61220, 32'she6b4a0bc, 32'she6b32f5b, 
               32'she6b1bdff, 32'she6b04ca6, 32'she6aedb51, 32'she6ad6a00, 32'she6abf8b3, 32'she6aa876a, 32'she6a91625, 32'she6a7a4e4, 
               32'she6a633a6, 32'she6a4c26d, 32'she6a35137, 32'she6a1e006, 32'she6a06ed8, 32'she69efdae, 32'she69d8c88, 32'she69c1b66, 
               32'she69aaa48, 32'she699392e, 32'she697c818, 32'she6965706, 32'she694e5f7, 32'she69374ed, 32'she69203e6, 32'she69092e4, 
               32'she68f21e5, 32'she68db0ea, 32'she68c3ff3, 32'she68acf00, 32'she6895e11, 32'she687ed26, 32'she6867c3f, 32'she6850b5c, 
               32'she6839a7c, 32'she68229a1, 32'she680b8ca, 32'she67f47f6, 32'she67dd727, 32'she67c665b, 32'she67af593, 32'she67984cf, 
               32'she6781410, 32'she676a354, 32'she675329c, 32'she673c1e8, 32'she6725138, 32'she670e08c, 32'she66f6fe3, 32'she66dff3f, 
               32'she66c8e9f, 32'she66b1e02, 32'she669ad6a, 32'she6683cd5, 32'she666cc45, 32'she6655bb8, 32'she663eb30, 32'she6627aab, 
               32'she6610a2a, 32'she65f99ae, 32'she65e2935, 32'she65cb8c0, 32'she65b484f, 32'she659d7e2, 32'she6586779, 32'she656f714, 
               32'she65586b3, 32'she6541656, 32'she652a5fc, 32'she65135a7, 32'she64fc556, 32'she64e5509, 32'she64ce4bf, 32'she64b747a, 
               32'she64a0438, 32'she64893fb, 32'she64723c2, 32'she645b38c, 32'she644435a, 32'she642d32d, 32'she6416303, 32'she63ff2de, 
               32'she63e82bc, 32'she63d129e, 32'she63ba285, 32'she63a326f, 32'she638c25d, 32'she637524f, 32'she635e245, 32'she6347240, 
               32'she633023e, 32'she6319240, 32'she6302246, 32'she62eb250, 32'she62d425e, 32'she62bd270, 32'she62a6286, 32'she628f2a0, 
               32'she62782be, 32'she62612e0, 32'she624a306, 32'she6233330, 32'she621c35e, 32'she6205390, 32'she61ee3c6, 32'she61d73ff, 
               32'she61c043d, 32'she61a947f, 32'she61924c5, 32'she617b50f, 32'she616455d, 32'she614d5af, 32'she6136605, 32'she611f65e, 
               32'she61086bc, 32'she60f171e, 32'she60da784, 32'she60c37ee, 32'she60ac85c, 32'she60958ce, 32'she607e944, 32'she60679bd, 
               32'she6050a3b, 32'she6039abd, 32'she6022b43, 32'she600bbcd, 32'she5ff4c5b, 32'she5fddced, 32'she5fc6d83, 32'she5fafe1d, 
               32'she5f98ebb, 32'she5f81f5d, 32'she5f6b003, 32'she5f540ad, 32'she5f3d15b, 32'she5f2620d, 32'she5f0f2c3, 32'she5ef837d, 
               32'she5ee143b, 32'she5eca4fd, 32'she5eb35c3, 32'she5e9c68d, 32'she5e8575b, 32'she5e6e82e, 32'she5e57904, 32'she5e409de, 
               32'she5e29abc, 32'she5e12b9f, 32'she5dfbc85, 32'she5de4d6f, 32'she5dcde5e, 32'she5db6f50, 32'she5da0047, 32'she5d89141, 
               32'she5d72240, 32'she5d5b342, 32'she5d44449, 32'she5d2d553, 32'she5d16662, 32'she5cff775, 32'she5ce888b, 32'she5cd19a6, 
               32'she5cbaac5, 32'she5ca3be8, 32'she5c8cd0f, 32'she5c75e3a, 32'she5c5ef69, 32'she5c4809c, 32'she5c311d3, 32'she5c1a30e, 
               32'she5c0344d, 32'she5bec590, 32'she5bd56d7, 32'she5bbe823, 32'she5ba7972, 32'she5b90ac6, 32'she5b79c1d, 32'she5b62d79, 
               32'she5b4bed8, 32'she5b3503c, 32'she5b1e1a3, 32'she5b0730f, 32'she5af047f, 32'she5ad95f3, 32'she5ac276b, 32'she5aab8e7, 
               32'she5a94a67, 32'she5a7dbeb, 32'she5a66d73, 32'she5a4feff, 32'she5a39090, 32'she5a22224, 32'she5a0b3bc, 32'she59f4559, 
               32'she59dd6f9, 32'she59c689e, 32'she59afa47, 32'she5998bf3, 32'she5981da4, 32'she596af59, 32'she5954112, 32'she593d2cf, 
               32'she5926490, 32'she590f656, 32'she58f881f, 32'she58e19ec, 32'she58cabbe, 32'she58b3d93, 32'she589cf6d, 32'she588614a, 
               32'she586f32c, 32'she5858512, 32'she58416fc, 32'she582a8ea, 32'she5813adc, 32'she57fccd2, 32'she57e5ecc, 32'she57cf0cb, 
               32'she57b82cd, 32'she57a14d4, 32'she578a6de, 32'she57738ed, 32'she575cb00, 32'she5745d17, 32'she572ef32, 32'she5718151, 
               32'she5701374, 32'she56ea59b, 32'she56d37c7, 32'she56bc9f6, 32'she56a5c2a, 32'she568ee61, 32'she567809d, 32'she56612dd, 
               32'she564a521, 32'she5633769, 32'she561c9b5, 32'she5605c06, 32'she55eee5a, 32'she55d80b2, 32'she55c130f, 32'she55aa570, 
               32'she55937d5, 32'she557ca3e, 32'she5565cab, 32'she554ef1c, 32'she5538191, 32'she552140a, 32'she550a688, 32'she54f3909, 
               32'she54dcb8f, 32'she54c5e19, 32'she54af0a7, 32'she5498339, 32'she54815cf, 32'she546a86a, 32'she5453b08, 32'she543cdab, 
               32'she5426051, 32'she540f2fc, 32'she53f85ab, 32'she53e185e, 32'she53cab15, 32'she53b3dd1, 32'she539d090, 32'she5386354, 
               32'she536f61b, 32'she53588e7, 32'she5341bb7, 32'she532ae8b, 32'she5314163, 32'she52fd440, 32'she52e6720, 32'she52cfa05, 
               32'she52b8cee, 32'she52a1fdb, 32'she528b2cc, 32'she52745c1, 32'she525d8ba, 32'she5246bb8, 32'she522feb9, 32'she52191bf, 
               32'she52024c9, 32'she51eb7d7, 32'she51d4ae9, 32'she51bddff, 32'she51a711a, 32'she5190438, 32'she517975b, 32'she5162a82, 
               32'she514bdad, 32'she51350dc, 32'she511e410, 32'she5107747, 32'she50f0a83, 32'she50d9dc3, 32'she50c3107, 32'she50ac44f, 
               32'she509579b, 32'she507eaec, 32'she5067e40, 32'she5051199, 32'she503a4f6, 32'she5023857, 32'she500cbbc, 32'she4ff5f26, 
               32'she4fdf294, 32'she4fc8605, 32'she4fb197b, 32'she4f9acf5, 32'she4f84074, 32'she4f6d3f6, 32'she4f5677d, 32'she4f3fb07, 
               32'she4f28e96, 32'she4f12229, 32'she4efb5c1, 32'she4ee495c, 32'she4ecdcfc, 32'she4eb70a0, 32'she4ea0448, 32'she4e897f4, 
               32'she4e72ba4, 32'she4e5bf59, 32'she4e45311, 32'she4e2e6ce, 32'she4e17a8f, 32'she4e00e54, 32'she4dea21e, 32'she4dd35eb, 
               32'she4dbc9bd, 32'she4da5d93, 32'she4d8f16d, 32'she4d7854c, 32'she4d6192e, 32'she4d4ad15, 32'she4d34100, 32'she4d1d4ef, 
               32'she4d068e2, 32'she4cefcda, 32'she4cd90d5, 32'she4cc24d5, 32'she4cab8d9, 32'she4c94ce2, 32'she4c7e0ee, 32'she4c674ff, 
               32'she4c50914, 32'she4c39d2d, 32'she4c2314a, 32'she4c0c56b, 32'she4bf5991, 32'she4bdedbb, 32'she4bc81e9, 32'she4bb161b, 
               32'she4b9aa52, 32'she4b83e8d, 32'she4b6d2cb, 32'she4b5670f, 32'she4b3fb56, 32'she4b28fa1, 32'she4b123f1, 32'she4afb845, 
               32'she4ae4c9d, 32'she4ace0fa, 32'she4ab755a, 32'she4aa09bf, 32'she4a89e28, 32'she4a73295, 32'she4a5c707, 32'she4a45b7c, 
               32'she4a2eff6, 32'she4a18474, 32'she4a018f7, 32'she49ead7d, 32'she49d4208, 32'she49bd697, 32'she49a6b2a, 32'she498ffc1, 
               32'she497945d, 32'she49628fd, 32'she494bda1, 32'she4935249, 32'she491e6f6, 32'she4907ba7, 32'she48f105c, 32'she48da515, 
               32'she48c39d3, 32'she48ace94, 32'she489635a, 32'she487f825, 32'she4868cf3, 32'she48521c6, 32'she483b69d, 32'she4824b78, 
               32'she480e057, 32'she47f753b, 32'she47e0a23, 32'she47c9f0f, 32'she47b33ff, 32'she479c8f4, 32'she4785ded, 32'she476f2ea, 
               32'she47587eb, 32'she4741cf1, 32'she472b1fa, 32'she4714709, 32'she46fdc1b, 32'she46e7131, 32'she46d064c, 32'she46b9b6b, 
               32'she46a308f, 32'she468c5b6, 32'she4675ae2, 32'she465f012, 32'she4648547, 32'she4631a7f, 32'she461afbc, 32'she46044fd, 
               32'she45eda43, 32'she45d6f8c, 32'she45c04da, 32'she45a9a2c, 32'she4592f83, 32'she457c4de, 32'she4565a3c, 32'she454efa0, 
               32'she4538507, 32'she4521a73, 32'she450afe3, 32'she44f4557, 32'she44ddad0, 32'she44c704d, 32'she44b05ce, 32'she4499b53, 
               32'she44830dd, 32'she446c66b, 32'she4455bfd, 32'she443f194, 32'she442872e, 32'she4411ccd, 32'she43fb271, 32'she43e4818, 
               32'she43cddc4, 32'she43b7374, 32'she43a0929, 32'she4389ee2, 32'she437349f, 32'she435ca60, 32'she4346026, 32'she432f5ef, 
               32'she4318bbe, 32'she4302190, 32'she42eb767, 32'she42d4d42, 32'she42be321, 32'she42a7905, 32'she4290eed, 32'she427a4d9, 
               32'she4263ac9, 32'she424d0be, 32'she42366b7, 32'she421fcb5, 32'she42092b6, 32'she41f28bc, 32'she41dbec7, 32'she41c54d5, 
               32'she41aeae8, 32'she41980ff, 32'she418171b, 32'she416ad3a, 32'she415435f, 32'she413d987, 32'she4126fb4, 32'she41105e5, 
               32'she40f9c1a, 32'she40e3254, 32'she40cc891, 32'she40b5ed4, 32'she409f51a, 32'she4088b65, 32'she40721b4, 32'she405b808, 
               32'she4044e60, 32'she402e4bc, 32'she4017b1c, 32'she4001181, 32'she3fea7ea, 32'she3fd3e57, 32'she3fbd4c9, 32'she3fa6b3f, 
               32'she3f901ba, 32'she3f79838, 32'she3f62ebb, 32'she3f4c542, 32'she3f35bce, 32'she3f1f25e, 32'she3f088f2, 32'she3ef1f8b, 
               32'she3edb628, 32'she3ec4cc9, 32'she3eae36f, 32'she3e97a19, 32'she3e810c7, 32'she3e6a77a, 32'she3e53e31, 32'she3e3d4ec, 
               32'she3e26bac, 32'she3e1026f, 32'she3df9938, 32'she3de3004, 32'she3dcc6d5, 32'she3db5dab, 32'she3d9f484, 32'she3d88b62, 
               32'she3d72245, 32'she3d5b92b, 32'she3d45016, 32'she3d2e706, 32'she3d17df9, 32'she3d014f1, 32'she3ceabee, 32'she3cd42ee, 
               32'she3cbd9f4, 32'she3ca70fd, 32'she3c9080b, 32'she3c79f1d, 32'she3c63633, 32'she3c4cd4e, 32'she3c3646d, 32'she3c1fb91, 
               32'she3c092b9, 32'she3bf29e5, 32'she3bdc116, 32'she3bc584b, 32'she3baef84, 32'she3b986c2, 32'she3b81e04, 32'she3b6b54a, 
               32'she3b54c95, 32'she3b3e3e4, 32'she3b27b38, 32'she3b1128f, 32'she3afa9ec, 32'she3ae414c, 32'she3acd8b1, 32'she3ab701b, 
               32'she3aa0788, 32'she3a89efa, 32'she3a73671, 32'she3a5cdec, 32'she3a4656b, 32'she3a2fcee, 32'she3a19476, 32'she3a02c03, 
               32'she39ec393, 32'she39d5b28, 32'she39bf2c2, 32'she39a8a60, 32'she3992202, 32'she397b9a8, 32'she3965153, 32'she394e903, 
               32'she39380b6, 32'she392186f, 32'she390b02b, 32'she38f47ec, 32'she38ddfb1, 32'she38c777b, 32'she38b0f49, 32'she389a71b, 
               32'she3883ef2, 32'she386d6cd, 32'she3856ead, 32'she3840691, 32'she3829e79, 32'she3813666, 32'she37fce57, 32'she37e664d, 
               32'she37cfe47, 32'she37b9645, 32'she37a2e48, 32'she378c64f, 32'she3775e5a, 32'she375f66a, 32'she3748e7f, 32'she3732697, 
               32'she371beb5, 32'she37056d6, 32'she36eeefc, 32'she36d8727, 32'she36c1f55, 32'she36ab788, 32'she3694fc0, 32'she367e7fc, 
               32'she366803c, 32'she3651881, 32'she363b0cb, 32'she3624918, 32'she360e16a, 32'she35f79c1, 32'she35e121c, 32'she35caa7b, 
               32'she35b42df, 32'she359db47, 32'she35873b3, 32'she3570c24, 32'she355a49a, 32'she3543d13, 32'she352d592, 32'she3516e14, 
               32'she350069b, 32'she34e9f27, 32'she34d37b7, 32'she34bd04b, 32'she34a68e4, 32'she3490181, 32'she3479a23, 32'she34632c9, 
               32'she344cb73, 32'she3436422, 32'she341fcd6, 32'she340958d, 32'she33f2e4a, 32'she33dc70a, 32'she33c5fcf, 32'she33af899, 
               32'she3399167, 32'she3382a39, 32'she336c310, 32'she3355beb, 32'she333f4cb, 32'she3328daf, 32'she3312698, 32'she32fbf85, 
               32'she32e5876, 32'she32cf16c, 32'she32b8a67, 32'she32a2365, 32'she328bc69, 32'she3275570, 32'she325ee7d, 32'she324878d, 
               32'she32320a2, 32'she321b9bc, 32'she32052da, 32'she31eebfc, 32'she31d8523, 32'she31c1e4e, 32'she31ab77e, 32'she31950b2, 
               32'she317e9eb, 32'she3168328, 32'she3151c6a, 32'she313b5b0, 32'she3124efa, 32'she310e849, 32'she30f819d, 32'she30e1af5, 
               32'she30cb451, 32'she30b4db2, 32'she309e717, 32'she3088081, 32'she30719ef, 32'she305b362, 32'she3044cd9, 32'she302e655, 
               32'she3017fd5, 32'she300195a, 32'she2feb2e3, 32'she2fd4c70, 32'she2fbe602, 32'she2fa7f99, 32'she2f91934, 32'she2f7b2d3, 
               32'she2f64c77, 32'she2f4e61f, 32'she2f37fcc, 32'she2f2197e, 32'she2f0b333, 32'she2ef4cee, 32'she2ede6ac, 32'she2ec8070, 
               32'she2eb1a37, 32'she2e9b404, 32'she2e84dd4, 32'she2e6e7aa, 32'she2e58183, 32'she2e41b62, 32'she2e2b544, 32'she2e14f2b, 
               32'she2dfe917, 32'she2de8307, 32'she2dd1cfc, 32'she2dbb6f5, 32'she2da50f3, 32'she2d8eaf5, 32'she2d784fb, 32'she2d61f07, 
               32'she2d4b916, 32'she2d3532a, 32'she2d1ed43, 32'she2d08760, 32'she2cf2182, 32'she2cdbba8, 32'she2cc55d2, 32'she2caf001, 
               32'she2c98a35, 32'she2c8246d, 32'she2c6beaa, 32'she2c558eb, 32'she2c3f331, 32'she2c28d7b, 32'she2c127c9, 32'she2bfc21d, 
               32'she2be5c74, 32'she2bcf6d1, 32'she2bb9131, 32'she2ba2b96, 32'she2b8c600, 32'she2b7606e, 32'she2b5fae1, 32'she2b49559, 
               32'she2b32fd4, 32'she2b1ca55, 32'she2b064da, 32'she2aeff63, 32'she2ad99f1, 32'she2ac3483, 32'she2aacf1a, 32'she2a969b6, 
               32'she2a80456, 32'she2a69efa, 32'she2a539a3, 32'she2a3d451, 32'she2a26f03, 32'she2a109b9, 32'she29fa474, 32'she29e3f34, 
               32'she29cd9f8, 32'she29b74c1, 32'she29a0f8e, 32'she298aa60, 32'she2974536, 32'she295e011, 32'she2947af1, 32'she29315d5, 
               32'she291b0bd, 32'she2904baa, 32'she28ee69c, 32'she28d8192, 32'she28c1c8c, 32'she28ab78c, 32'she289528f, 32'she287ed98, 
               32'she28688a4, 32'she28523b6, 32'she283becc, 32'she28259e6, 32'she280f505, 32'she27f9029, 32'she27e2b51, 32'she27cc67d, 
               32'she27b61af, 32'she279fce4, 32'she278981f, 32'she277335e, 32'she275cea1, 32'she27469e9, 32'she2730536, 32'she271a087, 
               32'she2703bdc, 32'she26ed736, 32'she26d7295, 32'she26c0df9, 32'she26aa960, 32'she26944cd, 32'she267e03e, 32'she2667bb3, 
               32'she265172e, 32'she263b2ac, 32'she2624e2f, 32'she260e9b7, 32'she25f8544, 32'she25e20d5, 32'she25cbc6a, 32'she25b5804, 
               32'she259f3a3, 32'she2588f46, 32'she2572aee, 32'she255c69b, 32'she254624b, 32'she252fe01, 32'she25199bb, 32'she250357a, 
               32'she24ed13d, 32'she24d6d05, 32'she24c08d1, 32'she24aa4a2, 32'she2494078, 32'she247dc52, 32'she2467831, 32'she2451414, 
               32'she243affc, 32'she2424be9, 32'she240e7da, 32'she23f83d0, 32'she23e1fca, 32'she23cbbc9, 32'she23b57cc, 32'she239f3d4, 
               32'she2388fe1, 32'she2372bf2, 32'she235c808, 32'she2346422, 32'she2330041, 32'she2319c65, 32'she230388d, 32'she22ed4ba, 
               32'she22d70eb, 32'she22c0d21, 32'she22aa95c, 32'she229459b, 32'she227e1df, 32'she2267e28, 32'she2251a75, 32'she223b6c6, 
               32'she222531c, 32'she220ef77, 32'she21f8bd7, 32'she21e283b, 32'she21cc4a3, 32'she21b6111, 32'she219fd82, 32'she21899f9, 
               32'she2173674, 32'she215d2f4, 32'she2146f78, 32'she2130c01, 32'she211a88f, 32'she2104521, 32'she20ee1b7, 32'she20d7e53, 
               32'she20c1af3, 32'she20ab798, 32'she2095441, 32'she207f0ef, 32'she2068da1, 32'she2052a58, 32'she203c714, 32'she20263d4, 
               32'she2010099, 32'she1ff9d63, 32'she1fe3a31, 32'she1fcd704, 32'she1fb73dc, 32'she1fa10b8, 32'she1f8ad98, 32'she1f74a7e, 
               32'she1f5e768, 32'she1f48457, 32'she1f3214a, 32'she1f1be42, 32'she1f05b3e, 32'she1eef83f, 32'she1ed9545, 32'she1ec3250, 
               32'she1eacf5f, 32'she1e96c73, 32'she1e8098b, 32'she1e6a6a8, 32'she1e543ca, 32'she1e3e0f0, 32'she1e27e1b, 32'she1e11b4b, 
               32'she1dfb87f, 32'she1de55b8, 32'she1dcf2f5, 32'she1db9037, 32'she1da2d7e, 32'she1d8caca, 32'she1d7681a, 32'she1d6056f, 
               32'she1d4a2c8, 32'she1d34026, 32'she1d1dd89, 32'she1d07af0, 32'she1cf185c, 32'she1cdb5cd, 32'she1cc5342, 32'she1caf0bc, 
               32'she1c98e3b, 32'she1c82bbe, 32'she1c6c946, 32'she1c566d3, 32'she1c40464, 32'she1c2a1fa, 32'she1c13f95, 32'she1bfdd34, 
               32'she1be7ad8, 32'she1bd1881, 32'she1bbb62e, 32'she1ba53e0, 32'she1b8f197, 32'she1b78f52, 32'she1b62d12, 32'she1b4cad7, 
               32'she1b368a0, 32'she1b2066e, 32'she1b0a441, 32'she1af4218, 32'she1addff4, 32'she1ac7dd5, 32'she1ab1bba, 32'she1a9b9a4, 
               32'she1a85793, 32'she1a6f586, 32'she1a5937e, 32'she1a4317b, 32'she1a2cf7c, 32'she1a16d83, 32'she1a00b8d, 32'she19ea99d, 
               32'she19d47b1, 32'she19be5ca, 32'she19a83e7, 32'she199220a, 32'she197c031, 32'she1965e5c, 32'she194fc8d, 32'she1939ac2, 
               32'she19238fb, 32'she190d73a, 32'she18f757d, 32'she18e13c4, 32'she18cb211, 32'she18b5062, 32'she189eeb8, 32'she1888d13, 
               32'she1872b72, 32'she185c9d6, 32'she184683e, 32'she18306ac, 32'she181a51e, 32'she1804395, 32'she17ee210, 32'she17d8090, 
               32'she17c1f15, 32'she17abd9f, 32'she1795c2d, 32'she177fac0, 32'she1769958, 32'she17537f4, 32'she173d695, 32'she172753b, 
               32'she17113e5, 32'she16fb295, 32'she16e5149, 32'she16cf001, 32'she16b8ebf, 32'she16a2d81, 32'she168cc48, 32'she1676b13, 
               32'she16609e3, 32'she164a8b8, 32'she1634792, 32'she161e671, 32'she1608554, 32'she15f243c, 32'she15dc328, 32'she15c621a, 
               32'she15b0110, 32'she159a00a, 32'she1583f0a, 32'she156de0e, 32'she1557d17, 32'she1541c25, 32'she152bb37, 32'she1515a4e, 
               32'she14ff96a, 32'she14e988b, 32'she14d37b0, 32'she14bd6da, 32'she14a7609, 32'she149153c, 32'she147b475, 32'she14653b2, 
               32'she144f2f3, 32'she143923a, 32'she1423185, 32'she140d0d5, 32'she13f702a, 32'she13e0f83, 32'she13caee1, 32'she13b4e44, 
               32'she139edac, 32'she1388d19, 32'she1372c8a, 32'she135cc00, 32'she1346b7a, 32'she1330afa, 32'she131aa7e, 32'she1304a07, 
               32'she12ee995, 32'she12d8927, 32'she12c28be, 32'she12ac85a, 32'she12967fb, 32'she12807a0, 32'she126a74a, 32'she12546f9, 
               32'she123e6ad, 32'she1228666, 32'she1212623, 32'she11fc5e5, 32'she11e65ac, 32'she11d0577, 32'she11ba547, 32'she11a451c, 
               32'she118e4f6, 32'she11784d5, 32'she11624b8, 32'she114c4a0, 32'she113648d, 32'she112047f, 32'she110a475, 32'she10f4470, 
               32'she10de470, 32'she10c8475, 32'she10b247f, 32'she109c48d, 32'she10864a0, 32'she10704b8, 32'she105a4d4, 32'she10444f6, 
               32'she102e51c, 32'she1018547, 32'she1002577, 32'she0fec5ab, 32'she0fd65e4, 32'she0fc0622, 32'she0faa665, 32'she0f946ad, 
               32'she0f7e6f9, 32'she0f6874a, 32'she0f527a0, 32'she0f3c7fb, 32'she0f2685b, 32'she0f108bf, 32'she0efa928, 32'she0ee4996, 
               32'she0ecea09, 32'she0eb8a80, 32'she0ea2afd, 32'she0e8cb7e, 32'she0e76c04, 32'she0e60c8e, 32'she0e4ad1e, 32'she0e34db2, 
               32'she0e1ee4b, 32'she0e08ee9, 32'she0df2f8c, 32'she0ddd033, 32'she0dc70e0, 32'she0db1191, 32'she0d9b247, 32'she0d85301, 
               32'she0d6f3c1, 32'she0d59485, 32'she0d4354e, 32'she0d2d61c, 32'she0d176ef, 32'she0d017c6, 32'she0ceb8a3, 32'she0cd5984, 
               32'she0cbfa6a, 32'she0ca9b55, 32'she0c93c44, 32'she0c7dd39, 32'she0c67e32, 32'she0c51f30, 32'she0c3c033, 32'she0c2613a, 
               32'she0c10247, 32'she0bfa358, 32'she0be446e, 32'she0bce589, 32'she0bb86a9, 32'she0ba27cd, 32'she0b8c8f7, 32'she0b76a25, 
               32'she0b60b58, 32'she0b4ac90, 32'she0b34dcd, 32'she0b1ef0e, 32'she0b09055, 32'she0af31a0, 32'she0add2f0, 32'she0ac7445, 
               32'she0ab159e, 32'she0a9b6fd, 32'she0a85860, 32'she0a6f9c8, 32'she0a59b35, 32'she0a43ca7, 32'she0a2de1e, 32'she0a17f99, 
               32'she0a0211a, 32'she09ec29f, 32'she09d6429, 32'she09c05b8, 32'she09aa74b, 32'she09948e4, 32'she097ea81, 32'she0968c24, 
               32'she0952dcb, 32'she093cf77, 32'she0927127, 32'she09112dd, 32'she08fb497, 32'she08e5657, 32'she08cf81b, 32'she08b99e4, 
               32'she08a3bb2, 32'she088dd85, 32'she0877f5c, 32'she0862139, 32'she084c31a, 32'she0836500, 32'she08206eb, 32'she080a8db, 
               32'she07f4acf, 32'she07decc9, 32'she07c8ec7, 32'she07b30cb, 32'she079d2d3, 32'she07874e0, 32'she07716f2, 32'she075b908, 
               32'she0745b24, 32'she072fd44, 32'she0719f6a, 32'she0704194, 32'she06ee3c3, 32'she06d85f7, 32'she06c2830, 32'she06aca6d, 
               32'she0696cb0, 32'she0680ef7, 32'she066b144, 32'she0655395, 32'she063f5eb, 32'she0629846, 32'she0613aa5, 32'she05fdd0a, 
               32'she05e7f74, 32'she05d21e2, 32'she05bc455, 32'she05a66cd, 32'she059094a, 32'she057abcc, 32'she0564e53, 32'she054f0df, 
               32'she053936f, 32'she0523605, 32'she050d89f, 32'she04f7b3e, 32'she04e1de3, 32'she04cc08c, 32'she04b6339, 32'she04a05ec, 
               32'she048a8a4, 32'she0474b60, 32'she045ee22, 32'she04490e8, 32'she04333b3, 32'she041d684, 32'she0407959, 32'she03f1c33, 
               32'she03dbf11, 32'she03c61f5, 32'she03b04de, 32'she039a7cb, 32'she0384abe, 32'she036edb5, 32'she03590b1, 32'she03433b2, 
               32'she032d6b8, 32'she03179c3, 32'she0301cd3, 32'she02ebfe8, 32'she02d6301, 32'she02c0620, 32'she02aa943, 32'she0294c6c, 
               32'she027ef99, 32'she02692cb, 32'she0253602, 32'she023d93e, 32'she0227c7f, 32'she0211fc5, 32'she01fc310, 32'she01e6660, 
               32'she01d09b4, 32'she01bad0e, 32'she01a506c, 32'she018f3cf, 32'she0179738, 32'she0163aa5, 32'she014de17, 32'she013818e, 
               32'she012250a, 32'she010c88b, 32'she00f6c11, 32'she00e0f9b, 32'she00cb32b, 32'she00b56bf, 32'she009fa59, 32'she0089df7, 
               32'she007419b, 32'she005e543, 32'she00488f0, 32'she0032ca2, 32'she001d05a, 32'she0007416, 32'shdfff17d7, 32'shdffdbb9c, 
               32'shdffc5f67, 32'shdffb0337, 32'shdff9a70c, 32'shdff84ae5, 32'shdff6eec4, 32'shdff592a7, 32'shdff43690, 32'shdff2da7d, 
               32'shdff17e70, 32'shdff02267, 32'shdfeec663, 32'shdfed6a64, 32'shdfec0e6a, 32'shdfeab276, 32'shdfe95686, 32'shdfe7fa9b, 
               32'shdfe69eb4, 32'shdfe542d3, 32'shdfe3e6f7, 32'shdfe28b20, 32'shdfe12f4e, 32'shdfdfd380, 32'shdfde77b8, 32'shdfdd1bf5, 
               32'shdfdbc036, 32'shdfda647d, 32'shdfd908c8, 32'shdfd7ad18, 32'shdfd6516e, 32'shdfd4f5c8, 32'shdfd39a27, 32'shdfd23e8c, 
               32'shdfd0e2f5, 32'shdfcf8763, 32'shdfce2bd6, 32'shdfccd04e, 32'shdfcb74cb, 32'shdfca194d, 32'shdfc8bdd4, 32'shdfc76260, 
               32'shdfc606f1, 32'shdfc4ab87, 32'shdfc35022, 32'shdfc1f4c2, 32'shdfc09967, 32'shdfbf3e11, 32'shdfbde2bf, 32'shdfbc8773, 
               32'shdfbb2c2c, 32'shdfb9d0ea, 32'shdfb875ac, 32'shdfb71a74, 32'shdfb5bf41, 32'shdfb46412, 32'shdfb308e9, 32'shdfb1adc4, 
               32'shdfb052a5, 32'shdfaef78b, 32'shdfad9c75, 32'shdfac4165, 32'shdfaae659, 32'shdfa98b53, 32'shdfa83051, 32'shdfa6d554, 
               32'shdfa57a5d, 32'shdfa41f6a, 32'shdfa2c47d, 32'shdfa16994, 32'shdfa00eb1, 32'shdf9eb3d2, 32'shdf9d58f8, 32'shdf9bfe24, 
               32'shdf9aa354, 32'shdf99488a, 32'shdf97edc4, 32'shdf969303, 32'shdf953848, 32'shdf93dd91, 32'shdf9282df, 32'shdf912833, 
               32'shdf8fcd8b, 32'shdf8e72e8, 32'shdf8d184b, 32'shdf8bbdb2, 32'shdf8a631f, 32'shdf890890, 32'shdf87ae06, 32'shdf865382, 
               32'shdf84f902, 32'shdf839e88, 32'shdf824412, 32'shdf80e9a2, 32'shdf7f8f36, 32'shdf7e34cf, 32'shdf7cda6e, 32'shdf7b8011, 
               32'shdf7a25ba, 32'shdf78cb67, 32'shdf77711a, 32'shdf7616d2, 32'shdf74bc8e, 32'shdf736250, 32'shdf720816, 32'shdf70ade2, 
               32'shdf6f53b3, 32'shdf6df988, 32'shdf6c9f63, 32'shdf6b4543, 32'shdf69eb27, 32'shdf689111, 32'shdf673700, 32'shdf65dcf4, 
               32'shdf6482ed, 32'shdf6328eb, 32'shdf61ceee, 32'shdf6074f5, 32'shdf5f1b02, 32'shdf5dc114, 32'shdf5c672b, 32'shdf5b0d48, 
               32'shdf59b369, 32'shdf58598f, 32'shdf56ffba, 32'shdf55a5ea, 32'shdf544c1f, 32'shdf52f25a, 32'shdf519899, 32'shdf503edd, 
               32'shdf4ee527, 32'shdf4d8b75, 32'shdf4c31c9, 32'shdf4ad821, 32'shdf497e7f, 32'shdf4824e1, 32'shdf46cb49, 32'shdf4571b6, 
               32'shdf441828, 32'shdf42be9e, 32'shdf41651a, 32'shdf400b9b, 32'shdf3eb221, 32'shdf3d58ac, 32'shdf3bff3c, 32'shdf3aa5d1, 
               32'shdf394c6b, 32'shdf37f30b, 32'shdf3699af, 32'shdf354058, 32'shdf33e707, 32'shdf328dba, 32'shdf313473, 32'shdf2fdb30, 
               32'shdf2e81f3, 32'shdf2d28bb, 32'shdf2bcf87, 32'shdf2a7659, 32'shdf291d30, 32'shdf27c40c, 32'shdf266aed, 32'shdf2511d3, 
               32'shdf23b8be, 32'shdf225fae, 32'shdf2106a4, 32'shdf1fad9e, 32'shdf1e549d, 32'shdf1cfba2, 32'shdf1ba2ab, 32'shdf1a49ba, 
               32'shdf18f0ce, 32'shdf1797e7, 32'shdf163f04, 32'shdf14e627, 32'shdf138d4f, 32'shdf12347c, 32'shdf10dbaf, 32'shdf0f82e6, 
               32'shdf0e2a22, 32'shdf0cd163, 32'shdf0b78aa, 32'shdf0a1ff5, 32'shdf08c746, 32'shdf076e9c, 32'shdf0615f7, 32'shdf04bd57, 
               32'shdf0364bc, 32'shdf020c26, 32'shdf00b395, 32'shdeff5b09, 32'shdefe0282, 32'shdefcaa01, 32'shdefb5184, 32'shdef9f90d, 
               32'shdef8a09b, 32'shdef7482d, 32'shdef5efc5, 32'shdef49762, 32'shdef33f04, 32'shdef1e6ab, 32'shdef08e58, 32'shdeef3609, 
               32'shdeedddc0, 32'shdeec857b, 32'shdeeb2d3c, 32'shdee9d502, 32'shdee87ccc, 32'shdee7249c, 32'shdee5cc72, 32'shdee4744c, 
               32'shdee31c2b, 32'shdee1c40f, 32'shdee06bf9, 32'shdedf13e8, 32'shdeddbbdb, 32'shdedc63d4, 32'shdedb0bd2, 32'shded9b3d5, 
               32'shded85bdd, 32'shded703eb, 32'shded5abfd, 32'shded45414, 32'shded2fc31, 32'shded1a453, 32'shded04c7a, 32'shdecef4a6, 
               32'shdecd9cd7, 32'shdecc450d, 32'shdecaed48, 32'shdec99589, 32'shdec83dce, 32'shdec6e619, 32'shdec58e69, 32'shdec436be, 
               32'shdec2df18, 32'shdec18777, 32'shdec02fdb, 32'shdebed845, 32'shdebd80b3, 32'shdebc2927, 32'shdebad1a0, 32'shdeb97a1e, 
               32'shdeb822a1, 32'shdeb6cb29, 32'shdeb573b7, 32'shdeb41c49, 32'shdeb2c4e1, 32'shdeb16d7d, 32'shdeb0161f, 32'shdeaebec6, 
               32'shdead6773, 32'shdeac1024, 32'shdeaab8da, 32'shdea96196, 32'shdea80a57, 32'shdea6b31d, 32'shdea55be8, 32'shdea404b8, 
               32'shdea2ad8d, 32'shdea15668, 32'shde9fff47, 32'shde9ea82c, 32'shde9d5116, 32'shde9bfa05, 32'shde9aa2f9, 32'shde994bf2, 
               32'shde97f4f1, 32'shde969df5, 32'shde9546fd, 32'shde93f00b, 32'shde92991e, 32'shde914237, 32'shde8feb54, 32'shde8e9477, 
               32'shde8d3d9e, 32'shde8be6cb, 32'shde8a8ffd, 32'shde893935, 32'shde87e271, 32'shde868bb2, 32'shde8534f9, 32'shde83de45, 
               32'shde828796, 32'shde8130ec, 32'shde7fda48, 32'shde7e83a8, 32'shde7d2d0e, 32'shde7bd679, 32'shde7a7fe9, 32'shde79295e, 
               32'shde77d2d8, 32'shde767c58, 32'shde7525dc, 32'shde73cf66, 32'shde7278f5, 32'shde71228a, 32'shde6fcc23, 32'shde6e75c2, 
               32'shde6d1f65, 32'shde6bc90e, 32'shde6a72bc, 32'shde691c70, 32'shde67c628, 32'shde666fe6, 32'shde6519a9, 32'shde63c371, 
               32'shde626d3e, 32'shde611710, 32'shde5fc0e8, 32'shde5e6ac4, 32'shde5d14a6, 32'shde5bbe8d, 32'shde5a687a, 32'shde59126b, 
               32'shde57bc62, 32'shde56665e, 32'shde55105f, 32'shde53ba65, 32'shde526471, 32'shde510e81, 32'shde4fb897, 32'shde4e62b2, 
               32'shde4d0cd2, 32'shde4bb6f8, 32'shde4a6122, 32'shde490b52, 32'shde47b587, 32'shde465fc2, 32'shde450a01, 32'shde43b446, 
               32'shde425e8f, 32'shde4108de, 32'shde3fb333, 32'shde3e5d8c, 32'shde3d07eb, 32'shde3bb24f, 32'shde3a5cb8, 32'shde390726, 
               32'shde37b199, 32'shde365c12, 32'shde350690, 32'shde33b113, 32'shde325b9b, 32'shde310629, 32'shde2fb0bc, 32'shde2e5b54, 
               32'shde2d05f1, 32'shde2bb093, 32'shde2a5b3b, 32'shde2905e8, 32'shde27b09a, 32'shde265b51, 32'shde25060e, 32'shde23b0cf, 
               32'shde225b96, 32'shde210662, 32'shde1fb134, 32'shde1e5c0a, 32'shde1d06e6, 32'shde1bb1c7, 32'shde1a5cad, 32'shde190799, 
               32'shde17b28a, 32'shde165d80, 32'shde15087b, 32'shde13b37b, 32'shde125e81, 32'shde11098c, 32'shde0fb49c, 32'shde0e5fb1, 
               32'shde0d0acc, 32'shde0bb5ec, 32'shde0a6111, 32'shde090c3b, 32'shde07b76b, 32'shde06629f, 32'shde050dd9, 32'shde03b919, 
               32'shde02645d, 32'shde010fa7, 32'shddffbaf6, 32'shddfe664a, 32'shddfd11a3, 32'shddfbbd02, 32'shddfa6866, 32'shddf913cf, 
               32'shddf7bf3e, 32'shddf66ab1, 32'shddf5162a, 32'shddf3c1a9, 32'shddf26d2c, 32'shddf118b5, 32'shddefc443, 32'shddee6fd6, 
               32'shdded1b6e, 32'shddebc70c, 32'shddea72af, 32'shdde91e57, 32'shdde7ca05, 32'shdde675b7, 32'shdde5216f, 32'shdde3cd2d, 
               32'shdde278ef, 32'shdde124b7, 32'shdddfd084, 32'shddde7c56, 32'shdddd282e, 32'shdddbd40b, 32'shddda7fed, 32'shddd92bd4, 
               32'shddd7d7c1, 32'shddd683b3, 32'shddd52faa, 32'shddd3dba6, 32'shddd287a8, 32'shddd133af, 32'shddcfdfbb, 32'shddce8bcd, 
               32'shddcd37e4, 32'shddcbe400, 32'shddca9021, 32'shddc93c48, 32'shddc7e873, 32'shddc694a5, 32'shddc540db, 32'shddc3ed17, 
               32'shddc29958, 32'shddc1459e, 32'shddbff1ea, 32'shddbe9e3a, 32'shddbd4a91, 32'shddbbf6ec, 32'shddbaa34d, 32'shddb94fb3, 
               32'shddb7fc1e, 32'shddb6a88f, 32'shddb55504, 32'shddb4017f, 32'shddb2ae00, 32'shddb15a86, 32'shddb00711, 32'shddaeb3a1, 
               32'shddad6036, 32'shddac0cd1, 32'shddaab972, 32'shdda96617, 32'shdda812c2, 32'shdda6bf72, 32'shdda56c27, 32'shdda418e2, 
               32'shdda2c5a2, 32'shdda17267, 32'shdda01f32, 32'shdd9ecc01, 32'shdd9d78d7, 32'shdd9c25b1, 32'shdd9ad291, 32'shdd997f76, 
               32'shdd982c60, 32'shdd96d950, 32'shdd958645, 32'shdd94333f, 32'shdd92e03f, 32'shdd918d44, 32'shdd903a4e, 32'shdd8ee75d, 
               32'shdd8d9472, 32'shdd8c418c, 32'shdd8aeeac, 32'shdd899bd1, 32'shdd8848fb, 32'shdd86f62a, 32'shdd85a35f, 32'shdd845099, 
               32'shdd82fdd8, 32'shdd81ab1d, 32'shdd805867, 32'shdd7f05b6, 32'shdd7db30b, 32'shdd7c6065, 32'shdd7b0dc4, 32'shdd79bb29, 
               32'shdd786892, 32'shdd771602, 32'shdd75c376, 32'shdd7470f0, 32'shdd731e6f, 32'shdd71cbf4, 32'shdd70797e, 32'shdd6f270d, 
               32'shdd6dd4a2, 32'shdd6c823b, 32'shdd6b2fdb, 32'shdd69dd7f, 32'shdd688b29, 32'shdd6738d8, 32'shdd65e68d, 32'shdd649447, 
               32'shdd634206, 32'shdd61efcb, 32'shdd609d94, 32'shdd5f4b64, 32'shdd5df938, 32'shdd5ca712, 32'shdd5b54f1, 32'shdd5a02d6, 
               32'shdd58b0c0, 32'shdd575eaf, 32'shdd560ca4, 32'shdd54ba9e, 32'shdd53689d, 32'shdd5216a2, 32'shdd50c4ac, 32'shdd4f72bb, 
               32'shdd4e20d0, 32'shdd4cceea, 32'shdd4b7d09, 32'shdd4a2b2e, 32'shdd48d958, 32'shdd478788, 32'shdd4635bd, 32'shdd44e3f7, 
               32'shdd439236, 32'shdd42407b, 32'shdd40eec5, 32'shdd3f9d15, 32'shdd3e4b6a, 32'shdd3cf9c4, 32'shdd3ba824, 32'shdd3a5689, 
               32'shdd3904f4, 32'shdd37b363, 32'shdd3661d8, 32'shdd351053, 32'shdd33bed3, 32'shdd326d58, 32'shdd311be3, 32'shdd2fca73, 
               32'shdd2e7908, 32'shdd2d27a3, 32'shdd2bd643, 32'shdd2a84e8, 32'shdd293393, 32'shdd27e243, 32'shdd2690f9, 32'shdd253fb4, 
               32'shdd23ee74, 32'shdd229d3a, 32'shdd214c05, 32'shdd1ffad5, 32'shdd1ea9ab, 32'shdd1d5886, 32'shdd1c0767, 32'shdd1ab64d, 
               32'shdd196538, 32'shdd181429, 32'shdd16c31f, 32'shdd15721b, 32'shdd14211b, 32'shdd12d022, 32'shdd117f2d, 32'shdd102e3e, 
               32'shdd0edd55, 32'shdd0d8c71, 32'shdd0c3b92, 32'shdd0aeab9, 32'shdd0999e4, 32'shdd084916, 32'shdd06f84d, 32'shdd05a789, 
               32'shdd0456ca, 32'shdd030611, 32'shdd01b55e, 32'shdd0064af, 32'shdcff1407, 32'shdcfdc363, 32'shdcfc72c5, 32'shdcfb222c, 
               32'shdcf9d199, 32'shdcf8810b, 32'shdcf73083, 32'shdcf5e000, 32'shdcf48f82, 32'shdcf33f0a, 32'shdcf1ee97, 32'shdcf09e2a, 
               32'shdcef4dc2, 32'shdcedfd5f, 32'shdcecad02, 32'shdceb5caa, 32'shdcea0c58, 32'shdce8bc0b, 32'shdce76bc3, 32'shdce61b81, 
               32'shdce4cb44, 32'shdce37b0d, 32'shdce22adb, 32'shdce0daae, 32'shdcdf8a87, 32'shdcde3a66, 32'shdcdcea49, 32'shdcdb9a32, 
               32'shdcda4a21, 32'shdcd8fa15, 32'shdcd7aa0e, 32'shdcd65a0d, 32'shdcd50a12, 32'shdcd3ba1b, 32'shdcd26a2a, 32'shdcd11a3f, 
               32'shdccfca59, 32'shdcce7a78, 32'shdccd2a9d, 32'shdccbdac7, 32'shdcca8af7, 32'shdcc93b2c, 32'shdcc7eb67, 32'shdcc69ba7, 
               32'shdcc54bec, 32'shdcc3fc37, 32'shdcc2ac87, 32'shdcc15cdd, 32'shdcc00d38, 32'shdcbebd99, 32'shdcbd6dff, 32'shdcbc1e6a, 
               32'shdcbacedb, 32'shdcb97f51, 32'shdcb82fcd, 32'shdcb6e04e, 32'shdcb590d5, 32'shdcb44161, 32'shdcb2f1f3, 32'shdcb1a28a, 
               32'shdcb05326, 32'shdcaf03c8, 32'shdcadb46f, 32'shdcac651c, 32'shdcab15ce, 32'shdca9c686, 32'shdca87743, 32'shdca72805, 
               32'shdca5d8cd, 32'shdca4899b, 32'shdca33a6e, 32'shdca1eb46, 32'shdca09c24, 32'shdc9f4d07, 32'shdc9dfdf0, 32'shdc9caede, 
               32'shdc9b5fd2, 32'shdc9a10cb, 32'shdc98c1ca, 32'shdc9772ce, 32'shdc9623d7, 32'shdc94d4e6, 32'shdc9385fa, 32'shdc923714, 
               32'shdc90e834, 32'shdc8f9958, 32'shdc8e4a83, 32'shdc8cfbb2, 32'shdc8bace8, 32'shdc8a5e22, 32'shdc890f62, 32'shdc87c0a8, 
               32'shdc8671f3, 32'shdc852344, 32'shdc83d49a, 32'shdc8285f5, 32'shdc813756, 32'shdc7fe8bc, 32'shdc7e9a28, 32'shdc7d4b9a, 
               32'shdc7bfd11, 32'shdc7aae8d, 32'shdc79600f, 32'shdc781196, 32'shdc76c323, 32'shdc7574b5, 32'shdc74264d, 32'shdc72d7ea, 
               32'shdc71898d, 32'shdc703b35, 32'shdc6eece2, 32'shdc6d9e96, 32'shdc6c504e, 32'shdc6b020c, 32'shdc69b3d0, 32'shdc686599, 
               32'shdc671768, 32'shdc65c93c, 32'shdc647b15, 32'shdc632cf4, 32'shdc61ded9, 32'shdc6090c3, 32'shdc5f42b2, 32'shdc5df4a7, 
               32'shdc5ca6a2, 32'shdc5b58a2, 32'shdc5a0aa8, 32'shdc58bcb3, 32'shdc576ec3, 32'shdc5620d9, 32'shdc54d2f5, 32'shdc538516, 
               32'shdc52373c, 32'shdc50e968, 32'shdc4f9b9a, 32'shdc4e4dd1, 32'shdc4d000d, 32'shdc4bb24f, 32'shdc4a6497, 32'shdc4916e4, 
               32'shdc47c936, 32'shdc467b8e, 32'shdc452dec, 32'shdc43e04f, 32'shdc4292b8, 32'shdc414526, 32'shdc3ff799, 32'shdc3eaa12, 
               32'shdc3d5c91, 32'shdc3c0f15, 32'shdc3ac19f, 32'shdc39742e, 32'shdc3826c3, 32'shdc36d95d, 32'shdc358bfd, 32'shdc343ea2, 
               32'shdc32f14d, 32'shdc31a3fd, 32'shdc3056b3, 32'shdc2f096e, 32'shdc2dbc2f, 32'shdc2c6ef5, 32'shdc2b21c1, 32'shdc29d493, 
               32'shdc28876a, 32'shdc273a46, 32'shdc25ed28, 32'shdc24a010, 32'shdc2352fd, 32'shdc2205f0, 32'shdc20b8e8, 32'shdc1f6be5, 
               32'shdc1e1ee9, 32'shdc1cd1f1, 32'shdc1b8500, 32'shdc1a3813, 32'shdc18eb2d, 32'shdc179e4c, 32'shdc165170, 32'shdc15049a, 
               32'shdc13b7c9, 32'shdc126afe, 32'shdc111e39, 32'shdc0fd179, 32'shdc0e84bf, 32'shdc0d380a, 32'shdc0beb5b, 32'shdc0a9eb1, 
               32'shdc09520d, 32'shdc08056e, 32'shdc06b8d5, 32'shdc056c42, 32'shdc041fb4, 32'shdc02d32b, 32'shdc0186a8, 32'shdc003a2b, 
               32'shdbfeedb3, 32'shdbfda141, 32'shdbfc54d4, 32'shdbfb086d, 32'shdbf9bc0c, 32'shdbf86fb0, 32'shdbf72359, 32'shdbf5d708, 
               32'shdbf48abd, 32'shdbf33e77, 32'shdbf1f237, 32'shdbf0a5fc, 32'shdbef59c7, 32'shdbee0d98, 32'shdbecc16e, 32'shdbeb7549, 
               32'shdbea292b, 32'shdbe8dd11, 32'shdbe790fe, 32'shdbe644ef, 32'shdbe4f8e7, 32'shdbe3ace4, 32'shdbe260e6, 32'shdbe114ef, 
               32'shdbdfc8fc, 32'shdbde7d10, 32'shdbdd3128, 32'shdbdbe547, 32'shdbda996b, 32'shdbd94d94, 32'shdbd801c3, 32'shdbd6b5f8, 
               32'shdbd56a32, 32'shdbd41e72, 32'shdbd2d2b8, 32'shdbd18703, 32'shdbd03b53, 32'shdbceefaa, 32'shdbcda405, 32'shdbcc5867, 
               32'shdbcb0cce, 32'shdbc9c13a, 32'shdbc875ac, 32'shdbc72a24, 32'shdbc5dea1, 32'shdbc49324, 32'shdbc347ac, 32'shdbc1fc3a, 
               32'shdbc0b0ce, 32'shdbbf6567, 32'shdbbe1a06, 32'shdbbcceaa, 32'shdbbb8354, 32'shdbba3804, 32'shdbb8ecb9, 32'shdbb7a174, 
               32'shdbb65634, 32'shdbb50afa, 32'shdbb3bfc6, 32'shdbb27497, 32'shdbb1296e, 32'shdbafde4a, 32'shdbae932c, 32'shdbad4814, 
               32'shdbabfd01, 32'shdbaab1f3, 32'shdba966ec, 32'shdba81bea, 32'shdba6d0ed, 32'shdba585f7, 32'shdba43b05, 32'shdba2f01a, 
               32'shdba1a534, 32'shdba05a53, 32'shdb9f0f78, 32'shdb9dc4a3, 32'shdb9c79d4, 32'shdb9b2f0a, 32'shdb99e445, 32'shdb989987, 
               32'shdb974ece, 32'shdb96041a, 32'shdb94b96c, 32'shdb936ec4, 32'shdb922421, 32'shdb90d984, 32'shdb8f8eed, 32'shdb8e445b, 
               32'shdb8cf9cf, 32'shdb8baf48, 32'shdb8a64c7, 32'shdb891a4c, 32'shdb87cfd6, 32'shdb868566, 32'shdb853afc, 32'shdb83f097, 
               32'shdb82a638, 32'shdb815bde, 32'shdb80118a, 32'shdb7ec73c, 32'shdb7d7cf3, 32'shdb7c32b0, 32'shdb7ae873, 32'shdb799e3b, 
               32'shdb785409, 32'shdb7709dc, 32'shdb75bfb5, 32'shdb747594, 32'shdb732b79, 32'shdb71e163, 32'shdb709752, 32'shdb6f4d48, 
               32'shdb6e0342, 32'shdb6cb943, 32'shdb6b6f49, 32'shdb6a2555, 32'shdb68db67, 32'shdb67917e, 32'shdb66479b, 32'shdb64fdbd, 
               32'shdb63b3e5, 32'shdb626a13, 32'shdb612046, 32'shdb5fd67f, 32'shdb5e8cbe, 32'shdb5d4302, 32'shdb5bf94c, 32'shdb5aaf9c, 
               32'shdb5965f1, 32'shdb581c4c, 32'shdb56d2ac, 32'shdb558913, 32'shdb543f7e, 32'shdb52f5f0, 32'shdb51ac67, 32'shdb5062e4, 
               32'shdb4f1967, 32'shdb4dcfef, 32'shdb4c867d, 32'shdb4b3d10, 32'shdb49f3a9, 32'shdb48aa48, 32'shdb4760ec, 32'shdb461797, 
               32'shdb44ce46, 32'shdb4384fc, 32'shdb423bb7, 32'shdb40f278, 32'shdb3fa93e, 32'shdb3e600a, 32'shdb3d16dc, 32'shdb3bcdb3, 
               32'shdb3a8491, 32'shdb393b73, 32'shdb37f25c, 32'shdb36a94a, 32'shdb35603e, 32'shdb341737, 32'shdb32ce36, 32'shdb31853b, 
               32'shdb303c46, 32'shdb2ef356, 32'shdb2daa6c, 32'shdb2c6187, 32'shdb2b18a9, 32'shdb29cfcf, 32'shdb2886fc, 32'shdb273e2e, 
               32'shdb25f566, 32'shdb24aca4, 32'shdb2363e7, 32'shdb221b30, 32'shdb20d27f, 32'shdb1f89d3, 32'shdb1e412d, 32'shdb1cf88d, 
               32'shdb1baff2, 32'shdb1a675e, 32'shdb191ece, 32'shdb17d645, 32'shdb168dc1, 32'shdb154543, 32'shdb13fccb, 32'shdb12b458, 
               32'shdb116beb, 32'shdb102383, 32'shdb0edb22, 32'shdb0d92c6, 32'shdb0c4a70, 32'shdb0b021f, 32'shdb09b9d4, 32'shdb08718f, 
               32'shdb072950, 32'shdb05e116, 32'shdb0498e2, 32'shdb0350b4, 32'shdb02088b, 32'shdb00c068, 32'shdaff784b, 32'shdafe3033, 
               32'shdafce821, 32'shdafba015, 32'shdafa580f, 32'shdaf9100e, 32'shdaf7c813, 32'shdaf6801e, 32'shdaf5382e, 32'shdaf3f045, 
               32'shdaf2a860, 32'shdaf16082, 32'shdaf018a9, 32'shdaeed0d6, 32'shdaed8909, 32'shdaec4141, 32'shdaeaf980, 32'shdae9b1c4, 
               32'shdae86a0d, 32'shdae7225c, 32'shdae5dab2, 32'shdae4930c, 32'shdae34b6d, 32'shdae203d3, 32'shdae0bc3f, 32'shdadf74b1, 
               32'shdade2d28, 32'shdadce5a5, 32'shdadb9e28, 32'shdada56b0, 32'shdad90f3f, 32'shdad7c7d3, 32'shdad6806d, 32'shdad5390c, 
               32'shdad3f1b1, 32'shdad2aa5c, 32'shdad1630d, 32'shdad01bc3, 32'shdaced47f, 32'shdacd8d41, 32'shdacc4609, 32'shdacafed6, 
               32'shdac9b7a9, 32'shdac87082, 32'shdac72961, 32'shdac5e245, 32'shdac49b2f, 32'shdac3541f, 32'shdac20d15, 32'shdac0c610, 
               32'shdabf7f11, 32'shdabe3818, 32'shdabcf124, 32'shdabbaa36, 32'shdaba634e, 32'shdab91c6c, 32'shdab7d590, 32'shdab68eb9, 
               32'shdab547e8, 32'shdab4011d, 32'shdab2ba57, 32'shdab17397, 32'shdab02cdd, 32'shdaaee629, 32'shdaad9f7b, 32'shdaac58d2, 
               32'shdaab122f, 32'shdaa9cb92, 32'shdaa884fa, 32'shdaa73e69, 32'shdaa5f7dd, 32'shdaa4b157, 32'shdaa36ad6, 32'shdaa2245c, 
               32'shdaa0dde7, 32'shda9f9778, 32'shda9e510e, 32'shda9d0aab, 32'shda9bc44d, 32'shda9a7df5, 32'shda9937a2, 32'shda97f156, 
               32'shda96ab0f, 32'shda9564ce, 32'shda941e93, 32'shda92d85d, 32'shda91922e, 32'shda904c04, 32'shda8f05e0, 32'shda8dbfc1, 
               32'shda8c79a9, 32'shda8b3396, 32'shda89ed89, 32'shda88a782, 32'shda876180, 32'shda861b84, 32'shda84d58f, 32'shda838f9e, 
               32'shda8249b4, 32'shda8103cf, 32'shda7fbdf1, 32'shda7e7818, 32'shda7d3244, 32'shda7bec77, 32'shda7aa6af, 32'shda7960ed, 
               32'shda781b31, 32'shda76d57b, 32'shda758fcb, 32'shda744a20, 32'shda73047b, 32'shda71bedc, 32'shda707942, 32'shda6f33af, 
               32'shda6dee21, 32'shda6ca899, 32'shda6b6317, 32'shda6a1d9b, 32'shda68d824, 32'shda6792b3, 32'shda664d48, 32'shda6507e3, 
               32'shda63c284, 32'shda627d2a, 32'shda6137d6, 32'shda5ff288, 32'shda5ead40, 32'shda5d67fe, 32'shda5c22c1, 32'shda5add8a, 
               32'shda599859, 32'shda58532e, 32'shda570e09, 32'shda55c8e9, 32'shda5483d0, 32'shda533ebc, 32'shda51f9ae, 32'shda50b4a5, 
               32'shda4f6fa3, 32'shda4e2aa6, 32'shda4ce5af, 32'shda4ba0be, 32'shda4a5bd3, 32'shda4916ed, 32'shda47d20e, 32'shda468d34, 
               32'shda454860, 32'shda440392, 32'shda42beca, 32'shda417a07, 32'shda40354a, 32'shda3ef093, 32'shda3dabe2, 32'shda3c6737, 
               32'shda3b2292, 32'shda39ddf2, 32'shda389958, 32'shda3754c4, 32'shda361036, 32'shda34cbae, 32'shda33872c, 32'shda3242af, 
               32'shda30fe38, 32'shda2fb9c7, 32'shda2e755c, 32'shda2d30f7, 32'shda2bec97, 32'shda2aa83e, 32'shda2963ea, 32'shda281f9c, 
               32'shda26db54, 32'shda259711, 32'shda2452d5, 32'shda230e9e, 32'shda21ca6e, 32'shda208643, 32'shda1f421e, 32'shda1dfdfe, 
               32'shda1cb9e5, 32'shda1b75d1, 32'shda1a31c4, 32'shda18edbc, 32'shda17a9ba, 32'shda1665be, 32'shda1521c7, 32'shda13ddd7, 
               32'shda1299ec, 32'shda115607, 32'shda101228, 32'shda0ece4f, 32'shda0d8a7c, 32'shda0c46af, 32'shda0b02e7, 32'shda09bf25, 
               32'shda087b69, 32'shda0737b3, 32'shda05f403, 32'shda04b059, 32'shda036cb5, 32'shda022916, 32'shda00e57d, 32'shd9ffa1eb, 
               32'shd9fe5e5e, 32'shd9fd1ad6, 32'shd9fbd755, 32'shd9fa93da, 32'shd9f95064, 32'shd9f80cf5, 32'shd9f6c98b, 32'shd9f58627, 
               32'shd9f442c9, 32'shd9f2ff71, 32'shd9f1bc1e, 32'shd9f078d2, 32'shd9ef358b, 32'shd9edf24b, 32'shd9ecaf10, 32'shd9eb6bdb, 
               32'shd9ea28ac, 32'shd9e8e582, 32'shd9e7a25f, 32'shd9e65f42, 32'shd9e51c2a, 32'shd9e3d918, 32'shd9e2960c, 32'shd9e15306, 
               32'shd9e01006, 32'shd9decd0c, 32'shd9dd8a18, 32'shd9dc4729, 32'shd9db0441, 32'shd9d9c15e, 32'shd9d87e81, 32'shd9d73baa, 
               32'shd9d5f8d9, 32'shd9d4b60e, 32'shd9d37349, 32'shd9d23089, 32'shd9d0edd0, 32'shd9cfab1c, 32'shd9ce686e, 32'shd9cd25c7, 
               32'shd9cbe325, 32'shd9caa089, 32'shd9c95df3, 32'shd9c81b62, 32'shd9c6d8d8, 32'shd9c59653, 32'shd9c453d5, 32'shd9c3115c, 
               32'shd9c1cee9, 32'shd9c08c7c, 32'shd9bf4a15, 32'shd9be07b4, 32'shd9bcc559, 32'shd9bb8304, 32'shd9ba40b5, 32'shd9b8fe6b, 
               32'shd9b7bc27, 32'shd9b679ea, 32'shd9b537b2, 32'shd9b3f580, 32'shd9b2b354, 32'shd9b1712e, 32'shd9b02f0e, 32'shd9aeecf4, 
               32'shd9adaadf, 32'shd9ac68d1, 32'shd9ab26c8, 32'shd9a9e4c6, 32'shd9a8a2c9, 32'shd9a760d2, 32'shd9a61ee1, 32'shd9a4dcf6, 
               32'shd9a39b11, 32'shd9a25932, 32'shd9a11759, 32'shd99fd586, 32'shd99e93b8, 32'shd99d51f1, 32'shd99c102f, 32'shd99ace74, 
               32'shd9998cbe, 32'shd9984b0e, 32'shd9970965, 32'shd995c7c1, 32'shd9948623, 32'shd993448b, 32'shd99202f8, 32'shd990c16c, 
               32'shd98f7fe6, 32'shd98e3e66, 32'shd98cfceb, 32'shd98bbb77, 32'shd98a7a08, 32'shd989389f, 32'shd987f73d, 32'shd986b5e0, 
               32'shd9857489, 32'shd9843338, 32'shd982f1ed, 32'shd981b0a8, 32'shd9806f69, 32'shd97f2e30, 32'shd97decfd, 32'shd97cabcf, 
               32'shd97b6aa8, 32'shd97a2986, 32'shd978e86b, 32'shd977a755, 32'shd9766646, 32'shd975253c, 32'shd973e438, 32'shd972a33b, 
               32'shd9716243, 32'shd9702151, 32'shd96ee065, 32'shd96d9f7f, 32'shd96c5e9f, 32'shd96b1dc5, 32'shd969dcf1, 32'shd9689c23, 
               32'shd9675b5a, 32'shd9661a98, 32'shd964d9dc, 32'shd9639926, 32'shd9625875, 32'shd96117cb, 32'shd95fd726, 32'shd95e9688, 
               32'shd95d55ef, 32'shd95c155c, 32'shd95ad4d0, 32'shd9599449, 32'shd95853c8, 32'shd957134d, 32'shd955d2d9, 32'shd954926a, 
               32'shd9535201, 32'shd952119e, 32'shd950d141, 32'shd94f90ea, 32'shd94e5099, 32'shd94d104e, 32'shd94bd009, 32'shd94a8fca, 
               32'shd9494f90, 32'shd9480f5d, 32'shd946cf30, 32'shd9458f09, 32'shd9444ee7, 32'shd9430ecc, 32'shd941ceb7, 32'shd9408ea7, 
               32'shd93f4e9e, 32'shd93e0e9b, 32'shd93cce9d, 32'shd93b8ea6, 32'shd93a4eb4, 32'shd9390ec9, 32'shd937cee3, 32'shd9368f04, 
               32'shd9354f2a, 32'shd9340f56, 32'shd932cf89, 32'shd9318fc1, 32'shd9305000, 32'shd92f1044, 32'shd92dd08e, 32'shd92c90df, 
               32'shd92b5135, 32'shd92a1191, 32'shd928d1f4, 32'shd927925c, 32'shd92652ca, 32'shd925133e, 32'shd923d3b9, 32'shd9229439, 
               32'shd92154bf, 32'shd920154b, 32'shd91ed5de, 32'shd91d9676, 32'shd91c5714, 32'shd91b17b8, 32'shd919d863, 32'shd9189913, 
               32'shd91759c9, 32'shd9161a85, 32'shd914db47, 32'shd9139c10, 32'shd9125cde, 32'shd9111db2, 32'shd90fde8c, 32'shd90e9f6d, 
               32'shd90d6053, 32'shd90c213f, 32'shd90ae231, 32'shd909a32a, 32'shd9086428, 32'shd907252c, 32'shd905e636, 32'shd904a747, 
               32'shd903685d, 32'shd9022979, 32'shd900ea9c, 32'shd8ffabc4, 32'shd8fe6cf2, 32'shd8fd2e27, 32'shd8fbef61, 32'shd8fab0a2, 
               32'shd8f971e8, 32'shd8f83335, 32'shd8f6f487, 32'shd8f5b5df, 32'shd8f4773e, 32'shd8f338a3, 32'shd8f1fa0d, 32'shd8f0bb7e, 
               32'shd8ef7cf4, 32'shd8ee3e71, 32'shd8ecfff4, 32'shd8ebc17c, 32'shd8ea830b, 32'shd8e944a0, 32'shd8e8063a, 32'shd8e6c7db, 
               32'shd8e58982, 32'shd8e44b2f, 32'shd8e30ce2, 32'shd8e1ce9b, 32'shd8e0905a, 32'shd8df521f, 32'shd8de13ea, 32'shd8dcd5bb, 
               32'shd8db9792, 32'shd8da596f, 32'shd8d91b52, 32'shd8d7dd3b, 32'shd8d69f2a, 32'shd8d56120, 32'shd8d4231b, 32'shd8d2e51c, 
               32'shd8d1a724, 32'shd8d06931, 32'shd8cf2b45, 32'shd8cded5e, 32'shd8ccaf7e, 32'shd8cb71a3, 32'shd8ca33cf, 32'shd8c8f601, 
               32'shd8c7b838, 32'shd8c67a76, 32'shd8c53cba, 32'shd8c3ff04, 32'shd8c2c154, 32'shd8c183aa, 32'shd8c04606, 32'shd8bf0868, 
               32'shd8bdcad0, 32'shd8bc8d3e, 32'shd8bb4fb3, 32'shd8ba122d, 32'shd8b8d4ad, 32'shd8b79734, 32'shd8b659c0, 32'shd8b51c53, 
               32'shd8b3deeb, 32'shd8b2a18a, 32'shd8b1642f, 32'shd8b026da, 32'shd8aee98a, 32'shd8adac41, 32'shd8ac6efe, 32'shd8ab31c1, 
               32'shd8a9f48a, 32'shd8a8b75a, 32'shd8a77a2f, 32'shd8a63d0a, 32'shd8a4ffec, 32'shd8a3c2d3, 32'shd8a285c0, 32'shd8a148b4, 
               32'shd8a00bae, 32'shd89ecead, 32'shd89d91b3, 32'shd89c54bf, 32'shd89b17d1, 32'shd899dae9, 32'shd8989e07, 32'shd897612b, 
               32'shd8962456, 32'shd894e786, 32'shd893aabc, 32'shd8926df9, 32'shd891313b, 32'shd88ff484, 32'shd88eb7d3, 32'shd88d7b28, 
               32'shd88c3e83, 32'shd88b01e4, 32'shd889c54b, 32'shd88888b8, 32'shd8874c2b, 32'shd8860fa4, 32'shd884d324, 32'shd88396a9, 
               32'shd8825a35, 32'shd8811dc7, 32'shd87fe15e, 32'shd87ea4fc, 32'shd87d68a0, 32'shd87c2c4a, 32'shd87aeffa, 32'shd879b3b1, 
               32'shd878776d, 32'shd8773b2f, 32'shd875fef8, 32'shd874c2c7, 32'shd873869b, 32'shd8724a76, 32'shd8710e57, 32'shd86fd23e, 
               32'shd86e962b, 32'shd86d5a1e, 32'shd86c1e18, 32'shd86ae217, 32'shd869a61d, 32'shd8686a28, 32'shd8672e3a, 32'shd865f252, 
               32'shd864b670, 32'shd8637a94, 32'shd8623ebe, 32'shd86102ee, 32'shd85fc725, 32'shd85e8b61, 32'shd85d4fa4, 32'shd85c13ed, 
               32'shd85ad83c, 32'shd8599c91, 32'shd85860ec, 32'shd857254d, 32'shd855e9b4, 32'shd854ae21, 32'shd8537295, 32'shd852370f, 
               32'shd850fb8e, 32'shd84fc014, 32'shd84e84a0, 32'shd84d4933, 32'shd84c0dcb, 32'shd84ad269, 32'shd849970e, 32'shd8485bb8, 
               32'shd8472069, 32'shd845e520, 32'shd844a9dd, 32'shd8436ea0, 32'shd8423369, 32'shd840f839, 32'shd83fbd0e, 32'shd83e81ea, 
               32'shd83d46cc, 32'shd83c0bb4, 32'shd83ad0a2, 32'shd8399596, 32'shd8385a90, 32'shd8371f91, 32'shd835e497, 32'shd834a9a4, 
               32'shd8336eb7, 32'shd83233d0, 32'shd830f8ef, 32'shd82fbe14, 32'shd82e833f, 32'shd82d4871, 32'shd82c0da9, 32'shd82ad2e7, 
               32'shd829982b, 32'shd8285d75, 32'shd82722c5, 32'shd825e81b, 32'shd824ad78, 32'shd82372db, 32'shd8223843, 32'shd820fdb2, 
               32'shd81fc328, 32'shd81e88a3, 32'shd81d4e24, 32'shd81c13ac, 32'shd81ad93a, 32'shd8199ecd, 32'shd8186468, 32'shd8172a08, 
               32'shd815efae, 32'shd814b55b, 32'shd8137b0d, 32'shd81240c6, 32'shd8110685, 32'shd80fcc4a, 32'shd80e9216, 32'shd80d57e7, 
               32'shd80c1dbf, 32'shd80ae39c, 32'shd809a980, 32'shd8086f6a, 32'shd807355b, 32'shd805fb51, 32'shd804c14e, 32'shd8038751, 
               32'shd8024d59, 32'shd8011369, 32'shd7ffd97e, 32'shd7fe9f99, 32'shd7fd65bb, 32'shd7fc2be3, 32'shd7faf211, 32'shd7f9b845, 
               32'shd7f87e7f, 32'shd7f744bf, 32'shd7f60b06, 32'shd7f4d153, 32'shd7f397a6, 32'shd7f25dff, 32'shd7f1245e, 32'shd7efeac4, 
               32'shd7eeb130, 32'shd7ed77a1, 32'shd7ec3e1a, 32'shd7eb0498, 32'shd7e9cb1c, 32'shd7e891a7, 32'shd7e75838, 32'shd7e61ece, 
               32'shd7e4e56c, 32'shd7e3ac0f, 32'shd7e272b8, 32'shd7e13968, 32'shd7e0001e, 32'shd7dec6da, 32'shd7dd8d9c, 32'shd7dc5465, 
               32'shd7db1b34, 32'shd7d9e208, 32'shd7d8a8e3, 32'shd7d76fc5, 32'shd7d636ac, 32'shd7d4fd9a, 32'shd7d3c48d, 32'shd7d28b87, 
               32'shd7d15288, 32'shd7d0198e, 32'shd7cee09b, 32'shd7cda7ad, 32'shd7cc6ec6, 32'shd7cb35e6, 32'shd7c9fd0b, 32'shd7c8c436, 
               32'shd7c78b68, 32'shd7c652a0, 32'shd7c519de, 32'shd7c3e123, 32'shd7c2a86d, 32'shd7c16fbe, 32'shd7c03715, 32'shd7befe72, 
               32'shd7bdc5d6, 32'shd7bc8d40, 32'shd7bb54af, 32'shd7ba1c25, 32'shd7b8e3a2, 32'shd7b7ab24, 32'shd7b672ad, 32'shd7b53a3c, 
               32'shd7b401d1, 32'shd7b2c96c, 32'shd7b1910e, 32'shd7b058b6, 32'shd7af2063, 32'shd7ade818, 32'shd7acafd2, 32'shd7ab7793, 
               32'shd7aa3f5a, 32'shd7a90727, 32'shd7a7cefa, 32'shd7a696d3, 32'shd7a55eb3, 32'shd7a42699, 32'shd7a2ee85, 32'shd7a1b678, 
               32'shd7a07e70, 32'shd79f466f, 32'shd79e0e74, 32'shd79cd680, 32'shd79b9e91, 32'shd79a66a9, 32'shd7992ec7, 32'shd797f6eb, 
               32'shd796bf16, 32'shd7958746, 32'shd7944f7d, 32'shd79317ba, 32'shd791dffe, 32'shd790a847, 32'shd78f7097, 32'shd78e38ed, 
               32'shd78d014a, 32'shd78bc9ac, 32'shd78a9215, 32'shd7895a84, 32'shd78822f9, 32'shd786eb75, 32'shd785b3f7, 32'shd7847c7f, 
               32'shd783450d, 32'shd7820da1, 32'shd780d63c, 32'shd77f9edd, 32'shd77e6784, 32'shd77d3032, 32'shd77bf8e6, 32'shd77ac1a0, 
               32'shd7798a60, 32'shd7785326, 32'shd7771bf3, 32'shd775e4c6, 32'shd774ad9f, 32'shd773767f, 32'shd7723f64, 32'shd7710850, 
               32'shd76fd143, 32'shd76e9a3b, 32'shd76d633a, 32'shd76c2c3f, 32'shd76af54a, 32'shd769be5c, 32'shd7688774, 32'shd7675092, 
               32'shd76619b6, 32'shd764e2e0, 32'shd763ac11, 32'shd7627548, 32'shd7613e86, 32'shd76007c9, 32'shd75ed113, 32'shd75d9a63, 
               32'shd75c63ba, 32'shd75b2d17, 32'shd759f679, 32'shd758bfe3, 32'shd7578952, 32'shd75652c8, 32'shd7551c44, 32'shd753e5c6, 
               32'shd752af4f, 32'shd75178de, 32'shd7504273, 32'shd74f0c0e, 32'shd74dd5b0, 32'shd74c9f58, 32'shd74b6906, 32'shd74a32bb, 
               32'shd748fc75, 32'shd747c636, 32'shd7468ffe, 32'shd74559cb, 32'shd744239f, 32'shd742ed79, 32'shd741b75a, 32'shd7408141, 
               32'shd73f4b2e, 32'shd73e1521, 32'shd73cdf1b, 32'shd73ba91a, 32'shd73a7321, 32'shd7393d2d, 32'shd7380740, 32'shd736d159, 
               32'shd7359b78, 32'shd734659e, 32'shd7332fca, 32'shd731f9fc, 32'shd730c434, 32'shd72f8e73, 32'shd72e58b8, 32'shd72d2304, 
               32'shd72bed55, 32'shd72ab7ad, 32'shd729820c, 32'shd7284c70, 32'shd72716db, 32'shd725e14c, 32'shd724abc4, 32'shd7237641, 
               32'shd72240c5, 32'shd7210b50, 32'shd71fd5e0, 32'shd71ea077, 32'shd71d6b15, 32'shd71c35b8, 32'shd71b0062, 32'shd719cb12, 
               32'shd71895c9, 32'shd7176086, 32'shd7162b49, 32'shd714f612, 32'shd713c0e2, 32'shd7128bb8, 32'shd7115694, 32'shd7102177, 
               32'shd70eec60, 32'shd70db74f, 32'shd70c8245, 32'shd70b4d41, 32'shd70a1843, 32'shd708e34c, 32'shd707ae5a, 32'shd7067970, 
               32'shd705448b, 32'shd7040fad, 32'shd702dad5, 32'shd701a604, 32'shd7007138, 32'shd6ff3c73, 32'shd6fe07b5, 32'shd6fcd2fd, 
               32'shd6fb9e4b, 32'shd6fa699f, 32'shd6f934fa, 32'shd6f8005b, 32'shd6f6cbc2, 32'shd6f59730, 32'shd6f462a4, 32'shd6f32e1f, 
               32'shd6f1f99f, 32'shd6f0c526, 32'shd6ef90b4, 32'shd6ee5c47, 32'shd6ed27e1, 32'shd6ebf382, 32'shd6eabf28, 32'shd6e98ad6, 
               32'shd6e85689, 32'shd6e72243, 32'shd6e5ee03, 32'shd6e4b9c9, 32'shd6e38596, 32'shd6e25169, 32'shd6e11d42, 32'shd6dfe922, 
               32'shd6deb508, 32'shd6dd80f5, 32'shd6dc4ce7, 32'shd6db18e0, 32'shd6d9e4e0, 32'shd6d8b0e6, 32'shd6d77cf2, 32'shd6d64904, 
               32'shd6d5151d, 32'shd6d3e13d, 32'shd6d2ad62, 32'shd6d1798e, 32'shd6d045c0, 32'shd6cf11f9, 32'shd6cdde38, 32'shd6ccaa7d, 
               32'shd6cb76c9, 32'shd6ca431b, 32'shd6c90f73, 32'shd6c7dbd2, 32'shd6c6a837, 32'shd6c574a2, 32'shd6c44114, 32'shd6c30d8c, 
               32'shd6c1da0b, 32'shd6c0a690, 32'shd6bf731b, 32'shd6be3fad, 32'shd6bd0c45, 32'shd6bbd8e3, 32'shd6baa588, 32'shd6b97233, 
               32'shd6b83ee4, 32'shd6b70b9c, 32'shd6b5d85a, 32'shd6b4a51f, 32'shd6b371ea, 32'shd6b23ebb, 32'shd6b10b92, 32'shd6afd870, 
               32'shd6aea555, 32'shd6ad7240, 32'shd6ac3f31, 32'shd6ab0c28, 32'shd6a9d926, 32'shd6a8a62a, 32'shd6a77335, 32'shd6a64046, 
               32'shd6a50d5d, 32'shd6a3da7b, 32'shd6a2a79f, 32'shd6a174ca, 32'shd6a041fa, 32'shd69f0f32, 32'shd69ddc6f, 32'shd69ca9b3, 
               32'shd69b76fe, 32'shd69a444f, 32'shd69911a6, 32'shd697df03, 32'shd696ac67, 32'shd69579d2, 32'shd6944742, 32'shd69314b9, 
               32'shd691e237, 32'shd690afbb, 32'shd68f7d45, 32'shd68e4ad6, 32'shd68d186d, 32'shd68be60a, 32'shd68ab3ae, 32'shd6898158, 
               32'shd6884f09, 32'shd6871cc0, 32'shd685ea7d, 32'shd684b841, 32'shd683860b, 32'shd68253dc, 32'shd68121b3, 32'shd67fef90, 
               32'shd67ebd74, 32'shd67d8b5e, 32'shd67c594f, 32'shd67b2746, 32'shd679f543, 32'shd678c347, 32'shd6779151, 32'shd6765f62, 
               32'shd6752d79, 32'shd673fb97, 32'shd672c9ba, 32'shd67197e5, 32'shd6706615, 32'shd66f344c, 32'shd66e028a, 32'shd66cd0ce, 
               32'shd66b9f18, 32'shd66a6d69, 32'shd6693bc0, 32'shd6680a1d, 32'shd666d881, 32'shd665a6ec, 32'shd664755c, 32'shd66343d4, 
               32'shd6621251, 32'shd660e0d5, 32'shd65faf60, 32'shd65e7df1, 32'shd65d4c88, 32'shd65c1b26, 32'shd65ae9ca, 32'shd659b874, 
               32'shd6588725, 32'shd65755dd, 32'shd656249b, 32'shd654f35f, 32'shd653c229, 32'shd65290fb, 32'shd6515fd2, 32'shd6502eb0, 
               32'shd64efd94, 32'shd64dcc7f, 32'shd64c9b71, 32'shd64b6a68, 32'shd64a3966, 32'shd649086b, 32'shd647d776, 32'shd646a687, 
               32'shd645759f, 32'shd64444bd, 32'shd64313e2, 32'shd641e30d, 32'shd640b23f, 32'shd63f8177, 32'shd63e50b5, 32'shd63d1ffa, 
               32'shd63bef46, 32'shd63abe97, 32'shd6398df0, 32'shd6385d4e, 32'shd6372cb3, 32'shd635fc1f, 32'shd634cb91, 32'shd6339b09, 
               32'shd6326a88, 32'shd6313a0e, 32'shd6300999, 32'shd62ed92c, 32'shd62da8c4, 32'shd62c7863, 32'shd62b4809, 32'shd62a17b5, 
               32'shd628e767, 32'shd627b720, 32'shd62686e0, 32'shd62556a6, 32'shd6242672, 32'shd622f645, 32'shd621c61e, 32'shd62095fe, 
               32'shd61f65e4, 32'shd61e35d0, 32'shd61d05c3, 32'shd61bd5bd, 32'shd61aa5bd, 32'shd61975c3, 32'shd61845d0, 32'shd61715e3, 
               32'shd615e5fd, 32'shd614b61d, 32'shd6138644, 32'shd6125671, 32'shd61126a5, 32'shd60ff6df, 32'shd60ec720, 32'shd60d9767, 
               32'shd60c67b4, 32'shd60b3808, 32'shd60a0863, 32'shd608d8c4, 32'shd607a92b, 32'shd6067999, 32'shd6054a0d, 32'shd6041a88, 
               32'shd602eb0a, 32'shd601bb91, 32'shd6008c20, 32'shd5ff5cb4, 32'shd5fe2d50, 32'shd5fcfdf1, 32'shd5fbce9a, 32'shd5fa9f48, 
               32'shd5f96ffd, 32'shd5f840b9, 32'shd5f7117b, 32'shd5f5e244, 32'shd5f4b313, 32'shd5f383e8, 32'shd5f254c4, 32'shd5f125a7, 
               32'shd5eff690, 32'shd5eec77f, 32'shd5ed9875, 32'shd5ec6972, 32'shd5eb3a75, 32'shd5ea0b7e, 32'shd5e8dc8e, 32'shd5e7ada4, 
               32'shd5e67ec1, 32'shd5e54fe5, 32'shd5e4210f, 32'shd5e2f23f, 32'shd5e1c376, 32'shd5e094b3, 32'shd5df65f7, 32'shd5de3742, 
               32'shd5dd0892, 32'shd5dbd9ea, 32'shd5daab48, 32'shd5d97cac, 32'shd5d84e17, 32'shd5d71f88, 32'shd5d5f100, 32'shd5d4c27e, 
               32'shd5d39403, 32'shd5d2658f, 32'shd5d13721, 32'shd5d008b9, 32'shd5ceda58, 32'shd5cdabfd, 32'shd5cc7da9, 32'shd5cb4f5c, 
               32'shd5ca2115, 32'shd5c8f2d4, 32'shd5c7c49a, 32'shd5c69666, 32'shd5c56839, 32'shd5c43a13, 32'shd5c30bf3, 32'shd5c1ddd9, 
               32'shd5c0afc6, 32'shd5bf81ba, 32'shd5be53b4, 32'shd5bd25b4, 32'shd5bbf7bc, 32'shd5bac9c9, 32'shd5b99bdd, 32'shd5b86df8, 
               32'shd5b74019, 32'shd5b61241, 32'shd5b4e46f, 32'shd5b3b6a4, 32'shd5b288df, 32'shd5b15b21, 32'shd5b02d69, 32'shd5aeffb8, 
               32'shd5add20d, 32'shd5aca469, 32'shd5ab76cb, 32'shd5aa4934, 32'shd5a91ba4, 32'shd5a7ee1a, 32'shd5a6c096, 32'shd5a59319, 
               32'shd5a465a3, 32'shd5a33833, 32'shd5a20aca, 32'shd5a0dd67, 32'shd59fb00b, 32'shd59e82b5, 32'shd59d5566, 32'shd59c281d, 
               32'shd59afadb, 32'shd599cd9f, 32'shd598a06a, 32'shd597733c, 32'shd5964614, 32'shd59518f2, 32'shd593ebd7, 32'shd592bec3, 
               32'shd59191b5, 32'shd59064ae, 32'shd58f37ad, 32'shd58e0ab3, 32'shd58cddbf, 32'shd58bb0d2, 32'shd58a83eb, 32'shd589570b, 
               32'shd5882a32, 32'shd586fd5f, 32'shd585d093, 32'shd584a3cd, 32'shd583770e, 32'shd5824a55, 32'shd5811da3, 32'shd57ff0f7, 
               32'shd57ec452, 32'shd57d97b4, 32'shd57c6b1c, 32'shd57b3e8a, 32'shd57a1200, 32'shd578e57b, 32'shd577b8fe, 32'shd5768c86, 
               32'shd5756016, 32'shd57433ac, 32'shd5730748, 32'shd571daeb, 32'shd570ae95, 32'shd56f8245, 32'shd56e55fc, 32'shd56d29b9, 
               32'shd56bfd7d, 32'shd56ad148, 32'shd569a519, 32'shd56878f1, 32'shd5674ccf, 32'shd56620b3, 32'shd564f49f, 32'shd563c891, 
               32'shd5629c89, 32'shd5617088, 32'shd560448e, 32'shd55f189a, 32'shd55decad, 32'shd55cc0c6, 32'shd55b94e6, 32'shd55a690c, 
               32'shd5593d3a, 32'shd558116d, 32'shd556e5a7, 32'shd555b9e8, 32'shd5548e30, 32'shd553627d, 32'shd55236d2, 32'shd5510b2d, 
               32'shd54fdf8f, 32'shd54eb3f7, 32'shd54d8866, 32'shd54c5cdb, 32'shd54b3157, 32'shd54a05da, 32'shd548da63, 32'shd547aef3, 
               32'shd5468389, 32'shd5455826, 32'shd5442cca, 32'shd5430174, 32'shd541d625, 32'shd540aadc, 32'shd53f7f9a, 32'shd53e545f, 
               32'shd53d292a, 32'shd53bfdfb, 32'shd53ad2d4, 32'shd539a7b3, 32'shd5387c98, 32'shd5375184, 32'shd5362677, 32'shd534fb70, 
               32'shd533d070, 32'shd532a577, 32'shd5317a84, 32'shd5304f97, 32'shd52f24b2, 32'shd52df9d3, 32'shd52ccefa, 32'shd52ba428, 
               32'shd52a795d, 32'shd5294e98, 32'shd52823da, 32'shd526f923, 32'shd525ce72, 32'shd524a3c7, 32'shd5237924, 32'shd5224e87, 
               32'shd52123f0, 32'shd51ff960, 32'shd51eced7, 32'shd51da455, 32'shd51c79d9, 32'shd51b4f63, 32'shd51a24f5, 32'shd518fa8c, 
               32'shd517d02b, 32'shd516a5d0, 32'shd5157b7c, 32'shd514512e, 32'shd51326e7, 32'shd511fca7, 32'shd510d26d, 32'shd50fa83a, 
               32'shd50e7e0d, 32'shd50d53e7, 32'shd50c29c8, 32'shd50affaf, 32'shd509d59d, 32'shd508ab91, 32'shd507818d, 32'shd506578e, 
               32'shd5052d97, 32'shd50403a6, 32'shd502d9bc, 32'shd501afd8, 32'shd50085fb, 32'shd4ff5c24, 32'shd4fe3255, 32'shd4fd088c, 
               32'shd4fbdec9, 32'shd4fab50d, 32'shd4f98b58, 32'shd4f861a9, 32'shd4f73801, 32'shd4f60e60, 32'shd4f4e4c5, 32'shd4f3bb31, 
               32'shd4f291a4, 32'shd4f1681d, 32'shd4f03e9d, 32'shd4ef1523, 32'shd4edebb0, 32'shd4ecc244, 32'shd4eb98de, 32'shd4ea6f80, 
               32'shd4e94627, 32'shd4e81cd6, 32'shd4e6f38b, 32'shd4e5ca46, 32'shd4e4a108, 32'shd4e377d1, 32'shd4e24ea1, 32'shd4e12577, 
               32'shd4dffc54, 32'shd4ded338, 32'shd4ddaa22, 32'shd4dc8113, 32'shd4db580a, 32'shd4da2f08, 32'shd4d9060d, 32'shd4d7dd18, 
               32'shd4d6b42b, 32'shd4d58b43, 32'shd4d46263, 32'shd4d33989, 32'shd4d210b5, 32'shd4d0e7e9, 32'shd4cfbf23, 32'shd4ce9664, 
               32'shd4cd6dab, 32'shd4cc44f9, 32'shd4cb1c4e, 32'shd4c9f3a9, 32'shd4c8cb0b, 32'shd4c7a274, 32'shd4c679e3, 32'shd4c55159, 
               32'shd4c428d6, 32'shd4c30059, 32'shd4c1d7e3, 32'shd4c0af74, 32'shd4bf870b, 32'shd4be5ea9, 32'shd4bd364e, 32'shd4bc0df9, 
               32'shd4bae5ab, 32'shd4b9bd64, 32'shd4b89523, 32'shd4b76ce9, 32'shd4b644b6, 32'shd4b51c8a, 32'shd4b3f464, 32'shd4b2cc44, 
               32'shd4b1a42c, 32'shd4b07c1a, 32'shd4af540f, 32'shd4ae2c0a, 32'shd4ad040c, 32'shd4abdc15, 32'shd4aab425, 32'shd4a98c3b, 
               32'shd4a86458, 32'shd4a73c7b, 32'shd4a614a6, 32'shd4a4ecd7, 32'shd4a3c50e, 32'shd4a29d4c, 32'shd4a17591, 32'shd4a04ddd, 
               32'shd49f2630, 32'shd49dfe89, 32'shd49cd6e8, 32'shd49baf4f, 32'shd49a87bc, 32'shd4996030, 32'shd49838aa, 32'shd497112b, 
               32'shd495e9b3, 32'shd494c242, 32'shd4939ad7, 32'shd4927373, 32'shd4914c16, 32'shd49024bf, 32'shd48efd6f, 32'shd48dd626, 
               32'shd48caee4, 32'shd48b87a8, 32'shd48a6073, 32'shd4893944, 32'shd488121d, 32'shd486eafc, 32'shd485c3e1, 32'shd4849cce, 
               32'shd48375c1, 32'shd4824ebb, 32'shd48127bb, 32'shd48000c2, 32'shd47ed9d0, 32'shd47db2e5, 32'shd47c8c00, 32'shd47b6523, 
               32'shd47a3e4b, 32'shd479177b, 32'shd477f0b1, 32'shd476c9ee, 32'shd475a332, 32'shd4747c7c, 32'shd47355cd, 32'shd4722f25, 
               32'shd4710883, 32'shd46fe1e8, 32'shd46ebb54, 32'shd46d94c7, 32'shd46c6e40, 32'shd46b47c0, 32'shd46a2147, 32'shd468fad5, 
               32'shd467d469, 32'shd466ae04, 32'shd46587a6, 32'shd464614e, 32'shd4633afd, 32'shd46214b3, 32'shd460ee70, 32'shd45fc833, 
               32'shd45ea1fd, 32'shd45d7bce, 32'shd45c55a5, 32'shd45b2f84, 32'shd45a0969, 32'shd458e354, 32'shd457bd47, 32'shd4569740, 
               32'shd4557140, 32'shd4544b46, 32'shd4532554, 32'shd451ff68, 32'shd450d983, 32'shd44fb3a4, 32'shd44e8dcd, 32'shd44d67fc, 
               32'shd44c4232, 32'shd44b1c6e, 32'shd449f6b1, 32'shd448d0fb, 32'shd447ab4c, 32'shd44685a4, 32'shd4456002, 32'shd4443a67, 
               32'shd44314d3, 32'shd441ef45, 32'shd440c9be, 32'shd43fa43e, 32'shd43e7ec5, 32'shd43d5952, 32'shd43c33e7, 32'shd43b0e81, 
               32'shd439e923, 32'shd438c3cc, 32'shd4379e7b, 32'shd4367931, 32'shd43553ee, 32'shd4342eb1, 32'shd433097b, 32'shd431e44c, 
               32'shd430bf24, 32'shd42f9a02, 32'shd42e74e8, 32'shd42d4fd4, 32'shd42c2ac6, 32'shd42b05c0, 32'shd429e0c0, 32'shd428bbc7, 
               32'shd42796d5, 32'shd42671ea, 32'shd4254d05, 32'shd4242827, 32'shd4230350, 32'shd421de7f, 32'shd420b9b6, 32'shd41f94f3, 
               32'shd41e7037, 32'shd41d4b81, 32'shd41c26d3, 32'shd41b022b, 32'shd419dd8a, 32'shd418b8f0, 32'shd417945c, 32'shd4166fd0, 
               32'shd4154b4a, 32'shd41426cb, 32'shd4130252, 32'shd411dde1, 32'shd410b976, 32'shd40f9512, 32'shd40e70b4, 32'shd40d4c5e, 
               32'shd40c280e, 32'shd40b03c5, 32'shd409df83, 32'shd408bb48, 32'shd4079713, 32'shd40672e5, 32'shd4054ebe, 32'shd4042a9e, 
               32'shd4030684, 32'shd401e271, 32'shd400be66, 32'shd3ff9a60, 32'shd3fe7662, 32'shd3fd526a, 32'shd3fc2e7a, 32'shd3fb0a90, 
               32'shd3f9e6ad, 32'shd3f8c2d0, 32'shd3f79efa, 32'shd3f67b2c, 32'shd3f55764, 32'shd3f433a2, 32'shd3f30fe8, 32'shd3f1ec34, 
               32'shd3f0c887, 32'shd3efa4e1, 32'shd3ee8142, 32'shd3ed5da9, 32'shd3ec3a18, 32'shd3eb168d, 32'shd3e9f309, 32'shd3e8cf8b, 
               32'shd3e7ac15, 32'shd3e688a5, 32'shd3e5653c, 32'shd3e441da, 32'shd3e31e7f, 32'shd3e1fb2a, 32'shd3e0d7dd, 32'shd3dfb496, 
               32'shd3de9156, 32'shd3dd6e1c, 32'shd3dc4aea, 32'shd3db27be, 32'shd3da049a, 32'shd3d8e17b, 32'shd3d7be64, 32'shd3d69b54, 
               32'shd3d5784a, 32'shd3d45547, 32'shd3d3324b, 32'shd3d20f56, 32'shd3d0ec68, 32'shd3cfc980, 32'shd3cea69f, 32'shd3cd83c6, 
               32'shd3cc60f2, 32'shd3cb3e26, 32'shd3ca1b61, 32'shd3c8f8a2, 32'shd3c7d5ea, 32'shd3c6b339, 32'shd3c5908f, 32'shd3c46dec, 
               32'shd3c34b4f, 32'shd3c228b9, 32'shd3c1062a, 32'shd3bfe3a2, 32'shd3bec121, 32'shd3bd9ea7, 32'shd3bc7c33, 32'shd3bb59c6, 
               32'shd3ba3760, 32'shd3b91501, 32'shd3b7f2a9, 32'shd3b6d057, 32'shd3b5ae0d, 32'shd3b48bc9, 32'shd3b3698c, 32'shd3b24756, 
               32'shd3b12526, 32'shd3b002fe, 32'shd3aee0dc, 32'shd3adbec1, 32'shd3ac9cad, 32'shd3ab7aa0, 32'shd3aa589a, 32'shd3a9369a, 
               32'shd3a814a2, 32'shd3a6f2b0, 32'shd3a5d0c5, 32'shd3a4aee1, 32'shd3a38d03, 32'shd3a26b2d, 32'shd3a1495d, 32'shd3a02795, 
               32'shd39f05d3, 32'shd39de418, 32'shd39cc263, 32'shd39ba0b6, 32'shd39a7f0f, 32'shd3995d70, 32'shd3983bd7, 32'shd3971a45, 
               32'shd395f8ba, 32'shd394d735, 32'shd393b5b8, 32'shd3929441, 32'shd39172d2, 32'shd3905169, 32'shd38f3007, 32'shd38e0eac, 
               32'shd38ced57, 32'shd38bcc0a, 32'shd38aaac3, 32'shd3898983, 32'shd388684a, 32'shd3874718, 32'shd38625ed, 32'shd38504c9, 
               32'shd383e3ab, 32'shd382c295, 32'shd381a185, 32'shd380807c, 32'shd37f5f7a, 32'shd37e3e7f, 32'shd37d1d8a, 32'shd37bfc9d, 
               32'shd37adbb6, 32'shd379bad7, 32'shd37899fe, 32'shd377792c, 32'shd3765861, 32'shd375379d, 32'shd37416df, 32'shd372f629, 
               32'shd371d579, 32'shd370b4d0, 32'shd36f942e, 32'shd36e7393, 32'shd36d52ff, 32'shd36c3272, 32'shd36b11eb, 32'shd369f16c, 
               32'shd368d0f3, 32'shd367b082, 32'shd3669017, 32'shd3656fb3, 32'shd3644f55, 32'shd3632eff, 32'shd3620eb0, 32'shd360ee67, 
               32'shd35fce26, 32'shd35eadeb, 32'shd35d8db7, 32'shd35c6d8a, 32'shd35b4d64, 32'shd35a2d45, 32'shd3590d2c, 32'shd357ed1b, 
               32'shd356cd11, 32'shd355ad0d, 32'shd3548d10, 32'shd3536d1a, 32'shd3524d2b, 32'shd3512d43, 32'shd3500d62, 32'shd34eed88, 
               32'shd34dcdb4, 32'shd34cade8, 32'shd34b8e22, 32'shd34a6e63, 32'shd3494eab, 32'shd3482efa, 32'shd3470f50, 32'shd345efad, 
               32'shd344d011, 32'shd343b07b, 32'shd34290ed, 32'shd3417165, 32'shd34051e5, 32'shd33f326b, 32'shd33e12f8, 32'shd33cf38c, 
               32'shd33bd427, 32'shd33ab4c9, 32'shd3399572, 32'shd3387621, 32'shd33756d8, 32'shd3363795, 32'shd335185a, 32'shd333f925, 
               32'shd332d9f7, 32'shd331bad0, 32'shd3309bb0, 32'shd32f7c97, 32'shd32e5d85, 32'shd32d3e7a, 32'shd32c1f75, 32'shd32b0078, 
               32'shd329e181, 32'shd328c292, 32'shd327a3a9, 32'shd32684c7, 32'shd32565ec, 32'shd3244718, 32'shd323284b, 32'shd3220985, 
               32'shd320eac6, 32'shd31fcc0e, 32'shd31ead5c, 32'shd31d8eb2, 32'shd31c700f, 32'shd31b5172, 32'shd31a32dc, 32'shd319144e, 
               32'shd317f5c6, 32'shd316d745, 32'shd315b8cb, 32'shd3149a58, 32'shd3137bec, 32'shd3125d86, 32'shd3113f28, 32'shd31020d1, 
               32'shd30f0280, 32'shd30de437, 32'shd30cc5f4, 32'shd30ba7b9, 32'shd30a8984, 32'shd3096b56, 32'shd3084d30, 32'shd3072f10, 
               32'shd30610f7, 32'shd304f2e5, 32'shd303d4da, 32'shd302b6d6, 32'shd30198d8, 32'shd3007ae2, 32'shd2ff5cf3, 32'shd2fe3f0b, 
               32'shd2fd2129, 32'shd2fc034f, 32'shd2fae57b, 32'shd2f9c7ae, 32'shd2f8a9e9, 32'shd2f78c2a, 32'shd2f66e72, 32'shd2f550c2, 
               32'shd2f43318, 32'shd2f31575, 32'shd2f1f7d9, 32'shd2f0da44, 32'shd2efbcb6, 32'shd2ee9f2e, 32'shd2ed81ae, 32'shd2ec6435, 
               32'shd2eb46c3, 32'shd2ea2957, 32'shd2e90bf3, 32'shd2e7ee96, 32'shd2e6d13f, 32'shd2e5b3f0, 32'shd2e496a7, 32'shd2e37965, 
               32'shd2e25c2b, 32'shd2e13ef7, 32'shd2e021ca, 32'shd2df04a5, 32'shd2dde786, 32'shd2dcca6e, 32'shd2dbad5d, 32'shd2da9053, 
               32'shd2d97350, 32'shd2d85654, 32'shd2d7395f, 32'shd2d61c71, 32'shd2d4ff8a, 32'shd2d3e2aa, 32'shd2d2c5d0, 32'shd2d1a8fe, 
               32'shd2d08c33, 32'shd2cf6f6f, 32'shd2ce52b1, 32'shd2cd35fb, 32'shd2cc194c, 32'shd2cafca3, 32'shd2c9e002, 32'shd2c8c367, 
               32'shd2c7a6d4, 32'shd2c68a47, 32'shd2c56dc2, 32'shd2c45143, 32'shd2c334cc, 32'shd2c2185b, 32'shd2c0fbf1, 32'shd2bfdf8f, 
               32'shd2bec333, 32'shd2bda6de, 32'shd2bc8a91, 32'shd2bb6e4a, 32'shd2ba520a, 32'shd2b935d1, 32'shd2b8199f, 32'shd2b6fd75, 
               32'shd2b5e151, 32'shd2b4c534, 32'shd2b3a91e, 32'shd2b28d0f, 32'shd2b17107, 32'shd2b05506, 32'shd2af390d, 32'shd2ae1d1a, 
               32'shd2ad012e, 32'shd2abe549, 32'shd2aac96b, 32'shd2a9ad94, 32'shd2a891c4, 32'shd2a775fb, 32'shd2a65a39, 32'shd2a53e7e, 
               32'shd2a422ca, 32'shd2a3071d, 32'shd2a1eb77, 32'shd2a0cfd8, 32'shd29fb440, 32'shd29e98af, 32'shd29d7d25, 32'shd29c61a2, 
               32'shd29b4626, 32'shd29a2ab1, 32'shd2990f43, 32'shd297f3dc, 32'shd296d87c, 32'shd295bd23, 32'shd294a1d0, 32'shd2938685, 
               32'shd2926b41, 32'shd2915004, 32'shd29034ce, 32'shd28f199f, 32'shd28dfe77, 32'shd28ce357, 32'shd28bc83d, 32'shd28aad2a, 
               32'shd289921e, 32'shd2887719, 32'shd2875c1b, 32'shd2864124, 32'shd2852634, 32'shd2840b4b, 32'shd282f069, 32'shd281d58e, 
               32'shd280babb, 32'shd27f9fee, 32'shd27e8528, 32'shd27d6a69, 32'shd27c4fb1, 32'shd27b3501, 32'shd27a1a57, 32'shd278ffb4, 
               32'shd277e518, 32'shd276ca84, 32'shd275aff6, 32'shd2749570, 32'shd2737af0, 32'shd2726077, 32'shd2714606, 32'shd2702b9b, 
               32'shd26f1138, 32'shd26df6db, 32'shd26cdc86, 32'shd26bc237, 32'shd26aa7f0, 32'shd2698db0, 32'shd2687376, 32'shd2675944, 
               32'shd2663f19, 32'shd26524f5, 32'shd2640ad7, 32'shd262f0c1, 32'shd261d6b2, 32'shd260bcaa, 32'shd25fa2a9, 32'shd25e88af, 
               32'shd25d6ebc, 32'shd25c54d0, 32'shd25b3aeb, 32'shd25a210d, 32'shd2590736, 32'shd257ed67, 32'shd256d39e, 32'shd255b9dc, 
               32'shd254a021, 32'shd253866e, 32'shd2526cc1, 32'shd251531c, 32'shd250397d, 32'shd24f1fe6, 32'shd24e0655, 32'shd24ceccc, 
               32'shd24bd34a, 32'shd24ab9ce, 32'shd249a05a, 32'shd24886ed, 32'shd2476d87, 32'shd2465428, 32'shd2453ad0, 32'shd244217f, 
               32'shd2430835, 32'shd241eef2, 32'shd240d5b6, 32'shd23fbc82, 32'shd23ea354, 32'shd23d8a2d, 32'shd23c710e, 32'shd23b57f5, 
               32'shd23a3ee4, 32'shd23925d9, 32'shd2380cd6, 32'shd236f3da, 32'shd235dae4, 32'shd234c1f6, 32'shd233a90f, 32'shd232902f, 
               32'shd2317756, 32'shd2305e84, 32'shd22f45b9, 32'shd22e2cf6, 32'shd22d1439, 32'shd22bfb83, 32'shd22ae2d5, 32'shd229ca2d, 
               32'shd228b18d, 32'shd22798f3, 32'shd2268061, 32'shd22567d6, 32'shd2244f52, 32'shd22336d5, 32'shd2221e5f, 32'shd22105f0, 
               32'shd21fed88, 32'shd21ed527, 32'shd21dbccd, 32'shd21ca47b, 32'shd21b8c2f, 32'shd21a73eb, 32'shd2195bad, 32'shd2184377, 
               32'shd2172b48, 32'shd216131f, 32'shd214fafe, 32'shd213e2e4, 32'shd212cad1, 32'shd211b2c5, 32'shd2109ac1, 32'shd20f82c3, 
               32'shd20e6acc, 32'shd20d52dd, 32'shd20c3af4, 32'shd20b2313, 32'shd20a0b39, 32'shd208f366, 32'shd207db9a, 32'shd206c3d5, 
               32'shd205ac17, 32'shd2049460, 32'shd2037cb0, 32'shd2026508, 32'shd2014d66, 32'shd20035cc, 32'shd1ff1e38, 32'shd1fe06ac, 
               32'shd1fcef27, 32'shd1fbd7a9, 32'shd1fac032, 32'shd1f9a8c2, 32'shd1f89159, 32'shd1f779f8, 32'shd1f6629d, 32'shd1f54b49, 
               32'shd1f433fd, 32'shd1f31cb8, 32'shd1f2057a, 32'shd1f0ee43, 32'shd1efd713, 32'shd1eebfea, 32'shd1eda8c8, 32'shd1ec91ad, 
               32'shd1eb7a9a, 32'shd1ea638d, 32'shd1e94c88, 32'shd1e8358a, 32'shd1e71e93, 32'shd1e607a3, 32'shd1e4f0ba, 32'shd1e3d9d8, 
               32'shd1e2c2fd, 32'shd1e1ac2a, 32'shd1e0955d, 32'shd1df7e98, 32'shd1de67da, 32'shd1dd5123, 32'shd1dc3a73, 32'shd1db23ca, 
               32'shd1da0d28, 32'shd1d8f68d, 32'shd1d7dffa, 32'shd1d6c96d, 32'shd1d5b2e8, 32'shd1d49c6a, 32'shd1d385f3, 32'shd1d26f83, 
               32'shd1d1591a, 32'shd1d042b8, 32'shd1cf2c5e, 32'shd1ce160a, 32'shd1ccffbe, 32'shd1cbe979, 32'shd1cad33b, 32'shd1c9bd04, 
               32'shd1c8a6d4, 32'shd1c790ab, 32'shd1c67a8a, 32'shd1c5646f, 32'shd1c44e5c, 32'shd1c33850, 32'shd1c2224b, 32'shd1c10c4d, 
               32'shd1bff656, 32'shd1bee066, 32'shd1bdca7e, 32'shd1bcb49c, 32'shd1bb9ec2, 32'shd1ba88ef, 32'shd1b97323, 32'shd1b85d5e, 
               32'shd1b747a0, 32'shd1b631ea, 32'shd1b51c3a, 32'shd1b40692, 32'shd1b2f0f1, 32'shd1b1db57, 32'shd1b0c5c4, 32'shd1afb038, 
               32'shd1ae9ab4, 32'shd1ad8536, 32'shd1ac6fc0, 32'shd1ab5a51, 32'shd1aa44e9, 32'shd1a92f88, 32'shd1a81a2e, 32'shd1a704dc, 
               32'shd1a5ef90, 32'shd1a4da4c, 32'shd1a3c50f, 32'shd1a2afd9, 32'shd1a19aaa, 32'shd1a08582, 32'shd19f7062, 32'shd19e5b48, 
               32'shd19d4636, 32'shd19c312b, 32'shd19b1c27, 32'shd19a072a, 32'shd198f235, 32'shd197dd46, 32'shd196c85f, 32'shd195b37f, 
               32'shd1949ea6, 32'shd19389d4, 32'shd1927509, 32'shd1916046, 32'shd1904b89, 32'shd18f36d4, 32'shd18e2226, 32'shd18d0d7f, 
               32'shd18bf8e0, 32'shd18ae447, 32'shd189cfb6, 32'shd188bb2b, 32'shd187a6a8, 32'shd186922d, 32'shd1857db8, 32'shd184694a, 
               32'shd18354e4, 32'shd1824085, 32'shd1812c2d, 32'shd18017dc, 32'shd17f0392, 32'shd17def50, 32'shd17cdb14, 32'shd17bc6e0, 
               32'shd17ab2b3, 32'shd1799e8d, 32'shd1788a6f, 32'shd1777657, 32'shd1766247, 32'shd1754e3e, 32'shd1743a3c, 32'shd1732641, 
               32'shd172124d, 32'shd170fe61, 32'shd16fea7c, 32'shd16ed69e, 32'shd16dc2c7, 32'shd16caef7, 32'shd16b9b2f, 32'shd16a876d, 
               32'shd16973b3, 32'shd1686000, 32'shd1674c54, 32'shd16638b0, 32'shd1652512, 32'shd164117c, 32'shd162fded, 32'shd161ea65, 
               32'shd160d6e5, 32'shd15fc36b, 32'shd15eaff9, 32'shd15d9c8e, 32'shd15c892a, 32'shd15b75cd, 32'shd15a6278, 32'shd1594f29, 
               32'shd1583be2, 32'shd15728a2, 32'shd156156a, 32'shd1550238, 32'shd153ef0e, 32'shd152dbeb, 32'shd151c8cf, 32'shd150b5ba, 
               32'shd14fa2ad, 32'shd14e8fa6, 32'shd14d7ca7, 32'shd14c69af, 32'shd14b56be, 32'shd14a43d5, 32'shd14930f3, 32'shd1481e17, 
               32'shd1470b44, 32'shd145f877, 32'shd144e5b1, 32'shd143d2f3, 32'shd142c03c, 32'shd141ad8c, 32'shd1409ae3, 32'shd13f8842, 
               32'shd13e75a8, 32'shd13d6315, 32'shd13c5089, 32'shd13b3e04, 32'shd13a2b87, 32'shd1391911, 32'shd13806a2, 32'shd136f43a, 
               32'shd135e1d9, 32'shd134cf80, 32'shd133bd2e, 32'shd132aae3, 32'shd131989f, 32'shd1308663, 32'shd12f742d, 32'shd12e61ff, 
               32'shd12d4fd9, 32'shd12c3db9, 32'shd12b2ba1, 32'shd12a198f, 32'shd1290786, 32'shd127f583, 32'shd126e387, 32'shd125d193, 
               32'shd124bfa6, 32'shd123adc0, 32'shd1229be2, 32'shd1218a0a, 32'shd120783a, 32'shd11f6671, 32'shd11e54b0, 32'shd11d42f5, 
               32'shd11c3142, 32'shd11b1f96, 32'shd11a0df1, 32'shd118fc54, 32'shd117eabd, 32'shd116d92e, 32'shd115c7a7, 32'shd114b626, 
               32'shd113a4ad, 32'shd112933b, 32'shd11181d0, 32'shd110706c, 32'shd10f5f10, 32'shd10e4dbb, 32'shd10d3c6d, 32'shd10c2b26, 
               32'shd10b19e7, 32'shd10a08ae, 32'shd108f77d, 32'shd107e654, 32'shd106d531, 32'shd105c416, 32'shd104b302, 32'shd103a1f5, 
               32'shd10290f0, 32'shd1017ff2, 32'shd1006efb, 32'shd0ff5e0b, 32'shd0fe4d22, 32'shd0fd3c41, 32'shd0fc2b67, 32'shd0fb1a94, 
               32'shd0fa09c9, 32'shd0f8f905, 32'shd0f7e848, 32'shd0f6d792, 32'shd0f5c6e3, 32'shd0f4b63c, 32'shd0f3a59c, 32'shd0f29503, 
               32'shd0f18472, 32'shd0f073e8, 32'shd0ef6365, 32'shd0ee52e9, 32'shd0ed4275, 32'shd0ec3208, 32'shd0eb21a2, 32'shd0ea1143, 
               32'shd0e900ec, 32'shd0e7f09b, 32'shd0e6e053, 32'shd0e5d011, 32'shd0e4bfd7, 32'shd0e3afa4, 32'shd0e29f78, 32'shd0e18f53, 
               32'shd0e07f36, 32'shd0df6f20, 32'shd0de5f11, 32'shd0dd4f0a, 32'shd0dc3f0a, 32'shd0db2f11, 32'shd0da1f1f, 32'shd0d90f35, 
               32'shd0d7ff51, 32'shd0d6ef76, 32'shd0d5dfa1, 32'shd0d4cfd4, 32'shd0d3c00e, 32'shd0d2b04f, 32'shd0d1a097, 32'shd0d090e7, 
               32'shd0cf813e, 32'shd0ce719d, 32'shd0cd6202, 32'shd0cc526f, 32'shd0cb42e3, 32'shd0ca335f, 32'shd0c923e1, 32'shd0c8146c, 
               32'shd0c704fd, 32'shd0c5f595, 32'shd0c4e635, 32'shd0c3d6dc, 32'shd0c2c78b, 32'shd0c1b841, 32'shd0c0a8fe, 32'shd0bf99c2, 
               32'shd0be8a8d, 32'shd0bd7b60, 32'shd0bc6c3a, 32'shd0bb5d1c, 32'shd0ba4e05, 32'shd0b93ef5, 32'shd0b82fec, 32'shd0b720eb, 
               32'shd0b611f1, 32'shd0b502fe, 32'shd0b3f412, 32'shd0b2e52e, 32'shd0b1d651, 32'shd0b0c77b, 32'shd0afb8ad, 32'shd0aea9e6, 
               32'shd0ad9b26, 32'shd0ac8c6e, 32'shd0ab7dbd, 32'shd0aa6f13, 32'shd0a96070, 32'shd0a851d5, 32'shd0a74341, 32'shd0a634b4, 
               32'shd0a5262f, 32'shd0a417b1, 32'shd0a3093a, 32'shd0a1facb, 32'shd0a0ec63, 32'shd09fde02, 32'shd09ecfa8, 32'shd09dc156, 
               32'shd09cb30b, 32'shd09ba4c8, 32'shd09a968b, 32'shd0998856, 32'shd0987a29, 32'shd0976c02, 32'shd0965de3, 32'shd0954fcc, 
               32'shd09441bb, 32'shd09333b2, 32'shd09225b0, 32'shd09117b6, 32'shd09009c3, 32'shd08efbd7, 32'shd08dedf2, 32'shd08ce015, 
               32'shd08bd23f, 32'shd08ac470, 32'shd089b6a9, 32'shd088a8e9, 32'shd0879b31, 32'shd0868d7f, 32'shd0857fd5, 32'shd0847233, 
               32'shd0836497, 32'shd0825703, 32'shd0814977, 32'shd0803bf1, 32'shd07f2e73, 32'shd07e20fc, 32'shd07d138d, 32'shd07c0625, 
               32'shd07af8c4, 32'shd079eb6b, 32'shd078de19, 32'shd077d0ce, 32'shd076c38b, 32'shd075b64f, 32'shd074a91a, 32'shd0739bec, 
               32'shd0728ec6, 32'shd07181a7, 32'shd0707490, 32'shd06f6780, 32'shd06e5a77, 32'shd06d4d76, 32'shd06c407c, 32'shd06b3389, 
               32'shd06a269d, 32'shd06919b9, 32'shd0680cdd, 32'shd0670007, 32'shd065f339, 32'shd064e673, 32'shd063d9b3, 32'shd062ccfb, 
               32'shd061c04a, 32'shd060b3a1, 32'shd05fa6ff, 32'shd05e9a64, 32'shd05d8dd1, 32'shd05c8145, 32'shd05b74c0, 32'shd05a6843, 
               32'shd0595bcd, 32'shd0584f5f, 32'shd05742f7, 32'shd0563698, 32'shd0552a3f, 32'shd0541dee, 32'shd05311a4, 32'shd0520562, 
               32'shd050f926, 32'shd04fecf3, 32'shd04ee0c6, 32'shd04dd4a1, 32'shd04cc884, 32'shd04bbc6d, 32'shd04ab05e, 32'shd049a457, 
               32'shd0489856, 32'shd0478c5d, 32'shd046806c, 32'shd0457482, 32'shd044689f, 32'shd0435cc3, 32'shd04250ef, 32'shd0414522, 
               32'shd040395d, 32'shd03f2d9f, 32'shd03e21e8, 32'shd03d1639, 32'shd03c0a91, 32'shd03afef1, 32'shd039f357, 32'shd038e7c5, 
               32'shd037dc3b, 32'shd036d0b8, 32'shd035c53c, 32'shd034b9c8, 32'shd033ae5b, 32'shd032a2f5, 32'shd0319797, 32'shd0308c40, 
               32'shd02f80f1, 32'shd02e75a8, 32'shd02d6a68, 32'shd02c5f2e, 32'shd02b53fc, 32'shd02a48d2, 32'shd0293dae, 32'shd0283293, 
               32'shd027277e, 32'shd0261c71, 32'shd025116b, 32'shd024066d, 32'shd022fb76, 32'shd021f086, 32'shd020e59e, 32'shd01fdabd, 
               32'shd01ecfe4, 32'shd01dc512, 32'shd01cba47, 32'shd01baf84, 32'shd01aa4c8, 32'shd0199a13, 32'shd0188f66, 32'shd01784c1, 
               32'shd0167a22, 32'shd0156f8b, 32'shd01464fc, 32'shd0135a73, 32'shd0124ff3, 32'shd0114579, 32'shd0103b07, 32'shd00f309d, 
               32'shd00e2639, 32'shd00d1bdd, 32'shd00c1189, 32'shd00b073c, 32'shd009fcf6, 32'shd008f2b8, 32'shd007e881, 32'shd006de52, 
               32'shd005d42a, 32'shd004ca09, 32'shd003bff0, 32'shd002b5de, 32'shd001abd3, 32'shd000a1d0, 32'shcfff97d5, 32'shcffe8de0, 
               32'shcffd83f4, 32'shcffc7a0e, 32'shcffb7030, 32'shcffa6659, 32'shcff95c8a, 32'shcff852c2, 32'shcff74902, 32'shcff63f49, 
               32'shcff53597, 32'shcff42bed, 32'shcff3224a, 32'shcff218af, 32'shcff10f1b, 32'shcff0058e, 32'shcfeefc09, 32'shcfedf28b, 
               32'shcfece915, 32'shcfebdfa6, 32'shcfead63f, 32'shcfe9ccdf, 32'shcfe8c386, 32'shcfe7ba35, 32'shcfe6b0eb, 32'shcfe5a7a8, 
               32'shcfe49e6d, 32'shcfe3953a, 32'shcfe28c0e, 32'shcfe182e9, 32'shcfe079cc, 32'shcfdf70b6, 32'shcfde67a7, 32'shcfdd5ea0, 
               32'shcfdc55a1, 32'shcfdb4ca8, 32'shcfda43b8, 32'shcfd93ace, 32'shcfd831ec, 32'shcfd72912, 32'shcfd6203f, 32'shcfd51773, 
               32'shcfd40eaf, 32'shcfd305f2, 32'shcfd1fd3d, 32'shcfd0f48f, 32'shcfcfebe8, 32'shcfcee349, 32'shcfcddab2, 32'shcfccd221, 
               32'shcfcbc999, 32'shcfcac117, 32'shcfc9b89d, 32'shcfc8b02b, 32'shcfc7a7c0, 32'shcfc69f5c, 32'shcfc59700, 32'shcfc48eab, 
               32'shcfc3865e, 32'shcfc27e18, 32'shcfc175da, 32'shcfc06da3, 32'shcfbf6573, 32'shcfbe5d4b, 32'shcfbd552b, 32'shcfbc4d11, 
               32'shcfbb4500, 32'shcfba3cf5, 32'shcfb934f2, 32'shcfb82cf7, 32'shcfb72503, 32'shcfb61d16, 32'shcfb51531, 32'shcfb40d54, 
               32'shcfb3057d, 32'shcfb1fdaf, 32'shcfb0f5e7, 32'shcfafee28, 32'shcfaee66f, 32'shcfaddebe, 32'shcfacd715, 32'shcfabcf73, 
               32'shcfaac7d8, 32'shcfa9c045, 32'shcfa8b8b9, 32'shcfa7b135, 32'shcfa6a9b8, 32'shcfa5a243, 32'shcfa49ad5, 32'shcfa3936f, 
               32'shcfa28c10, 32'shcfa184b8, 32'shcfa07d68, 32'shcf9f7620, 32'shcf9e6edf, 32'shcf9d67a5, 32'shcf9c6073, 32'shcf9b5948, 
               32'shcf9a5225, 32'shcf994b09, 32'shcf9843f5, 32'shcf973ce8, 32'shcf9635e2, 32'shcf952ee4, 32'shcf9427ee, 32'shcf9320ff, 
               32'shcf921a17, 32'shcf911337, 32'shcf900c5f, 32'shcf8f058e, 32'shcf8dfec4, 32'shcf8cf802, 32'shcf8bf147, 32'shcf8aea94, 
               32'shcf89e3e8, 32'shcf88dd44, 32'shcf87d6a7, 32'shcf86d012, 32'shcf85c984, 32'shcf84c2fd, 32'shcf83bc7e, 32'shcf82b607, 
               32'shcf81af97, 32'shcf80a92e, 32'shcf7fa2cd, 32'shcf7e9c74, 32'shcf7d9622, 32'shcf7c8fd7, 32'shcf7b8994, 32'shcf7a8359, 
               32'shcf797d24, 32'shcf7876f8, 32'shcf7770d3, 32'shcf766ab5, 32'shcf75649f, 32'shcf745e90, 32'shcf735889, 32'shcf725289, 
               32'shcf714c91, 32'shcf7046a0, 32'shcf6f40b7, 32'shcf6e3ad5, 32'shcf6d34fb, 32'shcf6c2f28, 32'shcf6b295d, 32'shcf6a2399, 
               32'shcf691ddd, 32'shcf681828, 32'shcf67127a, 32'shcf660cd5, 32'shcf650736, 32'shcf64019f, 32'shcf62fc10, 32'shcf61f688, 
               32'shcf60f108, 32'shcf5feb8f, 32'shcf5ee61e, 32'shcf5de0b4, 32'shcf5cdb51, 32'shcf5bd5f7, 32'shcf5ad0a3, 32'shcf59cb57, 
               32'shcf58c613, 32'shcf57c0d6, 32'shcf56bba1, 32'shcf55b673, 32'shcf54b14d, 32'shcf53ac2e, 32'shcf52a716, 32'shcf51a207, 
               32'shcf509cfe, 32'shcf4f97fe, 32'shcf4e9304, 32'shcf4d8e12, 32'shcf4c8928, 32'shcf4b8445, 32'shcf4a7f6a, 32'shcf497a96, 
               32'shcf4875ca, 32'shcf477105, 32'shcf466c48, 32'shcf456793, 32'shcf4462e4, 32'shcf435e3e, 32'shcf42599f, 32'shcf415507, 
               32'shcf405077, 32'shcf3f4bee, 32'shcf3e476d, 32'shcf3d42f4, 32'shcf3c3e82, 32'shcf3b3a17, 32'shcf3a35b4, 32'shcf393159, 
               32'shcf382d05, 32'shcf3728b8, 32'shcf362473, 32'shcf352036, 32'shcf341c00, 32'shcf3317d2, 32'shcf3213ab, 32'shcf310f8c, 
               32'shcf300b74, 32'shcf2f0764, 32'shcf2e035b, 32'shcf2cff5a, 32'shcf2bfb60, 32'shcf2af76e, 32'shcf29f383, 32'shcf28efa0, 
               32'shcf27ebc5, 32'shcf26e7f1, 32'shcf25e424, 32'shcf24e05f, 32'shcf23dca2, 32'shcf22d8ec, 32'shcf21d53e, 32'shcf20d197, 
               32'shcf1fcdf8, 32'shcf1eca60, 32'shcf1dc6d0, 32'shcf1cc347, 32'shcf1bbfc6, 32'shcf1abc4d, 32'shcf19b8db, 32'shcf18b570, 
               32'shcf17b20d, 32'shcf16aeb2, 32'shcf15ab5e, 32'shcf14a812, 32'shcf13a4cd, 32'shcf12a190, 32'shcf119e5a, 32'shcf109b2c, 
               32'shcf0f9805, 32'shcf0e94e6, 32'shcf0d91cf, 32'shcf0c8ebf, 32'shcf0b8bb7, 32'shcf0a88b6, 32'shcf0985bc, 32'shcf0882cb, 
               32'shcf077fe1, 32'shcf067cfe, 32'shcf057a23, 32'shcf04774f, 32'shcf037483, 32'shcf0271bf, 32'shcf016f02, 32'shcf006c4d, 
               32'shceff699f, 32'shcefe66f9, 32'shcefd645a, 32'shcefc61c3, 32'shcefb5f34, 32'shcefa5cac, 32'shcef95a2b, 32'shcef857b2, 
               32'shcef75541, 32'shcef652d7, 32'shcef55075, 32'shcef44e1b, 32'shcef34bc8, 32'shcef2497c, 32'shcef14738, 32'shcef044fc, 
               32'shceef42c7, 32'shceee409a, 32'shceed3e74, 32'shceec3c56, 32'shceeb3a40, 32'shceea3831, 32'shcee93629, 32'shcee8342a, 
               32'shcee73231, 32'shcee63041, 32'shcee52e58, 32'shcee42c76, 32'shcee32a9c, 32'shcee228ca, 32'shcee126ff, 32'shcee0253c, 
               32'shcedf2380, 32'shcede21cc, 32'shcedd2020, 32'shcedc1e7b, 32'shcedb1cde, 32'shceda1b48, 32'shced919ba, 32'shced81833, 
               32'shced716b4, 32'shced6153d, 32'shced513cd, 32'shced41265, 32'shced31104, 32'shced20fab, 32'shced10e59, 32'shced00d0f, 
               32'shcecf0bcd, 32'shcece0a92, 32'shcecd095f, 32'shcecc0833, 32'shcecb070f, 32'shceca05f3, 32'shcec904de, 32'shcec803d1, 
               32'shcec702cb, 32'shcec601cd, 32'shcec500d7, 32'shcec3ffe8, 32'shcec2ff01, 32'shcec1fe21, 32'shcec0fd49, 32'shcebffc79, 
               32'shcebefbb0, 32'shcebdfaee, 32'shcebcfa35, 32'shcebbf983, 32'shcebaf8d8, 32'shceb9f835, 32'shceb8f79a, 32'shceb7f706, 
               32'shceb6f67a, 32'shceb5f5f5, 32'shceb4f579, 32'shceb3f503, 32'shceb2f496, 32'shceb1f42f, 32'shceb0f3d1, 32'shceaff37a, 
               32'shceaef32b, 32'shceadf2e3, 32'shceacf2a3, 32'shceabf26b, 32'shceaaf23a, 32'shcea9f210, 32'shcea8f1ef, 32'shcea7f1d5, 
               32'shcea6f1c2, 32'shcea5f1b7, 32'shcea4f1b4, 32'shcea3f1b9, 32'shcea2f1c5, 32'shcea1f1d8, 32'shcea0f1f4, 32'shce9ff216, 
               32'shce9ef241, 32'shce9df273, 32'shce9cf2ad, 32'shce9bf2ee, 32'shce9af337, 32'shce99f387, 32'shce98f3e0, 32'shce97f43f, 
               32'shce96f4a7, 32'shce95f516, 32'shce94f58c, 32'shce93f60b, 32'shce92f691, 32'shce91f71e, 32'shce90f7b3, 32'shce8ff850, 
               32'shce8ef8f4, 32'shce8df9a0, 32'shce8cfa54, 32'shce8bfb0f, 32'shce8afbd2, 32'shce89fc9d, 32'shce88fd6f, 32'shce87fe48, 
               32'shce86ff2a, 32'shce860013, 32'shce850104, 32'shce8401fc, 32'shce8302fc, 32'shce820403, 32'shce810512, 32'shce800629, 
               32'shce7f0748, 32'shce7e086e, 32'shce7d099b, 32'shce7c0ad1, 32'shce7b0c0e, 32'shce7a0d52, 32'shce790e9f, 32'shce780ff3, 
               32'shce77114e, 32'shce7612b1, 32'shce75141c, 32'shce74158e, 32'shce731709, 32'shce72188a, 32'shce711a14, 32'shce701ba5, 
               32'shce6f1d3d, 32'shce6e1ede, 32'shce6d2086, 32'shce6c2235, 32'shce6b23ec, 32'shce6a25ab, 32'shce692772, 32'shce682940, 
               32'shce672b16, 32'shce662cf3, 32'shce652ed8, 32'shce6430c5, 32'shce6332ba, 32'shce6234b6, 32'shce6136b9, 32'shce6038c5, 
               32'shce5f3ad8, 32'shce5e3cf2, 32'shce5d3f15, 32'shce5c413f, 32'shce5b4370, 32'shce5a45aa, 32'shce5947eb, 32'shce584a33, 
               32'shce574c84, 32'shce564edc, 32'shce55513b, 32'shce5453a2, 32'shce535611, 32'shce525888, 32'shce515b06, 32'shce505d8c, 
               32'shce4f6019, 32'shce4e62af, 32'shce4d654c, 32'shce4c67f0, 32'shce4b6a9c, 32'shce4a6d50, 32'shce49700c, 32'shce4872cf, 
               32'shce47759a, 32'shce46786c, 32'shce457b47, 32'shce447e28, 32'shce438112, 32'shce428403, 32'shce4186fc, 32'shce4089fd, 
               32'shce3f8d05, 32'shce3e9015, 32'shce3d932c, 32'shce3c964c, 32'shce3b9973, 32'shce3a9ca1, 32'shce399fd7, 32'shce38a315, 
               32'shce37a65b, 32'shce36a9a8, 32'shce35acfd, 32'shce34b05a, 32'shce33b3be, 32'shce32b72a, 32'shce31ba9e, 32'shce30be19, 
               32'shce2fc19c, 32'shce2ec527, 32'shce2dc8ba, 32'shce2ccc54, 32'shce2bcff5, 32'shce2ad39f, 32'shce29d750, 32'shce28db09, 
               32'shce27dec9, 32'shce26e292, 32'shce25e662, 32'shce24ea39, 32'shce23ee18, 32'shce22f1ff, 32'shce21f5ee, 32'shce20f9e4, 
               32'shce1ffde2, 32'shce1f01e8, 32'shce1e05f6, 32'shce1d0a0b, 32'shce1c0e28, 32'shce1b124c, 32'shce1a1678, 32'shce191aac, 
               32'shce181ee8, 32'shce17232b, 32'shce162776, 32'shce152bc9, 32'shce143023, 32'shce133485, 32'shce1238ef, 32'shce113d60, 
               32'shce1041d9, 32'shce0f465a, 32'shce0e4ae3, 32'shce0d4f73, 32'shce0c540b, 32'shce0b58ab, 32'shce0a5d52, 32'shce096201, 
               32'shce0866b8, 32'shce076b77, 32'shce06703d, 32'shce05750b, 32'shce0479e0, 32'shce037ebe, 32'shce0283a3, 32'shce01888f, 
               32'shce008d84, 32'shcdff9280, 32'shcdfe9784, 32'shcdfd9c90, 32'shcdfca1a3, 32'shcdfba6be, 32'shcdfaabe1, 32'shcdf9b10b, 
               32'shcdf8b63d, 32'shcdf7bb77, 32'shcdf6c0b9, 32'shcdf5c602, 32'shcdf4cb53, 32'shcdf3d0ac, 32'shcdf2d60c, 32'shcdf1db74, 
               32'shcdf0e0e4, 32'shcdefe65c, 32'shcdeeebdb, 32'shcdedf162, 32'shcdecf6f1, 32'shcdebfc87, 32'shcdeb0226, 32'shcdea07cc, 
               32'shcde90d79, 32'shcde8132f, 32'shcde718ec, 32'shcde61eb1, 32'shcde5247d, 32'shcde42a52, 32'shcde3302e, 32'shcde23611, 
               32'shcde13bfd, 32'shcde041f0, 32'shcddf47eb, 32'shcdde4dee, 32'shcddd53f8, 32'shcddc5a0a, 32'shcddb6024, 32'shcdda6646, 
               32'shcdd96c6f, 32'shcdd872a0, 32'shcdd778d9, 32'shcdd67f19, 32'shcdd58562, 32'shcdd48bb2, 32'shcdd39209, 32'shcdd29869, 
               32'shcdd19ed0, 32'shcdd0a53f, 32'shcdcfabb6, 32'shcdceb234, 32'shcdcdb8ba, 32'shcdccbf48, 32'shcdcbc5de, 32'shcdcacc7b, 
               32'shcdc9d320, 32'shcdc8d9cd, 32'shcdc7e082, 32'shcdc6e73e, 32'shcdc5ee02, 32'shcdc4f4ce, 32'shcdc3fba2, 32'shcdc3027d, 
               32'shcdc20960, 32'shcdc1104b, 32'shcdc0173e, 32'shcdbf1e38, 32'shcdbe253a, 32'shcdbd2c44, 32'shcdbc3356, 32'shcdbb3a6f, 
               32'shcdba4190, 32'shcdb948b9, 32'shcdb84fea, 32'shcdb75722, 32'shcdb65e62, 32'shcdb565aa, 32'shcdb46cfa, 32'shcdb37451, 
               32'shcdb27bb0, 32'shcdb18317, 32'shcdb08a86, 32'shcdaf91fc, 32'shcdae997a, 32'shcdada100, 32'shcdaca88e, 32'shcdabb023, 
               32'shcdaab7c0, 32'shcda9bf65, 32'shcda8c712, 32'shcda7cec7, 32'shcda6d683, 32'shcda5de47, 32'shcda4e613, 32'shcda3ede6, 
               32'shcda2f5c2, 32'shcda1fda5, 32'shcda10590, 32'shcda00d82, 32'shcd9f157d, 32'shcd9e1d7f, 32'shcd9d2589, 32'shcd9c2d9a, 
               32'shcd9b35b4, 32'shcd9a3dd5, 32'shcd9945fe, 32'shcd984e2f, 32'shcd975668, 32'shcd965ea8, 32'shcd9566f0, 32'shcd946f40, 
               32'shcd937798, 32'shcd927ff7, 32'shcd91885e, 32'shcd9090cd, 32'shcd8f9944, 32'shcd8ea1c3, 32'shcd8daa49, 32'shcd8cb2d7, 
               32'shcd8bbb6d, 32'shcd8ac40b, 32'shcd89ccb0, 32'shcd88d55d, 32'shcd87de12, 32'shcd86e6cf, 32'shcd85ef94, 32'shcd84f860, 
               32'shcd840134, 32'shcd830a10, 32'shcd8212f4, 32'shcd811bdf, 32'shcd8024d3, 32'shcd7f2dce, 32'shcd7e36d1, 32'shcd7d3fdb, 
               32'shcd7c48ee, 32'shcd7b5208, 32'shcd7a5b2a, 32'shcd796454, 32'shcd786d85, 32'shcd7776bf, 32'shcd768000, 32'shcd758949, 
               32'shcd74929a, 32'shcd739bf2, 32'shcd72a553, 32'shcd71aebb, 32'shcd70b82b, 32'shcd6fc1a3, 32'shcd6ecb22, 32'shcd6dd4a9, 
               32'shcd6cde39, 32'shcd6be7d0, 32'shcd6af16e, 32'shcd69fb15, 32'shcd6904c3, 32'shcd680e79, 32'shcd671837, 32'shcd6621fd, 
               32'shcd652bcb, 32'shcd6435a0, 32'shcd633f7d, 32'shcd624962, 32'shcd61534f, 32'shcd605d44, 32'shcd5f6740, 32'shcd5e7144, 
               32'shcd5d7b50, 32'shcd5c8564, 32'shcd5b8f80, 32'shcd5a99a3, 32'shcd59a3ce, 32'shcd58ae01, 32'shcd57b83c, 32'shcd56c27f, 
               32'shcd55ccca, 32'shcd54d71c, 32'shcd53e176, 32'shcd52ebd8, 32'shcd51f642, 32'shcd5100b3, 32'shcd500b2d, 32'shcd4f15ae, 
               32'shcd4e2037, 32'shcd4d2ac8, 32'shcd4c3560, 32'shcd4b4001, 32'shcd4a4aa9, 32'shcd495559, 32'shcd486011, 32'shcd476ad1, 
               32'shcd467599, 32'shcd458068, 32'shcd448b3f, 32'shcd43961e, 32'shcd42a105, 32'shcd41abf4, 32'shcd40b6ea, 32'shcd3fc1e9, 
               32'shcd3eccef, 32'shcd3dd7fd, 32'shcd3ce313, 32'shcd3bee30, 32'shcd3af956, 32'shcd3a0483, 32'shcd390fb8, 32'shcd381af5, 
               32'shcd37263a, 32'shcd363187, 32'shcd353cdb, 32'shcd344837, 32'shcd33539c, 32'shcd325f08, 32'shcd316a7b, 32'shcd3075f7, 
               32'shcd2f817b, 32'shcd2e8d06, 32'shcd2d9899, 32'shcd2ca434, 32'shcd2bafd7, 32'shcd2abb81, 32'shcd29c734, 32'shcd28d2ee, 
               32'shcd27deb0, 32'shcd26ea7b, 32'shcd25f64c, 32'shcd250226, 32'shcd240e08, 32'shcd2319f1, 32'shcd2225e2, 32'shcd2131db, 
               32'shcd203ddc, 32'shcd1f49e5, 32'shcd1e55f6, 32'shcd1d620e, 32'shcd1c6e2e, 32'shcd1b7a57, 32'shcd1a8687, 32'shcd1992be, 
               32'shcd189efe, 32'shcd17ab46, 32'shcd16b795, 32'shcd15c3ec, 32'shcd14d04b, 32'shcd13dcb2, 32'shcd12e921, 32'shcd11f598, 
               32'shcd110216, 32'shcd100e9d, 32'shcd0f1b2b, 32'shcd0e27c1, 32'shcd0d345f, 32'shcd0c4105, 32'shcd0b4db3, 32'shcd0a5a68, 
               32'shcd096725, 32'shcd0873eb, 32'shcd0780b8, 32'shcd068d8d, 32'shcd059a6a, 32'shcd04a74e, 32'shcd03b43b, 32'shcd02c12f, 
               32'shcd01ce2b, 32'shcd00db30, 32'shccffe83c, 32'shccfef54f, 32'shccfe026b, 32'shccfd0f8f, 32'shccfc1cba, 32'shccfb29ed, 
               32'shccfa3729, 32'shccf9446c, 32'shccf851b7, 32'shccf75f09, 32'shccf66c64, 32'shccf579c7, 32'shccf48731, 32'shccf394a3, 
               32'shccf2a21d, 32'shccf1af9f, 32'shccf0bd29, 32'shccefcabb, 32'shcceed855, 32'shccede5f6, 32'shccecf3a0, 32'shccec0151, 
               32'shcceb0f0a, 32'shccea1ccb, 32'shcce92a94, 32'shcce83865, 32'shcce7463e, 32'shcce6541e, 32'shcce56206, 32'shcce46ff7, 
               32'shcce37def, 32'shcce28bef, 32'shcce199f7, 32'shcce0a807, 32'shccdfb61f, 32'shccdec43e, 32'shccddd266, 32'shccdce095, 
               32'shccdbeecc, 32'shccdafd0b, 32'shccda0b52, 32'shccd919a1, 32'shccd827f8, 32'shccd73657, 32'shccd644bd, 32'shccd5532c, 
               32'shccd461a2, 32'shccd37021, 32'shccd27ea7, 32'shccd18d35, 32'shccd09bcb, 32'shcccfaa69, 32'shccceb90e, 32'shcccdc7bc, 
               32'shccccd671, 32'shcccbe52f, 32'shcccaf3f4, 32'shccca02c1, 32'shccc91196, 32'shccc82073, 32'shccc72f58, 32'shccc63e45, 
               32'shccc54d3a, 32'shccc45c36, 32'shccc36b3b, 32'shccc27a47, 32'shccc1895c, 32'shccc09878, 32'shccbfa79c, 32'shccbeb6c8, 
               32'shccbdc5fc, 32'shccbcd538, 32'shccbbe47b, 32'shccbaf3c7, 32'shccba031a, 32'shccb91276, 32'shccb821d9, 32'shccb73144, 
               32'shccb640b8, 32'shccb55033, 32'shccb45fb6, 32'shccb36f41, 32'shccb27ed3, 32'shccb18e6e, 32'shccb09e11, 32'shccafadbb, 
               32'shccaebd6e, 32'shccadcd28, 32'shccacdcea, 32'shccabecb5, 32'shccaafc87, 32'shccaa0c61, 32'shcca91c43, 32'shcca82c2d, 
               32'shcca73c1e, 32'shcca64c18, 32'shcca55c1a, 32'shcca46c23, 32'shcca37c35, 32'shcca28c4e, 32'shcca19c6f, 32'shcca0ac99, 
               32'shcc9fbcca, 32'shcc9ecd03, 32'shcc9ddd44, 32'shcc9ced8d, 32'shcc9bfddd, 32'shcc9b0e36, 32'shcc9a1e97, 32'shcc992f00, 
               32'shcc983f70, 32'shcc974fe9, 32'shcc966069, 32'shcc9570f1, 32'shcc948182, 32'shcc93921a, 32'shcc92a2ba, 32'shcc91b362, 
               32'shcc90c412, 32'shcc8fd4ca, 32'shcc8ee58a, 32'shcc8df651, 32'shcc8d0721, 32'shcc8c17f9, 32'shcc8b28d8, 32'shcc8a39c0, 
               32'shcc894aaf, 32'shcc885ba7, 32'shcc876ca6, 32'shcc867dad, 32'shcc858ebc, 32'shcc849fd4, 32'shcc83b0f3, 32'shcc82c21a, 
               32'shcc81d349, 32'shcc80e47f, 32'shcc7ff5be, 32'shcc7f0705, 32'shcc7e1854, 32'shcc7d29aa, 32'shcc7c3b09, 32'shcc7b4c70, 
               32'shcc7a5dde, 32'shcc796f55, 32'shcc7880d3, 32'shcc779259, 32'shcc76a3e8, 32'shcc75b57e, 32'shcc74c71c, 32'shcc73d8c2, 
               32'shcc72ea70, 32'shcc71fc26, 32'shcc710de4, 32'shcc701faa, 32'shcc6f3178, 32'shcc6e434e, 32'shcc6d552c, 32'shcc6c6711, 
               32'shcc6b78ff, 32'shcc6a8af5, 32'shcc699cf2, 32'shcc68aef8, 32'shcc67c105, 32'shcc66d31b, 32'shcc65e538, 32'shcc64f75e, 
               32'shcc64098b, 32'shcc631bc0, 32'shcc622dfd, 32'shcc614043, 32'shcc605290, 32'shcc5f64e5, 32'shcc5e7742, 32'shcc5d89a7, 
               32'shcc5c9c14, 32'shcc5bae89, 32'shcc5ac106, 32'shcc59d38b, 32'shcc58e618, 32'shcc57f8ad, 32'shcc570b4a, 32'shcc561dee, 
               32'shcc55309b, 32'shcc544350, 32'shcc53560c, 32'shcc5268d1, 32'shcc517b9e, 32'shcc508e72, 32'shcc4fa14f, 32'shcc4eb433, 
               32'shcc4dc720, 32'shcc4cda14, 32'shcc4bed11, 32'shcc4b0015, 32'shcc4a1322, 32'shcc492636, 32'shcc483952, 32'shcc474c77, 
               32'shcc465fa3, 32'shcc4572d7, 32'shcc448614, 32'shcc439958, 32'shcc42aca4, 32'shcc41bff8, 32'shcc40d354, 32'shcc3fe6b8, 
               32'shcc3efa25, 32'shcc3e0d99, 32'shcc3d2115, 32'shcc3c3499, 32'shcc3b4825, 32'shcc3a5bb9, 32'shcc396f55, 32'shcc3882f9, 
               32'shcc3796a5, 32'shcc36aa59, 32'shcc35be15, 32'shcc34d1d9, 32'shcc33e5a5, 32'shcc32f979, 32'shcc320d55, 32'shcc312139, 
               32'shcc303524, 32'shcc2f4918, 32'shcc2e5d14, 32'shcc2d7118, 32'shcc2c8524, 32'shcc2b9938, 32'shcc2aad54, 32'shcc29c177, 
               32'shcc28d5a3, 32'shcc27e9d7, 32'shcc26fe13, 32'shcc261257, 32'shcc2526a2, 32'shcc243af6, 32'shcc234f52, 32'shcc2263b6, 
               32'shcc217822, 32'shcc208c95, 32'shcc1fa111, 32'shcc1eb595, 32'shcc1dca21, 32'shcc1cdeb5, 32'shcc1bf350, 32'shcc1b07f4, 
               32'shcc1a1ca0, 32'shcc193154, 32'shcc184610, 32'shcc175ad3, 32'shcc166f9f, 32'shcc158473, 32'shcc14994f, 32'shcc13ae33, 
               32'shcc12c31f, 32'shcc11d813, 32'shcc10ed0e, 32'shcc100212, 32'shcc0f171e, 32'shcc0e2c32, 32'shcc0d414e, 32'shcc0c5672, 
               32'shcc0b6b9e, 32'shcc0a80d2, 32'shcc09960e, 32'shcc08ab52, 32'shcc07c09e, 32'shcc06d5f2, 32'shcc05eb4e, 32'shcc0500b2, 
               32'shcc04161e, 32'shcc032b92, 32'shcc02410e, 32'shcc015692, 32'shcc006c1e, 32'shcbff81b2, 32'shcbfe974e, 32'shcbfdacf2, 
               32'shcbfcc29f, 32'shcbfbd853, 32'shcbfaee0f, 32'shcbfa03d3, 32'shcbf919a0, 32'shcbf82f74, 32'shcbf74550, 32'shcbf65b34, 
               32'shcbf57121, 32'shcbf48715, 32'shcbf39d12, 32'shcbf2b316, 32'shcbf1c923, 32'shcbf0df37, 32'shcbeff554, 32'shcbef0b78, 
               32'shcbee21a5, 32'shcbed37d9, 32'shcbec4e16, 32'shcbeb645b, 32'shcbea7aa7, 32'shcbe990fc, 32'shcbe8a759, 32'shcbe7bdbe, 
               32'shcbe6d42b, 32'shcbe5ea9f, 32'shcbe5011c, 32'shcbe417a1, 32'shcbe32e2e, 32'shcbe244c3, 32'shcbe15b60, 32'shcbe07205, 
               32'shcbdf88b3, 32'shcbde9f68, 32'shcbddb625, 32'shcbdcccea, 32'shcbdbe3b7, 32'shcbdafa8d, 32'shcbda116a, 32'shcbd92850, 
               32'shcbd83f3d, 32'shcbd75633, 32'shcbd66d30, 32'shcbd58436, 32'shcbd49b43, 32'shcbd3b259, 32'shcbd2c977, 32'shcbd1e09c, 
               32'shcbd0f7ca, 32'shcbd00f00, 32'shcbcf263e, 32'shcbce3d84, 32'shcbcd54d2, 32'shcbcc6c28, 32'shcbcb8386, 32'shcbca9aec, 
               32'shcbc9b25a, 32'shcbc8c9d1, 32'shcbc7e14f, 32'shcbc6f8d5, 32'shcbc61064, 32'shcbc527fa, 32'shcbc43f99, 32'shcbc3573f, 
               32'shcbc26eee, 32'shcbc186a5, 32'shcbc09e64, 32'shcbbfb62a, 32'shcbbecdf9, 32'shcbbde5d0, 32'shcbbcfdaf, 32'shcbbc1596, 
               32'shcbbb2d85, 32'shcbba457c, 32'shcbb95d7c, 32'shcbb87583, 32'shcbb78d92, 32'shcbb6a5aa, 32'shcbb5bdc9, 32'shcbb4d5f1, 
               32'shcbb3ee20, 32'shcbb30658, 32'shcbb21e98, 32'shcbb136df, 32'shcbb04f2f, 32'shcbaf6787, 32'shcbae7fe7, 32'shcbad984f, 
               32'shcbacb0bf, 32'shcbabc938, 32'shcbaae1b8, 32'shcba9fa40, 32'shcba912d1, 32'shcba82b69, 32'shcba7440a, 32'shcba65cb2, 
               32'shcba57563, 32'shcba48e1c, 32'shcba3a6dd, 32'shcba2bfa6, 32'shcba1d877, 32'shcba0f150, 32'shcba00a31, 32'shcb9f231a, 
               32'shcb9e3c0b, 32'shcb9d5505, 32'shcb9c6e06, 32'shcb9b8710, 32'shcb9aa021, 32'shcb99b93b, 32'shcb98d25d, 32'shcb97eb87, 
               32'shcb9704b9, 32'shcb961df3, 32'shcb953735, 32'shcb94507f, 32'shcb9369d1, 32'shcb92832c, 32'shcb919c8e, 32'shcb90b5f9, 
               32'shcb8fcf6b, 32'shcb8ee8e6, 32'shcb8e0269, 32'shcb8d1bf4, 32'shcb8c3587, 32'shcb8b4f22, 32'shcb8a68c5, 32'shcb898270, 
               32'shcb889c23, 32'shcb87b5df, 32'shcb86cfa2, 32'shcb85e96e, 32'shcb850342, 32'shcb841d1d, 32'shcb833701, 32'shcb8250ed, 
               32'shcb816ae1, 32'shcb8084de, 32'shcb7f9ee2, 32'shcb7eb8ee, 32'shcb7dd303, 32'shcb7ced1f, 32'shcb7c0744, 32'shcb7b2171, 
               32'shcb7a3ba5, 32'shcb7955e2, 32'shcb787027, 32'shcb778a75, 32'shcb76a4ca, 32'shcb75bf27, 32'shcb74d98d, 32'shcb73f3fa, 
               32'shcb730e70, 32'shcb7228ee, 32'shcb714373, 32'shcb705e01, 32'shcb6f7898, 32'shcb6e9336, 32'shcb6daddc, 32'shcb6cc88a, 
               32'shcb6be341, 32'shcb6afe00, 32'shcb6a18c6, 32'shcb693395, 32'shcb684e6c, 32'shcb67694b, 32'shcb668432, 32'shcb659f22, 
               32'shcb64ba19, 32'shcb63d518, 32'shcb62f020, 32'shcb620b30, 32'shcb612648, 32'shcb604168, 32'shcb5f5c90, 32'shcb5e77c0, 
               32'shcb5d92f8, 32'shcb5cae39, 32'shcb5bc981, 32'shcb5ae4d2, 32'shcb5a002b, 32'shcb591b8b, 32'shcb5836f4, 32'shcb575266, 
               32'shcb566ddf, 32'shcb558960, 32'shcb54a4ea, 32'shcb53c07b, 32'shcb52dc15, 32'shcb51f7b7, 32'shcb511361, 32'shcb502f13, 
               32'shcb4f4acd, 32'shcb4e6690, 32'shcb4d825a, 32'shcb4c9e2d, 32'shcb4bba08, 32'shcb4ad5ea, 32'shcb49f1d5, 32'shcb490dc9, 
               32'shcb4829c4, 32'shcb4745c7, 32'shcb4661d3, 32'shcb457de6, 32'shcb449a02, 32'shcb43b626, 32'shcb42d252, 32'shcb41ee86, 
               32'shcb410ac3, 32'shcb402707, 32'shcb3f4354, 32'shcb3e5fa8, 32'shcb3d7c05, 32'shcb3c986a, 32'shcb3bb4d7, 32'shcb3ad14d, 
               32'shcb39edca, 32'shcb390a50, 32'shcb3826dd, 32'shcb374373, 32'shcb366011, 32'shcb357cb7, 32'shcb349965, 32'shcb33b61c, 
               32'shcb32d2da, 32'shcb31efa1, 32'shcb310c70, 32'shcb302947, 32'shcb2f4626, 32'shcb2e630d, 32'shcb2d7ffc, 32'shcb2c9cf4, 
               32'shcb2bb9f4, 32'shcb2ad6fb, 32'shcb29f40b, 32'shcb291123, 32'shcb282e44, 32'shcb274b6c, 32'shcb26689d, 32'shcb2585d5, 
               32'shcb24a316, 32'shcb23c05f, 32'shcb22ddb1, 32'shcb21fb0a, 32'shcb21186b, 32'shcb2035d5, 32'shcb1f5347, 32'shcb1e70c1, 
               32'shcb1d8e43, 32'shcb1cabcd, 32'shcb1bc95f, 32'shcb1ae6fa, 32'shcb1a049d, 32'shcb192248, 32'shcb183ffb, 32'shcb175db6, 
               32'shcb167b79, 32'shcb159945, 32'shcb14b718, 32'shcb13d4f4, 32'shcb12f2d8, 32'shcb1210c4, 32'shcb112eb9, 32'shcb104cb5, 
               32'shcb0f6aba, 32'shcb0e88c7, 32'shcb0da6dc, 32'shcb0cc4f9, 32'shcb0be31e, 32'shcb0b014b, 32'shcb0a1f81, 32'shcb093dbf, 
               32'shcb085c05, 32'shcb077a53, 32'shcb0698a9, 32'shcb05b708, 32'shcb04d56e, 32'shcb03f3dd, 32'shcb031254, 32'shcb0230d3, 
               32'shcb014f5b, 32'shcb006dea, 32'shcaff8c82, 32'shcafeab22, 32'shcafdc9ca, 32'shcafce87a, 32'shcafc0732, 32'shcafb25f3, 
               32'shcafa44bc, 32'shcaf9638d, 32'shcaf88266, 32'shcaf7a147, 32'shcaf6c030, 32'shcaf5df22, 32'shcaf4fe1c, 32'shcaf41d1e, 
               32'shcaf33c28, 32'shcaf25b3a, 32'shcaf17a55, 32'shcaf09977, 32'shcaefb8a2, 32'shcaeed7d5, 32'shcaedf711, 32'shcaed1654, 
               32'shcaec35a0, 32'shcaeb54f3, 32'shcaea744f, 32'shcae993b4, 32'shcae8b320, 32'shcae7d295, 32'shcae6f211, 32'shcae61196, 
               32'shcae53123, 32'shcae450b9, 32'shcae37056, 32'shcae28ffc, 32'shcae1afaa, 32'shcae0cf60, 32'shcadfef1e, 32'shcadf0ee4, 
               32'shcade2eb3, 32'shcadd4e8a, 32'shcadc6e69, 32'shcadb8e50, 32'shcadaae40, 32'shcad9ce37, 32'shcad8ee37, 32'shcad80e3f, 
               32'shcad72e4f, 32'shcad64e68, 32'shcad56e88, 32'shcad48eb1, 32'shcad3aee2, 32'shcad2cf1b, 32'shcad1ef5d, 32'shcad10fa6, 
               32'shcad02ff8, 32'shcacf5052, 32'shcace70b4, 32'shcacd911f, 32'shcaccb191, 32'shcacbd20c, 32'shcacaf28f, 32'shcaca131a, 
               32'shcac933ae, 32'shcac8544a, 32'shcac774ed, 32'shcac69599, 32'shcac5b64e, 32'shcac4d70a, 32'shcac3f7cf, 32'shcac3189c, 
               32'shcac23971, 32'shcac15a4e, 32'shcac07b34, 32'shcabf9c21, 32'shcabebd17, 32'shcabdde16, 32'shcabcff1c, 32'shcabc202a, 
               32'shcabb4141, 32'shcaba6260, 32'shcab98388, 32'shcab8a4b7, 32'shcab7c5ef, 32'shcab6e72f, 32'shcab60877, 32'shcab529c7, 
               32'shcab44b1f, 32'shcab36c80, 32'shcab28de9, 32'shcab1af5a, 32'shcab0d0d4, 32'shcaaff255, 32'shcaaf13df, 32'shcaae3571, 
               32'shcaad570c, 32'shcaac78ae, 32'shcaab9a59, 32'shcaaabc0c, 32'shcaa9ddc7, 32'shcaa8ff8a, 32'shcaa82156, 32'shcaa7432a, 
               32'shcaa66506, 32'shcaa586ea, 32'shcaa4a8d7, 32'shcaa3cacc, 32'shcaa2ecc9, 32'shcaa20ece, 32'shcaa130db, 32'shcaa052f1, 
               32'shca9f750f, 32'shca9e9735, 32'shca9db964, 32'shca9cdb9a, 32'shca9bfdd9, 32'shca9b2020, 32'shca9a4270, 32'shca9964c7, 
               32'shca988727, 32'shca97a98f, 32'shca96cbff, 32'shca95ee78, 32'shca9510f8, 32'shca943381, 32'shca935613, 32'shca9278ac, 
               32'shca919b4e, 32'shca90bdf8, 32'shca8fe0aa, 32'shca8f0364, 32'shca8e2627, 32'shca8d48f2, 32'shca8c6bc5, 32'shca8b8ea0, 
               32'shca8ab184, 32'shca89d470, 32'shca88f764, 32'shca881a60, 32'shca873d65, 32'shca866072, 32'shca858387, 32'shca84a6a4, 
               32'shca83c9ca, 32'shca82ecf8, 32'shca82102e, 32'shca81336c, 32'shca8056b3, 32'shca7f7a02, 32'shca7e9d59, 32'shca7dc0b8, 
               32'shca7ce420, 32'shca7c078f, 32'shca7b2b08, 32'shca7a4e88, 32'shca797211, 32'shca7895a1, 32'shca77b93b, 32'shca76dcdc, 
               32'shca760086, 32'shca752437, 32'shca7447f2, 32'shca736bb4, 32'shca728f7f, 32'shca71b351, 32'shca70d72d, 32'shca6ffb10, 
               32'shca6f1efc, 32'shca6e42f0, 32'shca6d66ec, 32'shca6c8af0, 32'shca6baefd, 32'shca6ad312, 32'shca69f72f, 32'shca691b55, 
               32'shca683f83, 32'shca6763b9, 32'shca6687f7, 32'shca65ac3e, 32'shca64d08d, 32'shca63f4e4, 32'shca631943, 32'shca623dab, 
               32'shca61621b, 32'shca608693, 32'shca5fab13, 32'shca5ecf9c, 32'shca5df42d, 32'shca5d18c6, 32'shca5c3d68, 32'shca5b6212, 
               32'shca5a86c4, 32'shca59ab7e, 32'shca58d041, 32'shca57f50c, 32'shca5719df, 32'shca563eba, 32'shca55639e, 32'shca54888a, 
               32'shca53ad7e, 32'shca52d27b, 32'shca51f780, 32'shca511c8d, 32'shca5041a2, 32'shca4f66c0, 32'shca4e8be6, 32'shca4db114, 
               32'shca4cd64b, 32'shca4bfb89, 32'shca4b20d0, 32'shca4a4620, 32'shca496b77, 32'shca4890d7, 32'shca47b640, 32'shca46dbb0, 
               32'shca460129, 32'shca4526aa, 32'shca444c33, 32'shca4371c5, 32'shca42975f, 32'shca41bd01, 32'shca40e2ac, 32'shca40085e, 
               32'shca3f2e19, 32'shca3e53dd, 32'shca3d79a8, 32'shca3c9f7c, 32'shca3bc559, 32'shca3aeb3d, 32'shca3a112a, 32'shca39371f, 
               32'shca385d1d, 32'shca378322, 32'shca36a930, 32'shca35cf47, 32'shca34f565, 32'shca341b8c, 32'shca3341bb, 32'shca3267f3, 
               32'shca318e32, 32'shca30b47a, 32'shca2fdacb, 32'shca2f0123, 32'shca2e2784, 32'shca2d4dee, 32'shca2c745f, 32'shca2b9ad9, 
               32'shca2ac15b, 32'shca29e7e6, 32'shca290e79, 32'shca283514, 32'shca275bb7, 32'shca268263, 32'shca25a917, 32'shca24cfd3, 
               32'shca23f698, 32'shca231d64, 32'shca22443a, 32'shca216b17, 32'shca2091fd, 32'shca1fb8eb, 32'shca1edfe2, 32'shca1e06e0, 
               32'shca1d2de7, 32'shca1c54f7, 32'shca1b7c0e, 32'shca1aa32e, 32'shca19ca57, 32'shca18f187, 32'shca1818c0, 32'shca174001, 
               32'shca16674b, 32'shca158e9d, 32'shca14b5f7, 32'shca13dd59, 32'shca1304c4, 32'shca122c37, 32'shca1153b3, 32'shca107b37, 
               32'shca0fa2c3, 32'shca0eca57, 32'shca0df1f4, 32'shca0d1999, 32'shca0c4146, 32'shca0b68fc, 32'shca0a90ba, 32'shca09b880, 
               32'shca08e04f, 32'shca080826, 32'shca073005, 32'shca0657ed, 32'shca057fdd, 32'shca04a7d5, 32'shca03cfd5, 32'shca02f7de, 
               32'shca021fef, 32'shca014809, 32'shca00702b, 32'shc9ff9855, 32'shc9fec088, 32'shc9fde8c2, 32'shc9fd1106, 32'shc9fc3951, 
               32'shc9fb61a5, 32'shc9fa8a01, 32'shc9f9b266, 32'shc9f8dad3, 32'shc9f80348, 32'shc9f72bc5, 32'shc9f6544b, 32'shc9f57cd9, 
               32'shc9f4a570, 32'shc9f3ce0f, 32'shc9f2f6b6, 32'shc9f21f65, 32'shc9f1481d, 32'shc9f070dd, 32'shc9ef99a6, 32'shc9eec277, 
               32'shc9edeb50, 32'shc9ed1431, 32'shc9ec3d1b, 32'shc9eb660d, 32'shc9ea8f08, 32'shc9e9b80b, 32'shc9e8e116, 32'shc9e80a2a, 
               32'shc9e73346, 32'shc9e65c6a, 32'shc9e58596, 32'shc9e4aecb, 32'shc9e3d809, 32'shc9e3014e, 32'shc9e22a9c, 32'shc9e153f3, 
               32'shc9e07d51, 32'shc9dfa6b8, 32'shc9ded028, 32'shc9ddf99f, 32'shc9dd231f, 32'shc9dc4ca8, 32'shc9db7639, 32'shc9da9fd2, 
               32'shc9d9c973, 32'shc9d8f31d, 32'shc9d81ccf, 32'shc9d7468a, 32'shc9d6704c, 32'shc9d59a18, 32'shc9d4c3eb, 32'shc9d3edc7, 
               32'shc9d317ab, 32'shc9d24198, 32'shc9d16b8d, 32'shc9d0958a, 32'shc9cfbf90, 32'shc9cee99e, 32'shc9ce13b4, 32'shc9cd3dd3, 
               32'shc9cc67fa, 32'shc9cb922a, 32'shc9cabc62, 32'shc9c9e6a2, 32'shc9c910ea, 32'shc9c83b3b, 32'shc9c76595, 32'shc9c68ff6, 
               32'shc9c5ba60, 32'shc9c4e4d3, 32'shc9c40f4d, 32'shc9c339d0, 32'shc9c2645c, 32'shc9c18ef0, 32'shc9c0b98c, 32'shc9bfe430, 
               32'shc9bf0edd, 32'shc9be3993, 32'shc9bd6450, 32'shc9bc8f16, 32'shc9bbb9e5, 32'shc9bae4bc, 32'shc9ba0f9b, 32'shc9b93a82, 
               32'shc9b86572, 32'shc9b7906a, 32'shc9b6bb6b, 32'shc9b5e674, 32'shc9b51185, 32'shc9b43c9f, 32'shc9b367c1, 32'shc9b292eb, 
               32'shc9b1be1e, 32'shc9b0e95a, 32'shc9b0149d, 32'shc9af3fe9, 32'shc9ae6b3d, 32'shc9ad969a, 32'shc9acc1ff, 32'shc9abed6d, 
               32'shc9ab18e3, 32'shc9aa4461, 32'shc9a96fe7, 32'shc9a89b76, 32'shc9a7c70e, 32'shc9a6f2ae, 32'shc9a61e56, 32'shc9a54a06, 
               32'shc9a475bf, 32'shc9a3a180, 32'shc9a2cd4a, 32'shc9a1f91c, 32'shc9a124f7, 32'shc9a050d9, 32'shc99f7cc5, 32'shc99ea8b8, 
               32'shc99dd4b4, 32'shc99d00b8, 32'shc99c2cc5, 32'shc99b58da, 32'shc99a84f8, 32'shc999b11e, 32'shc998dd4c, 32'shc9980983, 
               32'shc99735c2, 32'shc9966209, 32'shc9958e59, 32'shc994bab1, 32'shc993e712, 32'shc993137b, 32'shc9923fed, 32'shc9916c66, 
               32'shc99098e9, 32'shc98fc573, 32'shc98ef206, 32'shc98e1ea2, 32'shc98d4b45, 32'shc98c77f2, 32'shc98ba4a6, 32'shc98ad163, 
               32'shc989fe29, 32'shc9892af6, 32'shc98857cd, 32'shc98784ab, 32'shc986b192, 32'shc985de82, 32'shc9850b79, 32'shc9843879, 
               32'shc9836582, 32'shc9829293, 32'shc981bfac, 32'shc980ecce, 32'shc98019f8, 32'shc97f472b, 32'shc97e7466, 32'shc97da1aa, 
               32'shc97ccef5, 32'shc97bfc4a, 32'shc97b29a6, 32'shc97a570b, 32'shc9798479, 32'shc978b1ef, 32'shc977df6d, 32'shc9770cf4, 
               32'shc9763a83, 32'shc975681a, 32'shc97495ba, 32'shc973c362, 32'shc972f113, 32'shc9721ecc, 32'shc9714c8e, 32'shc9707a58, 
               32'shc96fa82a, 32'shc96ed605, 32'shc96e03e8, 32'shc96d31d4, 32'shc96c5fc8, 32'shc96b8dc4, 32'shc96abbc9, 32'shc969e9d7, 
               32'shc96917ec, 32'shc968460a, 32'shc9677431, 32'shc966a260, 32'shc965d097, 32'shc964fed7, 32'shc9642d1f, 32'shc9635b70, 
               32'shc96289c9, 32'shc961b82b, 32'shc960e695, 32'shc9601507, 32'shc95f4382, 32'shc95e7205, 32'shc95da090, 32'shc95ccf25, 
               32'shc95bfdc1, 32'shc95b2c66, 32'shc95a5b13, 32'shc95989c9, 32'shc958b887, 32'shc957e74e, 32'shc957161d, 32'shc95644f4, 
               32'shc95573d4, 32'shc954a2bc, 32'shc953d1ad, 32'shc95300a6, 32'shc9522fa8, 32'shc9515eb2, 32'shc9508dc5, 32'shc94fbce0, 
               32'shc94eec03, 32'shc94e1b2f, 32'shc94d4a63, 32'shc94c79a0, 32'shc94ba8e5, 32'shc94ad832, 32'shc94a0788, 32'shc94936e7, 
               32'shc948664d, 32'shc94795bd, 32'shc946c534, 32'shc945f4b4, 32'shc945243d, 32'shc94453ce, 32'shc9438368, 32'shc942b30a, 
               32'shc941e2b4, 32'shc9411267, 32'shc9404222, 32'shc93f71e6, 32'shc93ea1b2, 32'shc93dd186, 32'shc93d0163, 32'shc93c3149, 
               32'shc93b6137, 32'shc93a912d, 32'shc939c12c, 32'shc938f133, 32'shc9382143, 32'shc937515b, 32'shc936817b, 32'shc935b1a5, 
               32'shc934e1d6, 32'shc9341210, 32'shc9334252, 32'shc932729d, 32'shc931a2f0, 32'shc930d34c, 32'shc93003b0, 32'shc92f341d, 
               32'shc92e6492, 32'shc92d9510, 32'shc92cc596, 32'shc92bf624, 32'shc92b26bb, 32'shc92a575a, 32'shc9298802, 32'shc928b8b3, 
               32'shc927e96b, 32'shc9271a2d, 32'shc9264af6, 32'shc9257bc8, 32'shc924aca3, 32'shc923dd86, 32'shc9230e71, 32'shc9223f65, 
               32'shc9217062, 32'shc920a167, 32'shc91fd274, 32'shc91f038a, 32'shc91e34a8, 32'shc91d65cf, 32'shc91c96fe, 32'shc91bc836, 
               32'shc91af976, 32'shc91a2abe, 32'shc9195c0f, 32'shc9188d69, 32'shc917becb, 32'shc916f035, 32'shc91621a8, 32'shc9155324, 
               32'shc91484a8, 32'shc913b634, 32'shc912e7c9, 32'shc9121966, 32'shc9114b0c, 32'shc9107cba, 32'shc90fae71, 32'shc90ee030, 
               32'shc90e11f7, 32'shc90d43c8, 32'shc90c75a0, 32'shc90ba781, 32'shc90ad96b, 32'shc90a0b5d, 32'shc9093d57, 32'shc9086f5a, 
               32'shc907a166, 32'shc906d379, 32'shc9060596, 32'shc90537bb, 32'shc90469e8, 32'shc9039c1e, 32'shc902ce5c, 32'shc90200a3, 
               32'shc90132f2, 32'shc900654a, 32'shc8ff97aa, 32'shc8feca13, 32'shc8fdfc84, 32'shc8fd2efe, 32'shc8fc6180, 32'shc8fb940b, 
               32'shc8fac69e, 32'shc8f9f939, 32'shc8f92bdd, 32'shc8f85e8a, 32'shc8f7913f, 32'shc8f6c3fd, 32'shc8f5f6c3, 32'shc8f52991, 
               32'shc8f45c68, 32'shc8f38f48, 32'shc8f2c230, 32'shc8f1f520, 32'shc8f12819, 32'shc8f05b1a, 32'shc8ef8e24, 32'shc8eec137, 
               32'shc8edf452, 32'shc8ed2775, 32'shc8ec5aa1, 32'shc8eb8dd6, 32'shc8eac112, 32'shc8e9f458, 32'shc8e927a6, 32'shc8e85afc, 
               32'shc8e78e5b, 32'shc8e6c1c2, 32'shc8e5f532, 32'shc8e528ab, 32'shc8e45c2c, 32'shc8e38fb5, 32'shc8e2c347, 32'shc8e1f6e1, 
               32'shc8e12a84, 32'shc8e05e2f, 32'shc8df91e3, 32'shc8dec5a0, 32'shc8ddf965, 32'shc8dd2d32, 32'shc8dc6108, 32'shc8db94e6, 
               32'shc8dac8cd, 32'shc8d9fcbd, 32'shc8d930b4, 32'shc8d864b5, 32'shc8d798be, 32'shc8d6cccf, 32'shc8d600e9, 32'shc8d5350c, 
               32'shc8d46936, 32'shc8d39d6a, 32'shc8d2d1a6, 32'shc8d205ea, 32'shc8d13a37, 32'shc8d06e8d, 32'shc8cfa2eb, 32'shc8ced751, 
               32'shc8ce0bc0, 32'shc8cd4038, 32'shc8cc74b8, 32'shc8cba940, 32'shc8caddd1, 32'shc8ca126b, 32'shc8c9470d, 32'shc8c87bb8, 
               32'shc8c7b06b, 32'shc8c6e527, 32'shc8c619eb, 32'shc8c54eb7, 32'shc8c4838d, 32'shc8c3b86a, 32'shc8c2ed50, 32'shc8c2223f, 
               32'shc8c15736, 32'shc8c08c36, 32'shc8bfc13f, 32'shc8bef64f, 32'shc8be2b69, 32'shc8bd608b, 32'shc8bc95b5, 32'shc8bbcae8, 
               32'shc8bb0023, 32'shc8ba3567, 32'shc8b96ab4, 32'shc8b8a009, 32'shc8b7d566, 32'shc8b70acc, 32'shc8b6403b, 32'shc8b575b2, 
               32'shc8b4ab32, 32'shc8b3e0ba, 32'shc8b3164a, 32'shc8b24be4, 32'shc8b18185, 32'shc8b0b730, 32'shc8afece2, 32'shc8af229e, 
               32'shc8ae5862, 32'shc8ad8e2e, 32'shc8acc403, 32'shc8abf9e0, 32'shc8ab2fc6, 32'shc8aa65b5, 32'shc8a99bac, 32'shc8a8d1ac, 
               32'shc8a807b4, 32'shc8a73dc4, 32'shc8a673dd, 32'shc8a5a9ff, 32'shc8a4e029, 32'shc8a4165c, 32'shc8a34c98, 32'shc8a282db, 
               32'shc8a1b928, 32'shc8a0ef7d, 32'shc8a025da, 32'shc89f5c40, 32'shc89e92af, 32'shc89dc926, 32'shc89cffa6, 32'shc89c362e, 
               32'shc89b6cbf, 32'shc89aa358, 32'shc899d9fa, 32'shc89910a4, 32'shc8984757, 32'shc8977e12, 32'shc896b4d6, 32'shc895eba3, 
               32'shc8952278, 32'shc8945956, 32'shc893903c, 32'shc892c72b, 32'shc891fe22, 32'shc8913522, 32'shc8906c2a, 32'shc88fa33b, 
               32'shc88eda54, 32'shc88e1176, 32'shc88d48a1, 32'shc88c7fd4, 32'shc88bb710, 32'shc88aee54, 32'shc88a25a1, 32'shc8895cf6, 
               32'shc8889454, 32'shc887cbba, 32'shc8870329, 32'shc8863aa1, 32'shc8857221, 32'shc884a9aa, 32'shc883e13b, 32'shc88318d5, 
               32'shc8825077, 32'shc8818822, 32'shc880bfd5, 32'shc87ff791, 32'shc87f2f56, 32'shc87e6723, 32'shc87d9ef8, 32'shc87cd6d7, 
               32'shc87c0ebd, 32'shc87b46ad, 32'shc87a7ea5, 32'shc879b6a5, 32'shc878eeae, 32'shc87826c0, 32'shc8775eda, 32'shc87696fd, 
               32'shc875cf28, 32'shc875075c, 32'shc8743f98, 32'shc87377dd, 32'shc872b02b, 32'shc871e881, 32'shc87120e0, 32'shc8705947, 
               32'shc86f91b7, 32'shc86eca2f, 32'shc86e02b0, 32'shc86d3b3a, 32'shc86c73cc, 32'shc86bac66, 32'shc86ae50a, 32'shc86a1db6, 
               32'shc869566a, 32'shc8688f27, 32'shc867c7ec, 32'shc86700ba, 32'shc8663991, 32'shc8657270, 32'shc864ab58, 32'shc863e449, 
               32'shc8631d42, 32'shc8625643, 32'shc8618f4d, 32'shc860c860, 32'shc860017b, 32'shc85f3a9f, 32'shc85e73cc, 32'shc85dad01, 
               32'shc85ce63e, 32'shc85c1f84, 32'shc85b58d3, 32'shc85a922b, 32'shc859cb8a, 32'shc85904f3, 32'shc8583e64, 32'shc85777de, 
               32'shc856b160, 32'shc855eaeb, 32'shc855247e, 32'shc8545e1a, 32'shc85397bf, 32'shc852d16c, 32'shc8520b22, 32'shc85144e0, 
               32'shc8507ea7, 32'shc84fb877, 32'shc84ef24f, 32'shc84e2c2f, 32'shc84d6619, 32'shc84ca00b, 32'shc84bda05, 32'shc84b1408, 
               32'shc84a4e14, 32'shc8498828, 32'shc848c245, 32'shc847fc6a, 32'shc8473698, 32'shc84670cf, 32'shc845ab0e, 32'shc844e556, 
               32'shc8441fa6, 32'shc84359ff, 32'shc8429461, 32'shc841cecb, 32'shc841093e, 32'shc84043b9, 32'shc83f7e3d, 32'shc83eb8ca, 
               32'shc83df35f, 32'shc83d2dfd, 32'shc83c68a3, 32'shc83ba352, 32'shc83ade0a, 32'shc83a18ca, 32'shc8395393, 32'shc8388e64, 
               32'shc837c93e, 32'shc8370420, 32'shc8363f0c, 32'shc83579ff, 32'shc834b4fc, 32'shc833f001, 32'shc8332b0e, 32'shc8326625, 
               32'shc831a143, 32'shc830dc6b, 32'shc830179b, 32'shc82f52d3, 32'shc82e8e15, 32'shc82dc95e, 32'shc82d04b1, 32'shc82c400c, 
               32'shc82b7b70, 32'shc82ab6dc, 32'shc829f251, 32'shc8292dce, 32'shc8286954, 32'shc827a4e3, 32'shc826e07a, 32'shc8261c1a, 
               32'shc82557c3, 32'shc8249374, 32'shc823cf2e, 32'shc8230af0, 32'shc82246bb, 32'shc821828f, 32'shc820be6b, 32'shc81ffa50, 
               32'shc81f363d, 32'shc81e7233, 32'shc81dae32, 32'shc81cea39, 32'shc81c2649, 32'shc81b6262, 32'shc81a9e83, 32'shc819daad, 
               32'shc81916df, 32'shc818531a, 32'shc8178f5e, 32'shc816cbaa, 32'shc81607ff, 32'shc815445d, 32'shc81480c3, 32'shc813bd32, 
               32'shc812f9a9, 32'shc8123629, 32'shc81172b2, 32'shc810af43, 32'shc80febdd, 32'shc80f287f, 32'shc80e652b, 32'shc80da1de, 
               32'shc80cde9b, 32'shc80c1b60, 32'shc80b582e, 32'shc80a9504, 32'shc809d1e3, 32'shc8090eca, 32'shc8084bba, 32'shc80788b3, 
               32'shc806c5b5, 32'shc80602bf, 32'shc8053fd2, 32'shc8047ced, 32'shc803ba11, 32'shc802f73d, 32'shc8023473, 32'shc80171b1, 
               32'shc800aef7, 32'shc7ffec46, 32'shc7ff299e, 32'shc7fe66fe, 32'shc7fda468, 32'shc7fce1d9, 32'shc7fc1f54, 32'shc7fb5cd7, 
               32'shc7fa9a62, 32'shc7f9d7f6, 32'shc7f91593, 32'shc7f85339, 32'shc7f790e7, 32'shc7f6ce9e, 32'shc7f60c5d, 32'shc7f54a25, 
               32'shc7f487f6, 32'shc7f3c5cf, 32'shc7f303b1, 32'shc7f2419c, 32'shc7f17f8f, 32'shc7f0bd8b, 32'shc7effb90, 32'shc7ef399d, 
               32'shc7ee77b3, 32'shc7edb5d2, 32'shc7ecf3f9, 32'shc7ec3229, 32'shc7eb7061, 32'shc7eaaea2, 32'shc7e9ecec, 32'shc7e92b3e, 
               32'shc7e8699a, 32'shc7e7a7fd, 32'shc7e6e66a, 32'shc7e624df, 32'shc7e5635c, 32'shc7e4a1e3, 32'shc7e3e072, 32'shc7e31f09, 
               32'shc7e25daa, 32'shc7e19c53, 32'shc7e0db04, 32'shc7e019be, 32'shc7df5881, 32'shc7de974d, 32'shc7ddd621, 32'shc7dd14fe, 
               32'shc7dc53e3, 32'shc7db92d2, 32'shc7dad1c9, 32'shc7da10c8, 32'shc7d94fd0, 32'shc7d88ee1, 32'shc7d7cdfb, 32'shc7d70d1d, 
               32'shc7d64c47, 32'shc7d58b7b, 32'shc7d4cab7, 32'shc7d409fc, 32'shc7d34949, 32'shc7d2889f, 32'shc7d1c7fe, 32'shc7d10766, 
               32'shc7d046d6, 32'shc7cf864e, 32'shc7cec5d0, 32'shc7ce055a, 32'shc7cd44ed, 32'shc7cc8488, 32'shc7cbc42c, 32'shc7cb03d9, 
               32'shc7ca438f, 32'shc7c9834d, 32'shc7c8c313, 32'shc7c802e3, 32'shc7c742bb, 32'shc7c6829c, 32'shc7c5c285, 32'shc7c50277, 
               32'shc7c44272, 32'shc7c38276, 32'shc7c2c282, 32'shc7c20297, 32'shc7c142b4, 32'shc7c082da, 32'shc7bfc309, 32'shc7bf0340, 
               32'shc7be4381, 32'shc7bd83ca, 32'shc7bcc41b, 32'shc7bc0475, 32'shc7bb44d8, 32'shc7ba8544, 32'shc7b9c5b8, 32'shc7b90635, 
               32'shc7b846ba, 32'shc7b78749, 32'shc7b6c7e0, 32'shc7b6087f, 32'shc7b54928, 32'shc7b489d9, 32'shc7b3ca92, 32'shc7b30b55, 
               32'shc7b24c20, 32'shc7b18cf3, 32'shc7b0cdd0, 32'shc7b00eb5, 32'shc7af4fa3, 32'shc7ae9099, 32'shc7add198, 32'shc7ad12a0, 
               32'shc7ac53b1, 32'shc7ab94ca, 32'shc7aad5ec, 32'shc7aa1716, 32'shc7a9584a, 32'shc7a89986, 32'shc7a7daca, 32'shc7a71c18, 
               32'shc7a65d6e, 32'shc7a59ecc, 32'shc7a4e034, 32'shc7a421a4, 32'shc7a3631d, 32'shc7a2a49e, 32'shc7a1e628, 32'shc7a127bb, 
               32'shc7a06957, 32'shc79faafb, 32'shc79eeca8, 32'shc79e2e5d, 32'shc79d701c, 32'shc79cb1e3, 32'shc79bf3b3, 32'shc79b358b, 
               32'shc79a776c, 32'shc799b956, 32'shc798fb48, 32'shc7983d44, 32'shc7977f48, 32'shc796c154, 32'shc7960369, 32'shc7954587, 
               32'shc79487ae, 32'shc793c9de, 32'shc7930c16, 32'shc7924e56, 32'shc79190a0, 32'shc790d2f2, 32'shc790154d, 32'shc78f57b1, 
               32'shc78e9a1d, 32'shc78ddc92, 32'shc78d1f10, 32'shc78c6196, 32'shc78ba425, 32'shc78ae6bd, 32'shc78a295e, 32'shc7896c07, 
               32'shc788aeb9, 32'shc787f174, 32'shc7873437, 32'shc7867703, 32'shc785b9d8, 32'shc784fcb5, 32'shc7843f9c, 32'shc783828b, 
               32'shc782c582, 32'shc7820883, 32'shc7814b8c, 32'shc7808e9d, 32'shc77fd1b8, 32'shc77f14db, 32'shc77e5807, 32'shc77d9b3c, 
               32'shc77cde79, 32'shc77c21bf, 32'shc77b650e, 32'shc77aa865, 32'shc779ebc5, 32'shc7792f2e, 32'shc77872a0, 32'shc777b61a, 
               32'shc776f99d, 32'shc7763d29, 32'shc77580be, 32'shc774c45b, 32'shc7740801, 32'shc7734bb0, 32'shc7728f67, 32'shc771d327, 
               32'shc77116f0, 32'shc7705ac2, 32'shc76f9e9c, 32'shc76ee27f, 32'shc76e266b, 32'shc76d6a5f, 32'shc76cae5c, 32'shc76bf262, 
               32'shc76b3671, 32'shc76a7a88, 32'shc769bea8, 32'shc76902d1, 32'shc7684702, 32'shc7678b3d, 32'shc766cf80, 32'shc76613cb, 
               32'shc7655820, 32'shc7649c7d, 32'shc763e0e3, 32'shc7632552, 32'shc76269c9, 32'shc761ae49, 32'shc760f2d2, 32'shc7603763, 
               32'shc75f7bfe, 32'shc75ec0a1, 32'shc75e054c, 32'shc75d4a01, 32'shc75c8ebe, 32'shc75bd384, 32'shc75b1853, 32'shc75a5d2a, 
               32'shc759a20a, 32'shc758e6f3, 32'shc7582be5, 32'shc75770df, 32'shc756b5e2, 32'shc755faee, 32'shc7554003, 32'shc7548520, 
               32'shc753ca46, 32'shc7530f75, 32'shc75254ac, 32'shc75199ed, 32'shc750df36, 32'shc7502488, 32'shc74f69e2, 32'shc74eaf45, 
               32'shc74df4b1, 32'shc74d3a26, 32'shc74c7fa4, 32'shc74bc52a, 32'shc74b0ab9, 32'shc74a5050, 32'shc74995f1, 32'shc748db9a, 
               32'shc748214c, 32'shc7476707, 32'shc746acca, 32'shc745f296, 32'shc745386b, 32'shc7447e49, 32'shc743c42f, 32'shc7430a1f, 
               32'shc7425016, 32'shc7419617, 32'shc740dc21, 32'shc7402233, 32'shc73f684e, 32'shc73eae71, 32'shc73df49e, 32'shc73d3ad3, 
               32'shc73c8111, 32'shc73bc758, 32'shc73b0da7, 32'shc73a53ff, 32'shc7399a60, 32'shc738e0ca, 32'shc738273d, 32'shc7376db8, 
               32'shc736b43c, 32'shc735fac8, 32'shc735415e, 32'shc73487fc, 32'shc733cea3, 32'shc7331553, 32'shc7325c0c, 32'shc731a2cd, 
               32'shc730e997, 32'shc730306a, 32'shc72f7745, 32'shc72ebe2a, 32'shc72e0517, 32'shc72d4c0d, 32'shc72c930b, 32'shc72bda13, 
               32'shc72b2123, 32'shc72a683c, 32'shc729af5d, 32'shc728f688, 32'shc7283dbb, 32'shc72784f7, 32'shc726cc3c, 32'shc7261389, 
               32'shc7255ae0, 32'shc724a23f, 32'shc723e9a6, 32'shc7233117, 32'shc7227890, 32'shc721c013, 32'shc721079d, 32'shc7204f31, 
               32'shc71f96ce, 32'shc71ede73, 32'shc71e2621, 32'shc71d6dd7, 32'shc71cb597, 32'shc71bfd5f, 32'shc71b4530, 32'shc71a8d0a, 
               32'shc719d4ed, 32'shc7191cd8, 32'shc71864cc, 32'shc717acc9, 32'shc716f4cf, 32'shc7163cdd, 32'shc71584f5, 32'shc714cd15, 
               32'shc714153e, 32'shc7135d6f, 32'shc712a5aa, 32'shc711eded, 32'shc7113639, 32'shc7107e8d, 32'shc70fc6eb, 32'shc70f0f51, 
               32'shc70e57c0, 32'shc70da038, 32'shc70ce8b9, 32'shc70c3142, 32'shc70b79d4, 32'shc70ac26f, 32'shc70a0b13, 32'shc70953c0, 
               32'shc7089c75, 32'shc707e533, 32'shc7072dfa, 32'shc70676ca, 32'shc705bfa2, 32'shc7050883, 32'shc704516d, 32'shc7039a60, 
               32'shc702e35c, 32'shc7022c60, 32'shc701756d, 32'shc700be83, 32'shc70007a2, 32'shc6ff50ca, 32'shc6fe99fa, 32'shc6fde333, 
               32'shc6fd2c75, 32'shc6fc75c0, 32'shc6fbbf13, 32'shc6fb0870, 32'shc6fa51d5, 32'shc6f99b43, 32'shc6f8e4b9, 32'shc6f82e39, 
               32'shc6f777c1, 32'shc6f6c152, 32'shc6f60aec, 32'shc6f5548f, 32'shc6f49e3a, 32'shc6f3e7ee, 32'shc6f331ab, 32'shc6f27b71, 
               32'shc6f1c540, 32'shc6f10f17, 32'shc6f058f8, 32'shc6efa2e1, 32'shc6eeecd3, 32'shc6ee36cd, 32'shc6ed80d1, 32'shc6eccadd, 
               32'shc6ec14f2, 32'shc6eb5f10, 32'shc6eaa936, 32'shc6e9f366, 32'shc6e93d9e, 32'shc6e887df, 32'shc6e7d229, 32'shc6e71c7c, 
               32'shc6e666d7, 32'shc6e5b13c, 32'shc6e4fba9, 32'shc6e4461f, 32'shc6e3909d, 32'shc6e2db25, 32'shc6e225b5, 32'shc6e1704e, 
               32'shc6e0baf0, 32'shc6e0059b, 32'shc6df504f, 32'shc6de9b0b, 32'shc6dde5d0, 32'shc6dd309e, 32'shc6dc7b75, 32'shc6dbc654, 
               32'shc6db113d, 32'shc6da5c2e, 32'shc6d9a728, 32'shc6d8f22b, 32'shc6d83d37, 32'shc6d7884b, 32'shc6d6d369, 32'shc6d61e8f, 
               32'shc6d569be, 32'shc6d4b4f5, 32'shc6d40036, 32'shc6d34b7f, 32'shc6d296d1, 32'shc6d1e22d, 32'shc6d12d90, 32'shc6d078fd, 
               32'shc6cfc472, 32'shc6cf0ff1, 32'shc6ce5b78, 32'shc6cda708, 32'shc6ccf2a1, 32'shc6cc3e42, 32'shc6cb89ed, 32'shc6cad5a0, 
               32'shc6ca215c, 32'shc6c96d21, 32'shc6c8b8ee, 32'shc6c804c5, 32'shc6c750a4, 32'shc6c69c8c, 32'shc6c5e87d, 32'shc6c53477, 
               32'shc6c4807a, 32'shc6c3cc85, 32'shc6c31899, 32'shc6c264b7, 32'shc6c1b0dd, 32'shc6c0fd0b, 32'shc6c04943, 32'shc6bf9583, 
               32'shc6bee1cd, 32'shc6be2e1f, 32'shc6bd7a7a, 32'shc6bcc6dd, 32'shc6bc134a, 32'shc6bb5fbf, 32'shc6baac3d, 32'shc6b9f8c5, 
               32'shc6b94554, 32'shc6b891ed, 32'shc6b7de8f, 32'shc6b72b39, 32'shc6b677ec, 32'shc6b5c4a8, 32'shc6b5116d, 32'shc6b45e3b, 
               32'shc6b3ab12, 32'shc6b2f7f1, 32'shc6b244d9, 32'shc6b191ca, 32'shc6b0dec4, 32'shc6b02bc7, 32'shc6af78d3, 32'shc6aec5e7, 
               32'shc6ae1304, 32'shc6ad602a, 32'shc6acad59, 32'shc6abfa91, 32'shc6ab47d2, 32'shc6aa951b, 32'shc6a9e26e, 32'shc6a92fc9, 
               32'shc6a87d2d, 32'shc6a7ca9a, 32'shc6a7180f, 32'shc6a6658e, 32'shc6a5b315, 32'shc6a500a5, 32'shc6a44e3e, 32'shc6a39be0, 
               32'shc6a2e98b, 32'shc6a2373f, 32'shc6a184fb, 32'shc6a0d2c0, 32'shc6a0208f, 32'shc69f6e66, 32'shc69ebc45, 32'shc69e0a2e, 
               32'shc69d5820, 32'shc69ca61a, 32'shc69bf41d, 32'shc69b4229, 32'shc69a903e, 32'shc699de5c, 32'shc6992c83, 32'shc6987ab2, 
               32'shc697c8eb, 32'shc697172c, 32'shc6966576, 32'shc695b3c9, 32'shc6950224, 32'shc6945089, 32'shc6939ef6, 32'shc692ed6d, 
               32'shc6923bec, 32'shc6918a74, 32'shc690d905, 32'shc690279f, 32'shc68f7641, 32'shc68ec4ed, 32'shc68e13a1, 32'shc68d625e, 
               32'shc68cb124, 32'shc68bfff3, 32'shc68b4ecb, 32'shc68a9dac, 32'shc689ec95, 32'shc6893b87, 32'shc6888a83, 32'shc687d987, 
               32'shc6872894, 32'shc68677a9, 32'shc685c6c8, 32'shc68515f0, 32'shc6846520, 32'shc683b459, 32'shc683039b, 32'shc68252e6, 
               32'shc681a23a, 32'shc680f197, 32'shc68040fc, 32'shc67f906b, 32'shc67edfe2, 32'shc67e2f62, 32'shc67d7eeb, 32'shc67cce7d, 
               32'shc67c1e18, 32'shc67b6dbc, 32'shc67abd68, 32'shc67a0d1e, 32'shc6795cdc, 32'shc678aca3, 32'shc677fc73, 32'shc6774c4c, 
               32'shc6769c2e, 32'shc675ec18, 32'shc6753c0c, 32'shc6748c08, 32'shc673dc0d, 32'shc6732c1b, 32'shc6727c32, 32'shc671cc52, 
               32'shc6711c7b, 32'shc6706cad, 32'shc66fbce7, 32'shc66f0d2b, 32'shc66e5d77, 32'shc66dadcc, 32'shc66cfe2a, 32'shc66c4e91, 
               32'shc66b9f01, 32'shc66aef79, 32'shc66a3ffb, 32'shc6699085, 32'shc668e119, 32'shc66831b5, 32'shc667825a, 32'shc666d308, 
               32'shc66623be, 32'shc665747e, 32'shc664c547, 32'shc6641618, 32'shc66366f3, 32'shc662b7d6, 32'shc66208c2, 32'shc66159b7, 
               32'shc660aab5, 32'shc65ffbbc, 32'shc65f4ccb, 32'shc65e9de4, 32'shc65def05, 32'shc65d4030, 32'shc65c9163, 32'shc65be29f, 
               32'shc65b33e4, 32'shc65a8532, 32'shc659d688, 32'shc65927e8, 32'shc6587951, 32'shc657cac2, 32'shc6571c3c, 32'shc6566dc0, 
               32'shc655bf4c, 32'shc65510e1, 32'shc654627f, 32'shc653b426, 32'shc65305d5, 32'shc652578e, 32'shc651a94f, 32'shc650fb1a, 
               32'shc6504ced, 32'shc64f9ec9, 32'shc64ef0ae, 32'shc64e429c, 32'shc64d9493, 32'shc64ce693, 32'shc64c389b, 32'shc64b8aad, 
               32'shc64adcc7, 32'shc64a2eeb, 32'shc6498117, 32'shc648d34c, 32'shc648258a, 32'shc64777d1, 32'shc646ca21, 32'shc6461c7a, 
               32'shc6456edb, 32'shc644c146, 32'shc64413b9, 32'shc6436636, 32'shc642b8bb, 32'shc6420b49, 32'shc6415de0, 32'shc640b080, 
               32'shc6400329, 32'shc63f55db, 32'shc63ea896, 32'shc63dfb59, 32'shc63d4e26, 32'shc63ca0fb, 32'shc63bf3d9, 32'shc63b46c1, 
               32'shc63a99b1, 32'shc639ecaa, 32'shc6393fac, 32'shc63892b7, 32'shc637e5ca, 32'shc63738e7, 32'shc6368c0d, 32'shc635df3b, 
               32'shc6353273, 32'shc63485b3, 32'shc633d8fc, 32'shc6332c4e, 32'shc6327faa, 32'shc631d30e, 32'shc631267a, 32'shc63079f0, 
               32'shc62fcd6f, 32'shc62f20f7, 32'shc62e7487, 32'shc62dc821, 32'shc62d1bc3, 32'shc62c6f6e, 32'shc62bc323, 32'shc62b16e0, 
               32'shc62a6aa6, 32'shc629be75, 32'shc629124d, 32'shc628662e, 32'shc627ba17, 32'shc6270e0a, 32'shc6266206, 32'shc625b60a, 
               32'shc6250a18, 32'shc6245e2e, 32'shc623b24d, 32'shc6230675, 32'shc6225aa6, 32'shc621aee1, 32'shc6210323, 32'shc620576f, 
               32'shc61fabc4, 32'shc61f0022, 32'shc61e5489, 32'shc61da8f8, 32'shc61cfd71, 32'shc61c51f2, 32'shc61ba67d, 32'shc61afb10, 
               32'shc61a4fac, 32'shc619a451, 32'shc618f8ff, 32'shc6184db6, 32'shc617a276, 32'shc616f73f, 32'shc6164c11, 32'shc615a0ec, 
               32'shc614f5cf, 32'shc6144abc, 32'shc6139fb2, 32'shc612f4b0, 32'shc61249b7, 32'shc6119ec8, 32'shc610f3e1, 32'shc6104903, 
               32'shc60f9e2e, 32'shc60ef362, 32'shc60e489f, 32'shc60d9de5, 32'shc60cf334, 32'shc60c488c, 32'shc60b9ded, 32'shc60af357, 
               32'shc60a48c9, 32'shc6099e45, 32'shc608f3c9, 32'shc6084957, 32'shc6079eed, 32'shc606f48c, 32'shc6064a35, 32'shc6059fe6, 
               32'shc604f5a0, 32'shc6044b63, 32'shc603a12f, 32'shc602f704, 32'shc6024ce2, 32'shc601a2c9, 32'shc600f8b9, 32'shc6004eb1, 
               32'shc5ffa4b3, 32'shc5fefabe, 32'shc5fe50d1, 32'shc5fda6ee, 32'shc5fcfd13, 32'shc5fc5342, 32'shc5fba979, 32'shc5faffb9, 
               32'shc5fa5603, 32'shc5f9ac55, 32'shc5f902b0, 32'shc5f85914, 32'shc5f7af81, 32'shc5f705f7, 32'shc5f65c76, 32'shc5f5b2fe, 
               32'shc5f5098f, 32'shc5f46029, 32'shc5f3b6cb, 32'shc5f30d77, 32'shc5f2642c, 32'shc5f1bae9, 32'shc5f111b0, 32'shc5f0687f, 
               32'shc5efbf58, 32'shc5ef1639, 32'shc5ee6d24, 32'shc5edc417, 32'shc5ed1b13, 32'shc5ec7218, 32'shc5ebc927, 32'shc5eb203e, 
               32'shc5ea775e, 32'shc5e9ce87, 32'shc5e925b9, 32'shc5e87cf4, 32'shc5e7d438, 32'shc5e72b85, 32'shc5e682db, 32'shc5e5da3a, 
               32'shc5e531a1, 32'shc5e48912, 32'shc5e3e08c, 32'shc5e3380e, 32'shc5e28f9a, 32'shc5e1e72f, 32'shc5e13ecc, 32'shc5e09673, 
               32'shc5dfee22, 32'shc5df45db, 32'shc5de9d9c, 32'shc5ddf566, 32'shc5dd4d3a, 32'shc5dca516, 32'shc5dbfcfb, 32'shc5db54e9, 
               32'shc5daace1, 32'shc5da04e1, 32'shc5d95cea, 32'shc5d8b4fc, 32'shc5d80d17, 32'shc5d7653b, 32'shc5d6bd68, 32'shc5d6159e, 
               32'shc5d56ddd, 32'shc5d4c625, 32'shc5d41e76, 32'shc5d376d0, 32'shc5d2cf33, 32'shc5d2279e, 32'shc5d18013, 32'shc5d0d891, 
               32'shc5d03118, 32'shc5cf89a7, 32'shc5cee240, 32'shc5ce3ae1, 32'shc5cd938c, 32'shc5ccec40, 32'shc5cc44fc, 32'shc5cb9dc2, 
               32'shc5caf690, 32'shc5ca4f68, 32'shc5c9a848, 32'shc5c90132, 32'shc5c85a24, 32'shc5c7b31f, 32'shc5c70c24, 32'shc5c66531, 
               32'shc5c5be47, 32'shc5c51767, 32'shc5c4708f, 32'shc5c3c9c0, 32'shc5c322fb, 32'shc5c27c3e, 32'shc5c1d58a, 32'shc5c12edf, 
               32'shc5c0883d, 32'shc5bfe1a5, 32'shc5bf3b15, 32'shc5be948e, 32'shc5bdee10, 32'shc5bd479b, 32'shc5bca12f, 32'shc5bbfacc, 
               32'shc5bb5472, 32'shc5baae21, 32'shc5ba07d9, 32'shc5b9619a, 32'shc5b8bb64, 32'shc5b81537, 32'shc5b76f13, 32'shc5b6c8f8, 
               32'shc5b622e6, 32'shc5b57cdd, 32'shc5b4d6dd, 32'shc5b430e6, 32'shc5b38af8, 32'shc5b2e513, 32'shc5b23f37, 32'shc5b19963, 
               32'shc5b0f399, 32'shc5b04dd8, 32'shc5afa820, 32'shc5af0271, 32'shc5ae5ccb, 32'shc5adb72d, 32'shc5ad1199, 32'shc5ac6c0e, 
               32'shc5abc68c, 32'shc5ab2113, 32'shc5aa7ba3, 32'shc5a9d63b, 32'shc5a930dd, 32'shc5a88b88, 32'shc5a7e63c, 32'shc5a740f8, 
               32'shc5a69bbe, 32'shc5a5f68d, 32'shc5a55165, 32'shc5a4ac46, 32'shc5a4072f, 32'shc5a36222, 32'shc5a2bd1e, 32'shc5a21823, 
               32'shc5a17330, 32'shc5a0ce47, 32'shc5a02967, 32'shc59f8490, 32'shc59edfc2, 32'shc59e3afc, 32'shc59d9640, 32'shc59cf18d, 
               32'shc59c4ce3, 32'shc59ba842, 32'shc59b03a9, 32'shc59a5f1a, 32'shc599ba94, 32'shc5991617, 32'shc59871a3, 32'shc597cd38, 
               32'shc59728d5, 32'shc596847c, 32'shc595e02c, 32'shc5953be5, 32'shc59497a7, 32'shc593f372, 32'shc5934f46, 32'shc592ab22, 
               32'shc5920708, 32'shc59162f7, 32'shc590beef, 32'shc5901af0, 32'shc58f76fa, 32'shc58ed30d, 32'shc58e2f29, 32'shc58d8b4e, 
               32'shc58ce77c, 32'shc58c43b3, 32'shc58b9ff3, 32'shc58afc3c, 32'shc58a588e, 32'shc589b4e9, 32'shc589114e, 32'shc5886dbb, 
               32'shc587ca31, 32'shc58726b0, 32'shc5868338, 32'shc585dfc9, 32'shc5853c63, 32'shc5849907, 32'shc583f5b3, 32'shc5835268, 
               32'shc582af26, 32'shc5820bee, 32'shc58168be, 32'shc580c597, 32'shc580227a, 32'shc57f7f65, 32'shc57edc5a, 32'shc57e3957, 
               32'shc57d965d, 32'shc57cf36d, 32'shc57c5085, 32'shc57bada7, 32'shc57b0ad1, 32'shc57a6805, 32'shc579c542, 32'shc5792287, 
               32'shc5787fd6, 32'shc577dd2d, 32'shc5773a8e, 32'shc57697f8, 32'shc575f56b, 32'shc57552e6, 32'shc574b06b, 32'shc5740df9, 
               32'shc5736b90, 32'shc572c930, 32'shc57226d9, 32'shc571848b, 32'shc570e246, 32'shc570400a, 32'shc56f9dd7, 32'shc56efbad, 
               32'shc56e598c, 32'shc56db774, 32'shc56d1565, 32'shc56c735f, 32'shc56bd163, 32'shc56b2f6f, 32'shc56a8d84, 32'shc569eba2, 
               32'shc56949ca, 32'shc568a7fa, 32'shc5680634, 32'shc5676476, 32'shc566c2c2, 32'shc5662116, 32'shc5657f74, 32'shc564ddda, 
               32'shc5643c4a, 32'shc5639ac3, 32'shc562f944, 32'shc56257cf, 32'shc561b663, 32'shc5611500, 32'shc56073a6, 32'shc55fd255, 
               32'shc55f310d, 32'shc55e8fce, 32'shc55dee98, 32'shc55d4d6b, 32'shc55cac47, 32'shc55c0b2c, 32'shc55b6a1a, 32'shc55ac912, 
               32'shc55a2812, 32'shc559871b, 32'shc558e62e, 32'shc5584549, 32'shc557a46e, 32'shc557039b, 32'shc55662d2, 32'shc555c211, 
               32'shc555215a, 32'shc55480ac, 32'shc553e007, 32'shc5533f6b, 32'shc5529ed7, 32'shc551fe4d, 32'shc5515dcc, 32'shc550bd54, 
               32'shc5501ce5, 32'shc54f7c7f, 32'shc54edc23, 32'shc54e3bcf, 32'shc54d9b84, 32'shc54cfb42, 32'shc54c5b0a, 32'shc54bbada, 
               32'shc54b1ab4, 32'shc54a7a96, 32'shc549da82, 32'shc5493a76, 32'shc5489a74, 32'shc547fa7b, 32'shc5475a8b, 32'shc546baa4, 
               32'shc5461ac6, 32'shc5457af1, 32'shc544db25, 32'shc5443b62, 32'shc5439ba8, 32'shc542fbf7, 32'shc5425c4f, 32'shc541bcb1, 
               32'shc5411d1b, 32'shc5407d8e, 32'shc53fde0b, 32'shc53f3e90, 32'shc53e9f1f, 32'shc53dffb7, 32'shc53d6057, 32'shc53cc101, 
               32'shc53c21b4, 32'shc53b8270, 32'shc53ae335, 32'shc53a4403, 32'shc539a4da, 32'shc53905ba, 32'shc53866a4, 32'shc537c796, 
               32'shc5372891, 32'shc5368996, 32'shc535eaa3, 32'shc5354bba, 32'shc534acd9, 32'shc5340e02, 32'shc5336f34, 32'shc532d06f, 
               32'shc53231b3, 32'shc5319300, 32'shc530f456, 32'shc53055b5, 32'shc52fb71d, 32'shc52f188e, 32'shc52e7a09, 32'shc52ddb8c, 
               32'shc52d3d18, 32'shc52c9eae, 32'shc52c004d, 32'shc52b61f4, 32'shc52ac3a5, 32'shc52a255f, 32'shc5298722, 32'shc528e8ee, 
               32'shc5284ac3, 32'shc527aca1, 32'shc5270e88, 32'shc5267078, 32'shc525d272, 32'shc5253474, 32'shc5249680, 32'shc523f894, 
               32'shc5235ab2, 32'shc522bcd9, 32'shc5221f08, 32'shc5218141, 32'shc520e383, 32'shc52045ce, 32'shc51fa822, 32'shc51f0a7f, 
               32'shc51e6ce6, 32'shc51dcf55, 32'shc51d31ce, 32'shc51c944f, 32'shc51bf6da, 32'shc51b596d, 32'shc51abc0a, 32'shc51a1eb0, 
               32'shc519815f, 32'shc518e417, 32'shc51846d8, 32'shc517a9a2, 32'shc5170c75, 32'shc5166f52, 32'shc515d237, 32'shc5153526, 
               32'shc514981d, 32'shc513fb1e, 32'shc5135e28, 32'shc512c13b, 32'shc5122457, 32'shc511877c, 32'shc510eaaa, 32'shc5104de1, 
               32'shc50fb121, 32'shc50f146b, 32'shc50e77bd, 32'shc50ddb19, 32'shc50d3e7d, 32'shc50ca1eb, 32'shc50c0562, 32'shc50b68e2, 
               32'shc50acc6b, 32'shc50a2ffd, 32'shc5099398, 32'shc508f73d, 32'shc5085aea, 32'shc507bea1, 32'shc5072260, 32'shc5068629, 
               32'shc505e9fb, 32'shc5054dd5, 32'shc504b1b9, 32'shc50415a6, 32'shc503799d, 32'shc502dd9c, 32'shc50241a4, 32'shc501a5b6, 
               32'shc50109d0, 32'shc5006df4, 32'shc4ffd221, 32'shc4ff3656, 32'shc4fe9a95, 32'shc4fdfedd, 32'shc4fd632f, 32'shc4fcc789, 
               32'shc4fc2bec, 32'shc4fb9059, 32'shc4faf4ce, 32'shc4fa594d, 32'shc4f9bdd4, 32'shc4f92265, 32'shc4f886ff, 32'shc4f7eba2, 
               32'shc4f7504e, 32'shc4f6b504, 32'shc4f619c2, 32'shc4f57e8a, 32'shc4f4e35a, 32'shc4f44834, 32'shc4f3ad17, 32'shc4f31202, 
               32'shc4f276f7, 32'shc4f1dbf6, 32'shc4f140fd, 32'shc4f0a60d, 32'shc4f00b27, 32'shc4ef7049, 32'shc4eed575, 32'shc4ee3aa9, 
               32'shc4ed9fe7, 32'shc4ed052e, 32'shc4ec6a7e, 32'shc4ebcfd8, 32'shc4eb353a, 32'shc4ea9aa5, 32'shc4ea001a, 32'shc4e96597, 
               32'shc4e8cb1e, 32'shc4e830ae, 32'shc4e79647, 32'shc4e6fbe9, 32'shc4e66194, 32'shc4e5c749, 32'shc4e52d06, 32'shc4e492cd, 
               32'shc4e3f89c, 32'shc4e35e75, 32'shc4e2c457, 32'shc4e22a42, 32'shc4e19036, 32'shc4e0f633, 32'shc4e05c3a, 32'shc4dfc249, 
               32'shc4df2862, 32'shc4de8e83, 32'shc4ddf4ae, 32'shc4dd5ae2, 32'shc4dcc11f, 32'shc4dc2765, 32'shc4db8db5, 32'shc4daf40d, 
               32'shc4da5a6f, 32'shc4d9c0d9, 32'shc4d9274d, 32'shc4d88dca, 32'shc4d7f450, 32'shc4d75adf, 32'shc4d6c177, 32'shc4d62819, 
               32'shc4d58ec3, 32'shc4d4f577, 32'shc4d45c34, 32'shc4d3c2fa, 32'shc4d329c9, 32'shc4d290a1, 32'shc4d1f782, 32'shc4d15e6d, 
               32'shc4d0c560, 32'shc4d02c5d, 32'shc4cf9363, 32'shc4cefa71, 32'shc4ce6189, 32'shc4cdc8ab, 32'shc4cd2fd5, 32'shc4cc9708, 
               32'shc4cbfe45, 32'shc4cb658b, 32'shc4caccd9, 32'shc4ca3431, 32'shc4c99b92, 32'shc4c902fd, 32'shc4c86a70, 32'shc4c7d1ec, 
               32'shc4c73972, 32'shc4c6a101, 32'shc4c60899, 32'shc4c5703a, 32'shc4c4d7e4, 32'shc4c43f97, 32'shc4c3a753, 32'shc4c30f19, 
               32'shc4c276e8, 32'shc4c1dec0, 32'shc4c146a0, 32'shc4c0ae8b, 32'shc4c0167e, 32'shc4bf7e7a, 32'shc4bee680, 32'shc4be4e8e, 
               32'shc4bdb6a6, 32'shc4bd1ec7, 32'shc4bc86f1, 32'shc4bbef24, 32'shc4bb5760, 32'shc4babfa6, 32'shc4ba27f5, 32'shc4b9904c, 
               32'shc4b8f8ad, 32'shc4b86117, 32'shc4b7c98a, 32'shc4b73207, 32'shc4b69a8c, 32'shc4b6031b, 32'shc4b56bb3, 32'shc4b4d453, 
               32'shc4b43cfd, 32'shc4b3a5b1, 32'shc4b30e6d, 32'shc4b27732, 32'shc4b1e001, 32'shc4b148d9, 32'shc4b0b1ba, 32'shc4b01aa4, 
               32'shc4af8397, 32'shc4aeec93, 32'shc4ae5599, 32'shc4adbea7, 32'shc4ad27bf, 32'shc4ac90e0, 32'shc4abfa0a, 32'shc4ab633d, 
               32'shc4aacc7a, 32'shc4aa35bf, 32'shc4a99f0e, 32'shc4a90866, 32'shc4a871c7, 32'shc4a7db31, 32'shc4a744a4, 32'shc4a6ae21, 
               32'shc4a617a6, 32'shc4a58135, 32'shc4a4eacd, 32'shc4a4546e, 32'shc4a3be18, 32'shc4a327cb, 32'shc4a29188, 32'shc4a1fb4e, 
               32'shc4a1651c, 32'shc4a0cef4, 32'shc4a038d6, 32'shc49fa2c0, 32'shc49f0cb3, 32'shc49e76b0, 32'shc49de0b6, 32'shc49d4ac5, 
               32'shc49cb4dd, 32'shc49c1efe, 32'shc49b8928, 32'shc49af35c, 32'shc49a5d98, 32'shc499c7de, 32'shc499322d, 32'shc4989c86, 
               32'shc49806e7, 32'shc4977151, 32'shc496dbc5, 32'shc4964642, 32'shc495b0c8, 32'shc4951b57, 32'shc49485ef, 32'shc493f091, 
               32'shc4935b3c, 32'shc492c5ef, 32'shc49230ac, 32'shc4919b72, 32'shc4910642, 32'shc490711a, 32'shc48fdbfc, 32'shc48f46e7, 
               32'shc48eb1db, 32'shc48e1cd8, 32'shc48d87de, 32'shc48cf2ee, 32'shc48c5e06, 32'shc48bc928, 32'shc48b3453, 32'shc48a9f87, 
               32'shc48a0ac4, 32'shc489760b, 32'shc488e15b, 32'shc4884cb3, 32'shc487b815, 32'shc4872381, 32'shc4868ef5, 32'shc485fa72, 
               32'shc48565f9, 32'shc484d189, 32'shc4843d22, 32'shc483a8c4, 32'shc4831470, 32'shc4828024, 32'shc481ebe2, 32'shc48157a9, 
               32'shc480c379, 32'shc4802f52, 32'shc47f9b34, 32'shc47f0720, 32'shc47e7315, 32'shc47ddf13, 32'shc47d4b1a, 32'shc47cb72a, 
               32'shc47c2344, 32'shc47b8f66, 32'shc47afb92, 32'shc47a67c7, 32'shc479d405, 32'shc479404d, 32'shc478ac9d, 32'shc47818f7, 
               32'shc477855a, 32'shc476f1c6, 32'shc4765e3b, 32'shc475caba, 32'shc4753741, 32'shc474a3d2, 32'shc474106c, 32'shc4737d10, 
               32'shc472e9bc, 32'shc4725671, 32'shc471c330, 32'shc4712ff8, 32'shc4709cc9, 32'shc47009a4, 32'shc46f7687, 32'shc46ee374, 
               32'shc46e5069, 32'shc46dbd69, 32'shc46d2a71, 32'shc46c9782, 32'shc46c049d, 32'shc46b71c1, 32'shc46adeee, 32'shc46a4c24, 
               32'shc469b963, 32'shc46926ac, 32'shc46893fd, 32'shc4680158, 32'shc4676ebc, 32'shc466dc2a, 32'shc46649a0, 32'shc465b720, 
               32'shc46524a9, 32'shc464923b, 32'shc463ffd6, 32'shc4636d7a, 32'shc462db28, 32'shc46248df, 32'shc461b69f, 32'shc4612468, 
               32'shc460923b, 32'shc4600016, 32'shc45f6dfb, 32'shc45edbe9, 32'shc45e49e0, 32'shc45db7e1, 32'shc45d25ea, 32'shc45c93fd, 
               32'shc45c0219, 32'shc45b703e, 32'shc45ade6c, 32'shc45a4ca4, 32'shc459bae5, 32'shc459292f, 32'shc4589782, 32'shc45805de, 
               32'shc4577444, 32'shc456e2b3, 32'shc456512b, 32'shc455bfac, 32'shc4552e36, 32'shc4549cca, 32'shc4540b67, 32'shc4537a0d, 
               32'shc452e8bc, 32'shc4525774, 32'shc451c636, 32'shc4513500, 32'shc450a3d4, 32'shc45012b2, 32'shc44f8198, 32'shc44ef088, 
               32'shc44e5f80, 32'shc44dce82, 32'shc44d3d8e, 32'shc44caca2, 32'shc44c1bc0, 32'shc44b8ae7, 32'shc44afa17, 32'shc44a6950, 
               32'shc449d892, 32'shc44947de, 32'shc448b733, 32'shc4482691, 32'shc44795f8, 32'shc4470569, 32'shc44674e3, 32'shc445e466, 
               32'shc44553f2, 32'shc444c387, 32'shc4443326, 32'shc443a2cd, 32'shc443127e, 32'shc4428239, 32'shc441f1fc, 32'shc44161c9, 
               32'shc440d19e, 32'shc440417d, 32'shc43fb166, 32'shc43f2157, 32'shc43e9152, 32'shc43e0156, 32'shc43d7163, 32'shc43ce179, 
               32'shc43c5199, 32'shc43bc1c2, 32'shc43b31f4, 32'shc43aa22f, 32'shc43a1273, 32'shc43982c1, 32'shc438f318, 32'shc4386378, 
               32'shc437d3e1, 32'shc4374454, 32'shc436b4cf, 32'shc4362554, 32'shc43595e3, 32'shc435067a, 32'shc434771b, 32'shc433e7c4, 
               32'shc4335877, 32'shc432c934, 32'shc43239f9, 32'shc431aac8, 32'shc4311ba0, 32'shc4308c81, 32'shc42ffd6b, 32'shc42f6e5f, 
               32'shc42edf5c, 32'shc42e5062, 32'shc42dc171, 32'shc42d328a, 32'shc42ca3ac, 32'shc42c14d7, 32'shc42b860b, 32'shc42af748, 
               32'shc42a688f, 32'shc429d9df, 32'shc4294b38, 32'shc428bc9a, 32'shc4282e06, 32'shc4279f7b, 32'shc42710f9, 32'shc4268280, 
               32'shc425f410, 32'shc42565aa, 32'shc424d74d, 32'shc42448f9, 32'shc423baae, 32'shc4232c6d, 32'shc4229e35, 32'shc4221006, 
               32'shc42181e0, 32'shc420f3c4, 32'shc42065b1, 32'shc41fd7a7, 32'shc41f49a6, 32'shc41ebbaf, 32'shc41e2dc0, 32'shc41d9fdb, 
               32'shc41d11ff, 32'shc41c842d, 32'shc41bf664, 32'shc41b68a3, 32'shc41adaed, 32'shc41a4d3f, 32'shc419bf9b, 32'shc41931ff, 
               32'shc418a46d, 32'shc41816e5, 32'shc4178965, 32'shc416fbef, 32'shc4166e82, 32'shc415e11f, 32'shc41553c4, 32'shc414c673, 
               32'shc414392b, 32'shc413abec, 32'shc4131eb7, 32'shc412918a, 32'shc4120467, 32'shc411774d, 32'shc410ea3d, 32'shc4105d36, 
               32'shc40fd037, 32'shc40f4343, 32'shc40eb657, 32'shc40e2975, 32'shc40d9c9c, 32'shc40d0fcc, 32'shc40c8305, 32'shc40bf648, 
               32'shc40b6994, 32'shc40adce9, 32'shc40a5047, 32'shc409c3af, 32'shc4093720, 32'shc408aa9a, 32'shc4081e1d, 32'shc40791aa, 
               32'shc4070540, 32'shc40678df, 32'shc405ec87, 32'shc4056039, 32'shc404d3f4, 32'shc40447b8, 32'shc403bb85, 32'shc4032f5c, 
               32'shc402a33c, 32'shc4021725, 32'shc4018b17, 32'shc400ff13, 32'shc4007318, 32'shc3ffe726, 32'shc3ff5b3d, 32'shc3fecf5e, 
               32'shc3fe4388, 32'shc3fdb7bb, 32'shc3fd2bf7, 32'shc3fca03d, 32'shc3fc148c, 32'shc3fb88e4, 32'shc3fafd45, 32'shc3fa71b0, 
               32'shc3f9e624, 32'shc3f95aa1, 32'shc3f8cf27, 32'shc3f843b7, 32'shc3f7b850, 32'shc3f72cf2, 32'shc3f6a19e, 32'shc3f61652, 
               32'shc3f58b10, 32'shc3f4ffd8, 32'shc3f474a8, 32'shc3f3e982, 32'shc3f35e65, 32'shc3f2d351, 32'shc3f24847, 32'shc3f1bd46, 
               32'shc3f1324e, 32'shc3f0a75f, 32'shc3f01c7a, 32'shc3ef919d, 32'shc3ef06cb, 32'shc3ee7c01, 32'shc3edf141, 32'shc3ed6689, 
               32'shc3ecdbdc, 32'shc3ec5137, 32'shc3ebc69c, 32'shc3eb3c0a, 32'shc3eab181, 32'shc3ea2701, 32'shc3e99c8b, 32'shc3e9121e, 
               32'shc3e887bb, 32'shc3e7fd60, 32'shc3e7730f, 32'shc3e6e8c7, 32'shc3e65e88, 32'shc3e5d453, 32'shc3e54a27, 32'shc3e4c004, 
               32'shc3e435ea, 32'shc3e3abda, 32'shc3e321d3, 32'shc3e297d5, 32'shc3e20de1, 32'shc3e183f6, 32'shc3e0fa14, 32'shc3e0703b, 
               32'shc3dfe66c, 32'shc3df5ca6, 32'shc3ded2e9, 32'shc3de4935, 32'shc3ddbf8b, 32'shc3dd35ea, 32'shc3dcac52, 32'shc3dc22c4, 
               32'shc3db993e, 32'shc3db0fc2, 32'shc3da8650, 32'shc3d9fce6, 32'shc3d97386, 32'shc3d8ea2f, 32'shc3d860e2, 32'shc3d7d79d, 
               32'shc3d74e62, 32'shc3d6c531, 32'shc3d63c08, 32'shc3d5b2e9, 32'shc3d529d3, 32'shc3d4a0c7, 32'shc3d417c3, 32'shc3d38ec9, 
               32'shc3d305d8, 32'shc3d27cf1, 32'shc3d1f413, 32'shc3d16b3e, 32'shc3d0e272, 32'shc3d059b0, 32'shc3cfd0f7, 32'shc3cf4847, 
               32'shc3cebfa0, 32'shc3ce3703, 32'shc3cdae6f, 32'shc3cd25e4, 32'shc3cc9d63, 32'shc3cc14eb, 32'shc3cb8c7c, 32'shc3cb0416, 
               32'shc3ca7bba, 32'shc3c9f367, 32'shc3c96b1e, 32'shc3c8e2dd, 32'shc3c85aa6, 32'shc3c7d278, 32'shc3c74a54, 32'shc3c6c238, 
               32'shc3c63a26, 32'shc3c5b21e, 32'shc3c52a1e, 32'shc3c4a228, 32'shc3c41a3b, 32'shc3c39258, 32'shc3c30a7e, 32'shc3c282ad, 
               32'shc3c1fae5, 32'shc3c17327, 32'shc3c0eb71, 32'shc3c063c6, 32'shc3bfdc23, 32'shc3bf548a, 32'shc3beccfa, 32'shc3be4573, 
               32'shc3bdbdf6, 32'shc3bd3682, 32'shc3bcaf17, 32'shc3bc27b6, 32'shc3bba05e, 32'shc3bb190f, 32'shc3ba91c9, 32'shc3ba0a8d, 
               32'shc3b9835a, 32'shc3b8fc30, 32'shc3b87510, 32'shc3b7edf9, 32'shc3b766eb, 32'shc3b6dfe6, 32'shc3b658eb, 32'shc3b5d1f9, 
               32'shc3b54b11, 32'shc3b4c431, 32'shc3b43d5b, 32'shc3b3b68f, 32'shc3b32fcb, 32'shc3b2a911, 32'shc3b22260, 32'shc3b19bb9, 
               32'shc3b1151b, 32'shc3b08e86, 32'shc3b007fa, 32'shc3af8178, 32'shc3aefaff, 32'shc3ae748f, 32'shc3adee28, 32'shc3ad67cb, 
               32'shc3ace178, 32'shc3ac5b2d, 32'shc3abd4ec, 32'shc3ab4eb4, 32'shc3aac885, 32'shc3aa4260, 32'shc3a9bc44, 32'shc3a93631, 
               32'shc3a8b028, 32'shc3a82a28, 32'shc3a7a431, 32'shc3a71e44, 32'shc3a6985f, 32'shc3a61285, 32'shc3a58cb3, 32'shc3a506eb, 
               32'shc3a4812c, 32'shc3a3fb76, 32'shc3a375ca, 32'shc3a2f027, 32'shc3a26a8d, 32'shc3a1e4fd, 32'shc3a15f76, 32'shc3a0d9f8, 
               32'shc3a05484, 32'shc39fcf18, 32'shc39f49b7, 32'shc39ec45e, 32'shc39e3f0f, 32'shc39db9c9, 32'shc39d348c, 32'shc39caf59, 
               32'shc39c2a2f, 32'shc39ba50e, 32'shc39b1ff7, 32'shc39a9ae9, 32'shc39a15e4, 32'shc39990e9, 32'shc3990bf7, 32'shc398870e, 
               32'shc398022f, 32'shc3977d59, 32'shc396f88c, 32'shc39673c8, 32'shc395ef0e, 32'shc3956a5d, 32'shc394e5b6, 32'shc3946117, 
               32'shc393dc82, 32'shc39357f7, 32'shc392d375, 32'shc3924efc, 32'shc391ca8c, 32'shc3914626, 32'shc390c1c9, 32'shc3903d75, 
               32'shc38fb92a, 32'shc38f34e9, 32'shc38eb0b2, 32'shc38e2c83, 32'shc38da85e, 32'shc38d2442, 32'shc38ca030, 32'shc38c1c27, 
               32'shc38b9827, 32'shc38b1431, 32'shc38a9043, 32'shc38a0c60, 32'shc3898885, 32'shc38904b4, 32'shc38880ec, 32'shc387fd2e, 
               32'shc3877978, 32'shc386f5cc, 32'shc386722a, 32'shc385ee91, 32'shc3856b01, 32'shc384e77a, 32'shc38463fd, 32'shc383e089, 
               32'shc3835d1e, 32'shc382d9bd, 32'shc3825665, 32'shc381d317, 32'shc3814fd1, 32'shc380cc95, 32'shc3804963, 32'shc37fc639, 
               32'shc37f4319, 32'shc37ec003, 32'shc37e3cf6, 32'shc37db9f2, 32'shc37d36f7, 32'shc37cb406, 32'shc37c311e, 32'shc37bae3f, 
               32'shc37b2b6a, 32'shc37aa89e, 32'shc37a25db, 32'shc379a322, 32'shc3792072, 32'shc3789dcb, 32'shc3781b2e, 32'shc377989a, 
               32'shc377160f, 32'shc376938e, 32'shc3761116, 32'shc3758ea7, 32'shc3750c42, 32'shc37489e6, 32'shc3740793, 32'shc373854a, 
               32'shc373030a, 32'shc37280d3, 32'shc371fea6, 32'shc3717c82, 32'shc370fa68, 32'shc3707856, 32'shc36ff64e, 32'shc36f7450, 
               32'shc36ef25b, 32'shc36e706f, 32'shc36dee8c, 32'shc36d6cb3, 32'shc36ceae3, 32'shc36c691d, 32'shc36be75f, 32'shc36b65ab, 
               32'shc36ae401, 32'shc36a6260, 32'shc369e0c8, 32'shc3695f3a, 32'shc368ddb4, 32'shc3685c39, 32'shc367dac6, 32'shc367595d, 
               32'shc366d7fd, 32'shc36656a7, 32'shc365d55a, 32'shc3655416, 32'shc364d2dc, 32'shc36451ab, 32'shc363d083, 32'shc3634f65, 
               32'shc362ce50, 32'shc3624d44, 32'shc361cc42, 32'shc3614b49, 32'shc360ca59, 32'shc3604973, 32'shc35fc896, 32'shc35f47c2, 
               32'shc35ec6f8, 32'shc35e4637, 32'shc35dc580, 32'shc35d44d2, 32'shc35cc42d, 32'shc35c4391, 32'shc35bc2ff, 32'shc35b4277, 
               32'shc35ac1f7, 32'shc35a4181, 32'shc359c114, 32'shc35940b1, 32'shc358c057, 32'shc3584006, 32'shc357bfbf, 32'shc3573f81, 
               32'shc356bf4d, 32'shc3563f21, 32'shc355bf00, 32'shc3553ee7, 32'shc354bed8, 32'shc3543ed2, 32'shc353bed6, 32'shc3533ee3, 
               32'shc352bef9, 32'shc3523f18, 32'shc351bf41, 32'shc3513f74, 32'shc350bfaf, 32'shc3503ff5, 32'shc34fc043, 32'shc34f409b, 
               32'shc34ec0fc, 32'shc34e4166, 32'shc34dc1da, 32'shc34d4257, 32'shc34cc2de, 32'shc34c436e, 32'shc34bc407, 32'shc34b44aa, 
               32'shc34ac556, 32'shc34a460b, 32'shc349c6ca, 32'shc3494792, 32'shc348c864, 32'shc348493f, 32'shc347ca23, 32'shc3474b10, 
               32'shc346cc07, 32'shc3464d07, 32'shc345ce11, 32'shc3454f24, 32'shc344d041, 32'shc3445166, 32'shc343d295, 32'shc34353ce, 
               32'shc342d510, 32'shc342565b, 32'shc341d7b0, 32'shc341590e, 32'shc340da75, 32'shc3405be6, 32'shc33fdd60, 32'shc33f5ee3, 
               32'shc33ee070, 32'shc33e6206, 32'shc33de3a5, 32'shc33d654e, 32'shc33ce701, 32'shc33c68bc, 32'shc33bea81, 32'shc33b6c50, 
               32'shc33aee27, 32'shc33a7009, 32'shc339f1f3, 32'shc33973e7, 32'shc338f5e4, 32'shc33877eb, 32'shc337f9fb, 32'shc3377c14, 
               32'shc336fe37, 32'shc3368063, 32'shc3360298, 32'shc33584d7, 32'shc3350720, 32'shc3348971, 32'shc3340bcc, 32'shc3338e30, 
               32'shc333109e, 32'shc3329315, 32'shc3321596, 32'shc3319820, 32'shc3311ab3, 32'shc3309d50, 32'shc3301ff5, 32'shc32fa2a5, 
               32'shc32f255e, 32'shc32ea820, 32'shc32e2aeb, 32'shc32dadc0, 32'shc32d309e, 32'shc32cb386, 32'shc32c3677, 32'shc32bb971, 
               32'shc32b3c75, 32'shc32abf82, 32'shc32a4299, 32'shc329c5b9, 32'shc32948e2, 32'shc328cc15, 32'shc3284f51, 32'shc327d296, 
               32'shc32755e5, 32'shc326d93e, 32'shc3265c9f, 32'shc325e00a, 32'shc325637f, 32'shc324e6fc, 32'shc3246a83, 32'shc323ee14, 
               32'shc32371ae, 32'shc322f551, 32'shc32278fe, 32'shc321fcb4, 32'shc3218073, 32'shc321043c, 32'shc320880e, 32'shc3200bea, 
               32'shc31f8fcf, 32'shc31f13bd, 32'shc31e97b5, 32'shc31e1bb6, 32'shc31d9fc1, 32'shc31d23d5, 32'shc31ca7f2, 32'shc31c2c19, 
               32'shc31bb049, 32'shc31b3483, 32'shc31ab8c6, 32'shc31a3d12, 32'shc319c168, 32'shc31945c7, 32'shc318ca2f, 32'shc3184ea1, 
               32'shc317d31c, 32'shc31757a1, 32'shc316dc2f, 32'shc31660c6, 32'shc315e567, 32'shc3156a11, 32'shc314eec5, 32'shc3147382, 
               32'shc313f848, 32'shc3137d18, 32'shc31301f1, 32'shc31286d4, 32'shc3120bc0, 32'shc31190b5, 32'shc31115b4, 32'shc3109abc, 
               32'shc3101fce, 32'shc30fa4e9, 32'shc30f2a0d, 32'shc30eaf3b, 32'shc30e3472, 32'shc30db9b3, 32'shc30d3efd, 32'shc30cc450, 
               32'shc30c49ad, 32'shc30bcf13, 32'shc30b5482, 32'shc30ad9fb, 32'shc30a5f7e, 32'shc309e509, 32'shc3096a9f, 32'shc308f03d, 
               32'shc30875e5, 32'shc307fb97, 32'shc3078151, 32'shc3070715, 32'shc3068ce3, 32'shc30612ba, 32'shc305989a, 32'shc3051e84, 
               32'shc304a477, 32'shc3042a74, 32'shc303b07a, 32'shc3033689, 32'shc302bca2, 32'shc30242c4, 32'shc301c8f0, 32'shc3014f25, 
               32'shc300d563, 32'shc3005bab, 32'shc2ffe1fc, 32'shc2ff6857, 32'shc2feeebb, 32'shc2fe7529, 32'shc2fdfb9f, 32'shc2fd8220, 
               32'shc2fd08a9, 32'shc2fc8f3c, 32'shc2fc15d9, 32'shc2fb9c7f, 32'shc2fb232e, 32'shc2faa9e7, 32'shc2fa30a9, 32'shc2f9b775, 
               32'shc2f93e4a, 32'shc2f8c528, 32'shc2f84c10, 32'shc2f7d301, 32'shc2f759fc, 32'shc2f6e100, 32'shc2f6680d, 32'shc2f5ef24, 
               32'shc2f57644, 32'shc2f4fd6e, 32'shc2f484a1, 32'shc2f40bdd, 32'shc2f39323, 32'shc2f31a73, 32'shc2f2a1cb, 32'shc2f2292e, 
               32'shc2f1b099, 32'shc2f1380e, 32'shc2f0bf8c, 32'shc2f04714, 32'shc2efcea6, 32'shc2ef5640, 32'shc2eedde4, 32'shc2ee6592, 
               32'shc2eded49, 32'shc2ed7509, 32'shc2ecfcd3, 32'shc2ec84a6, 32'shc2ec0c82, 32'shc2eb9468, 32'shc2eb1c58, 32'shc2eaa451, 
               32'shc2ea2c53, 32'shc2e9b45f, 32'shc2e93c74, 32'shc2e8c492, 32'shc2e84cba, 32'shc2e7d4ec, 32'shc2e75d26, 32'shc2e6e56b, 
               32'shc2e66db8, 32'shc2e5f60f, 32'shc2e57e70, 32'shc2e506da, 32'shc2e48f4d, 32'shc2e417ca, 32'shc2e3a050, 32'shc2e328df, 
               32'shc2e2b178, 32'shc2e23a1b, 32'shc2e1c2c7, 32'shc2e14b7c, 32'shc2e0d43b, 32'shc2e05d03, 32'shc2dfe5d4, 32'shc2df6eaf, 
               32'shc2def794, 32'shc2de8082, 32'shc2de0979, 32'shc2dd927a, 32'shc2dd1b84, 32'shc2dca497, 32'shc2dc2db4, 32'shc2dbb6db, 
               32'shc2db400a, 32'shc2dac944, 32'shc2da5286, 32'shc2d9dbd3, 32'shc2d96528, 32'shc2d8ee87, 32'shc2d877f0, 32'shc2d80161, 
               32'shc2d78add, 32'shc2d71461, 32'shc2d69df0, 32'shc2d62787, 32'shc2d5b128, 32'shc2d53ad3, 32'shc2d4c486, 32'shc2d44e44, 
               32'shc2d3d80a, 32'shc2d361db, 32'shc2d2ebb4, 32'shc2d27597, 32'shc2d1ff84, 32'shc2d1897a, 32'shc2d11379, 32'shc2d09d82, 
               32'shc2d02794, 32'shc2cfb1b0, 32'shc2cf3bd5, 32'shc2cec603, 32'shc2ce503b, 32'shc2cdda7d, 32'shc2cd64c7, 32'shc2ccef1c, 
               32'shc2cc7979, 32'shc2cc03e1, 32'shc2cb8e51, 32'shc2cb18cb, 32'shc2caa34f, 32'shc2ca2ddc, 32'shc2c9b872, 32'shc2c94312, 
               32'shc2c8cdbb, 32'shc2c8586e, 32'shc2c7e32a, 32'shc2c76def, 32'shc2c6f8be, 32'shc2c68397, 32'shc2c60e78, 32'shc2c59964, 
               32'shc2c52459, 32'shc2c4af57, 32'shc2c43a5e, 32'shc2c3c56f, 32'shc2c3508a, 32'shc2c2dbae, 32'shc2c266db, 32'shc2c1f212, 
               32'shc2c17d52, 32'shc2c1089c, 32'shc2c093ef, 32'shc2c01f4c, 32'shc2bfaab2, 32'shc2bf3622, 32'shc2bec19b, 32'shc2be4d1d, 
               32'shc2bdd8a9, 32'shc2bd643e, 32'shc2bcefdd, 32'shc2bc7b85, 32'shc2bc0737, 32'shc2bb92f2, 32'shc2bb1eb6, 32'shc2baaa84, 
               32'shc2ba365c, 32'shc2b9c23d, 32'shc2b94e27, 32'shc2b8da1b, 32'shc2b86618, 32'shc2b7f21f, 32'shc2b77e2f, 32'shc2b70a49, 
               32'shc2b6966c, 32'shc2b62298, 32'shc2b5aece, 32'shc2b53b0d, 32'shc2b4c756, 32'shc2b453a9, 32'shc2b3e004, 32'shc2b36c6a, 
               32'shc2b2f8d8, 32'shc2b28550, 32'shc2b211d2, 32'shc2b19e5d, 32'shc2b12af1, 32'shc2b0b78f, 32'shc2b04437, 32'shc2afd0e8, 
               32'shc2af5da2, 32'shc2aeea66, 32'shc2ae7733, 32'shc2ae0409, 32'shc2ad90ea, 32'shc2ad1dd3, 32'shc2acaac6, 32'shc2ac37c3, 
               32'shc2abc4c9, 32'shc2ab51d8, 32'shc2aadef1, 32'shc2aa6c13, 32'shc2a9f93f, 32'shc2a98674, 32'shc2a913b3, 32'shc2a8a0fb, 
               32'shc2a82e4d, 32'shc2a7bba8, 32'shc2a7490c, 32'shc2a6d67a, 32'shc2a663f2, 32'shc2a5f173, 32'shc2a57efd, 32'shc2a50c91, 
               32'shc2a49a2e, 32'shc2a427d5, 32'shc2a3b585, 32'shc2a3433f, 32'shc2a2d102, 32'shc2a25ecf, 32'shc2a1eca5, 32'shc2a17a84, 
               32'shc2a1086d, 32'shc2a09660, 32'shc2a0245c, 32'shc29fb261, 32'shc29f4070, 32'shc29ece88, 32'shc29e5caa, 32'shc29dead5, 
               32'shc29d790a, 32'shc29d0748, 32'shc29c9590, 32'shc29c23e1, 32'shc29bb23c, 32'shc29b40a0, 32'shc29acf0d, 32'shc29a5d84, 
               32'shc299ec05, 32'shc2997a8f, 32'shc2990922, 32'shc29897bf, 32'shc2982665, 32'shc297b515, 32'shc29743ce, 32'shc296d291, 
               32'shc296615d, 32'shc295f033, 32'shc2957f12, 32'shc2950dfb, 32'shc2949ced, 32'shc2942be8, 32'shc293baed, 32'shc29349fc, 
               32'shc292d914, 32'shc2926835, 32'shc291f760, 32'shc2918695, 32'shc29115d3, 32'shc290a51a, 32'shc290346b, 32'shc28fc3c5, 
               32'shc28f5329, 32'shc28ee296, 32'shc28e720d, 32'shc28e018d, 32'shc28d9117, 32'shc28d20aa, 32'shc28cb047, 32'shc28c3fed, 
               32'shc28bcf9c, 32'shc28b5f55, 32'shc28aef18, 32'shc28a7ee4, 32'shc28a0eb9, 32'shc2899e98, 32'shc2892e81, 32'shc288be73, 
               32'shc2884e6e, 32'shc287de73, 32'shc2876e82, 32'shc286fe99, 32'shc2868ebb, 32'shc2861ee6, 32'shc285af1a, 32'shc2853f58, 
               32'shc284cf9f, 32'shc2845ff0, 32'shc283f04a, 32'shc28380ad, 32'shc283111b, 32'shc282a191, 32'shc2823211, 32'shc281c29b, 
               32'shc281532e, 32'shc280e3cb, 32'shc2807471, 32'shc2800520, 32'shc27f95d9, 32'shc27f269c, 32'shc27eb768, 32'shc27e483d, 
               32'shc27dd91c, 32'shc27d6a05, 32'shc27cfaf7, 32'shc27c8bf2, 32'shc27c1cf7, 32'shc27bae06, 32'shc27b3f1e, 32'shc27ad03f, 
               32'shc27a616a, 32'shc279f29e, 32'shc27983dc, 32'shc2791523, 32'shc278a674, 32'shc27837ce, 32'shc277c932, 32'shc2775aa0, 
               32'shc276ec16, 32'shc2767d97, 32'shc2760f20, 32'shc275a0b4, 32'shc2753250, 32'shc274c3f7, 32'shc27455a6, 32'shc273e760, 
               32'shc2737922, 32'shc2730aee, 32'shc2729cc4, 32'shc2722ea3, 32'shc271c08c, 32'shc271527e, 32'shc270e47a, 32'shc270767f, 
               32'shc270088e, 32'shc26f9aa6, 32'shc26f2cc7, 32'shc26ebef2, 32'shc26e5127, 32'shc26de365, 32'shc26d75ad, 32'shc26d07fe, 
               32'shc26c9a58, 32'shc26c2cbd, 32'shc26bbf2a, 32'shc26b51a1, 32'shc26ae422, 32'shc26a76ac, 32'shc26a093f, 32'shc2699bdd, 
               32'shc2692e83, 32'shc268c133, 32'shc26853ed, 32'shc267e6b0, 32'shc267797c, 32'shc2670c52, 32'shc2669f32, 32'shc266321b, 
               32'shc265c50e, 32'shc265580a, 32'shc264eb0f, 32'shc2647e1e, 32'shc2641137, 32'shc263a459, 32'shc2633785, 32'shc262caba, 
               32'shc2625df8, 32'shc261f140, 32'shc2618492, 32'shc26117ed, 32'shc260ab51, 32'shc2603ec0, 32'shc25fd237, 32'shc25f65b8, 
               32'shc25ef943, 32'shc25e8cd7, 32'shc25e2074, 32'shc25db41c, 32'shc25d47cc, 32'shc25cdb86, 32'shc25c6f4a, 32'shc25c0317, 
               32'shc25b96ee, 32'shc25b2ace, 32'shc25abeb7, 32'shc25a52ab, 32'shc259e6a7, 32'shc2597aad, 32'shc2590ebd, 32'shc258a2d6, 
               32'shc25836f9, 32'shc257cb25, 32'shc2575f5b, 32'shc256f39a, 32'shc25687e3, 32'shc2561c35, 32'shc255b091, 32'shc25544f6, 
               32'shc254d965, 32'shc2546ddd, 32'shc254025f, 32'shc25396ea, 32'shc2532b7f, 32'shc252c01d, 32'shc25254c5, 32'shc251e976, 
               32'shc2517e31, 32'shc25112f6, 32'shc250a7c3, 32'shc2503c9b, 32'shc24fd17c, 32'shc24f6666, 32'shc24efb5a, 32'shc24e9057, 
               32'shc24e255e, 32'shc24dba6f, 32'shc24d4f89, 32'shc24ce4ac, 32'shc24c79d9, 32'shc24c0f10, 32'shc24ba450, 32'shc24b3999, 
               32'shc24aceed, 32'shc24a6449, 32'shc249f9af, 32'shc2498f1f, 32'shc2492498, 32'shc248ba1b, 32'shc2484fa7, 32'shc247e53c, 
               32'shc2477adc, 32'shc2471084, 32'shc246a637, 32'shc2463bf2, 32'shc245d1b8, 32'shc2456786, 32'shc244fd5f, 32'shc2449341, 
               32'shc244292c, 32'shc243bf21, 32'shc243551f, 32'shc242eb27, 32'shc2428139, 32'shc2421754, 32'shc241ad78, 32'shc24143a6, 
               32'shc240d9de, 32'shc240701f, 32'shc2400669, 32'shc23f9cbd, 32'shc23f331b, 32'shc23ec982, 32'shc23e5ff3, 32'shc23df66d, 
               32'shc23d8cf1, 32'shc23d237e, 32'shc23cba15, 32'shc23c50b5, 32'shc23be75f, 32'shc23b7e12, 32'shc23b14cf, 32'shc23aab95, 
               32'shc23a4265, 32'shc239d93f, 32'shc2397021, 32'shc239070e, 32'shc2389e04, 32'shc2383504, 32'shc237cc0d, 32'shc237631f, 
               32'shc236fa3b, 32'shc2369161, 32'shc2362890, 32'shc235bfc9, 32'shc235570b, 32'shc234ee57, 32'shc23485ac, 32'shc2341d0b, 
               32'shc233b473, 32'shc2334be5, 32'shc232e361, 32'shc2327ae6, 32'shc2321274, 32'shc231aa0c, 32'shc23141ae, 32'shc230d959, 
               32'shc230710d, 32'shc23008cb, 32'shc22fa093, 32'shc22f3864, 32'shc22ed03f, 32'shc22e6823, 32'shc22e0011, 32'shc22d9808, 
               32'shc22d3009, 32'shc22cc814, 32'shc22c6028, 32'shc22bf845, 32'shc22b906c, 32'shc22b289d, 32'shc22ac0d7, 32'shc22a591a, 
               32'shc229f167, 32'shc22989be, 32'shc229221e, 32'shc228ba88, 32'shc22852fb, 32'shc227eb78, 32'shc22783fe, 32'shc2271c8e, 
               32'shc226b528, 32'shc2264dcb, 32'shc225e677, 32'shc2257f2d, 32'shc22517ed, 32'shc224b0b6, 32'shc2244989, 32'shc223e265, 
               32'shc2237b4b, 32'shc223143a, 32'shc222ad33, 32'shc2224635, 32'shc221df41, 32'shc2217857, 32'shc2211176, 32'shc220aa9e, 
               32'shc22043d0, 32'shc21fdd0c, 32'shc21f7651, 32'shc21f0fa0, 32'shc21ea8f8, 32'shc21e425a, 32'shc21ddbc5, 32'shc21d753a, 
               32'shc21d0eb8, 32'shc21ca840, 32'shc21c41d2, 32'shc21bdb6d, 32'shc21b7511, 32'shc21b0ebf, 32'shc21aa877, 32'shc21a4238, 
               32'shc219dc03, 32'shc21975d7, 32'shc2190fb5, 32'shc218a99d, 32'shc218438e, 32'shc217dd88, 32'shc217778c, 32'shc217119a, 
               32'shc216abb1, 32'shc21645d2, 32'shc215dffc, 32'shc2157a30, 32'shc215146d, 32'shc214aeb4, 32'shc2144904, 32'shc213e35e, 
               32'shc2137dc2, 32'shc213182f, 32'shc212b2a5, 32'shc2124d26, 32'shc211e7af, 32'shc2118243, 32'shc2111cdf, 32'shc210b786, 
               32'shc2105236, 32'shc20fecef, 32'shc20f87b2, 32'shc20f227f, 32'shc20ebd55, 32'shc20e5835, 32'shc20df31e, 32'shc20d8e11, 
               32'shc20d290d, 32'shc20cc413, 32'shc20c5f22, 32'shc20bfa3b, 32'shc20b955e, 32'shc20b308a, 32'shc20acbc0, 32'shc20a66ff, 
               32'shc20a0248, 32'shc2099d9a, 32'shc20938f6, 32'shc208d45b, 32'shc2086fca, 32'shc2080b43, 32'shc207a6c5, 32'shc2074251, 
               32'shc206dde6, 32'shc2067985, 32'shc206152d, 32'shc205b0df, 32'shc2054c9b, 32'shc204e860, 32'shc204842e, 32'shc2042006, 
               32'shc203bbe8, 32'shc20357d3, 32'shc202f3c8, 32'shc2028fc6, 32'shc2022bce, 32'shc201c7e0, 32'shc20163fb, 32'shc201001f, 
               32'shc2009c4e, 32'shc2003885, 32'shc1ffd4c7, 32'shc1ff7111, 32'shc1ff0d66, 32'shc1fea9c4, 32'shc1fe462b, 32'shc1fde29c, 
               32'shc1fd7f17, 32'shc1fd1b9b, 32'shc1fcb829, 32'shc1fc54c0, 32'shc1fbf161, 32'shc1fb8e0c, 32'shc1fb2ac0, 32'shc1fac77e, 
               32'shc1fa6445, 32'shc1fa0115, 32'shc1f99df0, 32'shc1f93ad4, 32'shc1f8d7c1, 32'shc1f874b8, 32'shc1f811b9, 32'shc1f7aec3, 
               32'shc1f74bd6, 32'shc1f6e8f4, 32'shc1f6861a, 32'shc1f6234b, 32'shc1f5c085, 32'shc1f55dc8, 32'shc1f4fb15, 32'shc1f4986c, 
               32'shc1f435cc, 32'shc1f3d336, 32'shc1f370a9, 32'shc1f30e26, 32'shc1f2abad, 32'shc1f2493d, 32'shc1f1e6d7, 32'shc1f1847a, 
               32'shc1f12227, 32'shc1f0bfdd, 32'shc1f05d9d, 32'shc1effb66, 32'shc1ef9939, 32'shc1ef3716, 32'shc1eed4fc, 32'shc1ee72ec, 
               32'shc1ee10e5, 32'shc1edaee8, 32'shc1ed4cf5, 32'shc1eceb0b, 32'shc1ec892b, 32'shc1ec2754, 32'shc1ebc587, 32'shc1eb63c3, 
               32'shc1eb0209, 32'shc1eaa058, 32'shc1ea3eb1, 32'shc1e9dd14, 32'shc1e97b80, 32'shc1e919f6, 32'shc1e8b876, 32'shc1e856fe, 
               32'shc1e7f591, 32'shc1e7942d, 32'shc1e732d3, 32'shc1e6d182, 32'shc1e6703b, 32'shc1e60efd, 32'shc1e5adc9, 32'shc1e54c9f, 
               32'shc1e4eb7e, 32'shc1e48a67, 32'shc1e42959, 32'shc1e3c855, 32'shc1e3675a, 32'shc1e30669, 32'shc1e2a582, 32'shc1e244a4, 
               32'shc1e1e3d0, 32'shc1e18305, 32'shc1e12244, 32'shc1e0c18d, 32'shc1e060df, 32'shc1e0003a, 32'shc1df9fa0, 32'shc1df3f0f, 
               32'shc1dede87, 32'shc1de7e09, 32'shc1de1d94, 32'shc1ddbd2a, 32'shc1dd5cc8, 32'shc1dcfc71, 32'shc1dc9c23, 32'shc1dc3bde, 
               32'shc1dbdba3, 32'shc1db7b72, 32'shc1db1b4a, 32'shc1dabb2c, 32'shc1da5b17, 32'shc1d9fb0c, 32'shc1d99b0b, 32'shc1d93b13, 
               32'shc1d8db25, 32'shc1d87b40, 32'shc1d81b65, 32'shc1d7bb93, 32'shc1d75bcb, 32'shc1d6fc0d, 32'shc1d69c58, 32'shc1d63cad, 
               32'shc1d5dd0c, 32'shc1d57d74, 32'shc1d51de5, 32'shc1d4be60, 32'shc1d45ee5, 32'shc1d3ff73, 32'shc1d3a00b, 32'shc1d340ad, 
               32'shc1d2e158, 32'shc1d2820d, 32'shc1d222cb, 32'shc1d1c393, 32'shc1d16464, 32'shc1d1053f, 32'shc1d0a624, 32'shc1d04712, 
               32'shc1cfe80a, 32'shc1cf890c, 32'shc1cf2a17, 32'shc1cecb2b, 32'shc1ce6c49, 32'shc1ce0d71, 32'shc1cdaea3, 32'shc1cd4fde, 
               32'shc1ccf122, 32'shc1cc9270, 32'shc1cc33c8, 32'shc1cbd529, 32'shc1cb7694, 32'shc1cb1809, 32'shc1cab987, 32'shc1ca5b0f, 
               32'shc1c9fca0, 32'shc1c99e3b, 32'shc1c93fdf, 32'shc1c8e18d, 32'shc1c88345, 32'shc1c82506, 32'shc1c7c6d1, 32'shc1c768a6, 
               32'shc1c70a84, 32'shc1c6ac6b, 32'shc1c64e5d, 32'shc1c5f057, 32'shc1c5925c, 32'shc1c5346a, 32'shc1c4d682, 32'shc1c478a3, 
               32'shc1c41ace, 32'shc1c3bd02, 32'shc1c35f40, 32'shc1c30188, 32'shc1c2a3d9, 32'shc1c24634, 32'shc1c1e898, 32'shc1c18b06, 
               32'shc1c12d7e, 32'shc1c0cfff, 32'shc1c0728a, 32'shc1c0151e, 32'shc1bfb7bc, 32'shc1bf5a64, 32'shc1befd15, 32'shc1be9fd0, 
               32'shc1be4294, 32'shc1bde562, 32'shc1bd883a, 32'shc1bd2b1b, 32'shc1bcce06, 32'shc1bc70fa, 32'shc1bc13f8, 32'shc1bbb700, 
               32'shc1bb5a11, 32'shc1bafd2c, 32'shc1baa050, 32'shc1ba437e, 32'shc1b9e6b6, 32'shc1b989f7, 32'shc1b92d42, 32'shc1b8d097, 
               32'shc1b873f5, 32'shc1b8175c, 32'shc1b7bacd, 32'shc1b75e48, 32'shc1b701cd, 32'shc1b6a55b, 32'shc1b648f3, 32'shc1b5ec94, 
               32'shc1b5903f, 32'shc1b533f3, 32'shc1b4d7b1, 32'shc1b47b79, 32'shc1b41f4a, 32'shc1b3c325, 32'shc1b3670a, 32'shc1b30af8, 
               32'shc1b2aef0, 32'shc1b252f1, 32'shc1b1f6fc, 32'shc1b19b10, 32'shc1b13f2f, 32'shc1b0e356, 32'shc1b08788, 32'shc1b02bc3, 
               32'shc1afd007, 32'shc1af7456, 32'shc1af18ae, 32'shc1aebd0f, 32'shc1ae617a, 32'shc1ae05ef, 32'shc1adaa6d, 32'shc1ad4ef5, 
               32'shc1acf386, 32'shc1ac9821, 32'shc1ac3cc6, 32'shc1abe174, 32'shc1ab862c, 32'shc1ab2aee, 32'shc1aacfb9, 32'shc1aa748e, 
               32'shc1aa196c, 32'shc1a9be54, 32'shc1a96346, 32'shc1a90841, 32'shc1a8ad46, 32'shc1a85254, 32'shc1a7f76c, 32'shc1a79c8e, 
               32'shc1a741b9, 32'shc1a6e6ee, 32'shc1a68c2d, 32'shc1a63175, 32'shc1a5d6c7, 32'shc1a57c22, 32'shc1a52187, 32'shc1a4c6f6, 
               32'shc1a46c6e, 32'shc1a411f0, 32'shc1a3b77b, 32'shc1a35d10, 32'shc1a302af, 32'shc1a2a857, 32'shc1a24e09, 32'shc1a1f3c5, 
               32'shc1a1998a, 32'shc1a13f59, 32'shc1a0e531, 32'shc1a08b13, 32'shc1a030ff, 32'shc19fd6f4, 32'shc19f7cf3, 32'shc19f22fb, 
               32'shc19ec90d, 32'shc19e6f29, 32'shc19e154e, 32'shc19dbb7d, 32'shc19d61b6, 32'shc19d07f8, 32'shc19cae44, 32'shc19c549a, 
               32'shc19bfaf9, 32'shc19ba161, 32'shc19b47d4, 32'shc19aee50, 32'shc19a94d5, 32'shc19a3b64, 32'shc199e1fd, 32'shc199889f, 
               32'shc1992f4c, 32'shc198d601, 32'shc1987cc1, 32'shc1982389, 32'shc197ca5c, 32'shc1977138, 32'shc197181e, 32'shc196bf0d, 
               32'shc1966606, 32'shc1960d09, 32'shc195b415, 32'shc1955b2b, 32'shc195024b, 32'shc194a974, 32'shc19450a7, 32'shc193f7e3, 
               32'shc1939f29, 32'shc1934679, 32'shc192edd2, 32'shc1929535, 32'shc1923ca2, 32'shc191e418, 32'shc1918b98, 32'shc1913321, 
               32'shc190dab4, 32'shc1908251, 32'shc19029f7, 32'shc18fd1a7, 32'shc18f7961, 32'shc18f2124, 32'shc18ec8f1, 32'shc18e70c7, 
               32'shc18e18a7, 32'shc18dc091, 32'shc18d6884, 32'shc18d1081, 32'shc18cb888, 32'shc18c6098, 32'shc18c08b2, 32'shc18bb0d5, 
               32'shc18b5903, 32'shc18b0139, 32'shc18aa97a, 32'shc18a51c4, 32'shc189fa17, 32'shc189a275, 32'shc1894adc, 32'shc188f34c, 
               32'shc1889bc6, 32'shc188444a, 32'shc187ecd8, 32'shc187956f, 32'shc1873e10, 32'shc186e6ba, 32'shc1868f6e, 32'shc186382c, 
               32'shc185e0f3, 32'shc18589c4, 32'shc185329e, 32'shc184db82, 32'shc1848470, 32'shc1842d68, 32'shc183d669, 32'shc1837f73, 
               32'shc1832888, 32'shc182d1a6, 32'shc1827acd, 32'shc18223ff, 32'shc181cd3a, 32'shc181767e, 32'shc1811fcc, 32'shc180c924, 
               32'shc1807285, 32'shc1801bf1, 32'shc17fc565, 32'shc17f6ee4, 32'shc17f186c, 32'shc17ec1fd, 32'shc17e6b99, 32'shc17e153d, 
               32'shc17dbeec, 32'shc17d68a4, 32'shc17d1266, 32'shc17cbc32, 32'shc17c6607, 32'shc17c0fe5, 32'shc17bb9ce, 32'shc17b63c0, 
               32'shc17b0dbb, 32'shc17ab7c1, 32'shc17a61d0, 32'shc17a0be8, 32'shc179b60b, 32'shc1796036, 32'shc1790a6c, 32'shc178b4ab, 
               32'shc1785ef4, 32'shc1780946, 32'shc177b3a3, 32'shc1775e08, 32'shc1770878, 32'shc176b2f1, 32'shc1765d73, 32'shc1760800, 
               32'shc175b296, 32'shc1755d35, 32'shc17507df, 32'shc174b291, 32'shc1745d4e, 32'shc1740814, 32'shc173b2e4, 32'shc1735dbd, 
               32'shc17308a1, 32'shc172b38d, 32'shc1725e84, 32'shc1720984, 32'shc171b48e, 32'shc1715fa1, 32'shc1710abe, 32'shc170b5e5, 
               32'shc1706115, 32'shc1700c4f, 32'shc16fb792, 32'shc16f62e0, 32'shc16f0e36, 32'shc16eb997, 32'shc16e6501, 32'shc16e1075, 
               32'shc16dbbf3, 32'shc16d677a, 32'shc16d130a, 32'shc16cbea5, 32'shc16c6a49, 32'shc16c15f7, 32'shc16bc1ae, 32'shc16b6d6f, 
               32'shc16b193a, 32'shc16ac50e, 32'shc16a70ec, 32'shc16a1cd4, 32'shc169c8c5, 32'shc16974c0, 32'shc16920c5, 32'shc168ccd3, 
               32'shc16878eb, 32'shc168250c, 32'shc167d137, 32'shc1677d6c, 32'shc16729ab, 32'shc166d5f3, 32'shc1668245, 32'shc1662ea0, 
               32'shc165db05, 32'shc1658774, 32'shc16533ed, 32'shc164e06f, 32'shc1648cfa, 32'shc1643990, 32'shc163e62f, 32'shc16392d8, 
               32'shc1633f8a, 32'shc162ec46, 32'shc162990c, 32'shc16245db, 32'shc161f2b4, 32'shc1619f97, 32'shc1614c83, 32'shc160f979, 
               32'shc160a678, 32'shc1605382, 32'shc1600095, 32'shc15fadb1, 32'shc15f5ad7, 32'shc15f0807, 32'shc15eb541, 32'shc15e6284, 
               32'shc15e0fd1, 32'shc15dbd27, 32'shc15d6a88, 32'shc15d17f2, 32'shc15cc565, 32'shc15c72e2, 32'shc15c2069, 32'shc15bcdfa, 
               32'shc15b7b94, 32'shc15b2937, 32'shc15ad6e5, 32'shc15a849c, 32'shc15a325d, 32'shc159e027, 32'shc1598dfb, 32'shc1593bd9, 
               32'shc158e9c1, 32'shc15897b2, 32'shc15845ac, 32'shc157f3b1, 32'shc157a1bf, 32'shc1574fd7, 32'shc156fdf8, 32'shc156ac23, 
               32'shc1565a58, 32'shc1560896, 32'shc155b6de, 32'shc1556530, 32'shc155138c, 32'shc154c1f1, 32'shc154705f, 32'shc1541ed8, 
               32'shc153cd5a, 32'shc1537be5, 32'shc1532a7b, 32'shc152d91a, 32'shc15287c3, 32'shc1523675, 32'shc151e531, 32'shc15193f7, 
               32'shc15142c6, 32'shc150f19f, 32'shc150a082, 32'shc1504f6e, 32'shc14ffe64, 32'shc14fad64, 32'shc14f5c6d, 32'shc14f0b80, 
               32'shc14eba9d, 32'shc14e69c3, 32'shc14e18f3, 32'shc14dc82d, 32'shc14d7771, 32'shc14d26be, 32'shc14cd614, 32'shc14c8575, 
               32'shc14c34df, 32'shc14be453, 32'shc14b93d0, 32'shc14b4357, 32'shc14af2e8, 32'shc14aa282, 32'shc14a5226, 32'shc14a01d4, 
               32'shc149b18b, 32'shc149614c, 32'shc1491117, 32'shc148c0ec, 32'shc14870ca, 32'shc14820b2, 32'shc147d0a3, 32'shc147809e, 
               32'shc14730a3, 32'shc146e0b1, 32'shc14690ca, 32'shc14640eb, 32'shc145f117, 32'shc145a14c, 32'shc145518b, 32'shc14501d3, 
               32'shc144b225, 32'shc1446281, 32'shc14412e7, 32'shc143c356, 32'shc14373cf, 32'shc1432451, 32'shc142d4de, 32'shc1428574, 
               32'shc1423613, 32'shc141e6bc, 32'shc141976f, 32'shc141482c, 32'shc140f8f2, 32'shc140a9c2, 32'shc1405a9c, 32'shc1400b7f, 
               32'shc13fbc6c, 32'shc13f6d63, 32'shc13f1e63, 32'shc13ecf6d, 32'shc13e8081, 32'shc13e319e, 32'shc13de2c5, 32'shc13d93f6, 
               32'shc13d4530, 32'shc13cf674, 32'shc13ca7c2, 32'shc13c591a, 32'shc13c0a7b, 32'shc13bbbe6, 32'shc13b6d5a, 32'shc13b1ed8, 
               32'shc13ad060, 32'shc13a81f2, 32'shc13a338d, 32'shc139e532, 32'shc13996e0, 32'shc1394898, 32'shc138fa5a, 32'shc138ac26, 
               32'shc1385dfb, 32'shc1380fda, 32'shc137c1c3, 32'shc13773b5, 32'shc13725b1, 32'shc136d7b7, 32'shc13689c6, 32'shc1363bdf, 
               32'shc135ee02, 32'shc135a02f, 32'shc1355265, 32'shc13504a4, 32'shc134b6ee, 32'shc1346941, 32'shc1341b9e, 32'shc133ce04, 
               32'shc1338075, 32'shc13332ef, 32'shc132e572, 32'shc13297ff, 32'shc1324a96, 32'shc131fd37, 32'shc131afe1, 32'shc1316295, 
               32'shc1311553, 32'shc130c81a, 32'shc1307aeb, 32'shc1302dc6, 32'shc12fe0ab, 32'shc12f9399, 32'shc12f4690, 32'shc12ef992, 
               32'shc12eac9d, 32'shc12e5fb2, 32'shc12e12d1, 32'shc12dc5f9, 32'shc12d792b, 32'shc12d2c66, 32'shc12cdfac, 32'shc12c92fb, 
               32'shc12c4653, 32'shc12bf9b6, 32'shc12bad22, 32'shc12b6098, 32'shc12b1417, 32'shc12ac7a0, 32'shc12a7b33, 32'shc12a2ecf, 
               32'shc129e276, 32'shc1299626, 32'shc12949df, 32'shc128fda2, 32'shc128b16f, 32'shc1286546, 32'shc1281926, 32'shc127cd10, 
               32'shc1278104, 32'shc1273501, 32'shc126e909, 32'shc1269d19, 32'shc1265134, 32'shc1260558, 32'shc125b986, 32'shc1256dbe, 
               32'shc12521ff, 32'shc124d64a, 32'shc1248a9e, 32'shc1243efd, 32'shc123f365, 32'shc123a7d7, 32'shc1235c52, 32'shc12310d7, 
               32'shc122c566, 32'shc12279fe, 32'shc1222ea1, 32'shc121e34c, 32'shc1219802, 32'shc1214cc1, 32'shc121018a, 32'shc120b65d, 
               32'shc1206b39, 32'shc120201f, 32'shc11fd50f, 32'shc11f8a09, 32'shc11f3f0c, 32'shc11ef419, 32'shc11ea92f, 32'shc11e5e4f, 
               32'shc11e1379, 32'shc11dc8ad, 32'shc11d7dea, 32'shc11d3331, 32'shc11ce882, 32'shc11c9ddd, 32'shc11c5341, 32'shc11c08af, 
               32'shc11bbe26, 32'shc11b73a7, 32'shc11b2932, 32'shc11adec7, 32'shc11a9465, 32'shc11a4a0d, 32'shc119ffbf, 32'shc119b57a, 
               32'shc1196b3f, 32'shc119210e, 32'shc118d6e7, 32'shc1188cc9, 32'shc11842b5, 32'shc117f8ab, 32'shc117aeaa, 32'shc11764b3, 
               32'shc1171ac6, 32'shc116d0e2, 32'shc1168708, 32'shc1163d38, 32'shc115f372, 32'shc115a9b5, 32'shc1156002, 32'shc1151658, 
               32'shc114ccb9, 32'shc1148323, 32'shc1143997, 32'shc113f014, 32'shc113a69b, 32'shc1135d2c, 32'shc11313c7, 32'shc112ca6b, 
               32'shc1128119, 32'shc11237d0, 32'shc111ee92, 32'shc111a55d, 32'shc1115c32, 32'shc1111310, 32'shc110c9f8, 32'shc11080ea, 
               32'shc11037e6, 32'shc10feeeb, 32'shc10fa5fa, 32'shc10f5d13, 32'shc10f1435, 32'shc10ecb62, 32'shc10e8297, 32'shc10e39d7, 
               32'shc10df120, 32'shc10da873, 32'shc10d5fd0, 32'shc10d1736, 32'shc10ccea6, 32'shc10c8620, 32'shc10c3da4, 32'shc10bf531, 
               32'shc10bacc8, 32'shc10b6468, 32'shc10b1c13, 32'shc10ad3c7, 32'shc10a8b85, 32'shc10a434c, 32'shc109fb1d, 32'shc109b2f8, 
               32'shc1096add, 32'shc10922cb, 32'shc108dac3, 32'shc10892c5, 32'shc1084ad0, 32'shc10802e5, 32'shc107bb04, 32'shc107732d, 
               32'shc1072b5f, 32'shc106e39b, 32'shc1069be1, 32'shc1065430, 32'shc1060c89, 32'shc105c4ec, 32'shc1057d59, 32'shc10535cf, 
               32'shc104ee4f, 32'shc104a6d8, 32'shc1045f6c, 32'shc1041809, 32'shc103d0b0, 32'shc1038960, 32'shc103421b, 32'shc102fadf, 
               32'shc102b3ac, 32'shc1026c84, 32'shc1022565, 32'shc101de50, 32'shc1019744, 32'shc1015042, 32'shc101094a, 32'shc100c25c, 
               32'shc1007b77, 32'shc100349c, 32'shc0ffedcb, 32'shc0ffa704, 32'shc0ff6046, 32'shc0ff1992, 32'shc0fed2e8, 32'shc0fe8c47, 
               32'shc0fe45b0, 32'shc0fdff23, 32'shc0fdb8a0, 32'shc0fd7226, 32'shc0fd2bb6, 32'shc0fce54f, 32'shc0fc9ef3, 32'shc0fc58a0, 
               32'shc0fc1257, 32'shc0fbcc17, 32'shc0fb85e2, 32'shc0fb3fb6, 32'shc0faf993, 32'shc0fab37b, 32'shc0fa6d6c, 32'shc0fa2767, 
               32'shc0f9e16b, 32'shc0f99b7a, 32'shc0f95592, 32'shc0f90fb4, 32'shc0f8c9df, 32'shc0f88414, 32'shc0f83e53, 32'shc0f7f89c, 
               32'shc0f7b2ee, 32'shc0f76d4a, 32'shc0f727b0, 32'shc0f6e220, 32'shc0f69c99, 32'shc0f6571c, 32'shc0f611a8, 32'shc0f5cc3f, 
               32'shc0f586df, 32'shc0f54189, 32'shc0f4fc3c, 32'shc0f4b6fa, 32'shc0f471c1, 32'shc0f42c91, 32'shc0f3e76c, 32'shc0f3a250, 
               32'shc0f35d3e, 32'shc0f31836, 32'shc0f2d337, 32'shc0f28e42, 32'shc0f24957, 32'shc0f20475, 32'shc0f1bf9d, 32'shc0f17acf, 
               32'shc0f1360b, 32'shc0f0f151, 32'shc0f0aca0, 32'shc0f067f9, 32'shc0f0235b, 32'shc0efdec7, 32'shc0ef9a3d, 32'shc0ef55bd, 
               32'shc0ef1147, 32'shc0eeccda, 32'shc0ee8877, 32'shc0ee441e, 32'shc0edffce, 32'shc0edbb88, 32'shc0ed774c, 32'shc0ed3319, 
               32'shc0eceef1, 32'shc0ecaad2, 32'shc0ec66bc, 32'shc0ec22b1, 32'shc0ebdeaf, 32'shc0eb9ab7, 32'shc0eb56c9, 32'shc0eb12e4, 
               32'shc0eacf09, 32'shc0ea8b38, 32'shc0ea4771, 32'shc0ea03b3, 32'shc0e9bfff, 32'shc0e97c55, 32'shc0e938b4, 32'shc0e8f51d, 
               32'shc0e8b190, 32'shc0e86e0d, 32'shc0e82a93, 32'shc0e7e724, 32'shc0e7a3bd, 32'shc0e76061, 32'shc0e71d0e, 32'shc0e6d9c5, 
               32'shc0e69686, 32'shc0e65351, 32'shc0e61025, 32'shc0e5cd03, 32'shc0e589eb, 32'shc0e546dc, 32'shc0e503d7, 32'shc0e4c0dc, 
               32'shc0e47deb, 32'shc0e43b03, 32'shc0e3f825, 32'shc0e3b551, 32'shc0e37287, 32'shc0e32fc6, 32'shc0e2ed0f, 32'shc0e2aa62, 
               32'shc0e267be, 32'shc0e22525, 32'shc0e1e294, 32'shc0e1a00e, 32'shc0e15d92, 32'shc0e11b1f, 32'shc0e0d8b6, 32'shc0e09656, 
               32'shc0e05401, 32'shc0e011b5, 32'shc0dfcf73, 32'shc0df8d3a, 32'shc0df4b0b, 32'shc0df08e6, 32'shc0dec6cb, 32'shc0de84ba, 
               32'shc0de42b2, 32'shc0de00b4, 32'shc0ddbec0, 32'shc0dd7cd5, 32'shc0dd3af4, 32'shc0dcf91d, 32'shc0dcb750, 32'shc0dc758c, 
               32'shc0dc33d2, 32'shc0dbf222, 32'shc0dbb07c, 32'shc0db6edf, 32'shc0db2d4c, 32'shc0daebc3, 32'shc0daaa44, 32'shc0da68ce, 
               32'shc0da2762, 32'shc0d9e600, 32'shc0d9a4a7, 32'shc0d96359, 32'shc0d92214, 32'shc0d8e0d8, 32'shc0d89fa7, 32'shc0d85e7f, 
               32'shc0d81d61, 32'shc0d7dc4d, 32'shc0d79b42, 32'shc0d75a41, 32'shc0d7194a, 32'shc0d6d85d, 32'shc0d69779, 32'shc0d6569f, 
               32'shc0d615cf, 32'shc0d5d509, 32'shc0d5944c, 32'shc0d55399, 32'shc0d512f0, 32'shc0d4d251, 32'shc0d491bb, 32'shc0d4512f, 
               32'shc0d410ad, 32'shc0d3d034, 32'shc0d38fc6, 32'shc0d34f61, 32'shc0d30f05, 32'shc0d2ceb4, 32'shc0d28e6c, 32'shc0d24e2e, 
               32'shc0d20dfa, 32'shc0d1cdcf, 32'shc0d18dae, 32'shc0d14d97, 32'shc0d10d8a, 32'shc0d0cd87, 32'shc0d08d8d, 32'shc0d04d9d, 
               32'shc0d00db6, 32'shc0cfcdda, 32'shc0cf8e07, 32'shc0cf4e3e, 32'shc0cf0e7f, 32'shc0cecec9, 32'shc0ce8f1d, 32'shc0ce4f7b, 
               32'shc0ce0fe3, 32'shc0cdd054, 32'shc0cd90cf, 32'shc0cd5154, 32'shc0cd11e3, 32'shc0ccd27b, 32'shc0cc931d, 32'shc0cc53c9, 
               32'shc0cc147f, 32'shc0cbd53e, 32'shc0cb9607, 32'shc0cb56da, 32'shc0cb17b7, 32'shc0cad89d, 32'shc0ca998d, 32'shc0ca5a87, 
               32'shc0ca1b8a, 32'shc0c9dc98, 32'shc0c99daf, 32'shc0c95ed0, 32'shc0c91ffa, 32'shc0c8e12f, 32'shc0c8a26d, 32'shc0c863b4, 
               32'shc0c82506, 32'shc0c7e661, 32'shc0c7a7c6, 32'shc0c76935, 32'shc0c72aae, 32'shc0c6ec30, 32'shc0c6adbc, 32'shc0c66f52, 
               32'shc0c630f2, 32'shc0c5f29b, 32'shc0c5b44e, 32'shc0c5760b, 32'shc0c537d1, 32'shc0c4f9a2, 32'shc0c4bb7c, 32'shc0c47d60, 
               32'shc0c43f4d, 32'shc0c40144, 32'shc0c3c346, 32'shc0c38550, 32'shc0c34765, 32'shc0c30983, 32'shc0c2cbab, 32'shc0c28ddd, 
               32'shc0c25019, 32'shc0c2125e, 32'shc0c1d4ad, 32'shc0c19706, 32'shc0c15969, 32'shc0c11bd5, 32'shc0c0de4b, 32'shc0c0a0cb, 
               32'shc0c06355, 32'shc0c025e8, 32'shc0bfe885, 32'shc0bfab2c, 32'shc0bf6ddd, 32'shc0bf3097, 32'shc0bef35b, 32'shc0beb629, 
               32'shc0be7901, 32'shc0be3be2, 32'shc0bdfecd, 32'shc0bdc1c2, 32'shc0bd84c1, 32'shc0bd47c9, 32'shc0bd0adb, 32'shc0bccdf7, 
               32'shc0bc911d, 32'shc0bc544d, 32'shc0bc1786, 32'shc0bbdac9, 32'shc0bb9e15, 32'shc0bb616c, 32'shc0bb24cc, 32'shc0bae836, 
               32'shc0baabaa, 32'shc0ba6f27, 32'shc0ba32af, 32'shc0b9f640, 32'shc0b9b9da, 32'shc0b97d7f, 32'shc0b9412d, 32'shc0b904e5, 
               32'shc0b8c8a7, 32'shc0b88c73, 32'shc0b85048, 32'shc0b81427, 32'shc0b7d810, 32'shc0b79c02, 32'shc0b75fff, 32'shc0b72405, 
               32'shc0b6e815, 32'shc0b6ac2e, 32'shc0b67052, 32'shc0b6347f, 32'shc0b5f8b6, 32'shc0b5bcf7, 32'shc0b58141, 32'shc0b54595, 
               32'shc0b509f3, 32'shc0b4ce5b, 32'shc0b492cc, 32'shc0b45748, 32'shc0b41bcd, 32'shc0b3e05b, 32'shc0b3a4f4, 32'shc0b36996, 
               32'shc0b32e42, 32'shc0b2f2f8, 32'shc0b2b7b8, 32'shc0b27c81, 32'shc0b24154, 32'shc0b20631, 32'shc0b1cb17, 32'shc0b19008, 
               32'shc0b15502, 32'shc0b11a06, 32'shc0b0df13, 32'shc0b0a42b, 32'shc0b0694c, 32'shc0b02e77, 32'shc0aff3ac, 32'shc0afb8ea, 
               32'shc0af7e33, 32'shc0af4385, 32'shc0af08e0, 32'shc0aece46, 32'shc0ae93b5, 32'shc0ae592e, 32'shc0ae1eb1, 32'shc0ade43e, 
               32'shc0ada9d4, 32'shc0ad6f74, 32'shc0ad351e, 32'shc0acfad2, 32'shc0acc08f, 32'shc0ac8656, 32'shc0ac4c27, 32'shc0ac1202, 
               32'shc0abd7e6, 32'shc0ab9dd5, 32'shc0ab63cd, 32'shc0ab29ce, 32'shc0aaefda, 32'shc0aab5ef, 32'shc0aa7c0e, 32'shc0aa4237, 
               32'shc0aa086a, 32'shc0a9cea6, 32'shc0a994ec, 32'shc0a95b3c, 32'shc0a92196, 32'shc0a8e7f9, 32'shc0a8ae67, 32'shc0a874de, 
               32'shc0a83b5e, 32'shc0a801e9, 32'shc0a7c87d, 32'shc0a78f1b, 32'shc0a755c3, 32'shc0a71c75, 32'shc0a6e330, 32'shc0a6a9f5, 
               32'shc0a670c4, 32'shc0a6379d, 32'shc0a5fe7f, 32'shc0a5c56c, 32'shc0a58c62, 32'shc0a55361, 32'shc0a51a6b, 32'shc0a4e17e, 
               32'shc0a4a89b, 32'shc0a46fc2, 32'shc0a436f3, 32'shc0a3fe2d, 32'shc0a3c571, 32'shc0a38cbf, 32'shc0a35417, 32'shc0a31b78, 
               32'shc0a2e2e3, 32'shc0a2aa58, 32'shc0a271d7, 32'shc0a23960, 32'shc0a200f2, 32'shc0a1c88e, 32'shc0a19034, 32'shc0a157e4, 
               32'shc0a11f9d, 32'shc0a0e760, 32'shc0a0af2d, 32'shc0a07704, 32'shc0a03ee4, 32'shc0a006cf, 32'shc09fcec3, 32'shc09f96c1, 
               32'shc09f5ec8, 32'shc09f26da, 32'shc09eeef5, 32'shc09eb71a, 32'shc09e7f48, 32'shc09e4781, 32'shc09e0fc3, 32'shc09dd80f, 
               32'shc09da065, 32'shc09d68c4, 32'shc09d312e, 32'shc09cf9a1, 32'shc09cc21e, 32'shc09c8aa4, 32'shc09c5335, 32'shc09c1bcf, 
               32'shc09be473, 32'shc09bad21, 32'shc09b75d8, 32'shc09b3e9a, 32'shc09b0765, 32'shc09ad03a, 32'shc09a9918, 32'shc09a6201, 
               32'shc09a2af3, 32'shc099f3ef, 32'shc099bcf5, 32'shc0998604, 32'shc0994f1d, 32'shc0991840, 32'shc098e16d, 32'shc098aaa4, 
               32'shc09873e4, 32'shc0983d2f, 32'shc0980683, 32'shc097cfe0, 32'shc0979948, 32'shc09762b9, 32'shc0972c34, 32'shc096f5b9, 
               32'shc096bf48, 32'shc09688e0, 32'shc0965282, 32'shc0961c2e, 32'shc095e5e4, 32'shc095afa4, 32'shc095796d, 32'shc0954340, 
               32'shc0950d1d, 32'shc094d703, 32'shc094a0f4, 32'shc0946aee, 32'shc09434f2, 32'shc093ff00, 32'shc093c917, 32'shc0939339, 
               32'shc0935d64, 32'shc0932799, 32'shc092f1d7, 32'shc092bc20, 32'shc0928672, 32'shc09250ce, 32'shc0921b34, 32'shc091e5a4, 
               32'shc091b01d, 32'shc0917aa0, 32'shc091452d, 32'shc0910fc4, 32'shc090da64, 32'shc090a50e, 32'shc0906fc3, 32'shc0903a80, 
               32'shc0900548, 32'shc08fd019, 32'shc08f9af5, 32'shc08f65da, 32'shc08f30c8, 32'shc08efbc1, 32'shc08ec6c3, 32'shc08e91cf, 
               32'shc08e5ce5, 32'shc08e2805, 32'shc08df32e, 32'shc08dbe62, 32'shc08d899f, 32'shc08d54e5, 32'shc08d2036, 32'shc08ceb90, 
               32'shc08cb6f5, 32'shc08c8262, 32'shc08c4dda, 32'shc08c195c, 32'shc08be4e7, 32'shc08bb07c, 32'shc08b7c1b, 32'shc08b47c4, 
               32'shc08b1376, 32'shc08adf32, 32'shc08aaaf8, 32'shc08a76c8, 32'shc08a42a2, 32'shc08a0e85, 32'shc089da72, 32'shc089a669, 
               32'shc089726a, 32'shc0893e75, 32'shc0890a89, 32'shc088d6a7, 32'shc088a2cf, 32'shc0886f00, 32'shc0883b3c, 32'shc0880781, 
               32'shc087d3d0, 32'shc087a029, 32'shc0876c8c, 32'shc08738f8, 32'shc087056e, 32'shc086d1ee, 32'shc0869e78, 32'shc0866b0c, 
               32'shc08637a9, 32'shc0860450, 32'shc085d101, 32'shc0859dbc, 32'shc0856a80, 32'shc085374e, 32'shc0850426, 32'shc084d108, 
               32'shc0849df4, 32'shc0846ae9, 32'shc08437e9, 32'shc08404f2, 32'shc083d204, 32'shc0839f21, 32'shc0836c47, 32'shc0833978, 
               32'shc08306b2, 32'shc082d3f5, 32'shc082a143, 32'shc0826e9a, 32'shc0823bfb, 32'shc0820966, 32'shc081d6db, 32'shc081a45a, 
               32'shc08171e2, 32'shc0813f74, 32'shc0810d10, 32'shc080dab6, 32'shc080a865, 32'shc080761e, 32'shc08043e1, 32'shc08011ae, 
               32'shc07fdf85, 32'shc07fad65, 32'shc07f7b50, 32'shc07f4944, 32'shc07f1741, 32'shc07ee549, 32'shc07eb35a, 32'shc07e8176, 
               32'shc07e4f9b, 32'shc07e1dc9, 32'shc07dec02, 32'shc07dba44, 32'shc07d8890, 32'shc07d56e6, 32'shc07d2546, 32'shc07cf3b0, 
               32'shc07cc223, 32'shc07c90a0, 32'shc07c5f27, 32'shc07c2db8, 32'shc07bfc52, 32'shc07bcaf7, 32'shc07b99a5, 32'shc07b685d, 
               32'shc07b371e, 32'shc07b05ea, 32'shc07ad4bf, 32'shc07aa39e, 32'shc07a7287, 32'shc07a417a, 32'shc07a1076, 32'shc079df7c, 
               32'shc079ae8c, 32'shc0797da6, 32'shc0794cca, 32'shc0791bf7, 32'shc078eb2f, 32'shc078ba70, 32'shc07889bb, 32'shc078590f, 
               32'shc078286e, 32'shc077f7d6, 32'shc077c748, 32'shc07796c4, 32'shc0776649, 32'shc07735d9, 32'shc0770572, 32'shc076d515, 
               32'shc076a4c2, 32'shc0767478, 32'shc0764439, 32'shc0761403, 32'shc075e3d7, 32'shc075b3b5, 32'shc075839c, 32'shc075538e, 
               32'shc0752389, 32'shc074f38e, 32'shc074c39d, 32'shc07493b5, 32'shc07463d8, 32'shc0743404, 32'shc074043a, 32'shc073d47a, 
               32'shc073a4c3, 32'shc0737517, 32'shc0734574, 32'shc07315db, 32'shc072e64c, 32'shc072b6c6, 32'shc072874b, 32'shc07257d9, 
               32'shc0722871, 32'shc071f913, 32'shc071c9be, 32'shc0719a74, 32'shc0716b33, 32'shc0713bfc, 32'shc0710ccf, 32'shc070ddab, 
               32'shc070ae92, 32'shc0707f82, 32'shc070507c, 32'shc0702180, 32'shc06ff28e, 32'shc06fc3a5, 32'shc06f94c6, 32'shc06f65f1, 
               32'shc06f3726, 32'shc06f0865, 32'shc06ed9ad, 32'shc06eaaff, 32'shc06e7c5b, 32'shc06e4dc1, 32'shc06e1f31, 32'shc06df0aa, 
               32'shc06dc22e, 32'shc06d93bb, 32'shc06d6551, 32'shc06d36f2, 32'shc06d089d, 32'shc06cda51, 32'shc06cac0f, 32'shc06c7dd7, 
               32'shc06c4fa8, 32'shc06c2184, 32'shc06bf369, 32'shc06bc558, 32'shc06b9751, 32'shc06b6954, 32'shc06b3b60, 32'shc06b0d77, 
               32'shc06adf97, 32'shc06ab1c1, 32'shc06a83f5, 32'shc06a5632, 32'shc06a2879, 32'shc069facb, 32'shc069cd26, 32'shc0699f8a, 
               32'shc06971f9, 32'shc0694471, 32'shc06916f3, 32'shc068e97f, 32'shc068bc15, 32'shc0688eb5, 32'shc068615e, 32'shc0683411, 
               32'shc06806ce, 32'shc067d995, 32'shc067ac66, 32'shc0677f40, 32'shc0675225, 32'shc0672513, 32'shc066f80a, 32'shc066cb0c, 
               32'shc0669e18, 32'shc066712d, 32'shc066444c, 32'shc0661775, 32'shc065eaa8, 32'shc065bde4, 32'shc065912a, 32'shc065647b, 
               32'shc06537d4, 32'shc0650b38, 32'shc064dea6, 32'shc064b21d, 32'shc064859e, 32'shc0645929, 32'shc0642cbe, 32'shc064005d, 
               32'shc063d405, 32'shc063a7b7, 32'shc0637b73, 32'shc0634f39, 32'shc0632309, 32'shc062f6e2, 32'shc062cac6, 32'shc0629eb3, 
               32'shc06272aa, 32'shc06246aa, 32'shc0621ab5, 32'shc061eec9, 32'shc061c2e7, 32'shc061970f, 32'shc0616b41, 32'shc0613f7d, 
               32'shc06113c2, 32'shc060e811, 32'shc060bc6a, 32'shc06090cd, 32'shc060653a, 32'shc06039b0, 32'shc0600e30, 32'shc05fe2ba, 
               32'shc05fb74e, 32'shc05f8bec, 32'shc05f6093, 32'shc05f3545, 32'shc05f0a00, 32'shc05edec5, 32'shc05eb393, 32'shc05e886c, 
               32'shc05e5d4e, 32'shc05e323a, 32'shc05e0730, 32'shc05ddc30, 32'shc05db13a, 32'shc05d864d, 32'shc05d5b6b, 32'shc05d3092, 
               32'shc05d05c3, 32'shc05cdafd, 32'shc05cb042, 32'shc05c8590, 32'shc05c5ae8, 32'shc05c304a, 32'shc05c05b6, 32'shc05bdb2b, 
               32'shc05bb0ab, 32'shc05b8634, 32'shc05b5bc7, 32'shc05b3164, 32'shc05b070a, 32'shc05adcbb, 32'shc05ab275, 32'shc05a8839, 
               32'shc05a5e07, 32'shc05a33df, 32'shc05a09c0, 32'shc059dfac, 32'shc059b5a1, 32'shc0598ba0, 32'shc05961a9, 32'shc05937bb, 
               32'shc0590dd8, 32'shc058e3fe, 32'shc058ba2e, 32'shc0589068, 32'shc05866ac, 32'shc0583cf9, 32'shc0581350, 32'shc057e9b2, 
               32'shc057c01d, 32'shc0579691, 32'shc0576d10, 32'shc0574398, 32'shc0571a2b, 32'shc056f0c7, 32'shc056c76c, 32'shc0569e1c, 
               32'shc05674d6, 32'shc0564b99, 32'shc0562266, 32'shc055f93d, 32'shc055d01e, 32'shc055a708, 32'shc0557dfd, 32'shc05554fb, 
               32'shc0552c03, 32'shc0550315, 32'shc054da30, 32'shc054b156, 32'shc0548885, 32'shc0545fbe, 32'shc0543701, 32'shc0540e4e, 
               32'shc053e5a5, 32'shc053bd05, 32'shc053946f, 32'shc0536be3, 32'shc0534361, 32'shc0531ae9, 32'shc052f27a, 32'shc052ca16, 
               32'shc052a1bb, 32'shc052796a, 32'shc0525123, 32'shc05228e5, 32'shc05200b2, 32'shc051d888, 32'shc051b068, 32'shc0518852, 
               32'shc0516045, 32'shc0513843, 32'shc051104a, 32'shc050e85c, 32'shc050c077, 32'shc050989b, 32'shc05070ca, 32'shc0504902, 
               32'shc0502145, 32'shc04ff991, 32'shc04fd1e7, 32'shc04faa46, 32'shc04f82b0, 32'shc04f5b23, 32'shc04f33a1, 32'shc04f0c28, 
               32'shc04ee4b8, 32'shc04ebd53, 32'shc04e95f8, 32'shc04e6ea6, 32'shc04e475e, 32'shc04e2020, 32'shc04df8ec, 32'shc04dd1c1, 
               32'shc04daaa1, 32'shc04d838a, 32'shc04d5c7d, 32'shc04d357a, 32'shc04d0e81, 32'shc04ce791, 32'shc04cc0ac, 32'shc04c99d0, 
               32'shc04c72fe, 32'shc04c4c36, 32'shc04c2577, 32'shc04bfec3, 32'shc04bd818, 32'shc04bb177, 32'shc04b8ae0, 32'shc04b6453, 
               32'shc04b3dcf, 32'shc04b1756, 32'shc04af0e6, 32'shc04aca80, 32'shc04aa424, 32'shc04a7dd2, 32'shc04a5789, 32'shc04a314b, 
               32'shc04a0b16, 32'shc049e4eb, 32'shc049beca, 32'shc04998b2, 32'shc04972a5, 32'shc0494ca1, 32'shc04926a7, 32'shc04900b7, 
               32'shc048dad1, 32'shc048b4f5, 32'shc0488f22, 32'shc0486959, 32'shc048439b, 32'shc0481de5, 32'shc047f83a, 32'shc047d299, 
               32'shc047ad01, 32'shc0478773, 32'shc04761ef, 32'shc0473c75, 32'shc0471705, 32'shc046f19f, 32'shc046cc42, 32'shc046a6ef, 
               32'shc04681a6, 32'shc0465c67, 32'shc0463732, 32'shc0461206, 32'shc045ece5, 32'shc045c7cd, 32'shc045a2bf, 32'shc0457dba, 
               32'shc04558c0, 32'shc04533d0, 32'shc0450ee9, 32'shc044ea0c, 32'shc044c539, 32'shc044a070, 32'shc0447bb0, 32'shc04456fb, 
               32'shc044324f, 32'shc0440dad, 32'shc043e915, 32'shc043c487, 32'shc043a002, 32'shc0437b88, 32'shc0435717, 32'shc04332b0, 
               32'shc0430e53, 32'shc042ea00, 32'shc042c5b6, 32'shc042a177, 32'shc0427d41, 32'shc0425915, 32'shc04234f3, 32'shc04210da, 
               32'shc041eccc, 32'shc041c8c7, 32'shc041a4cd, 32'shc04180dc, 32'shc0415cf4, 32'shc0413917, 32'shc0411544, 32'shc040f17a, 
               32'shc040cdba, 32'shc040aa04, 32'shc0408658, 32'shc04062b6, 32'shc0403f1d, 32'shc0401b8e, 32'shc03ff80a, 32'shc03fd48f, 
               32'shc03fb11d, 32'shc03f8db6, 32'shc03f6a58, 32'shc03f4705, 32'shc03f23bb, 32'shc03f007b, 32'shc03edd45, 32'shc03eba18, 
               32'shc03e96f6, 32'shc03e73dd, 32'shc03e50ce, 32'shc03e2dc9, 32'shc03e0ace, 32'shc03de7dd, 32'shc03dc4f5, 32'shc03da217, 
               32'shc03d7f44, 32'shc03d5c79, 32'shc03d39b9, 32'shc03d1703, 32'shc03cf456, 32'shc03cd1b4, 32'shc03caf1b, 32'shc03c8c8c, 
               32'shc03c6a07, 32'shc03c478b, 32'shc03c251a, 32'shc03c02b2, 32'shc03be054, 32'shc03bbe00, 32'shc03b9bb6, 32'shc03b7975, 
               32'shc03b573f, 32'shc03b3512, 32'shc03b12ef, 32'shc03af0d6, 32'shc03acec7, 32'shc03aacc2, 32'shc03a8ac6, 32'shc03a68d4, 
               32'shc03a46ed, 32'shc03a250e, 32'shc03a033a, 32'shc039e170, 32'shc039bfaf, 32'shc0399df9, 32'shc0397c4c, 32'shc0395aa9, 
               32'shc0393910, 32'shc0391780, 32'shc038f5fb, 32'shc038d47f, 32'shc038b30d, 32'shc03891a5, 32'shc0387047, 32'shc0384ef3, 
               32'shc0382da8, 32'shc0380c68, 32'shc037eb31, 32'shc037ca04, 32'shc037a8e1, 32'shc03787c7, 32'shc03766b8, 32'shc03745b2, 
               32'shc03724b6, 32'shc03703c4, 32'shc036e2dc, 32'shc036c1fe, 32'shc036a129, 32'shc036805f, 32'shc0365f9e, 32'shc0363ee7, 
               32'shc0361e3a, 32'shc035fd96, 32'shc035dcfd, 32'shc035bc6d, 32'shc0359be8, 32'shc0357b6c, 32'shc0355afa, 32'shc0353a91, 
               32'shc0351a33, 32'shc034f9de, 32'shc034d994, 32'shc034b953, 32'shc034991c, 32'shc03478ee, 32'shc03458cb, 32'shc03438b1, 
               32'shc03418a2, 32'shc033f89c, 32'shc033d8a0, 32'shc033b8ad, 32'shc03398c5, 32'shc03378e7, 32'shc0335912, 32'shc0333947, 
               32'shc0331986, 32'shc032f9cf, 32'shc032da22, 32'shc032ba7e, 32'shc0329ae4, 32'shc0327b55, 32'shc0325bcf, 32'shc0323c52, 
               32'shc0321ce0, 32'shc031fd78, 32'shc031de19, 32'shc031bec4, 32'shc0319f79, 32'shc0318038, 32'shc0316101, 32'shc03141d3, 
               32'shc03122b0, 32'shc0310396, 32'shc030e486, 32'shc030c580, 32'shc030a684, 32'shc0308792, 32'shc03068a9, 32'shc03049ca, 
               32'shc0302af5, 32'shc0300c2a, 32'shc02fed69, 32'shc02fceb2, 32'shc02fb004, 32'shc02f9161, 32'shc02f72c7, 32'shc02f5437, 
               32'shc02f35b1, 32'shc02f1734, 32'shc02ef8c2, 32'shc02eda59, 32'shc02ebbfb, 32'shc02e9da6, 32'shc02e7f5b, 32'shc02e6119, 
               32'shc02e42e2, 32'shc02e24b4, 32'shc02e0691, 32'shc02de877, 32'shc02dca67, 32'shc02dac61, 32'shc02d8e64, 32'shc02d7072, 
               32'shc02d5289, 32'shc02d34aa, 32'shc02d16d5, 32'shc02cf90a, 32'shc02cdb49, 32'shc02cbd91, 32'shc02c9fe4, 32'shc02c8240, 
               32'shc02c64a6, 32'shc02c4716, 32'shc02c2990, 32'shc02c0c13, 32'shc02beea1, 32'shc02bd138, 32'shc02bb3d9, 32'shc02b9684, 
               32'shc02b7939, 32'shc02b5bf8, 32'shc02b3ec0, 32'shc02b2192, 32'shc02b046f, 32'shc02ae755, 32'shc02aca44, 32'shc02aad3e, 
               32'shc02a9042, 32'shc02a734f, 32'shc02a5666, 32'shc02a3988, 32'shc02a1cb2, 32'shc029ffe7, 32'shc029e326, 32'shc029c66e, 
               32'shc029a9c1, 32'shc0298d1d, 32'shc0297083, 32'shc02953f3, 32'shc029376c, 32'shc0291af0, 32'shc028fe7d, 32'shc028e215, 
               32'shc028c5b6, 32'shc028a961, 32'shc0288d15, 32'shc02870d4, 32'shc028549c, 32'shc028386f, 32'shc0281c4b, 32'shc0280031, 
               32'shc027e421, 32'shc027c81a, 32'shc027ac1e, 32'shc027902b, 32'shc0277442, 32'shc0275864, 32'shc0273c8e, 32'shc02720c3, 
               32'shc0270502, 32'shc026e94a, 32'shc026cd9d, 32'shc026b1f9, 32'shc026965f, 32'shc0267acf, 32'shc0265f48, 32'shc02643cc, 
               32'shc0262859, 32'shc0260cf0, 32'shc025f191, 32'shc025d63c, 32'shc025baf1, 32'shc0259fb0, 32'shc0258478, 32'shc025694a, 
               32'shc0254e27, 32'shc025330d, 32'shc02517fc, 32'shc024fcf6, 32'shc024e1fa, 32'shc024c707, 32'shc024ac1e, 32'shc024913f, 
               32'shc024766a, 32'shc0245b9f, 32'shc02440de, 32'shc0242626, 32'shc0240b78, 32'shc023f0d5, 32'shc023d63b, 32'shc023bbab, 
               32'shc023a124, 32'shc02386a8, 32'shc0236c35, 32'shc02351cc, 32'shc023376e, 32'shc0231d18, 32'shc02302cd, 32'shc022e88c, 
               32'shc022ce54, 32'shc022b427, 32'shc0229a03, 32'shc0227fe9, 32'shc02265d9, 32'shc0224bd3, 32'shc02231d6, 32'shc02217e4, 
               32'shc021fdfb, 32'shc021e41c, 32'shc021ca47, 32'shc021b07c, 32'shc02196bb, 32'shc0217d03, 32'shc0216356, 32'shc02149b2, 
               32'shc0213018, 32'shc0211688, 32'shc020fd02, 32'shc020e385, 32'shc020ca13, 32'shc020b0aa, 32'shc020974b, 32'shc0207df6, 
               32'shc02064ab, 32'shc0204b6a, 32'shc0203232, 32'shc0201905, 32'shc01fffe1, 32'shc01fe6c7, 32'shc01fcdb7, 32'shc01fb4b1, 
               32'shc01f9bb5, 32'shc01f82c2, 32'shc01f69da, 32'shc01f50fb, 32'shc01f3826, 32'shc01f1f5b, 32'shc01f069a, 32'shc01eede2, 
               32'shc01ed535, 32'shc01ebc91, 32'shc01ea3f7, 32'shc01e8b67, 32'shc01e72e1, 32'shc01e5a65, 32'shc01e41f3, 32'shc01e298a, 
               32'shc01e112b, 32'shc01df8d7, 32'shc01de08c, 32'shc01dc84a, 32'shc01db013, 32'shc01d97e6, 32'shc01d7fc2, 32'shc01d67a8, 
               32'shc01d4f99, 32'shc01d3792, 32'shc01d1f96, 32'shc01d07a4, 32'shc01cefbb, 32'shc01cd7dd, 32'shc01cc008, 32'shc01ca83d, 
               32'shc01c907c, 32'shc01c78c5, 32'shc01c6118, 32'shc01c4974, 32'shc01c31da, 32'shc01c1a4b, 32'shc01c02c5, 32'shc01beb48, 
               32'shc01bd3d6, 32'shc01bbc6e, 32'shc01ba50f, 32'shc01b8dbb, 32'shc01b7670, 32'shc01b5f2f, 32'shc01b47f8, 32'shc01b30ca, 
               32'shc01b19a7, 32'shc01b028d, 32'shc01aeb7e, 32'shc01ad478, 32'shc01abd7c, 32'shc01aa68a, 32'shc01a8fa1, 32'shc01a78c3, 
               32'shc01a61ee, 32'shc01a4b24, 32'shc01a3463, 32'shc01a1dac, 32'shc01a06fe, 32'shc019f05b, 32'shc019d9c2, 32'shc019c332, 
               32'shc019acac, 32'shc0199630, 32'shc0197fbe, 32'shc0196956, 32'shc01952f8, 32'shc0193ca3, 32'shc0192659, 32'shc0191018, 
               32'shc018f9e1, 32'shc018e3b4, 32'shc018cd91, 32'shc018b777, 32'shc018a168, 32'shc0188b62, 32'shc0187566, 32'shc0185f74, 
               32'shc018498c, 32'shc01833ae, 32'shc0181dda, 32'shc018080f, 32'shc017f24e, 32'shc017dc98, 32'shc017c6eb, 32'shc017b148, 
               32'shc0179bae, 32'shc017861f, 32'shc0177099, 32'shc0175b1e, 32'shc01745ac, 32'shc0173044, 32'shc0171ae6, 32'shc0170591, 
               32'shc016f047, 32'shc016db07, 32'shc016c5d0, 32'shc016b0a3, 32'shc0169b80, 32'shc0168667, 32'shc0167158, 32'shc0165c52, 
               32'shc0164757, 32'shc0163265, 32'shc0161d7d, 32'shc016089f, 32'shc015f3cb, 32'shc015df01, 32'shc015ca40, 32'shc015b58a, 
               32'shc015a0dd, 32'shc0158c3a, 32'shc01577a1, 32'shc0156312, 32'shc0154e8d, 32'shc0153a11, 32'shc01525a0, 32'shc0151138, 
               32'shc014fcda, 32'shc014e886, 32'shc014d43c, 32'shc014bffc, 32'shc014abc5, 32'shc0149799, 32'shc0148376, 32'shc0146f5d, 
               32'shc0145b4e, 32'shc0144749, 32'shc014334e, 32'shc0141f5c, 32'shc0140b75, 32'shc013f797, 32'shc013e3c3, 32'shc013cff9, 
               32'shc013bc39, 32'shc013a883, 32'shc01394d6, 32'shc0138134, 32'shc0136d9b, 32'shc0135a0c, 32'shc0134687, 32'shc013330c, 
               32'shc0131f9b, 32'shc0130c33, 32'shc012f8d6, 32'shc012e582, 32'shc012d238, 32'shc012bef8, 32'shc012abc2, 32'shc0129896, 
               32'shc0128574, 32'shc012725b, 32'shc0125f4c, 32'shc0124c47, 32'shc012394c, 32'shc012265b, 32'shc0121374, 32'shc0120097, 
               32'shc011edc3, 32'shc011daf9, 32'shc011c83a, 32'shc011b584, 32'shc011a2d8, 32'shc0119035, 32'shc0117d9d, 32'shc0116b0e, 
               32'shc011588a, 32'shc011460f, 32'shc011339e, 32'shc0112137, 32'shc0110eda, 32'shc010fc86, 32'shc010ea3d, 32'shc010d7fd, 
               32'shc010c5c7, 32'shc010b39b, 32'shc010a179, 32'shc0108f61, 32'shc0107d53, 32'shc0106b4e, 32'shc0105954, 32'shc0104763, 
               32'shc010357c, 32'shc010239f, 32'shc01011cc, 32'shc0100002, 32'shc00fee43, 32'shc00fdc8d, 32'shc00fcae2, 32'shc00fb940, 
               32'shc00fa7a8, 32'shc00f9619, 32'shc00f8495, 32'shc00f731b, 32'shc00f61aa, 32'shc00f5043, 32'shc00f3ee6, 32'shc00f2d93, 
               32'shc00f1c4a, 32'shc00f0b0b, 32'shc00ef9d6, 32'shc00ee8aa, 32'shc00ed788, 32'shc00ec670, 32'shc00eb562, 32'shc00ea45e, 
               32'shc00e9364, 32'shc00e8274, 32'shc00e718d, 32'shc00e60b0, 32'shc00e4fde, 32'shc00e3f15, 32'shc00e2e56, 32'shc00e1da0, 
               32'shc00e0cf5, 32'shc00dfc53, 32'shc00debbc, 32'shc00ddb2e, 32'shc00dcaaa, 32'shc00dba30, 32'shc00da9c0, 32'shc00d9959, 
               32'shc00d88fd, 32'shc00d78aa, 32'shc00d6861, 32'shc00d5823, 32'shc00d47ed, 32'shc00d37c2, 32'shc00d27a1, 32'shc00d178a, 
               32'shc00d077c, 32'shc00cf778, 32'shc00ce77e, 32'shc00cd78e, 32'shc00cc7a8, 32'shc00cb7cc, 32'shc00ca7f9, 32'shc00c9831, 
               32'shc00c8872, 32'shc00c78bd, 32'shc00c6912, 32'shc00c5971, 32'shc00c49da, 32'shc00c3a4d, 32'shc00c2ac9, 32'shc00c1b4f, 
               32'shc00c0be0, 32'shc00bfc7a, 32'shc00bed1e, 32'shc00bddcb, 32'shc00bce83, 32'shc00bbf44, 32'shc00bb010, 32'shc00ba0e5, 
               32'shc00b91c4, 32'shc00b82ad, 32'shc00b73a0, 32'shc00b649d, 32'shc00b55a3, 32'shc00b46b4, 32'shc00b37ce, 32'shc00b28f2, 
               32'shc00b1a20, 32'shc00b0b58, 32'shc00afc9a, 32'shc00aede5, 32'shc00adf3b, 32'shc00ad09a, 32'shc00ac203, 32'shc00ab376, 
               32'shc00aa4f3, 32'shc00a967a, 32'shc00a880a, 32'shc00a79a5, 32'shc00a6b49, 32'shc00a5cf8, 32'shc00a4eb0, 32'shc00a4072, 
               32'shc00a323d, 32'shc00a2413, 32'shc00a15f3, 32'shc00a07dc, 32'shc009f9cf, 32'shc009ebcc, 32'shc009ddd3, 32'shc009cfe4, 
               32'shc009c1ff, 32'shc009b423, 32'shc009a652, 32'shc009988a, 32'shc0098acc, 32'shc0097d18, 32'shc0096f6e, 32'shc00961ce, 
               32'shc0095438, 32'shc00946ab, 32'shc0093929, 32'shc0092bb0, 32'shc0091e41, 32'shc00910dc, 32'shc0090381, 32'shc008f62f, 
               32'shc008e8e8, 32'shc008dbaa, 32'shc008ce76, 32'shc008c14d, 32'shc008b42d, 32'shc008a716, 32'shc0089a0a, 32'shc0088d08, 
               32'shc008800f, 32'shc0087321, 32'shc008663c, 32'shc0085961, 32'shc0084c90, 32'shc0083fc8, 32'shc008330b, 32'shc0082658, 
               32'shc00819ae, 32'shc0080d0e, 32'shc0080078, 32'shc007f3ec, 32'shc007e76a, 32'shc007daf2, 32'shc007ce83, 32'shc007c21f, 
               32'shc007b5c4, 32'shc007a973, 32'shc0079d2c, 32'shc00790ef, 32'shc00784bc, 32'shc0077893, 32'shc0076c73, 32'shc007605d, 
               32'shc0075452, 32'shc0074850, 32'shc0073c58, 32'shc0073069, 32'shc0072485, 32'shc00718ab, 32'shc0070cda, 32'shc0070113, 
               32'shc006f556, 32'shc006e9a3, 32'shc006ddfa, 32'shc006d25b, 32'shc006c6c6, 32'shc006bb3a, 32'shc006afb8, 32'shc006a441, 
               32'shc00698d3, 32'shc0068d6f, 32'shc0068214, 32'shc00676c4, 32'shc0066b7d, 32'shc0066041, 32'shc006550e, 32'shc00649e5, 
               32'shc0063ec6, 32'shc00633b1, 32'shc00628a6, 32'shc0061da4, 32'shc00612ad, 32'shc00607bf, 32'shc005fcdb, 32'shc005f201, 
               32'shc005e731, 32'shc005dc6b, 32'shc005d1af, 32'shc005c6fc, 32'shc005bc54, 32'shc005b1b5, 32'shc005a720, 32'shc0059c95, 
               32'shc0059214, 32'shc005879c, 32'shc0057d2f, 32'shc00572cb, 32'shc0056872, 32'shc0055e22, 32'shc00553dc, 32'shc00549a0, 
               32'shc0053f6e, 32'shc0053545, 32'shc0052b27, 32'shc0052112, 32'shc0051707, 32'shc0050d06, 32'shc005030f, 32'shc004f922, 
               32'shc004ef3f, 32'shc004e566, 32'shc004db96, 32'shc004d1d0, 32'shc004c814, 32'shc004be62, 32'shc004b4ba, 32'shc004ab1c, 
               32'shc004a188, 32'shc00497fd, 32'shc0048e7d, 32'shc0048506, 32'shc0047b99, 32'shc0047236, 32'shc00468dd, 32'shc0045f8d, 
               32'shc0045648, 32'shc0044d0d, 32'shc00443db, 32'shc0043ab3, 32'shc0043195, 32'shc0042881, 32'shc0041f77, 32'shc0041676, 
               32'shc0040d80, 32'shc0040493, 32'shc003fbb0, 32'shc003f2d8, 32'shc003ea09, 32'shc003e143, 32'shc003d888, 32'shc003cfd7, 
               32'shc003c72f, 32'shc003be91, 32'shc003b5fe, 32'shc003ad74, 32'shc003a4f4, 32'shc0039c7d, 32'shc0039411, 32'shc0038baf, 
               32'shc0038356, 32'shc0037b07, 32'shc00372c2, 32'shc0036a87, 32'shc0036256, 32'shc0035a2f, 32'shc0035211, 32'shc00349fe, 
               32'shc00341f4, 32'shc00339f4, 32'shc00331fe, 32'shc0032a12, 32'shc0032230, 32'shc0031a58, 32'shc0031289, 32'shc0030ac5, 
               32'shc003030a, 32'shc002fb59, 32'shc002f3b2, 32'shc002ec15, 32'shc002e482, 32'shc002dcf8, 32'shc002d579, 32'shc002ce03, 
               32'shc002c697, 32'shc002bf35, 32'shc002b7dd, 32'shc002b08f, 32'shc002a94b, 32'shc002a210, 32'shc0029ae0, 32'shc00293b9, 
               32'shc0028c9c, 32'shc0028589, 32'shc0027e80, 32'shc0027781, 32'shc002708c, 32'shc00269a0, 32'shc00262be, 32'shc0025be7, 
               32'shc0025519, 32'shc0024e55, 32'shc002479b, 32'shc00240ea, 32'shc0023a44, 32'shc00233a7, 32'shc0022d15, 32'shc002268c, 
               32'shc002200d, 32'shc0021998, 32'shc002132d, 32'shc0020ccb, 32'shc0020674, 32'shc0020026, 32'shc001f9e2, 32'shc001f3a8, 
               32'shc001ed78, 32'shc001e752, 32'shc001e136, 32'shc001db24, 32'shc001d51b, 32'shc001cf1c, 32'shc001c928, 32'shc001c33d, 
               32'shc001bd5c, 32'shc001b784, 32'shc001b1b7, 32'shc001abf4, 32'shc001a63a, 32'shc001a08a, 32'shc0019ae5, 32'shc0019549, 
               32'shc0018fb6, 32'shc0018a2e, 32'shc00184b0, 32'shc0017f3b, 32'shc00179d1, 32'shc0017470, 32'shc0016f19, 32'shc00169cc, 
               32'shc0016489, 32'shc0015f50, 32'shc0015a20, 32'shc00154fb, 32'shc0014fdf, 32'shc0014acd, 32'shc00145c5, 32'shc00140c7, 
               32'shc0013bd3, 32'shc00136e8, 32'shc0013208, 32'shc0012d31, 32'shc0012865, 32'shc00123a2, 32'shc0011ee9, 32'shc0011a3a, 
               32'shc0011594, 32'shc00110f9, 32'shc0010c67, 32'shc00107e0, 32'shc0010362, 32'shc000feee, 32'shc000fa84, 32'shc000f624, 
               32'shc000f1ce, 32'shc000ed81, 32'shc000e93f, 32'shc000e506, 32'shc000e0d7, 32'shc000dcb2, 32'shc000d897, 32'shc000d486, 
               32'shc000d07e, 32'shc000cc81, 32'shc000c88d, 32'shc000c4a4, 32'shc000c0c4, 32'shc000bcee, 32'shc000b921, 32'shc000b55f, 
               32'shc000b1a7, 32'shc000adf8, 32'shc000aa54, 32'shc000a6b9, 32'shc000a328, 32'shc0009fa1, 32'shc0009c24, 32'shc00098b0, 
               32'shc0009547, 32'shc00091e7, 32'shc0008e92, 32'shc0008b46, 32'shc0008804, 32'shc00084cc, 32'shc000819d, 32'shc0007e79, 
               32'shc0007b5f, 32'shc000784e, 32'shc0007547, 32'shc000724a, 32'shc0006f57, 32'shc0006c6e, 32'shc000698f, 32'shc00066b9, 
               32'shc00063ee, 32'shc000612c, 32'shc0005e74, 32'shc0005bc7, 32'shc0005922, 32'shc0005688, 32'shc00053f8, 32'shc0005171, 
               32'shc0004ef5, 32'shc0004c82, 32'shc0004a19, 32'shc00047ba, 32'shc0004565, 32'shc000431a, 32'shc00040d9, 32'shc0003ea1, 
               32'shc0003c74, 32'shc0003a50, 32'shc0003836, 32'shc0003626, 32'shc0003420, 32'shc0003223, 32'shc0003031, 32'shc0002e48, 
               32'shc0002c6a, 32'shc0002a95, 32'shc00028ca, 32'shc0002709, 32'shc0002552, 32'shc00023a4, 32'shc0002201, 32'shc0002067, 
               32'shc0001ed8, 32'shc0001d52, 32'shc0001bd6, 32'shc0001a64, 32'shc00018fb, 32'shc000179d, 32'shc0001649, 32'shc00014fe, 
               32'shc00013bd, 32'shc0001286, 32'shc0001159, 32'shc0001036, 32'shc0000f1d, 32'shc0000e0d, 32'shc0000d08, 32'shc0000c0c, 
               32'shc0000b1a, 32'shc0000a33, 32'shc0000954, 32'shc0000880, 32'shc00007b6, 32'shc00006f5, 32'shc000063f, 32'shc0000592, 
               32'shc00004ef, 32'shc0000456, 32'shc00003c7, 32'shc0000342, 32'shc00002c7, 32'shc0000255, 32'shc00001ed, 32'shc0000190, 
               32'shc000013c, 32'shc00000f2, 32'shc00000b2, 32'shc000007b, 32'shc000004f, 32'shc000002c, 32'shc0000014, 32'shc0000005, 
               32'shc0000000, 32'shc0000005, 32'shc0000014, 32'shc000002c, 32'shc000004f, 32'shc000007b, 32'shc00000b2, 32'shc00000f2, 
               32'shc000013c, 32'shc0000190, 32'shc00001ed, 32'shc0000255, 32'shc00002c7, 32'shc0000342, 32'shc00003c7, 32'shc0000456, 
               32'shc00004ef, 32'shc0000592, 32'shc000063f, 32'shc00006f5, 32'shc00007b6, 32'shc0000880, 32'shc0000954, 32'shc0000a33, 
               32'shc0000b1a, 32'shc0000c0c, 32'shc0000d08, 32'shc0000e0d, 32'shc0000f1d, 32'shc0001036, 32'shc0001159, 32'shc0001286, 
               32'shc00013bd, 32'shc00014fe, 32'shc0001649, 32'shc000179d, 32'shc00018fb, 32'shc0001a64, 32'shc0001bd6, 32'shc0001d52, 
               32'shc0001ed8, 32'shc0002067, 32'shc0002201, 32'shc00023a4, 32'shc0002552, 32'shc0002709, 32'shc00028ca, 32'shc0002a95, 
               32'shc0002c6a, 32'shc0002e48, 32'shc0003031, 32'shc0003223, 32'shc0003420, 32'shc0003626, 32'shc0003836, 32'shc0003a50, 
               32'shc0003c74, 32'shc0003ea1, 32'shc00040d9, 32'shc000431a, 32'shc0004565, 32'shc00047ba, 32'shc0004a19, 32'shc0004c82, 
               32'shc0004ef5, 32'shc0005171, 32'shc00053f8, 32'shc0005688, 32'shc0005922, 32'shc0005bc7, 32'shc0005e74, 32'shc000612c, 
               32'shc00063ee, 32'shc00066b9, 32'shc000698f, 32'shc0006c6e, 32'shc0006f57, 32'shc000724a, 32'shc0007547, 32'shc000784e, 
               32'shc0007b5f, 32'shc0007e79, 32'shc000819d, 32'shc00084cc, 32'shc0008804, 32'shc0008b46, 32'shc0008e92, 32'shc00091e7, 
               32'shc0009547, 32'shc00098b0, 32'shc0009c24, 32'shc0009fa1, 32'shc000a328, 32'shc000a6b9, 32'shc000aa54, 32'shc000adf8, 
               32'shc000b1a7, 32'shc000b55f, 32'shc000b921, 32'shc000bcee, 32'shc000c0c4, 32'shc000c4a4, 32'shc000c88d, 32'shc000cc81, 
               32'shc000d07e, 32'shc000d486, 32'shc000d897, 32'shc000dcb2, 32'shc000e0d7, 32'shc000e506, 32'shc000e93f, 32'shc000ed81, 
               32'shc000f1ce, 32'shc000f624, 32'shc000fa84, 32'shc000feee, 32'shc0010362, 32'shc00107e0, 32'shc0010c67, 32'shc00110f9, 
               32'shc0011594, 32'shc0011a3a, 32'shc0011ee9, 32'shc00123a2, 32'shc0012865, 32'shc0012d31, 32'shc0013208, 32'shc00136e8, 
               32'shc0013bd3, 32'shc00140c7, 32'shc00145c5, 32'shc0014acd, 32'shc0014fdf, 32'shc00154fb, 32'shc0015a20, 32'shc0015f50, 
               32'shc0016489, 32'shc00169cc, 32'shc0016f19, 32'shc0017470, 32'shc00179d1, 32'shc0017f3b, 32'shc00184b0, 32'shc0018a2e, 
               32'shc0018fb6, 32'shc0019549, 32'shc0019ae5, 32'shc001a08a, 32'shc001a63a, 32'shc001abf4, 32'shc001b1b7, 32'shc001b784, 
               32'shc001bd5c, 32'shc001c33d, 32'shc001c928, 32'shc001cf1c, 32'shc001d51b, 32'shc001db24, 32'shc001e136, 32'shc001e752, 
               32'shc001ed78, 32'shc001f3a8, 32'shc001f9e2, 32'shc0020026, 32'shc0020674, 32'shc0020ccb, 32'shc002132d, 32'shc0021998, 
               32'shc002200d, 32'shc002268c, 32'shc0022d15, 32'shc00233a7, 32'shc0023a44, 32'shc00240ea, 32'shc002479b, 32'shc0024e55, 
               32'shc0025519, 32'shc0025be7, 32'shc00262be, 32'shc00269a0, 32'shc002708c, 32'shc0027781, 32'shc0027e80, 32'shc0028589, 
               32'shc0028c9c, 32'shc00293b9, 32'shc0029ae0, 32'shc002a210, 32'shc002a94b, 32'shc002b08f, 32'shc002b7dd, 32'shc002bf35, 
               32'shc002c697, 32'shc002ce03, 32'shc002d579, 32'shc002dcf8, 32'shc002e482, 32'shc002ec15, 32'shc002f3b2, 32'shc002fb59, 
               32'shc003030a, 32'shc0030ac5, 32'shc0031289, 32'shc0031a58, 32'shc0032230, 32'shc0032a12, 32'shc00331fe, 32'shc00339f4, 
               32'shc00341f4, 32'shc00349fe, 32'shc0035211, 32'shc0035a2f, 32'shc0036256, 32'shc0036a87, 32'shc00372c2, 32'shc0037b07, 
               32'shc0038356, 32'shc0038baf, 32'shc0039411, 32'shc0039c7d, 32'shc003a4f4, 32'shc003ad74, 32'shc003b5fe, 32'shc003be91, 
               32'shc003c72f, 32'shc003cfd7, 32'shc003d888, 32'shc003e143, 32'shc003ea09, 32'shc003f2d8, 32'shc003fbb0, 32'shc0040493, 
               32'shc0040d80, 32'shc0041676, 32'shc0041f77, 32'shc0042881, 32'shc0043195, 32'shc0043ab3, 32'shc00443db, 32'shc0044d0d, 
               32'shc0045648, 32'shc0045f8d, 32'shc00468dd, 32'shc0047236, 32'shc0047b99, 32'shc0048506, 32'shc0048e7d, 32'shc00497fd, 
               32'shc004a188, 32'shc004ab1c, 32'shc004b4ba, 32'shc004be62, 32'shc004c814, 32'shc004d1d0, 32'shc004db96, 32'shc004e566, 
               32'shc004ef3f, 32'shc004f922, 32'shc005030f, 32'shc0050d06, 32'shc0051707, 32'shc0052112, 32'shc0052b27, 32'shc0053545, 
               32'shc0053f6e, 32'shc00549a0, 32'shc00553dc, 32'shc0055e22, 32'shc0056872, 32'shc00572cb, 32'shc0057d2f, 32'shc005879c, 
               32'shc0059214, 32'shc0059c95, 32'shc005a720, 32'shc005b1b5, 32'shc005bc54, 32'shc005c6fc, 32'shc005d1af, 32'shc005dc6b, 
               32'shc005e731, 32'shc005f201, 32'shc005fcdb, 32'shc00607bf, 32'shc00612ad, 32'shc0061da4, 32'shc00628a6, 32'shc00633b1, 
               32'shc0063ec6, 32'shc00649e5, 32'shc006550e, 32'shc0066041, 32'shc0066b7d, 32'shc00676c4, 32'shc0068214, 32'shc0068d6f, 
               32'shc00698d3, 32'shc006a441, 32'shc006afb8, 32'shc006bb3a, 32'shc006c6c6, 32'shc006d25b, 32'shc006ddfa, 32'shc006e9a3, 
               32'shc006f556, 32'shc0070113, 32'shc0070cda, 32'shc00718ab, 32'shc0072485, 32'shc0073069, 32'shc0073c58, 32'shc0074850, 
               32'shc0075452, 32'shc007605d, 32'shc0076c73, 32'shc0077893, 32'shc00784bc, 32'shc00790ef, 32'shc0079d2c, 32'shc007a973, 
               32'shc007b5c4, 32'shc007c21f, 32'shc007ce83, 32'shc007daf2, 32'shc007e76a, 32'shc007f3ec, 32'shc0080078, 32'shc0080d0e, 
               32'shc00819ae, 32'shc0082658, 32'shc008330b, 32'shc0083fc8, 32'shc0084c90, 32'shc0085961, 32'shc008663c, 32'shc0087321, 
               32'shc008800f, 32'shc0088d08, 32'shc0089a0a, 32'shc008a716, 32'shc008b42d, 32'shc008c14d, 32'shc008ce76, 32'shc008dbaa, 
               32'shc008e8e8, 32'shc008f62f, 32'shc0090381, 32'shc00910dc, 32'shc0091e41, 32'shc0092bb0, 32'shc0093929, 32'shc00946ab, 
               32'shc0095438, 32'shc00961ce, 32'shc0096f6e, 32'shc0097d18, 32'shc0098acc, 32'shc009988a, 32'shc009a652, 32'shc009b423, 
               32'shc009c1ff, 32'shc009cfe4, 32'shc009ddd3, 32'shc009ebcc, 32'shc009f9cf, 32'shc00a07dc, 32'shc00a15f3, 32'shc00a2413, 
               32'shc00a323d, 32'shc00a4072, 32'shc00a4eb0, 32'shc00a5cf8, 32'shc00a6b49, 32'shc00a79a5, 32'shc00a880a, 32'shc00a967a, 
               32'shc00aa4f3, 32'shc00ab376, 32'shc00ac203, 32'shc00ad09a, 32'shc00adf3b, 32'shc00aede5, 32'shc00afc9a, 32'shc00b0b58, 
               32'shc00b1a20, 32'shc00b28f2, 32'shc00b37ce, 32'shc00b46b4, 32'shc00b55a3, 32'shc00b649d, 32'shc00b73a0, 32'shc00b82ad, 
               32'shc00b91c4, 32'shc00ba0e5, 32'shc00bb010, 32'shc00bbf44, 32'shc00bce83, 32'shc00bddcb, 32'shc00bed1e, 32'shc00bfc7a, 
               32'shc00c0be0, 32'shc00c1b4f, 32'shc00c2ac9, 32'shc00c3a4d, 32'shc00c49da, 32'shc00c5971, 32'shc00c6912, 32'shc00c78bd, 
               32'shc00c8872, 32'shc00c9831, 32'shc00ca7f9, 32'shc00cb7cc, 32'shc00cc7a8, 32'shc00cd78e, 32'shc00ce77e, 32'shc00cf778, 
               32'shc00d077c, 32'shc00d178a, 32'shc00d27a1, 32'shc00d37c2, 32'shc00d47ed, 32'shc00d5823, 32'shc00d6861, 32'shc00d78aa, 
               32'shc00d88fd, 32'shc00d9959, 32'shc00da9c0, 32'shc00dba30, 32'shc00dcaaa, 32'shc00ddb2e, 32'shc00debbc, 32'shc00dfc53, 
               32'shc00e0cf5, 32'shc00e1da0, 32'shc00e2e56, 32'shc00e3f15, 32'shc00e4fde, 32'shc00e60b0, 32'shc00e718d, 32'shc00e8274, 
               32'shc00e9364, 32'shc00ea45e, 32'shc00eb562, 32'shc00ec670, 32'shc00ed788, 32'shc00ee8aa, 32'shc00ef9d6, 32'shc00f0b0b, 
               32'shc00f1c4a, 32'shc00f2d93, 32'shc00f3ee6, 32'shc00f5043, 32'shc00f61aa, 32'shc00f731b, 32'shc00f8495, 32'shc00f9619, 
               32'shc00fa7a8, 32'shc00fb940, 32'shc00fcae2, 32'shc00fdc8d, 32'shc00fee43, 32'shc0100002, 32'shc01011cc, 32'shc010239f, 
               32'shc010357c, 32'shc0104763, 32'shc0105954, 32'shc0106b4e, 32'shc0107d53, 32'shc0108f61, 32'shc010a179, 32'shc010b39b, 
               32'shc010c5c7, 32'shc010d7fd, 32'shc010ea3d, 32'shc010fc86, 32'shc0110eda, 32'shc0112137, 32'shc011339e, 32'shc011460f, 
               32'shc011588a, 32'shc0116b0e, 32'shc0117d9d, 32'shc0119035, 32'shc011a2d8, 32'shc011b584, 32'shc011c83a, 32'shc011daf9, 
               32'shc011edc3, 32'shc0120097, 32'shc0121374, 32'shc012265b, 32'shc012394c, 32'shc0124c47, 32'shc0125f4c, 32'shc012725b, 
               32'shc0128574, 32'shc0129896, 32'shc012abc2, 32'shc012bef8, 32'shc012d238, 32'shc012e582, 32'shc012f8d6, 32'shc0130c33, 
               32'shc0131f9b, 32'shc013330c, 32'shc0134687, 32'shc0135a0c, 32'shc0136d9b, 32'shc0138134, 32'shc01394d6, 32'shc013a883, 
               32'shc013bc39, 32'shc013cff9, 32'shc013e3c3, 32'shc013f797, 32'shc0140b75, 32'shc0141f5c, 32'shc014334e, 32'shc0144749, 
               32'shc0145b4e, 32'shc0146f5d, 32'shc0148376, 32'shc0149799, 32'shc014abc5, 32'shc014bffc, 32'shc014d43c, 32'shc014e886, 
               32'shc014fcda, 32'shc0151138, 32'shc01525a0, 32'shc0153a11, 32'shc0154e8d, 32'shc0156312, 32'shc01577a1, 32'shc0158c3a, 
               32'shc015a0dd, 32'shc015b58a, 32'shc015ca40, 32'shc015df01, 32'shc015f3cb, 32'shc016089f, 32'shc0161d7d, 32'shc0163265, 
               32'shc0164757, 32'shc0165c52, 32'shc0167158, 32'shc0168667, 32'shc0169b80, 32'shc016b0a3, 32'shc016c5d0, 32'shc016db07, 
               32'shc016f047, 32'shc0170591, 32'shc0171ae6, 32'shc0173044, 32'shc01745ac, 32'shc0175b1e, 32'shc0177099, 32'shc017861f, 
               32'shc0179bae, 32'shc017b148, 32'shc017c6eb, 32'shc017dc98, 32'shc017f24e, 32'shc018080f, 32'shc0181dda, 32'shc01833ae, 
               32'shc018498c, 32'shc0185f74, 32'shc0187566, 32'shc0188b62, 32'shc018a168, 32'shc018b777, 32'shc018cd91, 32'shc018e3b4, 
               32'shc018f9e1, 32'shc0191018, 32'shc0192659, 32'shc0193ca3, 32'shc01952f8, 32'shc0196956, 32'shc0197fbe, 32'shc0199630, 
               32'shc019acac, 32'shc019c332, 32'shc019d9c2, 32'shc019f05b, 32'shc01a06fe, 32'shc01a1dac, 32'shc01a3463, 32'shc01a4b24, 
               32'shc01a61ee, 32'shc01a78c3, 32'shc01a8fa1, 32'shc01aa68a, 32'shc01abd7c, 32'shc01ad478, 32'shc01aeb7e, 32'shc01b028d, 
               32'shc01b19a7, 32'shc01b30ca, 32'shc01b47f8, 32'shc01b5f2f, 32'shc01b7670, 32'shc01b8dbb, 32'shc01ba50f, 32'shc01bbc6e, 
               32'shc01bd3d6, 32'shc01beb48, 32'shc01c02c5, 32'shc01c1a4b, 32'shc01c31da, 32'shc01c4974, 32'shc01c6118, 32'shc01c78c5, 
               32'shc01c907c, 32'shc01ca83d, 32'shc01cc008, 32'shc01cd7dd, 32'shc01cefbb, 32'shc01d07a4, 32'shc01d1f96, 32'shc01d3792, 
               32'shc01d4f99, 32'shc01d67a8, 32'shc01d7fc2, 32'shc01d97e6, 32'shc01db013, 32'shc01dc84a, 32'shc01de08c, 32'shc01df8d7, 
               32'shc01e112b, 32'shc01e298a, 32'shc01e41f3, 32'shc01e5a65, 32'shc01e72e1, 32'shc01e8b67, 32'shc01ea3f7, 32'shc01ebc91, 
               32'shc01ed535, 32'shc01eede2, 32'shc01f069a, 32'shc01f1f5b, 32'shc01f3826, 32'shc01f50fb, 32'shc01f69da, 32'shc01f82c2, 
               32'shc01f9bb5, 32'shc01fb4b1, 32'shc01fcdb7, 32'shc01fe6c7, 32'shc01fffe1, 32'shc0201905, 32'shc0203232, 32'shc0204b6a, 
               32'shc02064ab, 32'shc0207df6, 32'shc020974b, 32'shc020b0aa, 32'shc020ca13, 32'shc020e385, 32'shc020fd02, 32'shc0211688, 
               32'shc0213018, 32'shc02149b2, 32'shc0216356, 32'shc0217d03, 32'shc02196bb, 32'shc021b07c, 32'shc021ca47, 32'shc021e41c, 
               32'shc021fdfb, 32'shc02217e4, 32'shc02231d6, 32'shc0224bd3, 32'shc02265d9, 32'shc0227fe9, 32'shc0229a03, 32'shc022b427, 
               32'shc022ce54, 32'shc022e88c, 32'shc02302cd, 32'shc0231d18, 32'shc023376e, 32'shc02351cc, 32'shc0236c35, 32'shc02386a8, 
               32'shc023a124, 32'shc023bbab, 32'shc023d63b, 32'shc023f0d5, 32'shc0240b78, 32'shc0242626, 32'shc02440de, 32'shc0245b9f, 
               32'shc024766a, 32'shc024913f, 32'shc024ac1e, 32'shc024c707, 32'shc024e1fa, 32'shc024fcf6, 32'shc02517fc, 32'shc025330d, 
               32'shc0254e27, 32'shc025694a, 32'shc0258478, 32'shc0259fb0, 32'shc025baf1, 32'shc025d63c, 32'shc025f191, 32'shc0260cf0, 
               32'shc0262859, 32'shc02643cc, 32'shc0265f48, 32'shc0267acf, 32'shc026965f, 32'shc026b1f9, 32'shc026cd9d, 32'shc026e94a, 
               32'shc0270502, 32'shc02720c3, 32'shc0273c8e, 32'shc0275864, 32'shc0277442, 32'shc027902b, 32'shc027ac1e, 32'shc027c81a, 
               32'shc027e421, 32'shc0280031, 32'shc0281c4b, 32'shc028386f, 32'shc028549c, 32'shc02870d4, 32'shc0288d15, 32'shc028a961, 
               32'shc028c5b6, 32'shc028e215, 32'shc028fe7d, 32'shc0291af0, 32'shc029376c, 32'shc02953f3, 32'shc0297083, 32'shc0298d1d, 
               32'shc029a9c1, 32'shc029c66e, 32'shc029e326, 32'shc029ffe7, 32'shc02a1cb2, 32'shc02a3988, 32'shc02a5666, 32'shc02a734f, 
               32'shc02a9042, 32'shc02aad3e, 32'shc02aca44, 32'shc02ae755, 32'shc02b046f, 32'shc02b2192, 32'shc02b3ec0, 32'shc02b5bf8, 
               32'shc02b7939, 32'shc02b9684, 32'shc02bb3d9, 32'shc02bd138, 32'shc02beea1, 32'shc02c0c13, 32'shc02c2990, 32'shc02c4716, 
               32'shc02c64a6, 32'shc02c8240, 32'shc02c9fe4, 32'shc02cbd91, 32'shc02cdb49, 32'shc02cf90a, 32'shc02d16d5, 32'shc02d34aa, 
               32'shc02d5289, 32'shc02d7072, 32'shc02d8e64, 32'shc02dac61, 32'shc02dca67, 32'shc02de877, 32'shc02e0691, 32'shc02e24b4, 
               32'shc02e42e2, 32'shc02e6119, 32'shc02e7f5b, 32'shc02e9da6, 32'shc02ebbfb, 32'shc02eda59, 32'shc02ef8c2, 32'shc02f1734, 
               32'shc02f35b1, 32'shc02f5437, 32'shc02f72c7, 32'shc02f9161, 32'shc02fb004, 32'shc02fceb2, 32'shc02fed69, 32'shc0300c2a, 
               32'shc0302af5, 32'shc03049ca, 32'shc03068a9, 32'shc0308792, 32'shc030a684, 32'shc030c580, 32'shc030e486, 32'shc0310396, 
               32'shc03122b0, 32'shc03141d3, 32'shc0316101, 32'shc0318038, 32'shc0319f79, 32'shc031bec4, 32'shc031de19, 32'shc031fd78, 
               32'shc0321ce0, 32'shc0323c52, 32'shc0325bcf, 32'shc0327b55, 32'shc0329ae4, 32'shc032ba7e, 32'shc032da22, 32'shc032f9cf, 
               32'shc0331986, 32'shc0333947, 32'shc0335912, 32'shc03378e7, 32'shc03398c5, 32'shc033b8ad, 32'shc033d8a0, 32'shc033f89c, 
               32'shc03418a2, 32'shc03438b1, 32'shc03458cb, 32'shc03478ee, 32'shc034991c, 32'shc034b953, 32'shc034d994, 32'shc034f9de, 
               32'shc0351a33, 32'shc0353a91, 32'shc0355afa, 32'shc0357b6c, 32'shc0359be8, 32'shc035bc6d, 32'shc035dcfd, 32'shc035fd96, 
               32'shc0361e3a, 32'shc0363ee7, 32'shc0365f9e, 32'shc036805f, 32'shc036a129, 32'shc036c1fe, 32'shc036e2dc, 32'shc03703c4, 
               32'shc03724b6, 32'shc03745b2, 32'shc03766b8, 32'shc03787c7, 32'shc037a8e1, 32'shc037ca04, 32'shc037eb31, 32'shc0380c68, 
               32'shc0382da8, 32'shc0384ef3, 32'shc0387047, 32'shc03891a5, 32'shc038b30d, 32'shc038d47f, 32'shc038f5fb, 32'shc0391780, 
               32'shc0393910, 32'shc0395aa9, 32'shc0397c4c, 32'shc0399df9, 32'shc039bfaf, 32'shc039e170, 32'shc03a033a, 32'shc03a250e, 
               32'shc03a46ed, 32'shc03a68d4, 32'shc03a8ac6, 32'shc03aacc2, 32'shc03acec7, 32'shc03af0d6, 32'shc03b12ef, 32'shc03b3512, 
               32'shc03b573f, 32'shc03b7975, 32'shc03b9bb6, 32'shc03bbe00, 32'shc03be054, 32'shc03c02b2, 32'shc03c251a, 32'shc03c478b, 
               32'shc03c6a07, 32'shc03c8c8c, 32'shc03caf1b, 32'shc03cd1b4, 32'shc03cf456, 32'shc03d1703, 32'shc03d39b9, 32'shc03d5c79, 
               32'shc03d7f44, 32'shc03da217, 32'shc03dc4f5, 32'shc03de7dd, 32'shc03e0ace, 32'shc03e2dc9, 32'shc03e50ce, 32'shc03e73dd, 
               32'shc03e96f6, 32'shc03eba18, 32'shc03edd45, 32'shc03f007b, 32'shc03f23bb, 32'shc03f4705, 32'shc03f6a58, 32'shc03f8db6, 
               32'shc03fb11d, 32'shc03fd48f, 32'shc03ff80a, 32'shc0401b8e, 32'shc0403f1d, 32'shc04062b6, 32'shc0408658, 32'shc040aa04, 
               32'shc040cdba, 32'shc040f17a, 32'shc0411544, 32'shc0413917, 32'shc0415cf4, 32'shc04180dc, 32'shc041a4cd, 32'shc041c8c7, 
               32'shc041eccc, 32'shc04210da, 32'shc04234f3, 32'shc0425915, 32'shc0427d41, 32'shc042a177, 32'shc042c5b6, 32'shc042ea00, 
               32'shc0430e53, 32'shc04332b0, 32'shc0435717, 32'shc0437b88, 32'shc043a002, 32'shc043c487, 32'shc043e915, 32'shc0440dad, 
               32'shc044324f, 32'shc04456fb, 32'shc0447bb0, 32'shc044a070, 32'shc044c539, 32'shc044ea0c, 32'shc0450ee9, 32'shc04533d0, 
               32'shc04558c0, 32'shc0457dba, 32'shc045a2bf, 32'shc045c7cd, 32'shc045ece5, 32'shc0461206, 32'shc0463732, 32'shc0465c67, 
               32'shc04681a6, 32'shc046a6ef, 32'shc046cc42, 32'shc046f19f, 32'shc0471705, 32'shc0473c75, 32'shc04761ef, 32'shc0478773, 
               32'shc047ad01, 32'shc047d299, 32'shc047f83a, 32'shc0481de5, 32'shc048439b, 32'shc0486959, 32'shc0488f22, 32'shc048b4f5, 
               32'shc048dad1, 32'shc04900b7, 32'shc04926a7, 32'shc0494ca1, 32'shc04972a5, 32'shc04998b2, 32'shc049beca, 32'shc049e4eb, 
               32'shc04a0b16, 32'shc04a314b, 32'shc04a5789, 32'shc04a7dd2, 32'shc04aa424, 32'shc04aca80, 32'shc04af0e6, 32'shc04b1756, 
               32'shc04b3dcf, 32'shc04b6453, 32'shc04b8ae0, 32'shc04bb177, 32'shc04bd818, 32'shc04bfec3, 32'shc04c2577, 32'shc04c4c36, 
               32'shc04c72fe, 32'shc04c99d0, 32'shc04cc0ac, 32'shc04ce791, 32'shc04d0e81, 32'shc04d357a, 32'shc04d5c7d, 32'shc04d838a, 
               32'shc04daaa1, 32'shc04dd1c1, 32'shc04df8ec, 32'shc04e2020, 32'shc04e475e, 32'shc04e6ea6, 32'shc04e95f8, 32'shc04ebd53, 
               32'shc04ee4b8, 32'shc04f0c28, 32'shc04f33a1, 32'shc04f5b23, 32'shc04f82b0, 32'shc04faa46, 32'shc04fd1e7, 32'shc04ff991, 
               32'shc0502145, 32'shc0504902, 32'shc05070ca, 32'shc050989b, 32'shc050c077, 32'shc050e85c, 32'shc051104a, 32'shc0513843, 
               32'shc0516045, 32'shc0518852, 32'shc051b068, 32'shc051d888, 32'shc05200b2, 32'shc05228e5, 32'shc0525123, 32'shc052796a, 
               32'shc052a1bb, 32'shc052ca16, 32'shc052f27a, 32'shc0531ae9, 32'shc0534361, 32'shc0536be3, 32'shc053946f, 32'shc053bd05, 
               32'shc053e5a5, 32'shc0540e4e, 32'shc0543701, 32'shc0545fbe, 32'shc0548885, 32'shc054b156, 32'shc054da30, 32'shc0550315, 
               32'shc0552c03, 32'shc05554fb, 32'shc0557dfd, 32'shc055a708, 32'shc055d01e, 32'shc055f93d, 32'shc0562266, 32'shc0564b99, 
               32'shc05674d6, 32'shc0569e1c, 32'shc056c76c, 32'shc056f0c7, 32'shc0571a2b, 32'shc0574398, 32'shc0576d10, 32'shc0579691, 
               32'shc057c01d, 32'shc057e9b2, 32'shc0581350, 32'shc0583cf9, 32'shc05866ac, 32'shc0589068, 32'shc058ba2e, 32'shc058e3fe, 
               32'shc0590dd8, 32'shc05937bb, 32'shc05961a9, 32'shc0598ba0, 32'shc059b5a1, 32'shc059dfac, 32'shc05a09c0, 32'shc05a33df, 
               32'shc05a5e07, 32'shc05a8839, 32'shc05ab275, 32'shc05adcbb, 32'shc05b070a, 32'shc05b3164, 32'shc05b5bc7, 32'shc05b8634, 
               32'shc05bb0ab, 32'shc05bdb2b, 32'shc05c05b6, 32'shc05c304a, 32'shc05c5ae8, 32'shc05c8590, 32'shc05cb042, 32'shc05cdafd, 
               32'shc05d05c3, 32'shc05d3092, 32'shc05d5b6b, 32'shc05d864d, 32'shc05db13a, 32'shc05ddc30, 32'shc05e0730, 32'shc05e323a, 
               32'shc05e5d4e, 32'shc05e886c, 32'shc05eb393, 32'shc05edec5, 32'shc05f0a00, 32'shc05f3545, 32'shc05f6093, 32'shc05f8bec, 
               32'shc05fb74e, 32'shc05fe2ba, 32'shc0600e30, 32'shc06039b0, 32'shc060653a, 32'shc06090cd, 32'shc060bc6a, 32'shc060e811, 
               32'shc06113c2, 32'shc0613f7d, 32'shc0616b41, 32'shc061970f, 32'shc061c2e7, 32'shc061eec9, 32'shc0621ab5, 32'shc06246aa, 
               32'shc06272aa, 32'shc0629eb3, 32'shc062cac6, 32'shc062f6e2, 32'shc0632309, 32'shc0634f39, 32'shc0637b73, 32'shc063a7b7, 
               32'shc063d405, 32'shc064005d, 32'shc0642cbe, 32'shc0645929, 32'shc064859e, 32'shc064b21d, 32'shc064dea6, 32'shc0650b38, 
               32'shc06537d4, 32'shc065647b, 32'shc065912a, 32'shc065bde4, 32'shc065eaa8, 32'shc0661775, 32'shc066444c, 32'shc066712d, 
               32'shc0669e18, 32'shc066cb0c, 32'shc066f80a, 32'shc0672513, 32'shc0675225, 32'shc0677f40, 32'shc067ac66, 32'shc067d995, 
               32'shc06806ce, 32'shc0683411, 32'shc068615e, 32'shc0688eb5, 32'shc068bc15, 32'shc068e97f, 32'shc06916f3, 32'shc0694471, 
               32'shc06971f9, 32'shc0699f8a, 32'shc069cd26, 32'shc069facb, 32'shc06a2879, 32'shc06a5632, 32'shc06a83f5, 32'shc06ab1c1, 
               32'shc06adf97, 32'shc06b0d77, 32'shc06b3b60, 32'shc06b6954, 32'shc06b9751, 32'shc06bc558, 32'shc06bf369, 32'shc06c2184, 
               32'shc06c4fa8, 32'shc06c7dd7, 32'shc06cac0f, 32'shc06cda51, 32'shc06d089d, 32'shc06d36f2, 32'shc06d6551, 32'shc06d93bb, 
               32'shc06dc22e, 32'shc06df0aa, 32'shc06e1f31, 32'shc06e4dc1, 32'shc06e7c5b, 32'shc06eaaff, 32'shc06ed9ad, 32'shc06f0865, 
               32'shc06f3726, 32'shc06f65f1, 32'shc06f94c6, 32'shc06fc3a5, 32'shc06ff28e, 32'shc0702180, 32'shc070507c, 32'shc0707f82, 
               32'shc070ae92, 32'shc070ddab, 32'shc0710ccf, 32'shc0713bfc, 32'shc0716b33, 32'shc0719a74, 32'shc071c9be, 32'shc071f913, 
               32'shc0722871, 32'shc07257d9, 32'shc072874b, 32'shc072b6c6, 32'shc072e64c, 32'shc07315db, 32'shc0734574, 32'shc0737517, 
               32'shc073a4c3, 32'shc073d47a, 32'shc074043a, 32'shc0743404, 32'shc07463d8, 32'shc07493b5, 32'shc074c39d, 32'shc074f38e, 
               32'shc0752389, 32'shc075538e, 32'shc075839c, 32'shc075b3b5, 32'shc075e3d7, 32'shc0761403, 32'shc0764439, 32'shc0767478, 
               32'shc076a4c2, 32'shc076d515, 32'shc0770572, 32'shc07735d9, 32'shc0776649, 32'shc07796c4, 32'shc077c748, 32'shc077f7d6, 
               32'shc078286e, 32'shc078590f, 32'shc07889bb, 32'shc078ba70, 32'shc078eb2f, 32'shc0791bf7, 32'shc0794cca, 32'shc0797da6, 
               32'shc079ae8c, 32'shc079df7c, 32'shc07a1076, 32'shc07a417a, 32'shc07a7287, 32'shc07aa39e, 32'shc07ad4bf, 32'shc07b05ea, 
               32'shc07b371e, 32'shc07b685d, 32'shc07b99a5, 32'shc07bcaf7, 32'shc07bfc52, 32'shc07c2db8, 32'shc07c5f27, 32'shc07c90a0, 
               32'shc07cc223, 32'shc07cf3b0, 32'shc07d2546, 32'shc07d56e6, 32'shc07d8890, 32'shc07dba44, 32'shc07dec02, 32'shc07e1dc9, 
               32'shc07e4f9b, 32'shc07e8176, 32'shc07eb35a, 32'shc07ee549, 32'shc07f1741, 32'shc07f4944, 32'shc07f7b50, 32'shc07fad65, 
               32'shc07fdf85, 32'shc08011ae, 32'shc08043e1, 32'shc080761e, 32'shc080a865, 32'shc080dab6, 32'shc0810d10, 32'shc0813f74, 
               32'shc08171e2, 32'shc081a45a, 32'shc081d6db, 32'shc0820966, 32'shc0823bfb, 32'shc0826e9a, 32'shc082a143, 32'shc082d3f5, 
               32'shc08306b2, 32'shc0833978, 32'shc0836c47, 32'shc0839f21, 32'shc083d204, 32'shc08404f2, 32'shc08437e9, 32'shc0846ae9, 
               32'shc0849df4, 32'shc084d108, 32'shc0850426, 32'shc085374e, 32'shc0856a80, 32'shc0859dbc, 32'shc085d101, 32'shc0860450, 
               32'shc08637a9, 32'shc0866b0c, 32'shc0869e78, 32'shc086d1ee, 32'shc087056e, 32'shc08738f8, 32'shc0876c8c, 32'shc087a029, 
               32'shc087d3d0, 32'shc0880781, 32'shc0883b3c, 32'shc0886f00, 32'shc088a2cf, 32'shc088d6a7, 32'shc0890a89, 32'shc0893e75, 
               32'shc089726a, 32'shc089a669, 32'shc089da72, 32'shc08a0e85, 32'shc08a42a2, 32'shc08a76c8, 32'shc08aaaf8, 32'shc08adf32, 
               32'shc08b1376, 32'shc08b47c4, 32'shc08b7c1b, 32'shc08bb07c, 32'shc08be4e7, 32'shc08c195c, 32'shc08c4dda, 32'shc08c8262, 
               32'shc08cb6f5, 32'shc08ceb90, 32'shc08d2036, 32'shc08d54e5, 32'shc08d899f, 32'shc08dbe62, 32'shc08df32e, 32'shc08e2805, 
               32'shc08e5ce5, 32'shc08e91cf, 32'shc08ec6c3, 32'shc08efbc1, 32'shc08f30c8, 32'shc08f65da, 32'shc08f9af5, 32'shc08fd019, 
               32'shc0900548, 32'shc0903a80, 32'shc0906fc3, 32'shc090a50e, 32'shc090da64, 32'shc0910fc4, 32'shc091452d, 32'shc0917aa0, 
               32'shc091b01d, 32'shc091e5a4, 32'shc0921b34, 32'shc09250ce, 32'shc0928672, 32'shc092bc20, 32'shc092f1d7, 32'shc0932799, 
               32'shc0935d64, 32'shc0939339, 32'shc093c917, 32'shc093ff00, 32'shc09434f2, 32'shc0946aee, 32'shc094a0f4, 32'shc094d703, 
               32'shc0950d1d, 32'shc0954340, 32'shc095796d, 32'shc095afa4, 32'shc095e5e4, 32'shc0961c2e, 32'shc0965282, 32'shc09688e0, 
               32'shc096bf48, 32'shc096f5b9, 32'shc0972c34, 32'shc09762b9, 32'shc0979948, 32'shc097cfe0, 32'shc0980683, 32'shc0983d2f, 
               32'shc09873e4, 32'shc098aaa4, 32'shc098e16d, 32'shc0991840, 32'shc0994f1d, 32'shc0998604, 32'shc099bcf5, 32'shc099f3ef, 
               32'shc09a2af3, 32'shc09a6201, 32'shc09a9918, 32'shc09ad03a, 32'shc09b0765, 32'shc09b3e9a, 32'shc09b75d8, 32'shc09bad21, 
               32'shc09be473, 32'shc09c1bcf, 32'shc09c5335, 32'shc09c8aa4, 32'shc09cc21e, 32'shc09cf9a1, 32'shc09d312e, 32'shc09d68c4, 
               32'shc09da065, 32'shc09dd80f, 32'shc09e0fc3, 32'shc09e4781, 32'shc09e7f48, 32'shc09eb71a, 32'shc09eeef5, 32'shc09f26da, 
               32'shc09f5ec8, 32'shc09f96c1, 32'shc09fcec3, 32'shc0a006cf, 32'shc0a03ee4, 32'shc0a07704, 32'shc0a0af2d, 32'shc0a0e760, 
               32'shc0a11f9d, 32'shc0a157e4, 32'shc0a19034, 32'shc0a1c88e, 32'shc0a200f2, 32'shc0a23960, 32'shc0a271d7, 32'shc0a2aa58, 
               32'shc0a2e2e3, 32'shc0a31b78, 32'shc0a35417, 32'shc0a38cbf, 32'shc0a3c571, 32'shc0a3fe2d, 32'shc0a436f3, 32'shc0a46fc2, 
               32'shc0a4a89b, 32'shc0a4e17e, 32'shc0a51a6b, 32'shc0a55361, 32'shc0a58c62, 32'shc0a5c56c, 32'shc0a5fe7f, 32'shc0a6379d, 
               32'shc0a670c4, 32'shc0a6a9f5, 32'shc0a6e330, 32'shc0a71c75, 32'shc0a755c3, 32'shc0a78f1b, 32'shc0a7c87d, 32'shc0a801e9, 
               32'shc0a83b5e, 32'shc0a874de, 32'shc0a8ae67, 32'shc0a8e7f9, 32'shc0a92196, 32'shc0a95b3c, 32'shc0a994ec, 32'shc0a9cea6, 
               32'shc0aa086a, 32'shc0aa4237, 32'shc0aa7c0e, 32'shc0aab5ef, 32'shc0aaefda, 32'shc0ab29ce, 32'shc0ab63cd, 32'shc0ab9dd5, 
               32'shc0abd7e6, 32'shc0ac1202, 32'shc0ac4c27, 32'shc0ac8656, 32'shc0acc08f, 32'shc0acfad2, 32'shc0ad351e, 32'shc0ad6f74, 
               32'shc0ada9d4, 32'shc0ade43e, 32'shc0ae1eb1, 32'shc0ae592e, 32'shc0ae93b5, 32'shc0aece46, 32'shc0af08e0, 32'shc0af4385, 
               32'shc0af7e33, 32'shc0afb8ea, 32'shc0aff3ac, 32'shc0b02e77, 32'shc0b0694c, 32'shc0b0a42b, 32'shc0b0df13, 32'shc0b11a06, 
               32'shc0b15502, 32'shc0b19008, 32'shc0b1cb17, 32'shc0b20631, 32'shc0b24154, 32'shc0b27c81, 32'shc0b2b7b8, 32'shc0b2f2f8, 
               32'shc0b32e42, 32'shc0b36996, 32'shc0b3a4f4, 32'shc0b3e05b, 32'shc0b41bcd, 32'shc0b45748, 32'shc0b492cc, 32'shc0b4ce5b, 
               32'shc0b509f3, 32'shc0b54595, 32'shc0b58141, 32'shc0b5bcf7, 32'shc0b5f8b6, 32'shc0b6347f, 32'shc0b67052, 32'shc0b6ac2e, 
               32'shc0b6e815, 32'shc0b72405, 32'shc0b75fff, 32'shc0b79c02, 32'shc0b7d810, 32'shc0b81427, 32'shc0b85048, 32'shc0b88c73, 
               32'shc0b8c8a7, 32'shc0b904e5, 32'shc0b9412d, 32'shc0b97d7f, 32'shc0b9b9da, 32'shc0b9f640, 32'shc0ba32af, 32'shc0ba6f27, 
               32'shc0baabaa, 32'shc0bae836, 32'shc0bb24cc, 32'shc0bb616c, 32'shc0bb9e15, 32'shc0bbdac9, 32'shc0bc1786, 32'shc0bc544d, 
               32'shc0bc911d, 32'shc0bccdf7, 32'shc0bd0adb, 32'shc0bd47c9, 32'shc0bd84c1, 32'shc0bdc1c2, 32'shc0bdfecd, 32'shc0be3be2, 
               32'shc0be7901, 32'shc0beb629, 32'shc0bef35b, 32'shc0bf3097, 32'shc0bf6ddd, 32'shc0bfab2c, 32'shc0bfe885, 32'shc0c025e8, 
               32'shc0c06355, 32'shc0c0a0cb, 32'shc0c0de4b, 32'shc0c11bd5, 32'shc0c15969, 32'shc0c19706, 32'shc0c1d4ad, 32'shc0c2125e, 
               32'shc0c25019, 32'shc0c28ddd, 32'shc0c2cbab, 32'shc0c30983, 32'shc0c34765, 32'shc0c38550, 32'shc0c3c346, 32'shc0c40144, 
               32'shc0c43f4d, 32'shc0c47d60, 32'shc0c4bb7c, 32'shc0c4f9a2, 32'shc0c537d1, 32'shc0c5760b, 32'shc0c5b44e, 32'shc0c5f29b, 
               32'shc0c630f2, 32'shc0c66f52, 32'shc0c6adbc, 32'shc0c6ec30, 32'shc0c72aae, 32'shc0c76935, 32'shc0c7a7c6, 32'shc0c7e661, 
               32'shc0c82506, 32'shc0c863b4, 32'shc0c8a26d, 32'shc0c8e12f, 32'shc0c91ffa, 32'shc0c95ed0, 32'shc0c99daf, 32'shc0c9dc98, 
               32'shc0ca1b8a, 32'shc0ca5a87, 32'shc0ca998d, 32'shc0cad89d, 32'shc0cb17b7, 32'shc0cb56da, 32'shc0cb9607, 32'shc0cbd53e, 
               32'shc0cc147f, 32'shc0cc53c9, 32'shc0cc931d, 32'shc0ccd27b, 32'shc0cd11e3, 32'shc0cd5154, 32'shc0cd90cf, 32'shc0cdd054, 
               32'shc0ce0fe3, 32'shc0ce4f7b, 32'shc0ce8f1d, 32'shc0cecec9, 32'shc0cf0e7f, 32'shc0cf4e3e, 32'shc0cf8e07, 32'shc0cfcdda, 
               32'shc0d00db6, 32'shc0d04d9d, 32'shc0d08d8d, 32'shc0d0cd87, 32'shc0d10d8a, 32'shc0d14d97, 32'shc0d18dae, 32'shc0d1cdcf, 
               32'shc0d20dfa, 32'shc0d24e2e, 32'shc0d28e6c, 32'shc0d2ceb4, 32'shc0d30f05, 32'shc0d34f61, 32'shc0d38fc6, 32'shc0d3d034, 
               32'shc0d410ad, 32'shc0d4512f, 32'shc0d491bb, 32'shc0d4d251, 32'shc0d512f0, 32'shc0d55399, 32'shc0d5944c, 32'shc0d5d509, 
               32'shc0d615cf, 32'shc0d6569f, 32'shc0d69779, 32'shc0d6d85d, 32'shc0d7194a, 32'shc0d75a41, 32'shc0d79b42, 32'shc0d7dc4d, 
               32'shc0d81d61, 32'shc0d85e7f, 32'shc0d89fa7, 32'shc0d8e0d8, 32'shc0d92214, 32'shc0d96359, 32'shc0d9a4a7, 32'shc0d9e600, 
               32'shc0da2762, 32'shc0da68ce, 32'shc0daaa44, 32'shc0daebc3, 32'shc0db2d4c, 32'shc0db6edf, 32'shc0dbb07c, 32'shc0dbf222, 
               32'shc0dc33d2, 32'shc0dc758c, 32'shc0dcb750, 32'shc0dcf91d, 32'shc0dd3af4, 32'shc0dd7cd5, 32'shc0ddbec0, 32'shc0de00b4, 
               32'shc0de42b2, 32'shc0de84ba, 32'shc0dec6cb, 32'shc0df08e6, 32'shc0df4b0b, 32'shc0df8d3a, 32'shc0dfcf73, 32'shc0e011b5, 
               32'shc0e05401, 32'shc0e09656, 32'shc0e0d8b6, 32'shc0e11b1f, 32'shc0e15d92, 32'shc0e1a00e, 32'shc0e1e294, 32'shc0e22525, 
               32'shc0e267be, 32'shc0e2aa62, 32'shc0e2ed0f, 32'shc0e32fc6, 32'shc0e37287, 32'shc0e3b551, 32'shc0e3f825, 32'shc0e43b03, 
               32'shc0e47deb, 32'shc0e4c0dc, 32'shc0e503d7, 32'shc0e546dc, 32'shc0e589eb, 32'shc0e5cd03, 32'shc0e61025, 32'shc0e65351, 
               32'shc0e69686, 32'shc0e6d9c5, 32'shc0e71d0e, 32'shc0e76061, 32'shc0e7a3bd, 32'shc0e7e724, 32'shc0e82a93, 32'shc0e86e0d, 
               32'shc0e8b190, 32'shc0e8f51d, 32'shc0e938b4, 32'shc0e97c55, 32'shc0e9bfff, 32'shc0ea03b3, 32'shc0ea4771, 32'shc0ea8b38, 
               32'shc0eacf09, 32'shc0eb12e4, 32'shc0eb56c9, 32'shc0eb9ab7, 32'shc0ebdeaf, 32'shc0ec22b1, 32'shc0ec66bc, 32'shc0ecaad2, 
               32'shc0eceef1, 32'shc0ed3319, 32'shc0ed774c, 32'shc0edbb88, 32'shc0edffce, 32'shc0ee441e, 32'shc0ee8877, 32'shc0eeccda, 
               32'shc0ef1147, 32'shc0ef55bd, 32'shc0ef9a3d, 32'shc0efdec7, 32'shc0f0235b, 32'shc0f067f9, 32'shc0f0aca0, 32'shc0f0f151, 
               32'shc0f1360b, 32'shc0f17acf, 32'shc0f1bf9d, 32'shc0f20475, 32'shc0f24957, 32'shc0f28e42, 32'shc0f2d337, 32'shc0f31836, 
               32'shc0f35d3e, 32'shc0f3a250, 32'shc0f3e76c, 32'shc0f42c91, 32'shc0f471c1, 32'shc0f4b6fa, 32'shc0f4fc3c, 32'shc0f54189, 
               32'shc0f586df, 32'shc0f5cc3f, 32'shc0f611a8, 32'shc0f6571c, 32'shc0f69c99, 32'shc0f6e220, 32'shc0f727b0, 32'shc0f76d4a, 
               32'shc0f7b2ee, 32'shc0f7f89c, 32'shc0f83e53, 32'shc0f88414, 32'shc0f8c9df, 32'shc0f90fb4, 32'shc0f95592, 32'shc0f99b7a, 
               32'shc0f9e16b, 32'shc0fa2767, 32'shc0fa6d6c, 32'shc0fab37b, 32'shc0faf993, 32'shc0fb3fb6, 32'shc0fb85e2, 32'shc0fbcc17, 
               32'shc0fc1257, 32'shc0fc58a0, 32'shc0fc9ef3, 32'shc0fce54f, 32'shc0fd2bb6, 32'shc0fd7226, 32'shc0fdb8a0, 32'shc0fdff23, 
               32'shc0fe45b0, 32'shc0fe8c47, 32'shc0fed2e8, 32'shc0ff1992, 32'shc0ff6046, 32'shc0ffa704, 32'shc0ffedcb, 32'shc100349c, 
               32'shc1007b77, 32'shc100c25c, 32'shc101094a, 32'shc1015042, 32'shc1019744, 32'shc101de50, 32'shc1022565, 32'shc1026c84, 
               32'shc102b3ac, 32'shc102fadf, 32'shc103421b, 32'shc1038960, 32'shc103d0b0, 32'shc1041809, 32'shc1045f6c, 32'shc104a6d8, 
               32'shc104ee4f, 32'shc10535cf, 32'shc1057d59, 32'shc105c4ec, 32'shc1060c89, 32'shc1065430, 32'shc1069be1, 32'shc106e39b, 
               32'shc1072b5f, 32'shc107732d, 32'shc107bb04, 32'shc10802e5, 32'shc1084ad0, 32'shc10892c5, 32'shc108dac3, 32'shc10922cb, 
               32'shc1096add, 32'shc109b2f8, 32'shc109fb1d, 32'shc10a434c, 32'shc10a8b85, 32'shc10ad3c7, 32'shc10b1c13, 32'shc10b6468, 
               32'shc10bacc8, 32'shc10bf531, 32'shc10c3da4, 32'shc10c8620, 32'shc10ccea6, 32'shc10d1736, 32'shc10d5fd0, 32'shc10da873, 
               32'shc10df120, 32'shc10e39d7, 32'shc10e8297, 32'shc10ecb62, 32'shc10f1435, 32'shc10f5d13, 32'shc10fa5fa, 32'shc10feeeb, 
               32'shc11037e6, 32'shc11080ea, 32'shc110c9f8, 32'shc1111310, 32'shc1115c32, 32'shc111a55d, 32'shc111ee92, 32'shc11237d0, 
               32'shc1128119, 32'shc112ca6b, 32'shc11313c7, 32'shc1135d2c, 32'shc113a69b, 32'shc113f014, 32'shc1143997, 32'shc1148323, 
               32'shc114ccb9, 32'shc1151658, 32'shc1156002, 32'shc115a9b5, 32'shc115f372, 32'shc1163d38, 32'shc1168708, 32'shc116d0e2, 
               32'shc1171ac6, 32'shc11764b3, 32'shc117aeaa, 32'shc117f8ab, 32'shc11842b5, 32'shc1188cc9, 32'shc118d6e7, 32'shc119210e, 
               32'shc1196b3f, 32'shc119b57a, 32'shc119ffbf, 32'shc11a4a0d, 32'shc11a9465, 32'shc11adec7, 32'shc11b2932, 32'shc11b73a7, 
               32'shc11bbe26, 32'shc11c08af, 32'shc11c5341, 32'shc11c9ddd, 32'shc11ce882, 32'shc11d3331, 32'shc11d7dea, 32'shc11dc8ad, 
               32'shc11e1379, 32'shc11e5e4f, 32'shc11ea92f, 32'shc11ef419, 32'shc11f3f0c, 32'shc11f8a09, 32'shc11fd50f, 32'shc120201f, 
               32'shc1206b39, 32'shc120b65d, 32'shc121018a, 32'shc1214cc1, 32'shc1219802, 32'shc121e34c, 32'shc1222ea1, 32'shc12279fe, 
               32'shc122c566, 32'shc12310d7, 32'shc1235c52, 32'shc123a7d7, 32'shc123f365, 32'shc1243efd, 32'shc1248a9e, 32'shc124d64a, 
               32'shc12521ff, 32'shc1256dbe, 32'shc125b986, 32'shc1260558, 32'shc1265134, 32'shc1269d19, 32'shc126e909, 32'shc1273501, 
               32'shc1278104, 32'shc127cd10, 32'shc1281926, 32'shc1286546, 32'shc128b16f, 32'shc128fda2, 32'shc12949df, 32'shc1299626, 
               32'shc129e276, 32'shc12a2ecf, 32'shc12a7b33, 32'shc12ac7a0, 32'shc12b1417, 32'shc12b6098, 32'shc12bad22, 32'shc12bf9b6, 
               32'shc12c4653, 32'shc12c92fb, 32'shc12cdfac, 32'shc12d2c66, 32'shc12d792b, 32'shc12dc5f9, 32'shc12e12d1, 32'shc12e5fb2, 
               32'shc12eac9d, 32'shc12ef992, 32'shc12f4690, 32'shc12f9399, 32'shc12fe0ab, 32'shc1302dc6, 32'shc1307aeb, 32'shc130c81a, 
               32'shc1311553, 32'shc1316295, 32'shc131afe1, 32'shc131fd37, 32'shc1324a96, 32'shc13297ff, 32'shc132e572, 32'shc13332ef, 
               32'shc1338075, 32'shc133ce04, 32'shc1341b9e, 32'shc1346941, 32'shc134b6ee, 32'shc13504a4, 32'shc1355265, 32'shc135a02f, 
               32'shc135ee02, 32'shc1363bdf, 32'shc13689c6, 32'shc136d7b7, 32'shc13725b1, 32'shc13773b5, 32'shc137c1c3, 32'shc1380fda, 
               32'shc1385dfb, 32'shc138ac26, 32'shc138fa5a, 32'shc1394898, 32'shc13996e0, 32'shc139e532, 32'shc13a338d, 32'shc13a81f2, 
               32'shc13ad060, 32'shc13b1ed8, 32'shc13b6d5a, 32'shc13bbbe6, 32'shc13c0a7b, 32'shc13c591a, 32'shc13ca7c2, 32'shc13cf674, 
               32'shc13d4530, 32'shc13d93f6, 32'shc13de2c5, 32'shc13e319e, 32'shc13e8081, 32'shc13ecf6d, 32'shc13f1e63, 32'shc13f6d63, 
               32'shc13fbc6c, 32'shc1400b7f, 32'shc1405a9c, 32'shc140a9c2, 32'shc140f8f2, 32'shc141482c, 32'shc141976f, 32'shc141e6bc, 
               32'shc1423613, 32'shc1428574, 32'shc142d4de, 32'shc1432451, 32'shc14373cf, 32'shc143c356, 32'shc14412e7, 32'shc1446281, 
               32'shc144b225, 32'shc14501d3, 32'shc145518b, 32'shc145a14c, 32'shc145f117, 32'shc14640eb, 32'shc14690ca, 32'shc146e0b1, 
               32'shc14730a3, 32'shc147809e, 32'shc147d0a3, 32'shc14820b2, 32'shc14870ca, 32'shc148c0ec, 32'shc1491117, 32'shc149614c, 
               32'shc149b18b, 32'shc14a01d4, 32'shc14a5226, 32'shc14aa282, 32'shc14af2e8, 32'shc14b4357, 32'shc14b93d0, 32'shc14be453, 
               32'shc14c34df, 32'shc14c8575, 32'shc14cd614, 32'shc14d26be, 32'shc14d7771, 32'shc14dc82d, 32'shc14e18f3, 32'shc14e69c3, 
               32'shc14eba9d, 32'shc14f0b80, 32'shc14f5c6d, 32'shc14fad64, 32'shc14ffe64, 32'shc1504f6e, 32'shc150a082, 32'shc150f19f, 
               32'shc15142c6, 32'shc15193f7, 32'shc151e531, 32'shc1523675, 32'shc15287c3, 32'shc152d91a, 32'shc1532a7b, 32'shc1537be5, 
               32'shc153cd5a, 32'shc1541ed8, 32'shc154705f, 32'shc154c1f1, 32'shc155138c, 32'shc1556530, 32'shc155b6de, 32'shc1560896, 
               32'shc1565a58, 32'shc156ac23, 32'shc156fdf8, 32'shc1574fd7, 32'shc157a1bf, 32'shc157f3b1, 32'shc15845ac, 32'shc15897b2, 
               32'shc158e9c1, 32'shc1593bd9, 32'shc1598dfb, 32'shc159e027, 32'shc15a325d, 32'shc15a849c, 32'shc15ad6e5, 32'shc15b2937, 
               32'shc15b7b94, 32'shc15bcdfa, 32'shc15c2069, 32'shc15c72e2, 32'shc15cc565, 32'shc15d17f2, 32'shc15d6a88, 32'shc15dbd27, 
               32'shc15e0fd1, 32'shc15e6284, 32'shc15eb541, 32'shc15f0807, 32'shc15f5ad7, 32'shc15fadb1, 32'shc1600095, 32'shc1605382, 
               32'shc160a678, 32'shc160f979, 32'shc1614c83, 32'shc1619f97, 32'shc161f2b4, 32'shc16245db, 32'shc162990c, 32'shc162ec46, 
               32'shc1633f8a, 32'shc16392d8, 32'shc163e62f, 32'shc1643990, 32'shc1648cfa, 32'shc164e06f, 32'shc16533ed, 32'shc1658774, 
               32'shc165db05, 32'shc1662ea0, 32'shc1668245, 32'shc166d5f3, 32'shc16729ab, 32'shc1677d6c, 32'shc167d137, 32'shc168250c, 
               32'shc16878eb, 32'shc168ccd3, 32'shc16920c5, 32'shc16974c0, 32'shc169c8c5, 32'shc16a1cd4, 32'shc16a70ec, 32'shc16ac50e, 
               32'shc16b193a, 32'shc16b6d6f, 32'shc16bc1ae, 32'shc16c15f7, 32'shc16c6a49, 32'shc16cbea5, 32'shc16d130a, 32'shc16d677a, 
               32'shc16dbbf3, 32'shc16e1075, 32'shc16e6501, 32'shc16eb997, 32'shc16f0e36, 32'shc16f62e0, 32'shc16fb792, 32'shc1700c4f, 
               32'shc1706115, 32'shc170b5e5, 32'shc1710abe, 32'shc1715fa1, 32'shc171b48e, 32'shc1720984, 32'shc1725e84, 32'shc172b38d, 
               32'shc17308a1, 32'shc1735dbd, 32'shc173b2e4, 32'shc1740814, 32'shc1745d4e, 32'shc174b291, 32'shc17507df, 32'shc1755d35, 
               32'shc175b296, 32'shc1760800, 32'shc1765d73, 32'shc176b2f1, 32'shc1770878, 32'shc1775e08, 32'shc177b3a3, 32'shc1780946, 
               32'shc1785ef4, 32'shc178b4ab, 32'shc1790a6c, 32'shc1796036, 32'shc179b60b, 32'shc17a0be8, 32'shc17a61d0, 32'shc17ab7c1, 
               32'shc17b0dbb, 32'shc17b63c0, 32'shc17bb9ce, 32'shc17c0fe5, 32'shc17c6607, 32'shc17cbc32, 32'shc17d1266, 32'shc17d68a4, 
               32'shc17dbeec, 32'shc17e153d, 32'shc17e6b99, 32'shc17ec1fd, 32'shc17f186c, 32'shc17f6ee4, 32'shc17fc565, 32'shc1801bf1, 
               32'shc1807285, 32'shc180c924, 32'shc1811fcc, 32'shc181767e, 32'shc181cd3a, 32'shc18223ff, 32'shc1827acd, 32'shc182d1a6, 
               32'shc1832888, 32'shc1837f73, 32'shc183d669, 32'shc1842d68, 32'shc1848470, 32'shc184db82, 32'shc185329e, 32'shc18589c4, 
               32'shc185e0f3, 32'shc186382c, 32'shc1868f6e, 32'shc186e6ba, 32'shc1873e10, 32'shc187956f, 32'shc187ecd8, 32'shc188444a, 
               32'shc1889bc6, 32'shc188f34c, 32'shc1894adc, 32'shc189a275, 32'shc189fa17, 32'shc18a51c4, 32'shc18aa97a, 32'shc18b0139, 
               32'shc18b5903, 32'shc18bb0d5, 32'shc18c08b2, 32'shc18c6098, 32'shc18cb888, 32'shc18d1081, 32'shc18d6884, 32'shc18dc091, 
               32'shc18e18a7, 32'shc18e70c7, 32'shc18ec8f1, 32'shc18f2124, 32'shc18f7961, 32'shc18fd1a7, 32'shc19029f7, 32'shc1908251, 
               32'shc190dab4, 32'shc1913321, 32'shc1918b98, 32'shc191e418, 32'shc1923ca2, 32'shc1929535, 32'shc192edd2, 32'shc1934679, 
               32'shc1939f29, 32'shc193f7e3, 32'shc19450a7, 32'shc194a974, 32'shc195024b, 32'shc1955b2b, 32'shc195b415, 32'shc1960d09, 
               32'shc1966606, 32'shc196bf0d, 32'shc197181e, 32'shc1977138, 32'shc197ca5c, 32'shc1982389, 32'shc1987cc1, 32'shc198d601, 
               32'shc1992f4c, 32'shc199889f, 32'shc199e1fd, 32'shc19a3b64, 32'shc19a94d5, 32'shc19aee50, 32'shc19b47d4, 32'shc19ba161, 
               32'shc19bfaf9, 32'shc19c549a, 32'shc19cae44, 32'shc19d07f8, 32'shc19d61b6, 32'shc19dbb7d, 32'shc19e154e, 32'shc19e6f29, 
               32'shc19ec90d, 32'shc19f22fb, 32'shc19f7cf3, 32'shc19fd6f4, 32'shc1a030ff, 32'shc1a08b13, 32'shc1a0e531, 32'shc1a13f59, 
               32'shc1a1998a, 32'shc1a1f3c5, 32'shc1a24e09, 32'shc1a2a857, 32'shc1a302af, 32'shc1a35d10, 32'shc1a3b77b, 32'shc1a411f0, 
               32'shc1a46c6e, 32'shc1a4c6f6, 32'shc1a52187, 32'shc1a57c22, 32'shc1a5d6c7, 32'shc1a63175, 32'shc1a68c2d, 32'shc1a6e6ee, 
               32'shc1a741b9, 32'shc1a79c8e, 32'shc1a7f76c, 32'shc1a85254, 32'shc1a8ad46, 32'shc1a90841, 32'shc1a96346, 32'shc1a9be54, 
               32'shc1aa196c, 32'shc1aa748e, 32'shc1aacfb9, 32'shc1ab2aee, 32'shc1ab862c, 32'shc1abe174, 32'shc1ac3cc6, 32'shc1ac9821, 
               32'shc1acf386, 32'shc1ad4ef5, 32'shc1adaa6d, 32'shc1ae05ef, 32'shc1ae617a, 32'shc1aebd0f, 32'shc1af18ae, 32'shc1af7456, 
               32'shc1afd007, 32'shc1b02bc3, 32'shc1b08788, 32'shc1b0e356, 32'shc1b13f2f, 32'shc1b19b10, 32'shc1b1f6fc, 32'shc1b252f1, 
               32'shc1b2aef0, 32'shc1b30af8, 32'shc1b3670a, 32'shc1b3c325, 32'shc1b41f4a, 32'shc1b47b79, 32'shc1b4d7b1, 32'shc1b533f3, 
               32'shc1b5903f, 32'shc1b5ec94, 32'shc1b648f3, 32'shc1b6a55b, 32'shc1b701cd, 32'shc1b75e48, 32'shc1b7bacd, 32'shc1b8175c, 
               32'shc1b873f5, 32'shc1b8d097, 32'shc1b92d42, 32'shc1b989f7, 32'shc1b9e6b6, 32'shc1ba437e, 32'shc1baa050, 32'shc1bafd2c, 
               32'shc1bb5a11, 32'shc1bbb700, 32'shc1bc13f8, 32'shc1bc70fa, 32'shc1bcce06, 32'shc1bd2b1b, 32'shc1bd883a, 32'shc1bde562, 
               32'shc1be4294, 32'shc1be9fd0, 32'shc1befd15, 32'shc1bf5a64, 32'shc1bfb7bc, 32'shc1c0151e, 32'shc1c0728a, 32'shc1c0cfff, 
               32'shc1c12d7e, 32'shc1c18b06, 32'shc1c1e898, 32'shc1c24634, 32'shc1c2a3d9, 32'shc1c30188, 32'shc1c35f40, 32'shc1c3bd02, 
               32'shc1c41ace, 32'shc1c478a3, 32'shc1c4d682, 32'shc1c5346a, 32'shc1c5925c, 32'shc1c5f057, 32'shc1c64e5d, 32'shc1c6ac6b, 
               32'shc1c70a84, 32'shc1c768a6, 32'shc1c7c6d1, 32'shc1c82506, 32'shc1c88345, 32'shc1c8e18d, 32'shc1c93fdf, 32'shc1c99e3b, 
               32'shc1c9fca0, 32'shc1ca5b0f, 32'shc1cab987, 32'shc1cb1809, 32'shc1cb7694, 32'shc1cbd529, 32'shc1cc33c8, 32'shc1cc9270, 
               32'shc1ccf122, 32'shc1cd4fde, 32'shc1cdaea3, 32'shc1ce0d71, 32'shc1ce6c49, 32'shc1cecb2b, 32'shc1cf2a17, 32'shc1cf890c, 
               32'shc1cfe80a, 32'shc1d04712, 32'shc1d0a624, 32'shc1d1053f, 32'shc1d16464, 32'shc1d1c393, 32'shc1d222cb, 32'shc1d2820d, 
               32'shc1d2e158, 32'shc1d340ad, 32'shc1d3a00b, 32'shc1d3ff73, 32'shc1d45ee5, 32'shc1d4be60, 32'shc1d51de5, 32'shc1d57d74, 
               32'shc1d5dd0c, 32'shc1d63cad, 32'shc1d69c58, 32'shc1d6fc0d, 32'shc1d75bcb, 32'shc1d7bb93, 32'shc1d81b65, 32'shc1d87b40, 
               32'shc1d8db25, 32'shc1d93b13, 32'shc1d99b0b, 32'shc1d9fb0c, 32'shc1da5b17, 32'shc1dabb2c, 32'shc1db1b4a, 32'shc1db7b72, 
               32'shc1dbdba3, 32'shc1dc3bde, 32'shc1dc9c23, 32'shc1dcfc71, 32'shc1dd5cc8, 32'shc1ddbd2a, 32'shc1de1d94, 32'shc1de7e09, 
               32'shc1dede87, 32'shc1df3f0f, 32'shc1df9fa0, 32'shc1e0003a, 32'shc1e060df, 32'shc1e0c18d, 32'shc1e12244, 32'shc1e18305, 
               32'shc1e1e3d0, 32'shc1e244a4, 32'shc1e2a582, 32'shc1e30669, 32'shc1e3675a, 32'shc1e3c855, 32'shc1e42959, 32'shc1e48a67, 
               32'shc1e4eb7e, 32'shc1e54c9f, 32'shc1e5adc9, 32'shc1e60efd, 32'shc1e6703b, 32'shc1e6d182, 32'shc1e732d3, 32'shc1e7942d, 
               32'shc1e7f591, 32'shc1e856fe, 32'shc1e8b876, 32'shc1e919f6, 32'shc1e97b80, 32'shc1e9dd14, 32'shc1ea3eb1, 32'shc1eaa058, 
               32'shc1eb0209, 32'shc1eb63c3, 32'shc1ebc587, 32'shc1ec2754, 32'shc1ec892b, 32'shc1eceb0b, 32'shc1ed4cf5, 32'shc1edaee8, 
               32'shc1ee10e5, 32'shc1ee72ec, 32'shc1eed4fc, 32'shc1ef3716, 32'shc1ef9939, 32'shc1effb66, 32'shc1f05d9d, 32'shc1f0bfdd, 
               32'shc1f12227, 32'shc1f1847a, 32'shc1f1e6d7, 32'shc1f2493d, 32'shc1f2abad, 32'shc1f30e26, 32'shc1f370a9, 32'shc1f3d336, 
               32'shc1f435cc, 32'shc1f4986c, 32'shc1f4fb15, 32'shc1f55dc8, 32'shc1f5c085, 32'shc1f6234b, 32'shc1f6861a, 32'shc1f6e8f4, 
               32'shc1f74bd6, 32'shc1f7aec3, 32'shc1f811b9, 32'shc1f874b8, 32'shc1f8d7c1, 32'shc1f93ad4, 32'shc1f99df0, 32'shc1fa0115, 
               32'shc1fa6445, 32'shc1fac77e, 32'shc1fb2ac0, 32'shc1fb8e0c, 32'shc1fbf161, 32'shc1fc54c0, 32'shc1fcb829, 32'shc1fd1b9b, 
               32'shc1fd7f17, 32'shc1fde29c, 32'shc1fe462b, 32'shc1fea9c4, 32'shc1ff0d66, 32'shc1ff7111, 32'shc1ffd4c7, 32'shc2003885, 
               32'shc2009c4e, 32'shc201001f, 32'shc20163fb, 32'shc201c7e0, 32'shc2022bce, 32'shc2028fc6, 32'shc202f3c8, 32'shc20357d3, 
               32'shc203bbe8, 32'shc2042006, 32'shc204842e, 32'shc204e860, 32'shc2054c9b, 32'shc205b0df, 32'shc206152d, 32'shc2067985, 
               32'shc206dde6, 32'shc2074251, 32'shc207a6c5, 32'shc2080b43, 32'shc2086fca, 32'shc208d45b, 32'shc20938f6, 32'shc2099d9a, 
               32'shc20a0248, 32'shc20a66ff, 32'shc20acbc0, 32'shc20b308a, 32'shc20b955e, 32'shc20bfa3b, 32'shc20c5f22, 32'shc20cc413, 
               32'shc20d290d, 32'shc20d8e11, 32'shc20df31e, 32'shc20e5835, 32'shc20ebd55, 32'shc20f227f, 32'shc20f87b2, 32'shc20fecef, 
               32'shc2105236, 32'shc210b786, 32'shc2111cdf, 32'shc2118243, 32'shc211e7af, 32'shc2124d26, 32'shc212b2a5, 32'shc213182f, 
               32'shc2137dc2, 32'shc213e35e, 32'shc2144904, 32'shc214aeb4, 32'shc215146d, 32'shc2157a30, 32'shc215dffc, 32'shc21645d2, 
               32'shc216abb1, 32'shc217119a, 32'shc217778c, 32'shc217dd88, 32'shc218438e, 32'shc218a99d, 32'shc2190fb5, 32'shc21975d7, 
               32'shc219dc03, 32'shc21a4238, 32'shc21aa877, 32'shc21b0ebf, 32'shc21b7511, 32'shc21bdb6d, 32'shc21c41d2, 32'shc21ca840, 
               32'shc21d0eb8, 32'shc21d753a, 32'shc21ddbc5, 32'shc21e425a, 32'shc21ea8f8, 32'shc21f0fa0, 32'shc21f7651, 32'shc21fdd0c, 
               32'shc22043d0, 32'shc220aa9e, 32'shc2211176, 32'shc2217857, 32'shc221df41, 32'shc2224635, 32'shc222ad33, 32'shc223143a, 
               32'shc2237b4b, 32'shc223e265, 32'shc2244989, 32'shc224b0b6, 32'shc22517ed, 32'shc2257f2d, 32'shc225e677, 32'shc2264dcb, 
               32'shc226b528, 32'shc2271c8e, 32'shc22783fe, 32'shc227eb78, 32'shc22852fb, 32'shc228ba88, 32'shc229221e, 32'shc22989be, 
               32'shc229f167, 32'shc22a591a, 32'shc22ac0d7, 32'shc22b289d, 32'shc22b906c, 32'shc22bf845, 32'shc22c6028, 32'shc22cc814, 
               32'shc22d3009, 32'shc22d9808, 32'shc22e0011, 32'shc22e6823, 32'shc22ed03f, 32'shc22f3864, 32'shc22fa093, 32'shc23008cb, 
               32'shc230710d, 32'shc230d959, 32'shc23141ae, 32'shc231aa0c, 32'shc2321274, 32'shc2327ae6, 32'shc232e361, 32'shc2334be5, 
               32'shc233b473, 32'shc2341d0b, 32'shc23485ac, 32'shc234ee57, 32'shc235570b, 32'shc235bfc9, 32'shc2362890, 32'shc2369161, 
               32'shc236fa3b, 32'shc237631f, 32'shc237cc0d, 32'shc2383504, 32'shc2389e04, 32'shc239070e, 32'shc2397021, 32'shc239d93f, 
               32'shc23a4265, 32'shc23aab95, 32'shc23b14cf, 32'shc23b7e12, 32'shc23be75f, 32'shc23c50b5, 32'shc23cba15, 32'shc23d237e, 
               32'shc23d8cf1, 32'shc23df66d, 32'shc23e5ff3, 32'shc23ec982, 32'shc23f331b, 32'shc23f9cbd, 32'shc2400669, 32'shc240701f, 
               32'shc240d9de, 32'shc24143a6, 32'shc241ad78, 32'shc2421754, 32'shc2428139, 32'shc242eb27, 32'shc243551f, 32'shc243bf21, 
               32'shc244292c, 32'shc2449341, 32'shc244fd5f, 32'shc2456786, 32'shc245d1b8, 32'shc2463bf2, 32'shc246a637, 32'shc2471084, 
               32'shc2477adc, 32'shc247e53c, 32'shc2484fa7, 32'shc248ba1b, 32'shc2492498, 32'shc2498f1f, 32'shc249f9af, 32'shc24a6449, 
               32'shc24aceed, 32'shc24b3999, 32'shc24ba450, 32'shc24c0f10, 32'shc24c79d9, 32'shc24ce4ac, 32'shc24d4f89, 32'shc24dba6f, 
               32'shc24e255e, 32'shc24e9057, 32'shc24efb5a, 32'shc24f6666, 32'shc24fd17c, 32'shc2503c9b, 32'shc250a7c3, 32'shc25112f6, 
               32'shc2517e31, 32'shc251e976, 32'shc25254c5, 32'shc252c01d, 32'shc2532b7f, 32'shc25396ea, 32'shc254025f, 32'shc2546ddd, 
               32'shc254d965, 32'shc25544f6, 32'shc255b091, 32'shc2561c35, 32'shc25687e3, 32'shc256f39a, 32'shc2575f5b, 32'shc257cb25, 
               32'shc25836f9, 32'shc258a2d6, 32'shc2590ebd, 32'shc2597aad, 32'shc259e6a7, 32'shc25a52ab, 32'shc25abeb7, 32'shc25b2ace, 
               32'shc25b96ee, 32'shc25c0317, 32'shc25c6f4a, 32'shc25cdb86, 32'shc25d47cc, 32'shc25db41c, 32'shc25e2074, 32'shc25e8cd7, 
               32'shc25ef943, 32'shc25f65b8, 32'shc25fd237, 32'shc2603ec0, 32'shc260ab51, 32'shc26117ed, 32'shc2618492, 32'shc261f140, 
               32'shc2625df8, 32'shc262caba, 32'shc2633785, 32'shc263a459, 32'shc2641137, 32'shc2647e1e, 32'shc264eb0f, 32'shc265580a, 
               32'shc265c50e, 32'shc266321b, 32'shc2669f32, 32'shc2670c52, 32'shc267797c, 32'shc267e6b0, 32'shc26853ed, 32'shc268c133, 
               32'shc2692e83, 32'shc2699bdd, 32'shc26a093f, 32'shc26a76ac, 32'shc26ae422, 32'shc26b51a1, 32'shc26bbf2a, 32'shc26c2cbd, 
               32'shc26c9a58, 32'shc26d07fe, 32'shc26d75ad, 32'shc26de365, 32'shc26e5127, 32'shc26ebef2, 32'shc26f2cc7, 32'shc26f9aa6, 
               32'shc270088e, 32'shc270767f, 32'shc270e47a, 32'shc271527e, 32'shc271c08c, 32'shc2722ea3, 32'shc2729cc4, 32'shc2730aee, 
               32'shc2737922, 32'shc273e760, 32'shc27455a6, 32'shc274c3f7, 32'shc2753250, 32'shc275a0b4, 32'shc2760f20, 32'shc2767d97, 
               32'shc276ec16, 32'shc2775aa0, 32'shc277c932, 32'shc27837ce, 32'shc278a674, 32'shc2791523, 32'shc27983dc, 32'shc279f29e, 
               32'shc27a616a, 32'shc27ad03f, 32'shc27b3f1e, 32'shc27bae06, 32'shc27c1cf7, 32'shc27c8bf2, 32'shc27cfaf7, 32'shc27d6a05, 
               32'shc27dd91c, 32'shc27e483d, 32'shc27eb768, 32'shc27f269c, 32'shc27f95d9, 32'shc2800520, 32'shc2807471, 32'shc280e3cb, 
               32'shc281532e, 32'shc281c29b, 32'shc2823211, 32'shc282a191, 32'shc283111b, 32'shc28380ad, 32'shc283f04a, 32'shc2845ff0, 
               32'shc284cf9f, 32'shc2853f58, 32'shc285af1a, 32'shc2861ee6, 32'shc2868ebb, 32'shc286fe99, 32'shc2876e82, 32'shc287de73, 
               32'shc2884e6e, 32'shc288be73, 32'shc2892e81, 32'shc2899e98, 32'shc28a0eb9, 32'shc28a7ee4, 32'shc28aef18, 32'shc28b5f55, 
               32'shc28bcf9c, 32'shc28c3fed, 32'shc28cb047, 32'shc28d20aa, 32'shc28d9117, 32'shc28e018d, 32'shc28e720d, 32'shc28ee296, 
               32'shc28f5329, 32'shc28fc3c5, 32'shc290346b, 32'shc290a51a, 32'shc29115d3, 32'shc2918695, 32'shc291f760, 32'shc2926835, 
               32'shc292d914, 32'shc29349fc, 32'shc293baed, 32'shc2942be8, 32'shc2949ced, 32'shc2950dfb, 32'shc2957f12, 32'shc295f033, 
               32'shc296615d, 32'shc296d291, 32'shc29743ce, 32'shc297b515, 32'shc2982665, 32'shc29897bf, 32'shc2990922, 32'shc2997a8f, 
               32'shc299ec05, 32'shc29a5d84, 32'shc29acf0d, 32'shc29b40a0, 32'shc29bb23c, 32'shc29c23e1, 32'shc29c9590, 32'shc29d0748, 
               32'shc29d790a, 32'shc29dead5, 32'shc29e5caa, 32'shc29ece88, 32'shc29f4070, 32'shc29fb261, 32'shc2a0245c, 32'shc2a09660, 
               32'shc2a1086d, 32'shc2a17a84, 32'shc2a1eca5, 32'shc2a25ecf, 32'shc2a2d102, 32'shc2a3433f, 32'shc2a3b585, 32'shc2a427d5, 
               32'shc2a49a2e, 32'shc2a50c91, 32'shc2a57efd, 32'shc2a5f173, 32'shc2a663f2, 32'shc2a6d67a, 32'shc2a7490c, 32'shc2a7bba8, 
               32'shc2a82e4d, 32'shc2a8a0fb, 32'shc2a913b3, 32'shc2a98674, 32'shc2a9f93f, 32'shc2aa6c13, 32'shc2aadef1, 32'shc2ab51d8, 
               32'shc2abc4c9, 32'shc2ac37c3, 32'shc2acaac6, 32'shc2ad1dd3, 32'shc2ad90ea, 32'shc2ae0409, 32'shc2ae7733, 32'shc2aeea66, 
               32'shc2af5da2, 32'shc2afd0e8, 32'shc2b04437, 32'shc2b0b78f, 32'shc2b12af1, 32'shc2b19e5d, 32'shc2b211d2, 32'shc2b28550, 
               32'shc2b2f8d8, 32'shc2b36c6a, 32'shc2b3e004, 32'shc2b453a9, 32'shc2b4c756, 32'shc2b53b0d, 32'shc2b5aece, 32'shc2b62298, 
               32'shc2b6966c, 32'shc2b70a49, 32'shc2b77e2f, 32'shc2b7f21f, 32'shc2b86618, 32'shc2b8da1b, 32'shc2b94e27, 32'shc2b9c23d, 
               32'shc2ba365c, 32'shc2baaa84, 32'shc2bb1eb6, 32'shc2bb92f2, 32'shc2bc0737, 32'shc2bc7b85, 32'shc2bcefdd, 32'shc2bd643e, 
               32'shc2bdd8a9, 32'shc2be4d1d, 32'shc2bec19b, 32'shc2bf3622, 32'shc2bfaab2, 32'shc2c01f4c, 32'shc2c093ef, 32'shc2c1089c, 
               32'shc2c17d52, 32'shc2c1f212, 32'shc2c266db, 32'shc2c2dbae, 32'shc2c3508a, 32'shc2c3c56f, 32'shc2c43a5e, 32'shc2c4af57, 
               32'shc2c52459, 32'shc2c59964, 32'shc2c60e78, 32'shc2c68397, 32'shc2c6f8be, 32'shc2c76def, 32'shc2c7e32a, 32'shc2c8586e, 
               32'shc2c8cdbb, 32'shc2c94312, 32'shc2c9b872, 32'shc2ca2ddc, 32'shc2caa34f, 32'shc2cb18cb, 32'shc2cb8e51, 32'shc2cc03e1, 
               32'shc2cc7979, 32'shc2ccef1c, 32'shc2cd64c7, 32'shc2cdda7d, 32'shc2ce503b, 32'shc2cec603, 32'shc2cf3bd5, 32'shc2cfb1b0, 
               32'shc2d02794, 32'shc2d09d82, 32'shc2d11379, 32'shc2d1897a, 32'shc2d1ff84, 32'shc2d27597, 32'shc2d2ebb4, 32'shc2d361db, 
               32'shc2d3d80a, 32'shc2d44e44, 32'shc2d4c486, 32'shc2d53ad3, 32'shc2d5b128, 32'shc2d62787, 32'shc2d69df0, 32'shc2d71461, 
               32'shc2d78add, 32'shc2d80161, 32'shc2d877f0, 32'shc2d8ee87, 32'shc2d96528, 32'shc2d9dbd3, 32'shc2da5286, 32'shc2dac944, 
               32'shc2db400a, 32'shc2dbb6db, 32'shc2dc2db4, 32'shc2dca497, 32'shc2dd1b84, 32'shc2dd927a, 32'shc2de0979, 32'shc2de8082, 
               32'shc2def794, 32'shc2df6eaf, 32'shc2dfe5d4, 32'shc2e05d03, 32'shc2e0d43b, 32'shc2e14b7c, 32'shc2e1c2c7, 32'shc2e23a1b, 
               32'shc2e2b178, 32'shc2e328df, 32'shc2e3a050, 32'shc2e417ca, 32'shc2e48f4d, 32'shc2e506da, 32'shc2e57e70, 32'shc2e5f60f, 
               32'shc2e66db8, 32'shc2e6e56b, 32'shc2e75d26, 32'shc2e7d4ec, 32'shc2e84cba, 32'shc2e8c492, 32'shc2e93c74, 32'shc2e9b45f, 
               32'shc2ea2c53, 32'shc2eaa451, 32'shc2eb1c58, 32'shc2eb9468, 32'shc2ec0c82, 32'shc2ec84a6, 32'shc2ecfcd3, 32'shc2ed7509, 
               32'shc2eded49, 32'shc2ee6592, 32'shc2eedde4, 32'shc2ef5640, 32'shc2efcea6, 32'shc2f04714, 32'shc2f0bf8c, 32'shc2f1380e, 
               32'shc2f1b099, 32'shc2f2292e, 32'shc2f2a1cb, 32'shc2f31a73, 32'shc2f39323, 32'shc2f40bdd, 32'shc2f484a1, 32'shc2f4fd6e, 
               32'shc2f57644, 32'shc2f5ef24, 32'shc2f6680d, 32'shc2f6e100, 32'shc2f759fc, 32'shc2f7d301, 32'shc2f84c10, 32'shc2f8c528, 
               32'shc2f93e4a, 32'shc2f9b775, 32'shc2fa30a9, 32'shc2faa9e7, 32'shc2fb232e, 32'shc2fb9c7f, 32'shc2fc15d9, 32'shc2fc8f3c, 
               32'shc2fd08a9, 32'shc2fd8220, 32'shc2fdfb9f, 32'shc2fe7529, 32'shc2feeebb, 32'shc2ff6857, 32'shc2ffe1fc, 32'shc3005bab, 
               32'shc300d563, 32'shc3014f25, 32'shc301c8f0, 32'shc30242c4, 32'shc302bca2, 32'shc3033689, 32'shc303b07a, 32'shc3042a74, 
               32'shc304a477, 32'shc3051e84, 32'shc305989a, 32'shc30612ba, 32'shc3068ce3, 32'shc3070715, 32'shc3078151, 32'shc307fb97, 
               32'shc30875e5, 32'shc308f03d, 32'shc3096a9f, 32'shc309e509, 32'shc30a5f7e, 32'shc30ad9fb, 32'shc30b5482, 32'shc30bcf13, 
               32'shc30c49ad, 32'shc30cc450, 32'shc30d3efd, 32'shc30db9b3, 32'shc30e3472, 32'shc30eaf3b, 32'shc30f2a0d, 32'shc30fa4e9, 
               32'shc3101fce, 32'shc3109abc, 32'shc31115b4, 32'shc31190b5, 32'shc3120bc0, 32'shc31286d4, 32'shc31301f1, 32'shc3137d18, 
               32'shc313f848, 32'shc3147382, 32'shc314eec5, 32'shc3156a11, 32'shc315e567, 32'shc31660c6, 32'shc316dc2f, 32'shc31757a1, 
               32'shc317d31c, 32'shc3184ea1, 32'shc318ca2f, 32'shc31945c7, 32'shc319c168, 32'shc31a3d12, 32'shc31ab8c6, 32'shc31b3483, 
               32'shc31bb049, 32'shc31c2c19, 32'shc31ca7f2, 32'shc31d23d5, 32'shc31d9fc1, 32'shc31e1bb6, 32'shc31e97b5, 32'shc31f13bd, 
               32'shc31f8fcf, 32'shc3200bea, 32'shc320880e, 32'shc321043c, 32'shc3218073, 32'shc321fcb4, 32'shc32278fe, 32'shc322f551, 
               32'shc32371ae, 32'shc323ee14, 32'shc3246a83, 32'shc324e6fc, 32'shc325637f, 32'shc325e00a, 32'shc3265c9f, 32'shc326d93e, 
               32'shc32755e5, 32'shc327d296, 32'shc3284f51, 32'shc328cc15, 32'shc32948e2, 32'shc329c5b9, 32'shc32a4299, 32'shc32abf82, 
               32'shc32b3c75, 32'shc32bb971, 32'shc32c3677, 32'shc32cb386, 32'shc32d309e, 32'shc32dadc0, 32'shc32e2aeb, 32'shc32ea820, 
               32'shc32f255e, 32'shc32fa2a5, 32'shc3301ff5, 32'shc3309d50, 32'shc3311ab3, 32'shc3319820, 32'shc3321596, 32'shc3329315, 
               32'shc333109e, 32'shc3338e30, 32'shc3340bcc, 32'shc3348971, 32'shc3350720, 32'shc33584d7, 32'shc3360298, 32'shc3368063, 
               32'shc336fe37, 32'shc3377c14, 32'shc337f9fb, 32'shc33877eb, 32'shc338f5e4, 32'shc33973e7, 32'shc339f1f3, 32'shc33a7009, 
               32'shc33aee27, 32'shc33b6c50, 32'shc33bea81, 32'shc33c68bc, 32'shc33ce701, 32'shc33d654e, 32'shc33de3a5, 32'shc33e6206, 
               32'shc33ee070, 32'shc33f5ee3, 32'shc33fdd60, 32'shc3405be6, 32'shc340da75, 32'shc341590e, 32'shc341d7b0, 32'shc342565b, 
               32'shc342d510, 32'shc34353ce, 32'shc343d295, 32'shc3445166, 32'shc344d041, 32'shc3454f24, 32'shc345ce11, 32'shc3464d07, 
               32'shc346cc07, 32'shc3474b10, 32'shc347ca23, 32'shc348493f, 32'shc348c864, 32'shc3494792, 32'shc349c6ca, 32'shc34a460b, 
               32'shc34ac556, 32'shc34b44aa, 32'shc34bc407, 32'shc34c436e, 32'shc34cc2de, 32'shc34d4257, 32'shc34dc1da, 32'shc34e4166, 
               32'shc34ec0fc, 32'shc34f409b, 32'shc34fc043, 32'shc3503ff5, 32'shc350bfaf, 32'shc3513f74, 32'shc351bf41, 32'shc3523f18, 
               32'shc352bef9, 32'shc3533ee3, 32'shc353bed6, 32'shc3543ed2, 32'shc354bed8, 32'shc3553ee7, 32'shc355bf00, 32'shc3563f21, 
               32'shc356bf4d, 32'shc3573f81, 32'shc357bfbf, 32'shc3584006, 32'shc358c057, 32'shc35940b1, 32'shc359c114, 32'shc35a4181, 
               32'shc35ac1f7, 32'shc35b4277, 32'shc35bc2ff, 32'shc35c4391, 32'shc35cc42d, 32'shc35d44d2, 32'shc35dc580, 32'shc35e4637, 
               32'shc35ec6f8, 32'shc35f47c2, 32'shc35fc896, 32'shc3604973, 32'shc360ca59, 32'shc3614b49, 32'shc361cc42, 32'shc3624d44, 
               32'shc362ce50, 32'shc3634f65, 32'shc363d083, 32'shc36451ab, 32'shc364d2dc, 32'shc3655416, 32'shc365d55a, 32'shc36656a7, 
               32'shc366d7fd, 32'shc367595d, 32'shc367dac6, 32'shc3685c39, 32'shc368ddb4, 32'shc3695f3a, 32'shc369e0c8, 32'shc36a6260, 
               32'shc36ae401, 32'shc36b65ab, 32'shc36be75f, 32'shc36c691d, 32'shc36ceae3, 32'shc36d6cb3, 32'shc36dee8c, 32'shc36e706f, 
               32'shc36ef25b, 32'shc36f7450, 32'shc36ff64e, 32'shc3707856, 32'shc370fa68, 32'shc3717c82, 32'shc371fea6, 32'shc37280d3, 
               32'shc373030a, 32'shc373854a, 32'shc3740793, 32'shc37489e6, 32'shc3750c42, 32'shc3758ea7, 32'shc3761116, 32'shc376938e, 
               32'shc377160f, 32'shc377989a, 32'shc3781b2e, 32'shc3789dcb, 32'shc3792072, 32'shc379a322, 32'shc37a25db, 32'shc37aa89e, 
               32'shc37b2b6a, 32'shc37bae3f, 32'shc37c311e, 32'shc37cb406, 32'shc37d36f7, 32'shc37db9f2, 32'shc37e3cf6, 32'shc37ec003, 
               32'shc37f4319, 32'shc37fc639, 32'shc3804963, 32'shc380cc95, 32'shc3814fd1, 32'shc381d317, 32'shc3825665, 32'shc382d9bd, 
               32'shc3835d1e, 32'shc383e089, 32'shc38463fd, 32'shc384e77a, 32'shc3856b01, 32'shc385ee91, 32'shc386722a, 32'shc386f5cc, 
               32'shc3877978, 32'shc387fd2e, 32'shc38880ec, 32'shc38904b4, 32'shc3898885, 32'shc38a0c60, 32'shc38a9043, 32'shc38b1431, 
               32'shc38b9827, 32'shc38c1c27, 32'shc38ca030, 32'shc38d2442, 32'shc38da85e, 32'shc38e2c83, 32'shc38eb0b2, 32'shc38f34e9, 
               32'shc38fb92a, 32'shc3903d75, 32'shc390c1c9, 32'shc3914626, 32'shc391ca8c, 32'shc3924efc, 32'shc392d375, 32'shc39357f7, 
               32'shc393dc82, 32'shc3946117, 32'shc394e5b6, 32'shc3956a5d, 32'shc395ef0e, 32'shc39673c8, 32'shc396f88c, 32'shc3977d59, 
               32'shc398022f, 32'shc398870e, 32'shc3990bf7, 32'shc39990e9, 32'shc39a15e4, 32'shc39a9ae9, 32'shc39b1ff7, 32'shc39ba50e, 
               32'shc39c2a2f, 32'shc39caf59, 32'shc39d348c, 32'shc39db9c9, 32'shc39e3f0f, 32'shc39ec45e, 32'shc39f49b7, 32'shc39fcf18, 
               32'shc3a05484, 32'shc3a0d9f8, 32'shc3a15f76, 32'shc3a1e4fd, 32'shc3a26a8d, 32'shc3a2f027, 32'shc3a375ca, 32'shc3a3fb76, 
               32'shc3a4812c, 32'shc3a506eb, 32'shc3a58cb3, 32'shc3a61285, 32'shc3a6985f, 32'shc3a71e44, 32'shc3a7a431, 32'shc3a82a28, 
               32'shc3a8b028, 32'shc3a93631, 32'shc3a9bc44, 32'shc3aa4260, 32'shc3aac885, 32'shc3ab4eb4, 32'shc3abd4ec, 32'shc3ac5b2d, 
               32'shc3ace178, 32'shc3ad67cb, 32'shc3adee28, 32'shc3ae748f, 32'shc3aefaff, 32'shc3af8178, 32'shc3b007fa, 32'shc3b08e86, 
               32'shc3b1151b, 32'shc3b19bb9, 32'shc3b22260, 32'shc3b2a911, 32'shc3b32fcb, 32'shc3b3b68f, 32'shc3b43d5b, 32'shc3b4c431, 
               32'shc3b54b11, 32'shc3b5d1f9, 32'shc3b658eb, 32'shc3b6dfe6, 32'shc3b766eb, 32'shc3b7edf9, 32'shc3b87510, 32'shc3b8fc30, 
               32'shc3b9835a, 32'shc3ba0a8d, 32'shc3ba91c9, 32'shc3bb190f, 32'shc3bba05e, 32'shc3bc27b6, 32'shc3bcaf17, 32'shc3bd3682, 
               32'shc3bdbdf6, 32'shc3be4573, 32'shc3beccfa, 32'shc3bf548a, 32'shc3bfdc23, 32'shc3c063c6, 32'shc3c0eb71, 32'shc3c17327, 
               32'shc3c1fae5, 32'shc3c282ad, 32'shc3c30a7e, 32'shc3c39258, 32'shc3c41a3b, 32'shc3c4a228, 32'shc3c52a1e, 32'shc3c5b21e, 
               32'shc3c63a26, 32'shc3c6c238, 32'shc3c74a54, 32'shc3c7d278, 32'shc3c85aa6, 32'shc3c8e2dd, 32'shc3c96b1e, 32'shc3c9f367, 
               32'shc3ca7bba, 32'shc3cb0416, 32'shc3cb8c7c, 32'shc3cc14eb, 32'shc3cc9d63, 32'shc3cd25e4, 32'shc3cdae6f, 32'shc3ce3703, 
               32'shc3cebfa0, 32'shc3cf4847, 32'shc3cfd0f7, 32'shc3d059b0, 32'shc3d0e272, 32'shc3d16b3e, 32'shc3d1f413, 32'shc3d27cf1, 
               32'shc3d305d8, 32'shc3d38ec9, 32'shc3d417c3, 32'shc3d4a0c7, 32'shc3d529d3, 32'shc3d5b2e9, 32'shc3d63c08, 32'shc3d6c531, 
               32'shc3d74e62, 32'shc3d7d79d, 32'shc3d860e2, 32'shc3d8ea2f, 32'shc3d97386, 32'shc3d9fce6, 32'shc3da8650, 32'shc3db0fc2, 
               32'shc3db993e, 32'shc3dc22c4, 32'shc3dcac52, 32'shc3dd35ea, 32'shc3ddbf8b, 32'shc3de4935, 32'shc3ded2e9, 32'shc3df5ca6, 
               32'shc3dfe66c, 32'shc3e0703b, 32'shc3e0fa14, 32'shc3e183f6, 32'shc3e20de1, 32'shc3e297d5, 32'shc3e321d3, 32'shc3e3abda, 
               32'shc3e435ea, 32'shc3e4c004, 32'shc3e54a27, 32'shc3e5d453, 32'shc3e65e88, 32'shc3e6e8c7, 32'shc3e7730f, 32'shc3e7fd60, 
               32'shc3e887bb, 32'shc3e9121e, 32'shc3e99c8b, 32'shc3ea2701, 32'shc3eab181, 32'shc3eb3c0a, 32'shc3ebc69c, 32'shc3ec5137, 
               32'shc3ecdbdc, 32'shc3ed6689, 32'shc3edf141, 32'shc3ee7c01, 32'shc3ef06cb, 32'shc3ef919d, 32'shc3f01c7a, 32'shc3f0a75f, 
               32'shc3f1324e, 32'shc3f1bd46, 32'shc3f24847, 32'shc3f2d351, 32'shc3f35e65, 32'shc3f3e982, 32'shc3f474a8, 32'shc3f4ffd8, 
               32'shc3f58b10, 32'shc3f61652, 32'shc3f6a19e, 32'shc3f72cf2, 32'shc3f7b850, 32'shc3f843b7, 32'shc3f8cf27, 32'shc3f95aa1, 
               32'shc3f9e624, 32'shc3fa71b0, 32'shc3fafd45, 32'shc3fb88e4, 32'shc3fc148c, 32'shc3fca03d, 32'shc3fd2bf7, 32'shc3fdb7bb, 
               32'shc3fe4388, 32'shc3fecf5e, 32'shc3ff5b3d, 32'shc3ffe726, 32'shc4007318, 32'shc400ff13, 32'shc4018b17, 32'shc4021725, 
               32'shc402a33c, 32'shc4032f5c, 32'shc403bb85, 32'shc40447b8, 32'shc404d3f4, 32'shc4056039, 32'shc405ec87, 32'shc40678df, 
               32'shc4070540, 32'shc40791aa, 32'shc4081e1d, 32'shc408aa9a, 32'shc4093720, 32'shc409c3af, 32'shc40a5047, 32'shc40adce9, 
               32'shc40b6994, 32'shc40bf648, 32'shc40c8305, 32'shc40d0fcc, 32'shc40d9c9c, 32'shc40e2975, 32'shc40eb657, 32'shc40f4343, 
               32'shc40fd037, 32'shc4105d36, 32'shc410ea3d, 32'shc411774d, 32'shc4120467, 32'shc412918a, 32'shc4131eb7, 32'shc413abec, 
               32'shc414392b, 32'shc414c673, 32'shc41553c4, 32'shc415e11f, 32'shc4166e82, 32'shc416fbef, 32'shc4178965, 32'shc41816e5, 
               32'shc418a46d, 32'shc41931ff, 32'shc419bf9b, 32'shc41a4d3f, 32'shc41adaed, 32'shc41b68a3, 32'shc41bf664, 32'shc41c842d, 
               32'shc41d11ff, 32'shc41d9fdb, 32'shc41e2dc0, 32'shc41ebbaf, 32'shc41f49a6, 32'shc41fd7a7, 32'shc42065b1, 32'shc420f3c4, 
               32'shc42181e0, 32'shc4221006, 32'shc4229e35, 32'shc4232c6d, 32'shc423baae, 32'shc42448f9, 32'shc424d74d, 32'shc42565aa, 
               32'shc425f410, 32'shc4268280, 32'shc42710f9, 32'shc4279f7b, 32'shc4282e06, 32'shc428bc9a, 32'shc4294b38, 32'shc429d9df, 
               32'shc42a688f, 32'shc42af748, 32'shc42b860b, 32'shc42c14d7, 32'shc42ca3ac, 32'shc42d328a, 32'shc42dc171, 32'shc42e5062, 
               32'shc42edf5c, 32'shc42f6e5f, 32'shc42ffd6b, 32'shc4308c81, 32'shc4311ba0, 32'shc431aac8, 32'shc43239f9, 32'shc432c934, 
               32'shc4335877, 32'shc433e7c4, 32'shc434771b, 32'shc435067a, 32'shc43595e3, 32'shc4362554, 32'shc436b4cf, 32'shc4374454, 
               32'shc437d3e1, 32'shc4386378, 32'shc438f318, 32'shc43982c1, 32'shc43a1273, 32'shc43aa22f, 32'shc43b31f4, 32'shc43bc1c2, 
               32'shc43c5199, 32'shc43ce179, 32'shc43d7163, 32'shc43e0156, 32'shc43e9152, 32'shc43f2157, 32'shc43fb166, 32'shc440417d, 
               32'shc440d19e, 32'shc44161c9, 32'shc441f1fc, 32'shc4428239, 32'shc443127e, 32'shc443a2cd, 32'shc4443326, 32'shc444c387, 
               32'shc44553f2, 32'shc445e466, 32'shc44674e3, 32'shc4470569, 32'shc44795f8, 32'shc4482691, 32'shc448b733, 32'shc44947de, 
               32'shc449d892, 32'shc44a6950, 32'shc44afa17, 32'shc44b8ae7, 32'shc44c1bc0, 32'shc44caca2, 32'shc44d3d8e, 32'shc44dce82, 
               32'shc44e5f80, 32'shc44ef088, 32'shc44f8198, 32'shc45012b2, 32'shc450a3d4, 32'shc4513500, 32'shc451c636, 32'shc4525774, 
               32'shc452e8bc, 32'shc4537a0d, 32'shc4540b67, 32'shc4549cca, 32'shc4552e36, 32'shc455bfac, 32'shc456512b, 32'shc456e2b3, 
               32'shc4577444, 32'shc45805de, 32'shc4589782, 32'shc459292f, 32'shc459bae5, 32'shc45a4ca4, 32'shc45ade6c, 32'shc45b703e, 
               32'shc45c0219, 32'shc45c93fd, 32'shc45d25ea, 32'shc45db7e1, 32'shc45e49e0, 32'shc45edbe9, 32'shc45f6dfb, 32'shc4600016, 
               32'shc460923b, 32'shc4612468, 32'shc461b69f, 32'shc46248df, 32'shc462db28, 32'shc4636d7a, 32'shc463ffd6, 32'shc464923b, 
               32'shc46524a9, 32'shc465b720, 32'shc46649a0, 32'shc466dc2a, 32'shc4676ebc, 32'shc4680158, 32'shc46893fd, 32'shc46926ac, 
               32'shc469b963, 32'shc46a4c24, 32'shc46adeee, 32'shc46b71c1, 32'shc46c049d, 32'shc46c9782, 32'shc46d2a71, 32'shc46dbd69, 
               32'shc46e5069, 32'shc46ee374, 32'shc46f7687, 32'shc47009a4, 32'shc4709cc9, 32'shc4712ff8, 32'shc471c330, 32'shc4725671, 
               32'shc472e9bc, 32'shc4737d10, 32'shc474106c, 32'shc474a3d2, 32'shc4753741, 32'shc475caba, 32'shc4765e3b, 32'shc476f1c6, 
               32'shc477855a, 32'shc47818f7, 32'shc478ac9d, 32'shc479404d, 32'shc479d405, 32'shc47a67c7, 32'shc47afb92, 32'shc47b8f66, 
               32'shc47c2344, 32'shc47cb72a, 32'shc47d4b1a, 32'shc47ddf13, 32'shc47e7315, 32'shc47f0720, 32'shc47f9b34, 32'shc4802f52, 
               32'shc480c379, 32'shc48157a9, 32'shc481ebe2, 32'shc4828024, 32'shc4831470, 32'shc483a8c4, 32'shc4843d22, 32'shc484d189, 
               32'shc48565f9, 32'shc485fa72, 32'shc4868ef5, 32'shc4872381, 32'shc487b815, 32'shc4884cb3, 32'shc488e15b, 32'shc489760b, 
               32'shc48a0ac4, 32'shc48a9f87, 32'shc48b3453, 32'shc48bc928, 32'shc48c5e06, 32'shc48cf2ee, 32'shc48d87de, 32'shc48e1cd8, 
               32'shc48eb1db, 32'shc48f46e7, 32'shc48fdbfc, 32'shc490711a, 32'shc4910642, 32'shc4919b72, 32'shc49230ac, 32'shc492c5ef, 
               32'shc4935b3c, 32'shc493f091, 32'shc49485ef, 32'shc4951b57, 32'shc495b0c8, 32'shc4964642, 32'shc496dbc5, 32'shc4977151, 
               32'shc49806e7, 32'shc4989c86, 32'shc499322d, 32'shc499c7de, 32'shc49a5d98, 32'shc49af35c, 32'shc49b8928, 32'shc49c1efe, 
               32'shc49cb4dd, 32'shc49d4ac5, 32'shc49de0b6, 32'shc49e76b0, 32'shc49f0cb3, 32'shc49fa2c0, 32'shc4a038d6, 32'shc4a0cef4, 
               32'shc4a1651c, 32'shc4a1fb4e, 32'shc4a29188, 32'shc4a327cb, 32'shc4a3be18, 32'shc4a4546e, 32'shc4a4eacd, 32'shc4a58135, 
               32'shc4a617a6, 32'shc4a6ae21, 32'shc4a744a4, 32'shc4a7db31, 32'shc4a871c7, 32'shc4a90866, 32'shc4a99f0e, 32'shc4aa35bf, 
               32'shc4aacc7a, 32'shc4ab633d, 32'shc4abfa0a, 32'shc4ac90e0, 32'shc4ad27bf, 32'shc4adbea7, 32'shc4ae5599, 32'shc4aeec93, 
               32'shc4af8397, 32'shc4b01aa4, 32'shc4b0b1ba, 32'shc4b148d9, 32'shc4b1e001, 32'shc4b27732, 32'shc4b30e6d, 32'shc4b3a5b1, 
               32'shc4b43cfd, 32'shc4b4d453, 32'shc4b56bb3, 32'shc4b6031b, 32'shc4b69a8c, 32'shc4b73207, 32'shc4b7c98a, 32'shc4b86117, 
               32'shc4b8f8ad, 32'shc4b9904c, 32'shc4ba27f5, 32'shc4babfa6, 32'shc4bb5760, 32'shc4bbef24, 32'shc4bc86f1, 32'shc4bd1ec7, 
               32'shc4bdb6a6, 32'shc4be4e8e, 32'shc4bee680, 32'shc4bf7e7a, 32'shc4c0167e, 32'shc4c0ae8b, 32'shc4c146a0, 32'shc4c1dec0, 
               32'shc4c276e8, 32'shc4c30f19, 32'shc4c3a753, 32'shc4c43f97, 32'shc4c4d7e4, 32'shc4c5703a, 32'shc4c60899, 32'shc4c6a101, 
               32'shc4c73972, 32'shc4c7d1ec, 32'shc4c86a70, 32'shc4c902fd, 32'shc4c99b92, 32'shc4ca3431, 32'shc4caccd9, 32'shc4cb658b, 
               32'shc4cbfe45, 32'shc4cc9708, 32'shc4cd2fd5, 32'shc4cdc8ab, 32'shc4ce6189, 32'shc4cefa71, 32'shc4cf9363, 32'shc4d02c5d, 
               32'shc4d0c560, 32'shc4d15e6d, 32'shc4d1f782, 32'shc4d290a1, 32'shc4d329c9, 32'shc4d3c2fa, 32'shc4d45c34, 32'shc4d4f577, 
               32'shc4d58ec3, 32'shc4d62819, 32'shc4d6c177, 32'shc4d75adf, 32'shc4d7f450, 32'shc4d88dca, 32'shc4d9274d, 32'shc4d9c0d9, 
               32'shc4da5a6f, 32'shc4daf40d, 32'shc4db8db5, 32'shc4dc2765, 32'shc4dcc11f, 32'shc4dd5ae2, 32'shc4ddf4ae, 32'shc4de8e83, 
               32'shc4df2862, 32'shc4dfc249, 32'shc4e05c3a, 32'shc4e0f633, 32'shc4e19036, 32'shc4e22a42, 32'shc4e2c457, 32'shc4e35e75, 
               32'shc4e3f89c, 32'shc4e492cd, 32'shc4e52d06, 32'shc4e5c749, 32'shc4e66194, 32'shc4e6fbe9, 32'shc4e79647, 32'shc4e830ae, 
               32'shc4e8cb1e, 32'shc4e96597, 32'shc4ea001a, 32'shc4ea9aa5, 32'shc4eb353a, 32'shc4ebcfd8, 32'shc4ec6a7e, 32'shc4ed052e, 
               32'shc4ed9fe7, 32'shc4ee3aa9, 32'shc4eed575, 32'shc4ef7049, 32'shc4f00b27, 32'shc4f0a60d, 32'shc4f140fd, 32'shc4f1dbf6, 
               32'shc4f276f7, 32'shc4f31202, 32'shc4f3ad17, 32'shc4f44834, 32'shc4f4e35a, 32'shc4f57e8a, 32'shc4f619c2, 32'shc4f6b504, 
               32'shc4f7504e, 32'shc4f7eba2, 32'shc4f886ff, 32'shc4f92265, 32'shc4f9bdd4, 32'shc4fa594d, 32'shc4faf4ce, 32'shc4fb9059, 
               32'shc4fc2bec, 32'shc4fcc789, 32'shc4fd632f, 32'shc4fdfedd, 32'shc4fe9a95, 32'shc4ff3656, 32'shc4ffd221, 32'shc5006df4, 
               32'shc50109d0, 32'shc501a5b6, 32'shc50241a4, 32'shc502dd9c, 32'shc503799d, 32'shc50415a6, 32'shc504b1b9, 32'shc5054dd5, 
               32'shc505e9fb, 32'shc5068629, 32'shc5072260, 32'shc507bea1, 32'shc5085aea, 32'shc508f73d, 32'shc5099398, 32'shc50a2ffd, 
               32'shc50acc6b, 32'shc50b68e2, 32'shc50c0562, 32'shc50ca1eb, 32'shc50d3e7d, 32'shc50ddb19, 32'shc50e77bd, 32'shc50f146b, 
               32'shc50fb121, 32'shc5104de1, 32'shc510eaaa, 32'shc511877c, 32'shc5122457, 32'shc512c13b, 32'shc5135e28, 32'shc513fb1e, 
               32'shc514981d, 32'shc5153526, 32'shc515d237, 32'shc5166f52, 32'shc5170c75, 32'shc517a9a2, 32'shc51846d8, 32'shc518e417, 
               32'shc519815f, 32'shc51a1eb0, 32'shc51abc0a, 32'shc51b596d, 32'shc51bf6da, 32'shc51c944f, 32'shc51d31ce, 32'shc51dcf55, 
               32'shc51e6ce6, 32'shc51f0a7f, 32'shc51fa822, 32'shc52045ce, 32'shc520e383, 32'shc5218141, 32'shc5221f08, 32'shc522bcd9, 
               32'shc5235ab2, 32'shc523f894, 32'shc5249680, 32'shc5253474, 32'shc525d272, 32'shc5267078, 32'shc5270e88, 32'shc527aca1, 
               32'shc5284ac3, 32'shc528e8ee, 32'shc5298722, 32'shc52a255f, 32'shc52ac3a5, 32'shc52b61f4, 32'shc52c004d, 32'shc52c9eae, 
               32'shc52d3d18, 32'shc52ddb8c, 32'shc52e7a09, 32'shc52f188e, 32'shc52fb71d, 32'shc53055b5, 32'shc530f456, 32'shc5319300, 
               32'shc53231b3, 32'shc532d06f, 32'shc5336f34, 32'shc5340e02, 32'shc534acd9, 32'shc5354bba, 32'shc535eaa3, 32'shc5368996, 
               32'shc5372891, 32'shc537c796, 32'shc53866a4, 32'shc53905ba, 32'shc539a4da, 32'shc53a4403, 32'shc53ae335, 32'shc53b8270, 
               32'shc53c21b4, 32'shc53cc101, 32'shc53d6057, 32'shc53dffb7, 32'shc53e9f1f, 32'shc53f3e90, 32'shc53fde0b, 32'shc5407d8e, 
               32'shc5411d1b, 32'shc541bcb1, 32'shc5425c4f, 32'shc542fbf7, 32'shc5439ba8, 32'shc5443b62, 32'shc544db25, 32'shc5457af1, 
               32'shc5461ac6, 32'shc546baa4, 32'shc5475a8b, 32'shc547fa7b, 32'shc5489a74, 32'shc5493a76, 32'shc549da82, 32'shc54a7a96, 
               32'shc54b1ab4, 32'shc54bbada, 32'shc54c5b0a, 32'shc54cfb42, 32'shc54d9b84, 32'shc54e3bcf, 32'shc54edc23, 32'shc54f7c7f, 
               32'shc5501ce5, 32'shc550bd54, 32'shc5515dcc, 32'shc551fe4d, 32'shc5529ed7, 32'shc5533f6b, 32'shc553e007, 32'shc55480ac, 
               32'shc555215a, 32'shc555c211, 32'shc55662d2, 32'shc557039b, 32'shc557a46e, 32'shc5584549, 32'shc558e62e, 32'shc559871b, 
               32'shc55a2812, 32'shc55ac912, 32'shc55b6a1a, 32'shc55c0b2c, 32'shc55cac47, 32'shc55d4d6b, 32'shc55dee98, 32'shc55e8fce, 
               32'shc55f310d, 32'shc55fd255, 32'shc56073a6, 32'shc5611500, 32'shc561b663, 32'shc56257cf, 32'shc562f944, 32'shc5639ac3, 
               32'shc5643c4a, 32'shc564ddda, 32'shc5657f74, 32'shc5662116, 32'shc566c2c2, 32'shc5676476, 32'shc5680634, 32'shc568a7fa, 
               32'shc56949ca, 32'shc569eba2, 32'shc56a8d84, 32'shc56b2f6f, 32'shc56bd163, 32'shc56c735f, 32'shc56d1565, 32'shc56db774, 
               32'shc56e598c, 32'shc56efbad, 32'shc56f9dd7, 32'shc570400a, 32'shc570e246, 32'shc571848b, 32'shc57226d9, 32'shc572c930, 
               32'shc5736b90, 32'shc5740df9, 32'shc574b06b, 32'shc57552e6, 32'shc575f56b, 32'shc57697f8, 32'shc5773a8e, 32'shc577dd2d, 
               32'shc5787fd6, 32'shc5792287, 32'shc579c542, 32'shc57a6805, 32'shc57b0ad1, 32'shc57bada7, 32'shc57c5085, 32'shc57cf36d, 
               32'shc57d965d, 32'shc57e3957, 32'shc57edc5a, 32'shc57f7f65, 32'shc580227a, 32'shc580c597, 32'shc58168be, 32'shc5820bee, 
               32'shc582af26, 32'shc5835268, 32'shc583f5b3, 32'shc5849907, 32'shc5853c63, 32'shc585dfc9, 32'shc5868338, 32'shc58726b0, 
               32'shc587ca31, 32'shc5886dbb, 32'shc589114e, 32'shc589b4e9, 32'shc58a588e, 32'shc58afc3c, 32'shc58b9ff3, 32'shc58c43b3, 
               32'shc58ce77c, 32'shc58d8b4e, 32'shc58e2f29, 32'shc58ed30d, 32'shc58f76fa, 32'shc5901af0, 32'shc590beef, 32'shc59162f7, 
               32'shc5920708, 32'shc592ab22, 32'shc5934f46, 32'shc593f372, 32'shc59497a7, 32'shc5953be5, 32'shc595e02c, 32'shc596847c, 
               32'shc59728d5, 32'shc597cd38, 32'shc59871a3, 32'shc5991617, 32'shc599ba94, 32'shc59a5f1a, 32'shc59b03a9, 32'shc59ba842, 
               32'shc59c4ce3, 32'shc59cf18d, 32'shc59d9640, 32'shc59e3afc, 32'shc59edfc2, 32'shc59f8490, 32'shc5a02967, 32'shc5a0ce47, 
               32'shc5a17330, 32'shc5a21823, 32'shc5a2bd1e, 32'shc5a36222, 32'shc5a4072f, 32'shc5a4ac46, 32'shc5a55165, 32'shc5a5f68d, 
               32'shc5a69bbe, 32'shc5a740f8, 32'shc5a7e63c, 32'shc5a88b88, 32'shc5a930dd, 32'shc5a9d63b, 32'shc5aa7ba3, 32'shc5ab2113, 
               32'shc5abc68c, 32'shc5ac6c0e, 32'shc5ad1199, 32'shc5adb72d, 32'shc5ae5ccb, 32'shc5af0271, 32'shc5afa820, 32'shc5b04dd8, 
               32'shc5b0f399, 32'shc5b19963, 32'shc5b23f37, 32'shc5b2e513, 32'shc5b38af8, 32'shc5b430e6, 32'shc5b4d6dd, 32'shc5b57cdd, 
               32'shc5b622e6, 32'shc5b6c8f8, 32'shc5b76f13, 32'shc5b81537, 32'shc5b8bb64, 32'shc5b9619a, 32'shc5ba07d9, 32'shc5baae21, 
               32'shc5bb5472, 32'shc5bbfacc, 32'shc5bca12f, 32'shc5bd479b, 32'shc5bdee10, 32'shc5be948e, 32'shc5bf3b15, 32'shc5bfe1a5, 
               32'shc5c0883d, 32'shc5c12edf, 32'shc5c1d58a, 32'shc5c27c3e, 32'shc5c322fb, 32'shc5c3c9c0, 32'shc5c4708f, 32'shc5c51767, 
               32'shc5c5be47, 32'shc5c66531, 32'shc5c70c24, 32'shc5c7b31f, 32'shc5c85a24, 32'shc5c90132, 32'shc5c9a848, 32'shc5ca4f68, 
               32'shc5caf690, 32'shc5cb9dc2, 32'shc5cc44fc, 32'shc5ccec40, 32'shc5cd938c, 32'shc5ce3ae1, 32'shc5cee240, 32'shc5cf89a7, 
               32'shc5d03118, 32'shc5d0d891, 32'shc5d18013, 32'shc5d2279e, 32'shc5d2cf33, 32'shc5d376d0, 32'shc5d41e76, 32'shc5d4c625, 
               32'shc5d56ddd, 32'shc5d6159e, 32'shc5d6bd68, 32'shc5d7653b, 32'shc5d80d17, 32'shc5d8b4fc, 32'shc5d95cea, 32'shc5da04e1, 
               32'shc5daace1, 32'shc5db54e9, 32'shc5dbfcfb, 32'shc5dca516, 32'shc5dd4d3a, 32'shc5ddf566, 32'shc5de9d9c, 32'shc5df45db, 
               32'shc5dfee22, 32'shc5e09673, 32'shc5e13ecc, 32'shc5e1e72f, 32'shc5e28f9a, 32'shc5e3380e, 32'shc5e3e08c, 32'shc5e48912, 
               32'shc5e531a1, 32'shc5e5da3a, 32'shc5e682db, 32'shc5e72b85, 32'shc5e7d438, 32'shc5e87cf4, 32'shc5e925b9, 32'shc5e9ce87, 
               32'shc5ea775e, 32'shc5eb203e, 32'shc5ebc927, 32'shc5ec7218, 32'shc5ed1b13, 32'shc5edc417, 32'shc5ee6d24, 32'shc5ef1639, 
               32'shc5efbf58, 32'shc5f0687f, 32'shc5f111b0, 32'shc5f1bae9, 32'shc5f2642c, 32'shc5f30d77, 32'shc5f3b6cb, 32'shc5f46029, 
               32'shc5f5098f, 32'shc5f5b2fe, 32'shc5f65c76, 32'shc5f705f7, 32'shc5f7af81, 32'shc5f85914, 32'shc5f902b0, 32'shc5f9ac55, 
               32'shc5fa5603, 32'shc5faffb9, 32'shc5fba979, 32'shc5fc5342, 32'shc5fcfd13, 32'shc5fda6ee, 32'shc5fe50d1, 32'shc5fefabe, 
               32'shc5ffa4b3, 32'shc6004eb1, 32'shc600f8b9, 32'shc601a2c9, 32'shc6024ce2, 32'shc602f704, 32'shc603a12f, 32'shc6044b63, 
               32'shc604f5a0, 32'shc6059fe6, 32'shc6064a35, 32'shc606f48c, 32'shc6079eed, 32'shc6084957, 32'shc608f3c9, 32'shc6099e45, 
               32'shc60a48c9, 32'shc60af357, 32'shc60b9ded, 32'shc60c488c, 32'shc60cf334, 32'shc60d9de5, 32'shc60e489f, 32'shc60ef362, 
               32'shc60f9e2e, 32'shc6104903, 32'shc610f3e1, 32'shc6119ec8, 32'shc61249b7, 32'shc612f4b0, 32'shc6139fb2, 32'shc6144abc, 
               32'shc614f5cf, 32'shc615a0ec, 32'shc6164c11, 32'shc616f73f, 32'shc617a276, 32'shc6184db6, 32'shc618f8ff, 32'shc619a451, 
               32'shc61a4fac, 32'shc61afb10, 32'shc61ba67d, 32'shc61c51f2, 32'shc61cfd71, 32'shc61da8f8, 32'shc61e5489, 32'shc61f0022, 
               32'shc61fabc4, 32'shc620576f, 32'shc6210323, 32'shc621aee1, 32'shc6225aa6, 32'shc6230675, 32'shc623b24d, 32'shc6245e2e, 
               32'shc6250a18, 32'shc625b60a, 32'shc6266206, 32'shc6270e0a, 32'shc627ba17, 32'shc628662e, 32'shc629124d, 32'shc629be75, 
               32'shc62a6aa6, 32'shc62b16e0, 32'shc62bc323, 32'shc62c6f6e, 32'shc62d1bc3, 32'shc62dc821, 32'shc62e7487, 32'shc62f20f7, 
               32'shc62fcd6f, 32'shc63079f0, 32'shc631267a, 32'shc631d30e, 32'shc6327faa, 32'shc6332c4e, 32'shc633d8fc, 32'shc63485b3, 
               32'shc6353273, 32'shc635df3b, 32'shc6368c0d, 32'shc63738e7, 32'shc637e5ca, 32'shc63892b7, 32'shc6393fac, 32'shc639ecaa, 
               32'shc63a99b1, 32'shc63b46c1, 32'shc63bf3d9, 32'shc63ca0fb, 32'shc63d4e26, 32'shc63dfb59, 32'shc63ea896, 32'shc63f55db, 
               32'shc6400329, 32'shc640b080, 32'shc6415de0, 32'shc6420b49, 32'shc642b8bb, 32'shc6436636, 32'shc64413b9, 32'shc644c146, 
               32'shc6456edb, 32'shc6461c7a, 32'shc646ca21, 32'shc64777d1, 32'shc648258a, 32'shc648d34c, 32'shc6498117, 32'shc64a2eeb, 
               32'shc64adcc7, 32'shc64b8aad, 32'shc64c389b, 32'shc64ce693, 32'shc64d9493, 32'shc64e429c, 32'shc64ef0ae, 32'shc64f9ec9, 
               32'shc6504ced, 32'shc650fb1a, 32'shc651a94f, 32'shc652578e, 32'shc65305d5, 32'shc653b426, 32'shc654627f, 32'shc65510e1, 
               32'shc655bf4c, 32'shc6566dc0, 32'shc6571c3c, 32'shc657cac2, 32'shc6587951, 32'shc65927e8, 32'shc659d688, 32'shc65a8532, 
               32'shc65b33e4, 32'shc65be29f, 32'shc65c9163, 32'shc65d4030, 32'shc65def05, 32'shc65e9de4, 32'shc65f4ccb, 32'shc65ffbbc, 
               32'shc660aab5, 32'shc66159b7, 32'shc66208c2, 32'shc662b7d6, 32'shc66366f3, 32'shc6641618, 32'shc664c547, 32'shc665747e, 
               32'shc66623be, 32'shc666d308, 32'shc667825a, 32'shc66831b5, 32'shc668e119, 32'shc6699085, 32'shc66a3ffb, 32'shc66aef79, 
               32'shc66b9f01, 32'shc66c4e91, 32'shc66cfe2a, 32'shc66dadcc, 32'shc66e5d77, 32'shc66f0d2b, 32'shc66fbce7, 32'shc6706cad, 
               32'shc6711c7b, 32'shc671cc52, 32'shc6727c32, 32'shc6732c1b, 32'shc673dc0d, 32'shc6748c08, 32'shc6753c0c, 32'shc675ec18, 
               32'shc6769c2e, 32'shc6774c4c, 32'shc677fc73, 32'shc678aca3, 32'shc6795cdc, 32'shc67a0d1e, 32'shc67abd68, 32'shc67b6dbc, 
               32'shc67c1e18, 32'shc67cce7d, 32'shc67d7eeb, 32'shc67e2f62, 32'shc67edfe2, 32'shc67f906b, 32'shc68040fc, 32'shc680f197, 
               32'shc681a23a, 32'shc68252e6, 32'shc683039b, 32'shc683b459, 32'shc6846520, 32'shc68515f0, 32'shc685c6c8, 32'shc68677a9, 
               32'shc6872894, 32'shc687d987, 32'shc6888a83, 32'shc6893b87, 32'shc689ec95, 32'shc68a9dac, 32'shc68b4ecb, 32'shc68bfff3, 
               32'shc68cb124, 32'shc68d625e, 32'shc68e13a1, 32'shc68ec4ed, 32'shc68f7641, 32'shc690279f, 32'shc690d905, 32'shc6918a74, 
               32'shc6923bec, 32'shc692ed6d, 32'shc6939ef6, 32'shc6945089, 32'shc6950224, 32'shc695b3c9, 32'shc6966576, 32'shc697172c, 
               32'shc697c8eb, 32'shc6987ab2, 32'shc6992c83, 32'shc699de5c, 32'shc69a903e, 32'shc69b4229, 32'shc69bf41d, 32'shc69ca61a, 
               32'shc69d5820, 32'shc69e0a2e, 32'shc69ebc45, 32'shc69f6e66, 32'shc6a0208f, 32'shc6a0d2c0, 32'shc6a184fb, 32'shc6a2373f, 
               32'shc6a2e98b, 32'shc6a39be0, 32'shc6a44e3e, 32'shc6a500a5, 32'shc6a5b315, 32'shc6a6658e, 32'shc6a7180f, 32'shc6a7ca9a, 
               32'shc6a87d2d, 32'shc6a92fc9, 32'shc6a9e26e, 32'shc6aa951b, 32'shc6ab47d2, 32'shc6abfa91, 32'shc6acad59, 32'shc6ad602a, 
               32'shc6ae1304, 32'shc6aec5e7, 32'shc6af78d3, 32'shc6b02bc7, 32'shc6b0dec4, 32'shc6b191ca, 32'shc6b244d9, 32'shc6b2f7f1, 
               32'shc6b3ab12, 32'shc6b45e3b, 32'shc6b5116d, 32'shc6b5c4a8, 32'shc6b677ec, 32'shc6b72b39, 32'shc6b7de8f, 32'shc6b891ed, 
               32'shc6b94554, 32'shc6b9f8c5, 32'shc6baac3d, 32'shc6bb5fbf, 32'shc6bc134a, 32'shc6bcc6dd, 32'shc6bd7a7a, 32'shc6be2e1f, 
               32'shc6bee1cd, 32'shc6bf9583, 32'shc6c04943, 32'shc6c0fd0b, 32'shc6c1b0dd, 32'shc6c264b7, 32'shc6c31899, 32'shc6c3cc85, 
               32'shc6c4807a, 32'shc6c53477, 32'shc6c5e87d, 32'shc6c69c8c, 32'shc6c750a4, 32'shc6c804c5, 32'shc6c8b8ee, 32'shc6c96d21, 
               32'shc6ca215c, 32'shc6cad5a0, 32'shc6cb89ed, 32'shc6cc3e42, 32'shc6ccf2a1, 32'shc6cda708, 32'shc6ce5b78, 32'shc6cf0ff1, 
               32'shc6cfc472, 32'shc6d078fd, 32'shc6d12d90, 32'shc6d1e22d, 32'shc6d296d1, 32'shc6d34b7f, 32'shc6d40036, 32'shc6d4b4f5, 
               32'shc6d569be, 32'shc6d61e8f, 32'shc6d6d369, 32'shc6d7884b, 32'shc6d83d37, 32'shc6d8f22b, 32'shc6d9a728, 32'shc6da5c2e, 
               32'shc6db113d, 32'shc6dbc654, 32'shc6dc7b75, 32'shc6dd309e, 32'shc6dde5d0, 32'shc6de9b0b, 32'shc6df504f, 32'shc6e0059b, 
               32'shc6e0baf0, 32'shc6e1704e, 32'shc6e225b5, 32'shc6e2db25, 32'shc6e3909d, 32'shc6e4461f, 32'shc6e4fba9, 32'shc6e5b13c, 
               32'shc6e666d7, 32'shc6e71c7c, 32'shc6e7d229, 32'shc6e887df, 32'shc6e93d9e, 32'shc6e9f366, 32'shc6eaa936, 32'shc6eb5f10, 
               32'shc6ec14f2, 32'shc6eccadd, 32'shc6ed80d1, 32'shc6ee36cd, 32'shc6eeecd3, 32'shc6efa2e1, 32'shc6f058f8, 32'shc6f10f17, 
               32'shc6f1c540, 32'shc6f27b71, 32'shc6f331ab, 32'shc6f3e7ee, 32'shc6f49e3a, 32'shc6f5548f, 32'shc6f60aec, 32'shc6f6c152, 
               32'shc6f777c1, 32'shc6f82e39, 32'shc6f8e4b9, 32'shc6f99b43, 32'shc6fa51d5, 32'shc6fb0870, 32'shc6fbbf13, 32'shc6fc75c0, 
               32'shc6fd2c75, 32'shc6fde333, 32'shc6fe99fa, 32'shc6ff50ca, 32'shc70007a2, 32'shc700be83, 32'shc701756d, 32'shc7022c60, 
               32'shc702e35c, 32'shc7039a60, 32'shc704516d, 32'shc7050883, 32'shc705bfa2, 32'shc70676ca, 32'shc7072dfa, 32'shc707e533, 
               32'shc7089c75, 32'shc70953c0, 32'shc70a0b13, 32'shc70ac26f, 32'shc70b79d4, 32'shc70c3142, 32'shc70ce8b9, 32'shc70da038, 
               32'shc70e57c0, 32'shc70f0f51, 32'shc70fc6eb, 32'shc7107e8d, 32'shc7113639, 32'shc711eded, 32'shc712a5aa, 32'shc7135d6f, 
               32'shc714153e, 32'shc714cd15, 32'shc71584f5, 32'shc7163cdd, 32'shc716f4cf, 32'shc717acc9, 32'shc71864cc, 32'shc7191cd8, 
               32'shc719d4ed, 32'shc71a8d0a, 32'shc71b4530, 32'shc71bfd5f, 32'shc71cb597, 32'shc71d6dd7, 32'shc71e2621, 32'shc71ede73, 
               32'shc71f96ce, 32'shc7204f31, 32'shc721079d, 32'shc721c013, 32'shc7227890, 32'shc7233117, 32'shc723e9a6, 32'shc724a23f, 
               32'shc7255ae0, 32'shc7261389, 32'shc726cc3c, 32'shc72784f7, 32'shc7283dbb, 32'shc728f688, 32'shc729af5d, 32'shc72a683c, 
               32'shc72b2123, 32'shc72bda13, 32'shc72c930b, 32'shc72d4c0d, 32'shc72e0517, 32'shc72ebe2a, 32'shc72f7745, 32'shc730306a, 
               32'shc730e997, 32'shc731a2cd, 32'shc7325c0c, 32'shc7331553, 32'shc733cea3, 32'shc73487fc, 32'shc735415e, 32'shc735fac8, 
               32'shc736b43c, 32'shc7376db8, 32'shc738273d, 32'shc738e0ca, 32'shc7399a60, 32'shc73a53ff, 32'shc73b0da7, 32'shc73bc758, 
               32'shc73c8111, 32'shc73d3ad3, 32'shc73df49e, 32'shc73eae71, 32'shc73f684e, 32'shc7402233, 32'shc740dc21, 32'shc7419617, 
               32'shc7425016, 32'shc7430a1f, 32'shc743c42f, 32'shc7447e49, 32'shc745386b, 32'shc745f296, 32'shc746acca, 32'shc7476707, 
               32'shc748214c, 32'shc748db9a, 32'shc74995f1, 32'shc74a5050, 32'shc74b0ab9, 32'shc74bc52a, 32'shc74c7fa4, 32'shc74d3a26, 
               32'shc74df4b1, 32'shc74eaf45, 32'shc74f69e2, 32'shc7502488, 32'shc750df36, 32'shc75199ed, 32'shc75254ac, 32'shc7530f75, 
               32'shc753ca46, 32'shc7548520, 32'shc7554003, 32'shc755faee, 32'shc756b5e2, 32'shc75770df, 32'shc7582be5, 32'shc758e6f3, 
               32'shc759a20a, 32'shc75a5d2a, 32'shc75b1853, 32'shc75bd384, 32'shc75c8ebe, 32'shc75d4a01, 32'shc75e054c, 32'shc75ec0a1, 
               32'shc75f7bfe, 32'shc7603763, 32'shc760f2d2, 32'shc761ae49, 32'shc76269c9, 32'shc7632552, 32'shc763e0e3, 32'shc7649c7d, 
               32'shc7655820, 32'shc76613cb, 32'shc766cf80, 32'shc7678b3d, 32'shc7684702, 32'shc76902d1, 32'shc769bea8, 32'shc76a7a88, 
               32'shc76b3671, 32'shc76bf262, 32'shc76cae5c, 32'shc76d6a5f, 32'shc76e266b, 32'shc76ee27f, 32'shc76f9e9c, 32'shc7705ac2, 
               32'shc77116f0, 32'shc771d327, 32'shc7728f67, 32'shc7734bb0, 32'shc7740801, 32'shc774c45b, 32'shc77580be, 32'shc7763d29, 
               32'shc776f99d, 32'shc777b61a, 32'shc77872a0, 32'shc7792f2e, 32'shc779ebc5, 32'shc77aa865, 32'shc77b650e, 32'shc77c21bf, 
               32'shc77cde79, 32'shc77d9b3c, 32'shc77e5807, 32'shc77f14db, 32'shc77fd1b8, 32'shc7808e9d, 32'shc7814b8c, 32'shc7820883, 
               32'shc782c582, 32'shc783828b, 32'shc7843f9c, 32'shc784fcb5, 32'shc785b9d8, 32'shc7867703, 32'shc7873437, 32'shc787f174, 
               32'shc788aeb9, 32'shc7896c07, 32'shc78a295e, 32'shc78ae6bd, 32'shc78ba425, 32'shc78c6196, 32'shc78d1f10, 32'shc78ddc92, 
               32'shc78e9a1d, 32'shc78f57b1, 32'shc790154d, 32'shc790d2f2, 32'shc79190a0, 32'shc7924e56, 32'shc7930c16, 32'shc793c9de, 
               32'shc79487ae, 32'shc7954587, 32'shc7960369, 32'shc796c154, 32'shc7977f48, 32'shc7983d44, 32'shc798fb48, 32'shc799b956, 
               32'shc79a776c, 32'shc79b358b, 32'shc79bf3b3, 32'shc79cb1e3, 32'shc79d701c, 32'shc79e2e5d, 32'shc79eeca8, 32'shc79faafb, 
               32'shc7a06957, 32'shc7a127bb, 32'shc7a1e628, 32'shc7a2a49e, 32'shc7a3631d, 32'shc7a421a4, 32'shc7a4e034, 32'shc7a59ecc, 
               32'shc7a65d6e, 32'shc7a71c18, 32'shc7a7daca, 32'shc7a89986, 32'shc7a9584a, 32'shc7aa1716, 32'shc7aad5ec, 32'shc7ab94ca, 
               32'shc7ac53b1, 32'shc7ad12a0, 32'shc7add198, 32'shc7ae9099, 32'shc7af4fa3, 32'shc7b00eb5, 32'shc7b0cdd0, 32'shc7b18cf3, 
               32'shc7b24c20, 32'shc7b30b55, 32'shc7b3ca92, 32'shc7b489d9, 32'shc7b54928, 32'shc7b6087f, 32'shc7b6c7e0, 32'shc7b78749, 
               32'shc7b846ba, 32'shc7b90635, 32'shc7b9c5b8, 32'shc7ba8544, 32'shc7bb44d8, 32'shc7bc0475, 32'shc7bcc41b, 32'shc7bd83ca, 
               32'shc7be4381, 32'shc7bf0340, 32'shc7bfc309, 32'shc7c082da, 32'shc7c142b4, 32'shc7c20297, 32'shc7c2c282, 32'shc7c38276, 
               32'shc7c44272, 32'shc7c50277, 32'shc7c5c285, 32'shc7c6829c, 32'shc7c742bb, 32'shc7c802e3, 32'shc7c8c313, 32'shc7c9834d, 
               32'shc7ca438f, 32'shc7cb03d9, 32'shc7cbc42c, 32'shc7cc8488, 32'shc7cd44ed, 32'shc7ce055a, 32'shc7cec5d0, 32'shc7cf864e, 
               32'shc7d046d6, 32'shc7d10766, 32'shc7d1c7fe, 32'shc7d2889f, 32'shc7d34949, 32'shc7d409fc, 32'shc7d4cab7, 32'shc7d58b7b, 
               32'shc7d64c47, 32'shc7d70d1d, 32'shc7d7cdfb, 32'shc7d88ee1, 32'shc7d94fd0, 32'shc7da10c8, 32'shc7dad1c9, 32'shc7db92d2, 
               32'shc7dc53e3, 32'shc7dd14fe, 32'shc7ddd621, 32'shc7de974d, 32'shc7df5881, 32'shc7e019be, 32'shc7e0db04, 32'shc7e19c53, 
               32'shc7e25daa, 32'shc7e31f09, 32'shc7e3e072, 32'shc7e4a1e3, 32'shc7e5635c, 32'shc7e624df, 32'shc7e6e66a, 32'shc7e7a7fd, 
               32'shc7e8699a, 32'shc7e92b3e, 32'shc7e9ecec, 32'shc7eaaea2, 32'shc7eb7061, 32'shc7ec3229, 32'shc7ecf3f9, 32'shc7edb5d2, 
               32'shc7ee77b3, 32'shc7ef399d, 32'shc7effb90, 32'shc7f0bd8b, 32'shc7f17f8f, 32'shc7f2419c, 32'shc7f303b1, 32'shc7f3c5cf, 
               32'shc7f487f6, 32'shc7f54a25, 32'shc7f60c5d, 32'shc7f6ce9e, 32'shc7f790e7, 32'shc7f85339, 32'shc7f91593, 32'shc7f9d7f6, 
               32'shc7fa9a62, 32'shc7fb5cd7, 32'shc7fc1f54, 32'shc7fce1d9, 32'shc7fda468, 32'shc7fe66fe, 32'shc7ff299e, 32'shc7ffec46, 
               32'shc800aef7, 32'shc80171b1, 32'shc8023473, 32'shc802f73d, 32'shc803ba11, 32'shc8047ced, 32'shc8053fd2, 32'shc80602bf, 
               32'shc806c5b5, 32'shc80788b3, 32'shc8084bba, 32'shc8090eca, 32'shc809d1e3, 32'shc80a9504, 32'shc80b582e, 32'shc80c1b60, 
               32'shc80cde9b, 32'shc80da1de, 32'shc80e652b, 32'shc80f287f, 32'shc80febdd, 32'shc810af43, 32'shc81172b2, 32'shc8123629, 
               32'shc812f9a9, 32'shc813bd32, 32'shc81480c3, 32'shc815445d, 32'shc81607ff, 32'shc816cbaa, 32'shc8178f5e, 32'shc818531a, 
               32'shc81916df, 32'shc819daad, 32'shc81a9e83, 32'shc81b6262, 32'shc81c2649, 32'shc81cea39, 32'shc81dae32, 32'shc81e7233, 
               32'shc81f363d, 32'shc81ffa50, 32'shc820be6b, 32'shc821828f, 32'shc82246bb, 32'shc8230af0, 32'shc823cf2e, 32'shc8249374, 
               32'shc82557c3, 32'shc8261c1a, 32'shc826e07a, 32'shc827a4e3, 32'shc8286954, 32'shc8292dce, 32'shc829f251, 32'shc82ab6dc, 
               32'shc82b7b70, 32'shc82c400c, 32'shc82d04b1, 32'shc82dc95e, 32'shc82e8e15, 32'shc82f52d3, 32'shc830179b, 32'shc830dc6b, 
               32'shc831a143, 32'shc8326625, 32'shc8332b0e, 32'shc833f001, 32'shc834b4fc, 32'shc83579ff, 32'shc8363f0c, 32'shc8370420, 
               32'shc837c93e, 32'shc8388e64, 32'shc8395393, 32'shc83a18ca, 32'shc83ade0a, 32'shc83ba352, 32'shc83c68a3, 32'shc83d2dfd, 
               32'shc83df35f, 32'shc83eb8ca, 32'shc83f7e3d, 32'shc84043b9, 32'shc841093e, 32'shc841cecb, 32'shc8429461, 32'shc84359ff, 
               32'shc8441fa6, 32'shc844e556, 32'shc845ab0e, 32'shc84670cf, 32'shc8473698, 32'shc847fc6a, 32'shc848c245, 32'shc8498828, 
               32'shc84a4e14, 32'shc84b1408, 32'shc84bda05, 32'shc84ca00b, 32'shc84d6619, 32'shc84e2c2f, 32'shc84ef24f, 32'shc84fb877, 
               32'shc8507ea7, 32'shc85144e0, 32'shc8520b22, 32'shc852d16c, 32'shc85397bf, 32'shc8545e1a, 32'shc855247e, 32'shc855eaeb, 
               32'shc856b160, 32'shc85777de, 32'shc8583e64, 32'shc85904f3, 32'shc859cb8a, 32'shc85a922b, 32'shc85b58d3, 32'shc85c1f84, 
               32'shc85ce63e, 32'shc85dad01, 32'shc85e73cc, 32'shc85f3a9f, 32'shc860017b, 32'shc860c860, 32'shc8618f4d, 32'shc8625643, 
               32'shc8631d42, 32'shc863e449, 32'shc864ab58, 32'shc8657270, 32'shc8663991, 32'shc86700ba, 32'shc867c7ec, 32'shc8688f27, 
               32'shc869566a, 32'shc86a1db6, 32'shc86ae50a, 32'shc86bac66, 32'shc86c73cc, 32'shc86d3b3a, 32'shc86e02b0, 32'shc86eca2f, 
               32'shc86f91b7, 32'shc8705947, 32'shc87120e0, 32'shc871e881, 32'shc872b02b, 32'shc87377dd, 32'shc8743f98, 32'shc875075c, 
               32'shc875cf28, 32'shc87696fd, 32'shc8775eda, 32'shc87826c0, 32'shc878eeae, 32'shc879b6a5, 32'shc87a7ea5, 32'shc87b46ad, 
               32'shc87c0ebd, 32'shc87cd6d7, 32'shc87d9ef8, 32'shc87e6723, 32'shc87f2f56, 32'shc87ff791, 32'shc880bfd5, 32'shc8818822, 
               32'shc8825077, 32'shc88318d5, 32'shc883e13b, 32'shc884a9aa, 32'shc8857221, 32'shc8863aa1, 32'shc8870329, 32'shc887cbba, 
               32'shc8889454, 32'shc8895cf6, 32'shc88a25a1, 32'shc88aee54, 32'shc88bb710, 32'shc88c7fd4, 32'shc88d48a1, 32'shc88e1176, 
               32'shc88eda54, 32'shc88fa33b, 32'shc8906c2a, 32'shc8913522, 32'shc891fe22, 32'shc892c72b, 32'shc893903c, 32'shc8945956, 
               32'shc8952278, 32'shc895eba3, 32'shc896b4d6, 32'shc8977e12, 32'shc8984757, 32'shc89910a4, 32'shc899d9fa, 32'shc89aa358, 
               32'shc89b6cbf, 32'shc89c362e, 32'shc89cffa6, 32'shc89dc926, 32'shc89e92af, 32'shc89f5c40, 32'shc8a025da, 32'shc8a0ef7d, 
               32'shc8a1b928, 32'shc8a282db, 32'shc8a34c98, 32'shc8a4165c, 32'shc8a4e029, 32'shc8a5a9ff, 32'shc8a673dd, 32'shc8a73dc4, 
               32'shc8a807b4, 32'shc8a8d1ac, 32'shc8a99bac, 32'shc8aa65b5, 32'shc8ab2fc6, 32'shc8abf9e0, 32'shc8acc403, 32'shc8ad8e2e, 
               32'shc8ae5862, 32'shc8af229e, 32'shc8afece2, 32'shc8b0b730, 32'shc8b18185, 32'shc8b24be4, 32'shc8b3164a, 32'shc8b3e0ba, 
               32'shc8b4ab32, 32'shc8b575b2, 32'shc8b6403b, 32'shc8b70acc, 32'shc8b7d566, 32'shc8b8a009, 32'shc8b96ab4, 32'shc8ba3567, 
               32'shc8bb0023, 32'shc8bbcae8, 32'shc8bc95b5, 32'shc8bd608b, 32'shc8be2b69, 32'shc8bef64f, 32'shc8bfc13f, 32'shc8c08c36, 
               32'shc8c15736, 32'shc8c2223f, 32'shc8c2ed50, 32'shc8c3b86a, 32'shc8c4838d, 32'shc8c54eb7, 32'shc8c619eb, 32'shc8c6e527, 
               32'shc8c7b06b, 32'shc8c87bb8, 32'shc8c9470d, 32'shc8ca126b, 32'shc8caddd1, 32'shc8cba940, 32'shc8cc74b8, 32'shc8cd4038, 
               32'shc8ce0bc0, 32'shc8ced751, 32'shc8cfa2eb, 32'shc8d06e8d, 32'shc8d13a37, 32'shc8d205ea, 32'shc8d2d1a6, 32'shc8d39d6a, 
               32'shc8d46936, 32'shc8d5350c, 32'shc8d600e9, 32'shc8d6cccf, 32'shc8d798be, 32'shc8d864b5, 32'shc8d930b4, 32'shc8d9fcbd, 
               32'shc8dac8cd, 32'shc8db94e6, 32'shc8dc6108, 32'shc8dd2d32, 32'shc8ddf965, 32'shc8dec5a0, 32'shc8df91e3, 32'shc8e05e2f, 
               32'shc8e12a84, 32'shc8e1f6e1, 32'shc8e2c347, 32'shc8e38fb5, 32'shc8e45c2c, 32'shc8e528ab, 32'shc8e5f532, 32'shc8e6c1c2, 
               32'shc8e78e5b, 32'shc8e85afc, 32'shc8e927a6, 32'shc8e9f458, 32'shc8eac112, 32'shc8eb8dd6, 32'shc8ec5aa1, 32'shc8ed2775, 
               32'shc8edf452, 32'shc8eec137, 32'shc8ef8e24, 32'shc8f05b1a, 32'shc8f12819, 32'shc8f1f520, 32'shc8f2c230, 32'shc8f38f48, 
               32'shc8f45c68, 32'shc8f52991, 32'shc8f5f6c3, 32'shc8f6c3fd, 32'shc8f7913f, 32'shc8f85e8a, 32'shc8f92bdd, 32'shc8f9f939, 
               32'shc8fac69e, 32'shc8fb940b, 32'shc8fc6180, 32'shc8fd2efe, 32'shc8fdfc84, 32'shc8feca13, 32'shc8ff97aa, 32'shc900654a, 
               32'shc90132f2, 32'shc90200a3, 32'shc902ce5c, 32'shc9039c1e, 32'shc90469e8, 32'shc90537bb, 32'shc9060596, 32'shc906d379, 
               32'shc907a166, 32'shc9086f5a, 32'shc9093d57, 32'shc90a0b5d, 32'shc90ad96b, 32'shc90ba781, 32'shc90c75a0, 32'shc90d43c8, 
               32'shc90e11f7, 32'shc90ee030, 32'shc90fae71, 32'shc9107cba, 32'shc9114b0c, 32'shc9121966, 32'shc912e7c9, 32'shc913b634, 
               32'shc91484a8, 32'shc9155324, 32'shc91621a8, 32'shc916f035, 32'shc917becb, 32'shc9188d69, 32'shc9195c0f, 32'shc91a2abe, 
               32'shc91af976, 32'shc91bc836, 32'shc91c96fe, 32'shc91d65cf, 32'shc91e34a8, 32'shc91f038a, 32'shc91fd274, 32'shc920a167, 
               32'shc9217062, 32'shc9223f65, 32'shc9230e71, 32'shc923dd86, 32'shc924aca3, 32'shc9257bc8, 32'shc9264af6, 32'shc9271a2d, 
               32'shc927e96b, 32'shc928b8b3, 32'shc9298802, 32'shc92a575a, 32'shc92b26bb, 32'shc92bf624, 32'shc92cc596, 32'shc92d9510, 
               32'shc92e6492, 32'shc92f341d, 32'shc93003b0, 32'shc930d34c, 32'shc931a2f0, 32'shc932729d, 32'shc9334252, 32'shc9341210, 
               32'shc934e1d6, 32'shc935b1a5, 32'shc936817b, 32'shc937515b, 32'shc9382143, 32'shc938f133, 32'shc939c12c, 32'shc93a912d, 
               32'shc93b6137, 32'shc93c3149, 32'shc93d0163, 32'shc93dd186, 32'shc93ea1b2, 32'shc93f71e6, 32'shc9404222, 32'shc9411267, 
               32'shc941e2b4, 32'shc942b30a, 32'shc9438368, 32'shc94453ce, 32'shc945243d, 32'shc945f4b4, 32'shc946c534, 32'shc94795bd, 
               32'shc948664d, 32'shc94936e7, 32'shc94a0788, 32'shc94ad832, 32'shc94ba8e5, 32'shc94c79a0, 32'shc94d4a63, 32'shc94e1b2f, 
               32'shc94eec03, 32'shc94fbce0, 32'shc9508dc5, 32'shc9515eb2, 32'shc9522fa8, 32'shc95300a6, 32'shc953d1ad, 32'shc954a2bc, 
               32'shc95573d4, 32'shc95644f4, 32'shc957161d, 32'shc957e74e, 32'shc958b887, 32'shc95989c9, 32'shc95a5b13, 32'shc95b2c66, 
               32'shc95bfdc1, 32'shc95ccf25, 32'shc95da090, 32'shc95e7205, 32'shc95f4382, 32'shc9601507, 32'shc960e695, 32'shc961b82b, 
               32'shc96289c9, 32'shc9635b70, 32'shc9642d1f, 32'shc964fed7, 32'shc965d097, 32'shc966a260, 32'shc9677431, 32'shc968460a, 
               32'shc96917ec, 32'shc969e9d7, 32'shc96abbc9, 32'shc96b8dc4, 32'shc96c5fc8, 32'shc96d31d4, 32'shc96e03e8, 32'shc96ed605, 
               32'shc96fa82a, 32'shc9707a58, 32'shc9714c8e, 32'shc9721ecc, 32'shc972f113, 32'shc973c362, 32'shc97495ba, 32'shc975681a, 
               32'shc9763a83, 32'shc9770cf4, 32'shc977df6d, 32'shc978b1ef, 32'shc9798479, 32'shc97a570b, 32'shc97b29a6, 32'shc97bfc4a, 
               32'shc97ccef5, 32'shc97da1aa, 32'shc97e7466, 32'shc97f472b, 32'shc98019f8, 32'shc980ecce, 32'shc981bfac, 32'shc9829293, 
               32'shc9836582, 32'shc9843879, 32'shc9850b79, 32'shc985de82, 32'shc986b192, 32'shc98784ab, 32'shc98857cd, 32'shc9892af6, 
               32'shc989fe29, 32'shc98ad163, 32'shc98ba4a6, 32'shc98c77f2, 32'shc98d4b45, 32'shc98e1ea2, 32'shc98ef206, 32'shc98fc573, 
               32'shc99098e9, 32'shc9916c66, 32'shc9923fed, 32'shc993137b, 32'shc993e712, 32'shc994bab1, 32'shc9958e59, 32'shc9966209, 
               32'shc99735c2, 32'shc9980983, 32'shc998dd4c, 32'shc999b11e, 32'shc99a84f8, 32'shc99b58da, 32'shc99c2cc5, 32'shc99d00b8, 
               32'shc99dd4b4, 32'shc99ea8b8, 32'shc99f7cc5, 32'shc9a050d9, 32'shc9a124f7, 32'shc9a1f91c, 32'shc9a2cd4a, 32'shc9a3a180, 
               32'shc9a475bf, 32'shc9a54a06, 32'shc9a61e56, 32'shc9a6f2ae, 32'shc9a7c70e, 32'shc9a89b76, 32'shc9a96fe7, 32'shc9aa4461, 
               32'shc9ab18e3, 32'shc9abed6d, 32'shc9acc1ff, 32'shc9ad969a, 32'shc9ae6b3d, 32'shc9af3fe9, 32'shc9b0149d, 32'shc9b0e95a, 
               32'shc9b1be1e, 32'shc9b292eb, 32'shc9b367c1, 32'shc9b43c9f, 32'shc9b51185, 32'shc9b5e674, 32'shc9b6bb6b, 32'shc9b7906a, 
               32'shc9b86572, 32'shc9b93a82, 32'shc9ba0f9b, 32'shc9bae4bc, 32'shc9bbb9e5, 32'shc9bc8f16, 32'shc9bd6450, 32'shc9be3993, 
               32'shc9bf0edd, 32'shc9bfe430, 32'shc9c0b98c, 32'shc9c18ef0, 32'shc9c2645c, 32'shc9c339d0, 32'shc9c40f4d, 32'shc9c4e4d3, 
               32'shc9c5ba60, 32'shc9c68ff6, 32'shc9c76595, 32'shc9c83b3b, 32'shc9c910ea, 32'shc9c9e6a2, 32'shc9cabc62, 32'shc9cb922a, 
               32'shc9cc67fa, 32'shc9cd3dd3, 32'shc9ce13b4, 32'shc9cee99e, 32'shc9cfbf90, 32'shc9d0958a, 32'shc9d16b8d, 32'shc9d24198, 
               32'shc9d317ab, 32'shc9d3edc7, 32'shc9d4c3eb, 32'shc9d59a18, 32'shc9d6704c, 32'shc9d7468a, 32'shc9d81ccf, 32'shc9d8f31d, 
               32'shc9d9c973, 32'shc9da9fd2, 32'shc9db7639, 32'shc9dc4ca8, 32'shc9dd231f, 32'shc9ddf99f, 32'shc9ded028, 32'shc9dfa6b8, 
               32'shc9e07d51, 32'shc9e153f3, 32'shc9e22a9c, 32'shc9e3014e, 32'shc9e3d809, 32'shc9e4aecb, 32'shc9e58596, 32'shc9e65c6a, 
               32'shc9e73346, 32'shc9e80a2a, 32'shc9e8e116, 32'shc9e9b80b, 32'shc9ea8f08, 32'shc9eb660d, 32'shc9ec3d1b, 32'shc9ed1431, 
               32'shc9edeb50, 32'shc9eec277, 32'shc9ef99a6, 32'shc9f070dd, 32'shc9f1481d, 32'shc9f21f65, 32'shc9f2f6b6, 32'shc9f3ce0f, 
               32'shc9f4a570, 32'shc9f57cd9, 32'shc9f6544b, 32'shc9f72bc5, 32'shc9f80348, 32'shc9f8dad3, 32'shc9f9b266, 32'shc9fa8a01, 
               32'shc9fb61a5, 32'shc9fc3951, 32'shc9fd1106, 32'shc9fde8c2, 32'shc9fec088, 32'shc9ff9855, 32'shca00702b, 32'shca014809, 
               32'shca021fef, 32'shca02f7de, 32'shca03cfd5, 32'shca04a7d5, 32'shca057fdd, 32'shca0657ed, 32'shca073005, 32'shca080826, 
               32'shca08e04f, 32'shca09b880, 32'shca0a90ba, 32'shca0b68fc, 32'shca0c4146, 32'shca0d1999, 32'shca0df1f4, 32'shca0eca57, 
               32'shca0fa2c3, 32'shca107b37, 32'shca1153b3, 32'shca122c37, 32'shca1304c4, 32'shca13dd59, 32'shca14b5f7, 32'shca158e9d, 
               32'shca16674b, 32'shca174001, 32'shca1818c0, 32'shca18f187, 32'shca19ca57, 32'shca1aa32e, 32'shca1b7c0e, 32'shca1c54f7, 
               32'shca1d2de7, 32'shca1e06e0, 32'shca1edfe2, 32'shca1fb8eb, 32'shca2091fd, 32'shca216b17, 32'shca22443a, 32'shca231d64, 
               32'shca23f698, 32'shca24cfd3, 32'shca25a917, 32'shca268263, 32'shca275bb7, 32'shca283514, 32'shca290e79, 32'shca29e7e6, 
               32'shca2ac15b, 32'shca2b9ad9, 32'shca2c745f, 32'shca2d4dee, 32'shca2e2784, 32'shca2f0123, 32'shca2fdacb, 32'shca30b47a, 
               32'shca318e32, 32'shca3267f3, 32'shca3341bb, 32'shca341b8c, 32'shca34f565, 32'shca35cf47, 32'shca36a930, 32'shca378322, 
               32'shca385d1d, 32'shca39371f, 32'shca3a112a, 32'shca3aeb3d, 32'shca3bc559, 32'shca3c9f7c, 32'shca3d79a8, 32'shca3e53dd, 
               32'shca3f2e19, 32'shca40085e, 32'shca40e2ac, 32'shca41bd01, 32'shca42975f, 32'shca4371c5, 32'shca444c33, 32'shca4526aa, 
               32'shca460129, 32'shca46dbb0, 32'shca47b640, 32'shca4890d7, 32'shca496b77, 32'shca4a4620, 32'shca4b20d0, 32'shca4bfb89, 
               32'shca4cd64b, 32'shca4db114, 32'shca4e8be6, 32'shca4f66c0, 32'shca5041a2, 32'shca511c8d, 32'shca51f780, 32'shca52d27b, 
               32'shca53ad7e, 32'shca54888a, 32'shca55639e, 32'shca563eba, 32'shca5719df, 32'shca57f50c, 32'shca58d041, 32'shca59ab7e, 
               32'shca5a86c4, 32'shca5b6212, 32'shca5c3d68, 32'shca5d18c6, 32'shca5df42d, 32'shca5ecf9c, 32'shca5fab13, 32'shca608693, 
               32'shca61621b, 32'shca623dab, 32'shca631943, 32'shca63f4e4, 32'shca64d08d, 32'shca65ac3e, 32'shca6687f7, 32'shca6763b9, 
               32'shca683f83, 32'shca691b55, 32'shca69f72f, 32'shca6ad312, 32'shca6baefd, 32'shca6c8af0, 32'shca6d66ec, 32'shca6e42f0, 
               32'shca6f1efc, 32'shca6ffb10, 32'shca70d72d, 32'shca71b351, 32'shca728f7f, 32'shca736bb4, 32'shca7447f2, 32'shca752437, 
               32'shca760086, 32'shca76dcdc, 32'shca77b93b, 32'shca7895a1, 32'shca797211, 32'shca7a4e88, 32'shca7b2b08, 32'shca7c078f, 
               32'shca7ce420, 32'shca7dc0b8, 32'shca7e9d59, 32'shca7f7a02, 32'shca8056b3, 32'shca81336c, 32'shca82102e, 32'shca82ecf8, 
               32'shca83c9ca, 32'shca84a6a4, 32'shca858387, 32'shca866072, 32'shca873d65, 32'shca881a60, 32'shca88f764, 32'shca89d470, 
               32'shca8ab184, 32'shca8b8ea0, 32'shca8c6bc5, 32'shca8d48f2, 32'shca8e2627, 32'shca8f0364, 32'shca8fe0aa, 32'shca90bdf8, 
               32'shca919b4e, 32'shca9278ac, 32'shca935613, 32'shca943381, 32'shca9510f8, 32'shca95ee78, 32'shca96cbff, 32'shca97a98f, 
               32'shca988727, 32'shca9964c7, 32'shca9a4270, 32'shca9b2020, 32'shca9bfdd9, 32'shca9cdb9a, 32'shca9db964, 32'shca9e9735, 
               32'shca9f750f, 32'shcaa052f1, 32'shcaa130db, 32'shcaa20ece, 32'shcaa2ecc9, 32'shcaa3cacc, 32'shcaa4a8d7, 32'shcaa586ea, 
               32'shcaa66506, 32'shcaa7432a, 32'shcaa82156, 32'shcaa8ff8a, 32'shcaa9ddc7, 32'shcaaabc0c, 32'shcaab9a59, 32'shcaac78ae, 
               32'shcaad570c, 32'shcaae3571, 32'shcaaf13df, 32'shcaaff255, 32'shcab0d0d4, 32'shcab1af5a, 32'shcab28de9, 32'shcab36c80, 
               32'shcab44b1f, 32'shcab529c7, 32'shcab60877, 32'shcab6e72f, 32'shcab7c5ef, 32'shcab8a4b7, 32'shcab98388, 32'shcaba6260, 
               32'shcabb4141, 32'shcabc202a, 32'shcabcff1c, 32'shcabdde16, 32'shcabebd17, 32'shcabf9c21, 32'shcac07b34, 32'shcac15a4e, 
               32'shcac23971, 32'shcac3189c, 32'shcac3f7cf, 32'shcac4d70a, 32'shcac5b64e, 32'shcac69599, 32'shcac774ed, 32'shcac8544a, 
               32'shcac933ae, 32'shcaca131a, 32'shcacaf28f, 32'shcacbd20c, 32'shcaccb191, 32'shcacd911f, 32'shcace70b4, 32'shcacf5052, 
               32'shcad02ff8, 32'shcad10fa6, 32'shcad1ef5d, 32'shcad2cf1b, 32'shcad3aee2, 32'shcad48eb1, 32'shcad56e88, 32'shcad64e68, 
               32'shcad72e4f, 32'shcad80e3f, 32'shcad8ee37, 32'shcad9ce37, 32'shcadaae40, 32'shcadb8e50, 32'shcadc6e69, 32'shcadd4e8a, 
               32'shcade2eb3, 32'shcadf0ee4, 32'shcadfef1e, 32'shcae0cf60, 32'shcae1afaa, 32'shcae28ffc, 32'shcae37056, 32'shcae450b9, 
               32'shcae53123, 32'shcae61196, 32'shcae6f211, 32'shcae7d295, 32'shcae8b320, 32'shcae993b4, 32'shcaea744f, 32'shcaeb54f3, 
               32'shcaec35a0, 32'shcaed1654, 32'shcaedf711, 32'shcaeed7d5, 32'shcaefb8a2, 32'shcaf09977, 32'shcaf17a55, 32'shcaf25b3a, 
               32'shcaf33c28, 32'shcaf41d1e, 32'shcaf4fe1c, 32'shcaf5df22, 32'shcaf6c030, 32'shcaf7a147, 32'shcaf88266, 32'shcaf9638d, 
               32'shcafa44bc, 32'shcafb25f3, 32'shcafc0732, 32'shcafce87a, 32'shcafdc9ca, 32'shcafeab22, 32'shcaff8c82, 32'shcb006dea, 
               32'shcb014f5b, 32'shcb0230d3, 32'shcb031254, 32'shcb03f3dd, 32'shcb04d56e, 32'shcb05b708, 32'shcb0698a9, 32'shcb077a53, 
               32'shcb085c05, 32'shcb093dbf, 32'shcb0a1f81, 32'shcb0b014b, 32'shcb0be31e, 32'shcb0cc4f9, 32'shcb0da6dc, 32'shcb0e88c7, 
               32'shcb0f6aba, 32'shcb104cb5, 32'shcb112eb9, 32'shcb1210c4, 32'shcb12f2d8, 32'shcb13d4f4, 32'shcb14b718, 32'shcb159945, 
               32'shcb167b79, 32'shcb175db6, 32'shcb183ffb, 32'shcb192248, 32'shcb1a049d, 32'shcb1ae6fa, 32'shcb1bc95f, 32'shcb1cabcd, 
               32'shcb1d8e43, 32'shcb1e70c1, 32'shcb1f5347, 32'shcb2035d5, 32'shcb21186b, 32'shcb21fb0a, 32'shcb22ddb1, 32'shcb23c05f, 
               32'shcb24a316, 32'shcb2585d5, 32'shcb26689d, 32'shcb274b6c, 32'shcb282e44, 32'shcb291123, 32'shcb29f40b, 32'shcb2ad6fb, 
               32'shcb2bb9f4, 32'shcb2c9cf4, 32'shcb2d7ffc, 32'shcb2e630d, 32'shcb2f4626, 32'shcb302947, 32'shcb310c70, 32'shcb31efa1, 
               32'shcb32d2da, 32'shcb33b61c, 32'shcb349965, 32'shcb357cb7, 32'shcb366011, 32'shcb374373, 32'shcb3826dd, 32'shcb390a50, 
               32'shcb39edca, 32'shcb3ad14d, 32'shcb3bb4d7, 32'shcb3c986a, 32'shcb3d7c05, 32'shcb3e5fa8, 32'shcb3f4354, 32'shcb402707, 
               32'shcb410ac3, 32'shcb41ee86, 32'shcb42d252, 32'shcb43b626, 32'shcb449a02, 32'shcb457de6, 32'shcb4661d3, 32'shcb4745c7, 
               32'shcb4829c4, 32'shcb490dc9, 32'shcb49f1d5, 32'shcb4ad5ea, 32'shcb4bba08, 32'shcb4c9e2d, 32'shcb4d825a, 32'shcb4e6690, 
               32'shcb4f4acd, 32'shcb502f13, 32'shcb511361, 32'shcb51f7b7, 32'shcb52dc15, 32'shcb53c07b, 32'shcb54a4ea, 32'shcb558960, 
               32'shcb566ddf, 32'shcb575266, 32'shcb5836f4, 32'shcb591b8b, 32'shcb5a002b, 32'shcb5ae4d2, 32'shcb5bc981, 32'shcb5cae39, 
               32'shcb5d92f8, 32'shcb5e77c0, 32'shcb5f5c90, 32'shcb604168, 32'shcb612648, 32'shcb620b30, 32'shcb62f020, 32'shcb63d518, 
               32'shcb64ba19, 32'shcb659f22, 32'shcb668432, 32'shcb67694b, 32'shcb684e6c, 32'shcb693395, 32'shcb6a18c6, 32'shcb6afe00, 
               32'shcb6be341, 32'shcb6cc88a, 32'shcb6daddc, 32'shcb6e9336, 32'shcb6f7898, 32'shcb705e01, 32'shcb714373, 32'shcb7228ee, 
               32'shcb730e70, 32'shcb73f3fa, 32'shcb74d98d, 32'shcb75bf27, 32'shcb76a4ca, 32'shcb778a75, 32'shcb787027, 32'shcb7955e2, 
               32'shcb7a3ba5, 32'shcb7b2171, 32'shcb7c0744, 32'shcb7ced1f, 32'shcb7dd303, 32'shcb7eb8ee, 32'shcb7f9ee2, 32'shcb8084de, 
               32'shcb816ae1, 32'shcb8250ed, 32'shcb833701, 32'shcb841d1d, 32'shcb850342, 32'shcb85e96e, 32'shcb86cfa2, 32'shcb87b5df, 
               32'shcb889c23, 32'shcb898270, 32'shcb8a68c5, 32'shcb8b4f22, 32'shcb8c3587, 32'shcb8d1bf4, 32'shcb8e0269, 32'shcb8ee8e6, 
               32'shcb8fcf6b, 32'shcb90b5f9, 32'shcb919c8e, 32'shcb92832c, 32'shcb9369d1, 32'shcb94507f, 32'shcb953735, 32'shcb961df3, 
               32'shcb9704b9, 32'shcb97eb87, 32'shcb98d25d, 32'shcb99b93b, 32'shcb9aa021, 32'shcb9b8710, 32'shcb9c6e06, 32'shcb9d5505, 
               32'shcb9e3c0b, 32'shcb9f231a, 32'shcba00a31, 32'shcba0f150, 32'shcba1d877, 32'shcba2bfa6, 32'shcba3a6dd, 32'shcba48e1c, 
               32'shcba57563, 32'shcba65cb2, 32'shcba7440a, 32'shcba82b69, 32'shcba912d1, 32'shcba9fa40, 32'shcbaae1b8, 32'shcbabc938, 
               32'shcbacb0bf, 32'shcbad984f, 32'shcbae7fe7, 32'shcbaf6787, 32'shcbb04f2f, 32'shcbb136df, 32'shcbb21e98, 32'shcbb30658, 
               32'shcbb3ee20, 32'shcbb4d5f1, 32'shcbb5bdc9, 32'shcbb6a5aa, 32'shcbb78d92, 32'shcbb87583, 32'shcbb95d7c, 32'shcbba457c, 
               32'shcbbb2d85, 32'shcbbc1596, 32'shcbbcfdaf, 32'shcbbde5d0, 32'shcbbecdf9, 32'shcbbfb62a, 32'shcbc09e64, 32'shcbc186a5, 
               32'shcbc26eee, 32'shcbc3573f, 32'shcbc43f99, 32'shcbc527fa, 32'shcbc61064, 32'shcbc6f8d5, 32'shcbc7e14f, 32'shcbc8c9d1, 
               32'shcbc9b25a, 32'shcbca9aec, 32'shcbcb8386, 32'shcbcc6c28, 32'shcbcd54d2, 32'shcbce3d84, 32'shcbcf263e, 32'shcbd00f00, 
               32'shcbd0f7ca, 32'shcbd1e09c, 32'shcbd2c977, 32'shcbd3b259, 32'shcbd49b43, 32'shcbd58436, 32'shcbd66d30, 32'shcbd75633, 
               32'shcbd83f3d, 32'shcbd92850, 32'shcbda116a, 32'shcbdafa8d, 32'shcbdbe3b7, 32'shcbdcccea, 32'shcbddb625, 32'shcbde9f68, 
               32'shcbdf88b3, 32'shcbe07205, 32'shcbe15b60, 32'shcbe244c3, 32'shcbe32e2e, 32'shcbe417a1, 32'shcbe5011c, 32'shcbe5ea9f, 
               32'shcbe6d42b, 32'shcbe7bdbe, 32'shcbe8a759, 32'shcbe990fc, 32'shcbea7aa7, 32'shcbeb645b, 32'shcbec4e16, 32'shcbed37d9, 
               32'shcbee21a5, 32'shcbef0b78, 32'shcbeff554, 32'shcbf0df37, 32'shcbf1c923, 32'shcbf2b316, 32'shcbf39d12, 32'shcbf48715, 
               32'shcbf57121, 32'shcbf65b34, 32'shcbf74550, 32'shcbf82f74, 32'shcbf919a0, 32'shcbfa03d3, 32'shcbfaee0f, 32'shcbfbd853, 
               32'shcbfcc29f, 32'shcbfdacf2, 32'shcbfe974e, 32'shcbff81b2, 32'shcc006c1e, 32'shcc015692, 32'shcc02410e, 32'shcc032b92, 
               32'shcc04161e, 32'shcc0500b2, 32'shcc05eb4e, 32'shcc06d5f2, 32'shcc07c09e, 32'shcc08ab52, 32'shcc09960e, 32'shcc0a80d2, 
               32'shcc0b6b9e, 32'shcc0c5672, 32'shcc0d414e, 32'shcc0e2c32, 32'shcc0f171e, 32'shcc100212, 32'shcc10ed0e, 32'shcc11d813, 
               32'shcc12c31f, 32'shcc13ae33, 32'shcc14994f, 32'shcc158473, 32'shcc166f9f, 32'shcc175ad3, 32'shcc184610, 32'shcc193154, 
               32'shcc1a1ca0, 32'shcc1b07f4, 32'shcc1bf350, 32'shcc1cdeb5, 32'shcc1dca21, 32'shcc1eb595, 32'shcc1fa111, 32'shcc208c95, 
               32'shcc217822, 32'shcc2263b6, 32'shcc234f52, 32'shcc243af6, 32'shcc2526a2, 32'shcc261257, 32'shcc26fe13, 32'shcc27e9d7, 
               32'shcc28d5a3, 32'shcc29c177, 32'shcc2aad54, 32'shcc2b9938, 32'shcc2c8524, 32'shcc2d7118, 32'shcc2e5d14, 32'shcc2f4918, 
               32'shcc303524, 32'shcc312139, 32'shcc320d55, 32'shcc32f979, 32'shcc33e5a5, 32'shcc34d1d9, 32'shcc35be15, 32'shcc36aa59, 
               32'shcc3796a5, 32'shcc3882f9, 32'shcc396f55, 32'shcc3a5bb9, 32'shcc3b4825, 32'shcc3c3499, 32'shcc3d2115, 32'shcc3e0d99, 
               32'shcc3efa25, 32'shcc3fe6b8, 32'shcc40d354, 32'shcc41bff8, 32'shcc42aca4, 32'shcc439958, 32'shcc448614, 32'shcc4572d7, 
               32'shcc465fa3, 32'shcc474c77, 32'shcc483952, 32'shcc492636, 32'shcc4a1322, 32'shcc4b0015, 32'shcc4bed11, 32'shcc4cda14, 
               32'shcc4dc720, 32'shcc4eb433, 32'shcc4fa14f, 32'shcc508e72, 32'shcc517b9e, 32'shcc5268d1, 32'shcc53560c, 32'shcc544350, 
               32'shcc55309b, 32'shcc561dee, 32'shcc570b4a, 32'shcc57f8ad, 32'shcc58e618, 32'shcc59d38b, 32'shcc5ac106, 32'shcc5bae89, 
               32'shcc5c9c14, 32'shcc5d89a7, 32'shcc5e7742, 32'shcc5f64e5, 32'shcc605290, 32'shcc614043, 32'shcc622dfd, 32'shcc631bc0, 
               32'shcc64098b, 32'shcc64f75e, 32'shcc65e538, 32'shcc66d31b, 32'shcc67c105, 32'shcc68aef8, 32'shcc699cf2, 32'shcc6a8af5, 
               32'shcc6b78ff, 32'shcc6c6711, 32'shcc6d552c, 32'shcc6e434e, 32'shcc6f3178, 32'shcc701faa, 32'shcc710de4, 32'shcc71fc26, 
               32'shcc72ea70, 32'shcc73d8c2, 32'shcc74c71c, 32'shcc75b57e, 32'shcc76a3e8, 32'shcc779259, 32'shcc7880d3, 32'shcc796f55, 
               32'shcc7a5dde, 32'shcc7b4c70, 32'shcc7c3b09, 32'shcc7d29aa, 32'shcc7e1854, 32'shcc7f0705, 32'shcc7ff5be, 32'shcc80e47f, 
               32'shcc81d349, 32'shcc82c21a, 32'shcc83b0f3, 32'shcc849fd4, 32'shcc858ebc, 32'shcc867dad, 32'shcc876ca6, 32'shcc885ba7, 
               32'shcc894aaf, 32'shcc8a39c0, 32'shcc8b28d8, 32'shcc8c17f9, 32'shcc8d0721, 32'shcc8df651, 32'shcc8ee58a, 32'shcc8fd4ca, 
               32'shcc90c412, 32'shcc91b362, 32'shcc92a2ba, 32'shcc93921a, 32'shcc948182, 32'shcc9570f1, 32'shcc966069, 32'shcc974fe9, 
               32'shcc983f70, 32'shcc992f00, 32'shcc9a1e97, 32'shcc9b0e36, 32'shcc9bfddd, 32'shcc9ced8d, 32'shcc9ddd44, 32'shcc9ecd03, 
               32'shcc9fbcca, 32'shcca0ac99, 32'shcca19c6f, 32'shcca28c4e, 32'shcca37c35, 32'shcca46c23, 32'shcca55c1a, 32'shcca64c18, 
               32'shcca73c1e, 32'shcca82c2d, 32'shcca91c43, 32'shccaa0c61, 32'shccaafc87, 32'shccabecb5, 32'shccacdcea, 32'shccadcd28, 
               32'shccaebd6e, 32'shccafadbb, 32'shccb09e11, 32'shccb18e6e, 32'shccb27ed3, 32'shccb36f41, 32'shccb45fb6, 32'shccb55033, 
               32'shccb640b8, 32'shccb73144, 32'shccb821d9, 32'shccb91276, 32'shccba031a, 32'shccbaf3c7, 32'shccbbe47b, 32'shccbcd538, 
               32'shccbdc5fc, 32'shccbeb6c8, 32'shccbfa79c, 32'shccc09878, 32'shccc1895c, 32'shccc27a47, 32'shccc36b3b, 32'shccc45c36, 
               32'shccc54d3a, 32'shccc63e45, 32'shccc72f58, 32'shccc82073, 32'shccc91196, 32'shccca02c1, 32'shcccaf3f4, 32'shcccbe52f, 
               32'shccccd671, 32'shcccdc7bc, 32'shccceb90e, 32'shcccfaa69, 32'shccd09bcb, 32'shccd18d35, 32'shccd27ea7, 32'shccd37021, 
               32'shccd461a2, 32'shccd5532c, 32'shccd644bd, 32'shccd73657, 32'shccd827f8, 32'shccd919a1, 32'shccda0b52, 32'shccdafd0b, 
               32'shccdbeecc, 32'shccdce095, 32'shccddd266, 32'shccdec43e, 32'shccdfb61f, 32'shcce0a807, 32'shcce199f7, 32'shcce28bef, 
               32'shcce37def, 32'shcce46ff7, 32'shcce56206, 32'shcce6541e, 32'shcce7463e, 32'shcce83865, 32'shcce92a94, 32'shccea1ccb, 
               32'shcceb0f0a, 32'shccec0151, 32'shccecf3a0, 32'shccede5f6, 32'shcceed855, 32'shccefcabb, 32'shccf0bd29, 32'shccf1af9f, 
               32'shccf2a21d, 32'shccf394a3, 32'shccf48731, 32'shccf579c7, 32'shccf66c64, 32'shccf75f09, 32'shccf851b7, 32'shccf9446c, 
               32'shccfa3729, 32'shccfb29ed, 32'shccfc1cba, 32'shccfd0f8f, 32'shccfe026b, 32'shccfef54f, 32'shccffe83c, 32'shcd00db30, 
               32'shcd01ce2b, 32'shcd02c12f, 32'shcd03b43b, 32'shcd04a74e, 32'shcd059a6a, 32'shcd068d8d, 32'shcd0780b8, 32'shcd0873eb, 
               32'shcd096725, 32'shcd0a5a68, 32'shcd0b4db3, 32'shcd0c4105, 32'shcd0d345f, 32'shcd0e27c1, 32'shcd0f1b2b, 32'shcd100e9d, 
               32'shcd110216, 32'shcd11f598, 32'shcd12e921, 32'shcd13dcb2, 32'shcd14d04b, 32'shcd15c3ec, 32'shcd16b795, 32'shcd17ab46, 
               32'shcd189efe, 32'shcd1992be, 32'shcd1a8687, 32'shcd1b7a57, 32'shcd1c6e2e, 32'shcd1d620e, 32'shcd1e55f6, 32'shcd1f49e5, 
               32'shcd203ddc, 32'shcd2131db, 32'shcd2225e2, 32'shcd2319f1, 32'shcd240e08, 32'shcd250226, 32'shcd25f64c, 32'shcd26ea7b, 
               32'shcd27deb0, 32'shcd28d2ee, 32'shcd29c734, 32'shcd2abb81, 32'shcd2bafd7, 32'shcd2ca434, 32'shcd2d9899, 32'shcd2e8d06, 
               32'shcd2f817b, 32'shcd3075f7, 32'shcd316a7b, 32'shcd325f08, 32'shcd33539c, 32'shcd344837, 32'shcd353cdb, 32'shcd363187, 
               32'shcd37263a, 32'shcd381af5, 32'shcd390fb8, 32'shcd3a0483, 32'shcd3af956, 32'shcd3bee30, 32'shcd3ce313, 32'shcd3dd7fd, 
               32'shcd3eccef, 32'shcd3fc1e9, 32'shcd40b6ea, 32'shcd41abf4, 32'shcd42a105, 32'shcd43961e, 32'shcd448b3f, 32'shcd458068, 
               32'shcd467599, 32'shcd476ad1, 32'shcd486011, 32'shcd495559, 32'shcd4a4aa9, 32'shcd4b4001, 32'shcd4c3560, 32'shcd4d2ac8, 
               32'shcd4e2037, 32'shcd4f15ae, 32'shcd500b2d, 32'shcd5100b3, 32'shcd51f642, 32'shcd52ebd8, 32'shcd53e176, 32'shcd54d71c, 
               32'shcd55ccca, 32'shcd56c27f, 32'shcd57b83c, 32'shcd58ae01, 32'shcd59a3ce, 32'shcd5a99a3, 32'shcd5b8f80, 32'shcd5c8564, 
               32'shcd5d7b50, 32'shcd5e7144, 32'shcd5f6740, 32'shcd605d44, 32'shcd61534f, 32'shcd624962, 32'shcd633f7d, 32'shcd6435a0, 
               32'shcd652bcb, 32'shcd6621fd, 32'shcd671837, 32'shcd680e79, 32'shcd6904c3, 32'shcd69fb15, 32'shcd6af16e, 32'shcd6be7d0, 
               32'shcd6cde39, 32'shcd6dd4a9, 32'shcd6ecb22, 32'shcd6fc1a3, 32'shcd70b82b, 32'shcd71aebb, 32'shcd72a553, 32'shcd739bf2, 
               32'shcd74929a, 32'shcd758949, 32'shcd768000, 32'shcd7776bf, 32'shcd786d85, 32'shcd796454, 32'shcd7a5b2a, 32'shcd7b5208, 
               32'shcd7c48ee, 32'shcd7d3fdb, 32'shcd7e36d1, 32'shcd7f2dce, 32'shcd8024d3, 32'shcd811bdf, 32'shcd8212f4, 32'shcd830a10, 
               32'shcd840134, 32'shcd84f860, 32'shcd85ef94, 32'shcd86e6cf, 32'shcd87de12, 32'shcd88d55d, 32'shcd89ccb0, 32'shcd8ac40b, 
               32'shcd8bbb6d, 32'shcd8cb2d7, 32'shcd8daa49, 32'shcd8ea1c3, 32'shcd8f9944, 32'shcd9090cd, 32'shcd91885e, 32'shcd927ff7, 
               32'shcd937798, 32'shcd946f40, 32'shcd9566f0, 32'shcd965ea8, 32'shcd975668, 32'shcd984e2f, 32'shcd9945fe, 32'shcd9a3dd5, 
               32'shcd9b35b4, 32'shcd9c2d9a, 32'shcd9d2589, 32'shcd9e1d7f, 32'shcd9f157d, 32'shcda00d82, 32'shcda10590, 32'shcda1fda5, 
               32'shcda2f5c2, 32'shcda3ede6, 32'shcda4e613, 32'shcda5de47, 32'shcda6d683, 32'shcda7cec7, 32'shcda8c712, 32'shcda9bf65, 
               32'shcdaab7c0, 32'shcdabb023, 32'shcdaca88e, 32'shcdada100, 32'shcdae997a, 32'shcdaf91fc, 32'shcdb08a86, 32'shcdb18317, 
               32'shcdb27bb0, 32'shcdb37451, 32'shcdb46cfa, 32'shcdb565aa, 32'shcdb65e62, 32'shcdb75722, 32'shcdb84fea, 32'shcdb948b9, 
               32'shcdba4190, 32'shcdbb3a6f, 32'shcdbc3356, 32'shcdbd2c44, 32'shcdbe253a, 32'shcdbf1e38, 32'shcdc0173e, 32'shcdc1104b, 
               32'shcdc20960, 32'shcdc3027d, 32'shcdc3fba2, 32'shcdc4f4ce, 32'shcdc5ee02, 32'shcdc6e73e, 32'shcdc7e082, 32'shcdc8d9cd, 
               32'shcdc9d320, 32'shcdcacc7b, 32'shcdcbc5de, 32'shcdccbf48, 32'shcdcdb8ba, 32'shcdceb234, 32'shcdcfabb6, 32'shcdd0a53f, 
               32'shcdd19ed0, 32'shcdd29869, 32'shcdd39209, 32'shcdd48bb2, 32'shcdd58562, 32'shcdd67f19, 32'shcdd778d9, 32'shcdd872a0, 
               32'shcdd96c6f, 32'shcdda6646, 32'shcddb6024, 32'shcddc5a0a, 32'shcddd53f8, 32'shcdde4dee, 32'shcddf47eb, 32'shcde041f0, 
               32'shcde13bfd, 32'shcde23611, 32'shcde3302e, 32'shcde42a52, 32'shcde5247d, 32'shcde61eb1, 32'shcde718ec, 32'shcde8132f, 
               32'shcde90d79, 32'shcdea07cc, 32'shcdeb0226, 32'shcdebfc87, 32'shcdecf6f1, 32'shcdedf162, 32'shcdeeebdb, 32'shcdefe65c, 
               32'shcdf0e0e4, 32'shcdf1db74, 32'shcdf2d60c, 32'shcdf3d0ac, 32'shcdf4cb53, 32'shcdf5c602, 32'shcdf6c0b9, 32'shcdf7bb77, 
               32'shcdf8b63d, 32'shcdf9b10b, 32'shcdfaabe1, 32'shcdfba6be, 32'shcdfca1a3, 32'shcdfd9c90, 32'shcdfe9784, 32'shcdff9280, 
               32'shce008d84, 32'shce01888f, 32'shce0283a3, 32'shce037ebe, 32'shce0479e0, 32'shce05750b, 32'shce06703d, 32'shce076b77, 
               32'shce0866b8, 32'shce096201, 32'shce0a5d52, 32'shce0b58ab, 32'shce0c540b, 32'shce0d4f73, 32'shce0e4ae3, 32'shce0f465a, 
               32'shce1041d9, 32'shce113d60, 32'shce1238ef, 32'shce133485, 32'shce143023, 32'shce152bc9, 32'shce162776, 32'shce17232b, 
               32'shce181ee8, 32'shce191aac, 32'shce1a1678, 32'shce1b124c, 32'shce1c0e28, 32'shce1d0a0b, 32'shce1e05f6, 32'shce1f01e8, 
               32'shce1ffde2, 32'shce20f9e4, 32'shce21f5ee, 32'shce22f1ff, 32'shce23ee18, 32'shce24ea39, 32'shce25e662, 32'shce26e292, 
               32'shce27dec9, 32'shce28db09, 32'shce29d750, 32'shce2ad39f, 32'shce2bcff5, 32'shce2ccc54, 32'shce2dc8ba, 32'shce2ec527, 
               32'shce2fc19c, 32'shce30be19, 32'shce31ba9e, 32'shce32b72a, 32'shce33b3be, 32'shce34b05a, 32'shce35acfd, 32'shce36a9a8, 
               32'shce37a65b, 32'shce38a315, 32'shce399fd7, 32'shce3a9ca1, 32'shce3b9973, 32'shce3c964c, 32'shce3d932c, 32'shce3e9015, 
               32'shce3f8d05, 32'shce4089fd, 32'shce4186fc, 32'shce428403, 32'shce438112, 32'shce447e28, 32'shce457b47, 32'shce46786c, 
               32'shce47759a, 32'shce4872cf, 32'shce49700c, 32'shce4a6d50, 32'shce4b6a9c, 32'shce4c67f0, 32'shce4d654c, 32'shce4e62af, 
               32'shce4f6019, 32'shce505d8c, 32'shce515b06, 32'shce525888, 32'shce535611, 32'shce5453a2, 32'shce55513b, 32'shce564edc, 
               32'shce574c84, 32'shce584a33, 32'shce5947eb, 32'shce5a45aa, 32'shce5b4370, 32'shce5c413f, 32'shce5d3f15, 32'shce5e3cf2, 
               32'shce5f3ad8, 32'shce6038c5, 32'shce6136b9, 32'shce6234b6, 32'shce6332ba, 32'shce6430c5, 32'shce652ed8, 32'shce662cf3, 
               32'shce672b16, 32'shce682940, 32'shce692772, 32'shce6a25ab, 32'shce6b23ec, 32'shce6c2235, 32'shce6d2086, 32'shce6e1ede, 
               32'shce6f1d3d, 32'shce701ba5, 32'shce711a14, 32'shce72188a, 32'shce731709, 32'shce74158e, 32'shce75141c, 32'shce7612b1, 
               32'shce77114e, 32'shce780ff3, 32'shce790e9f, 32'shce7a0d52, 32'shce7b0c0e, 32'shce7c0ad1, 32'shce7d099b, 32'shce7e086e, 
               32'shce7f0748, 32'shce800629, 32'shce810512, 32'shce820403, 32'shce8302fc, 32'shce8401fc, 32'shce850104, 32'shce860013, 
               32'shce86ff2a, 32'shce87fe48, 32'shce88fd6f, 32'shce89fc9d, 32'shce8afbd2, 32'shce8bfb0f, 32'shce8cfa54, 32'shce8df9a0, 
               32'shce8ef8f4, 32'shce8ff850, 32'shce90f7b3, 32'shce91f71e, 32'shce92f691, 32'shce93f60b, 32'shce94f58c, 32'shce95f516, 
               32'shce96f4a7, 32'shce97f43f, 32'shce98f3e0, 32'shce99f387, 32'shce9af337, 32'shce9bf2ee, 32'shce9cf2ad, 32'shce9df273, 
               32'shce9ef241, 32'shce9ff216, 32'shcea0f1f4, 32'shcea1f1d8, 32'shcea2f1c5, 32'shcea3f1b9, 32'shcea4f1b4, 32'shcea5f1b7, 
               32'shcea6f1c2, 32'shcea7f1d5, 32'shcea8f1ef, 32'shcea9f210, 32'shceaaf23a, 32'shceabf26b, 32'shceacf2a3, 32'shceadf2e3, 
               32'shceaef32b, 32'shceaff37a, 32'shceb0f3d1, 32'shceb1f42f, 32'shceb2f496, 32'shceb3f503, 32'shceb4f579, 32'shceb5f5f5, 
               32'shceb6f67a, 32'shceb7f706, 32'shceb8f79a, 32'shceb9f835, 32'shcebaf8d8, 32'shcebbf983, 32'shcebcfa35, 32'shcebdfaee, 
               32'shcebefbb0, 32'shcebffc79, 32'shcec0fd49, 32'shcec1fe21, 32'shcec2ff01, 32'shcec3ffe8, 32'shcec500d7, 32'shcec601cd, 
               32'shcec702cb, 32'shcec803d1, 32'shcec904de, 32'shceca05f3, 32'shcecb070f, 32'shcecc0833, 32'shcecd095f, 32'shcece0a92, 
               32'shcecf0bcd, 32'shced00d0f, 32'shced10e59, 32'shced20fab, 32'shced31104, 32'shced41265, 32'shced513cd, 32'shced6153d, 
               32'shced716b4, 32'shced81833, 32'shced919ba, 32'shceda1b48, 32'shcedb1cde, 32'shcedc1e7b, 32'shcedd2020, 32'shcede21cc, 
               32'shcedf2380, 32'shcee0253c, 32'shcee126ff, 32'shcee228ca, 32'shcee32a9c, 32'shcee42c76, 32'shcee52e58, 32'shcee63041, 
               32'shcee73231, 32'shcee8342a, 32'shcee93629, 32'shceea3831, 32'shceeb3a40, 32'shceec3c56, 32'shceed3e74, 32'shceee409a, 
               32'shceef42c7, 32'shcef044fc, 32'shcef14738, 32'shcef2497c, 32'shcef34bc8, 32'shcef44e1b, 32'shcef55075, 32'shcef652d7, 
               32'shcef75541, 32'shcef857b2, 32'shcef95a2b, 32'shcefa5cac, 32'shcefb5f34, 32'shcefc61c3, 32'shcefd645a, 32'shcefe66f9, 
               32'shceff699f, 32'shcf006c4d, 32'shcf016f02, 32'shcf0271bf, 32'shcf037483, 32'shcf04774f, 32'shcf057a23, 32'shcf067cfe, 
               32'shcf077fe1, 32'shcf0882cb, 32'shcf0985bc, 32'shcf0a88b6, 32'shcf0b8bb7, 32'shcf0c8ebf, 32'shcf0d91cf, 32'shcf0e94e6, 
               32'shcf0f9805, 32'shcf109b2c, 32'shcf119e5a, 32'shcf12a190, 32'shcf13a4cd, 32'shcf14a812, 32'shcf15ab5e, 32'shcf16aeb2, 
               32'shcf17b20d, 32'shcf18b570, 32'shcf19b8db, 32'shcf1abc4d, 32'shcf1bbfc6, 32'shcf1cc347, 32'shcf1dc6d0, 32'shcf1eca60, 
               32'shcf1fcdf8, 32'shcf20d197, 32'shcf21d53e, 32'shcf22d8ec, 32'shcf23dca2, 32'shcf24e05f, 32'shcf25e424, 32'shcf26e7f1, 
               32'shcf27ebc5, 32'shcf28efa0, 32'shcf29f383, 32'shcf2af76e, 32'shcf2bfb60, 32'shcf2cff5a, 32'shcf2e035b, 32'shcf2f0764, 
               32'shcf300b74, 32'shcf310f8c, 32'shcf3213ab, 32'shcf3317d2, 32'shcf341c00, 32'shcf352036, 32'shcf362473, 32'shcf3728b8, 
               32'shcf382d05, 32'shcf393159, 32'shcf3a35b4, 32'shcf3b3a17, 32'shcf3c3e82, 32'shcf3d42f4, 32'shcf3e476d, 32'shcf3f4bee, 
               32'shcf405077, 32'shcf415507, 32'shcf42599f, 32'shcf435e3e, 32'shcf4462e4, 32'shcf456793, 32'shcf466c48, 32'shcf477105, 
               32'shcf4875ca, 32'shcf497a96, 32'shcf4a7f6a, 32'shcf4b8445, 32'shcf4c8928, 32'shcf4d8e12, 32'shcf4e9304, 32'shcf4f97fe, 
               32'shcf509cfe, 32'shcf51a207, 32'shcf52a716, 32'shcf53ac2e, 32'shcf54b14d, 32'shcf55b673, 32'shcf56bba1, 32'shcf57c0d6, 
               32'shcf58c613, 32'shcf59cb57, 32'shcf5ad0a3, 32'shcf5bd5f7, 32'shcf5cdb51, 32'shcf5de0b4, 32'shcf5ee61e, 32'shcf5feb8f, 
               32'shcf60f108, 32'shcf61f688, 32'shcf62fc10, 32'shcf64019f, 32'shcf650736, 32'shcf660cd5, 32'shcf67127a, 32'shcf681828, 
               32'shcf691ddd, 32'shcf6a2399, 32'shcf6b295d, 32'shcf6c2f28, 32'shcf6d34fb, 32'shcf6e3ad5, 32'shcf6f40b7, 32'shcf7046a0, 
               32'shcf714c91, 32'shcf725289, 32'shcf735889, 32'shcf745e90, 32'shcf75649f, 32'shcf766ab5, 32'shcf7770d3, 32'shcf7876f8, 
               32'shcf797d24, 32'shcf7a8359, 32'shcf7b8994, 32'shcf7c8fd7, 32'shcf7d9622, 32'shcf7e9c74, 32'shcf7fa2cd, 32'shcf80a92e, 
               32'shcf81af97, 32'shcf82b607, 32'shcf83bc7e, 32'shcf84c2fd, 32'shcf85c984, 32'shcf86d012, 32'shcf87d6a7, 32'shcf88dd44, 
               32'shcf89e3e8, 32'shcf8aea94, 32'shcf8bf147, 32'shcf8cf802, 32'shcf8dfec4, 32'shcf8f058e, 32'shcf900c5f, 32'shcf911337, 
               32'shcf921a17, 32'shcf9320ff, 32'shcf9427ee, 32'shcf952ee4, 32'shcf9635e2, 32'shcf973ce8, 32'shcf9843f5, 32'shcf994b09, 
               32'shcf9a5225, 32'shcf9b5948, 32'shcf9c6073, 32'shcf9d67a5, 32'shcf9e6edf, 32'shcf9f7620, 32'shcfa07d68, 32'shcfa184b8, 
               32'shcfa28c10, 32'shcfa3936f, 32'shcfa49ad5, 32'shcfa5a243, 32'shcfa6a9b8, 32'shcfa7b135, 32'shcfa8b8b9, 32'shcfa9c045, 
               32'shcfaac7d8, 32'shcfabcf73, 32'shcfacd715, 32'shcfaddebe, 32'shcfaee66f, 32'shcfafee28, 32'shcfb0f5e7, 32'shcfb1fdaf, 
               32'shcfb3057d, 32'shcfb40d54, 32'shcfb51531, 32'shcfb61d16, 32'shcfb72503, 32'shcfb82cf7, 32'shcfb934f2, 32'shcfba3cf5, 
               32'shcfbb4500, 32'shcfbc4d11, 32'shcfbd552b, 32'shcfbe5d4b, 32'shcfbf6573, 32'shcfc06da3, 32'shcfc175da, 32'shcfc27e18, 
               32'shcfc3865e, 32'shcfc48eab, 32'shcfc59700, 32'shcfc69f5c, 32'shcfc7a7c0, 32'shcfc8b02b, 32'shcfc9b89d, 32'shcfcac117, 
               32'shcfcbc999, 32'shcfccd221, 32'shcfcddab2, 32'shcfcee349, 32'shcfcfebe8, 32'shcfd0f48f, 32'shcfd1fd3d, 32'shcfd305f2, 
               32'shcfd40eaf, 32'shcfd51773, 32'shcfd6203f, 32'shcfd72912, 32'shcfd831ec, 32'shcfd93ace, 32'shcfda43b8, 32'shcfdb4ca8, 
               32'shcfdc55a1, 32'shcfdd5ea0, 32'shcfde67a7, 32'shcfdf70b6, 32'shcfe079cc, 32'shcfe182e9, 32'shcfe28c0e, 32'shcfe3953a, 
               32'shcfe49e6d, 32'shcfe5a7a8, 32'shcfe6b0eb, 32'shcfe7ba35, 32'shcfe8c386, 32'shcfe9ccdf, 32'shcfead63f, 32'shcfebdfa6, 
               32'shcfece915, 32'shcfedf28b, 32'shcfeefc09, 32'shcff0058e, 32'shcff10f1b, 32'shcff218af, 32'shcff3224a, 32'shcff42bed, 
               32'shcff53597, 32'shcff63f49, 32'shcff74902, 32'shcff852c2, 32'shcff95c8a, 32'shcffa6659, 32'shcffb7030, 32'shcffc7a0e, 
               32'shcffd83f4, 32'shcffe8de0, 32'shcfff97d5, 32'shd000a1d0, 32'shd001abd3, 32'shd002b5de, 32'shd003bff0, 32'shd004ca09, 
               32'shd005d42a, 32'shd006de52, 32'shd007e881, 32'shd008f2b8, 32'shd009fcf6, 32'shd00b073c, 32'shd00c1189, 32'shd00d1bdd, 
               32'shd00e2639, 32'shd00f309d, 32'shd0103b07, 32'shd0114579, 32'shd0124ff3, 32'shd0135a73, 32'shd01464fc, 32'shd0156f8b, 
               32'shd0167a22, 32'shd01784c1, 32'shd0188f66, 32'shd0199a13, 32'shd01aa4c8, 32'shd01baf84, 32'shd01cba47, 32'shd01dc512, 
               32'shd01ecfe4, 32'shd01fdabd, 32'shd020e59e, 32'shd021f086, 32'shd022fb76, 32'shd024066d, 32'shd025116b, 32'shd0261c71, 
               32'shd027277e, 32'shd0283293, 32'shd0293dae, 32'shd02a48d2, 32'shd02b53fc, 32'shd02c5f2e, 32'shd02d6a68, 32'shd02e75a8, 
               32'shd02f80f1, 32'shd0308c40, 32'shd0319797, 32'shd032a2f5, 32'shd033ae5b, 32'shd034b9c8, 32'shd035c53c, 32'shd036d0b8, 
               32'shd037dc3b, 32'shd038e7c5, 32'shd039f357, 32'shd03afef1, 32'shd03c0a91, 32'shd03d1639, 32'shd03e21e8, 32'shd03f2d9f, 
               32'shd040395d, 32'shd0414522, 32'shd04250ef, 32'shd0435cc3, 32'shd044689f, 32'shd0457482, 32'shd046806c, 32'shd0478c5d, 
               32'shd0489856, 32'shd049a457, 32'shd04ab05e, 32'shd04bbc6d, 32'shd04cc884, 32'shd04dd4a1, 32'shd04ee0c6, 32'shd04fecf3, 
               32'shd050f926, 32'shd0520562, 32'shd05311a4, 32'shd0541dee, 32'shd0552a3f, 32'shd0563698, 32'shd05742f7, 32'shd0584f5f, 
               32'shd0595bcd, 32'shd05a6843, 32'shd05b74c0, 32'shd05c8145, 32'shd05d8dd1, 32'shd05e9a64, 32'shd05fa6ff, 32'shd060b3a1, 
               32'shd061c04a, 32'shd062ccfb, 32'shd063d9b3, 32'shd064e673, 32'shd065f339, 32'shd0670007, 32'shd0680cdd, 32'shd06919b9, 
               32'shd06a269d, 32'shd06b3389, 32'shd06c407c, 32'shd06d4d76, 32'shd06e5a77, 32'shd06f6780, 32'shd0707490, 32'shd07181a7, 
               32'shd0728ec6, 32'shd0739bec, 32'shd074a91a, 32'shd075b64f, 32'shd076c38b, 32'shd077d0ce, 32'shd078de19, 32'shd079eb6b, 
               32'shd07af8c4, 32'shd07c0625, 32'shd07d138d, 32'shd07e20fc, 32'shd07f2e73, 32'shd0803bf1, 32'shd0814977, 32'shd0825703, 
               32'shd0836497, 32'shd0847233, 32'shd0857fd5, 32'shd0868d7f, 32'shd0879b31, 32'shd088a8e9, 32'shd089b6a9, 32'shd08ac470, 
               32'shd08bd23f, 32'shd08ce015, 32'shd08dedf2, 32'shd08efbd7, 32'shd09009c3, 32'shd09117b6, 32'shd09225b0, 32'shd09333b2, 
               32'shd09441bb, 32'shd0954fcc, 32'shd0965de3, 32'shd0976c02, 32'shd0987a29, 32'shd0998856, 32'shd09a968b, 32'shd09ba4c8, 
               32'shd09cb30b, 32'shd09dc156, 32'shd09ecfa8, 32'shd09fde02, 32'shd0a0ec63, 32'shd0a1facb, 32'shd0a3093a, 32'shd0a417b1, 
               32'shd0a5262f, 32'shd0a634b4, 32'shd0a74341, 32'shd0a851d5, 32'shd0a96070, 32'shd0aa6f13, 32'shd0ab7dbd, 32'shd0ac8c6e, 
               32'shd0ad9b26, 32'shd0aea9e6, 32'shd0afb8ad, 32'shd0b0c77b, 32'shd0b1d651, 32'shd0b2e52e, 32'shd0b3f412, 32'shd0b502fe, 
               32'shd0b611f1, 32'shd0b720eb, 32'shd0b82fec, 32'shd0b93ef5, 32'shd0ba4e05, 32'shd0bb5d1c, 32'shd0bc6c3a, 32'shd0bd7b60, 
               32'shd0be8a8d, 32'shd0bf99c2, 32'shd0c0a8fe, 32'shd0c1b841, 32'shd0c2c78b, 32'shd0c3d6dc, 32'shd0c4e635, 32'shd0c5f595, 
               32'shd0c704fd, 32'shd0c8146c, 32'shd0c923e1, 32'shd0ca335f, 32'shd0cb42e3, 32'shd0cc526f, 32'shd0cd6202, 32'shd0ce719d, 
               32'shd0cf813e, 32'shd0d090e7, 32'shd0d1a097, 32'shd0d2b04f, 32'shd0d3c00e, 32'shd0d4cfd4, 32'shd0d5dfa1, 32'shd0d6ef76, 
               32'shd0d7ff51, 32'shd0d90f35, 32'shd0da1f1f, 32'shd0db2f11, 32'shd0dc3f0a, 32'shd0dd4f0a, 32'shd0de5f11, 32'shd0df6f20, 
               32'shd0e07f36, 32'shd0e18f53, 32'shd0e29f78, 32'shd0e3afa4, 32'shd0e4bfd7, 32'shd0e5d011, 32'shd0e6e053, 32'shd0e7f09b, 
               32'shd0e900ec, 32'shd0ea1143, 32'shd0eb21a2, 32'shd0ec3208, 32'shd0ed4275, 32'shd0ee52e9, 32'shd0ef6365, 32'shd0f073e8, 
               32'shd0f18472, 32'shd0f29503, 32'shd0f3a59c, 32'shd0f4b63c, 32'shd0f5c6e3, 32'shd0f6d792, 32'shd0f7e848, 32'shd0f8f905, 
               32'shd0fa09c9, 32'shd0fb1a94, 32'shd0fc2b67, 32'shd0fd3c41, 32'shd0fe4d22, 32'shd0ff5e0b, 32'shd1006efb, 32'shd1017ff2, 
               32'shd10290f0, 32'shd103a1f5, 32'shd104b302, 32'shd105c416, 32'shd106d531, 32'shd107e654, 32'shd108f77d, 32'shd10a08ae, 
               32'shd10b19e7, 32'shd10c2b26, 32'shd10d3c6d, 32'shd10e4dbb, 32'shd10f5f10, 32'shd110706c, 32'shd11181d0, 32'shd112933b, 
               32'shd113a4ad, 32'shd114b626, 32'shd115c7a7, 32'shd116d92e, 32'shd117eabd, 32'shd118fc54, 32'shd11a0df1, 32'shd11b1f96, 
               32'shd11c3142, 32'shd11d42f5, 32'shd11e54b0, 32'shd11f6671, 32'shd120783a, 32'shd1218a0a, 32'shd1229be2, 32'shd123adc0, 
               32'shd124bfa6, 32'shd125d193, 32'shd126e387, 32'shd127f583, 32'shd1290786, 32'shd12a198f, 32'shd12b2ba1, 32'shd12c3db9, 
               32'shd12d4fd9, 32'shd12e61ff, 32'shd12f742d, 32'shd1308663, 32'shd131989f, 32'shd132aae3, 32'shd133bd2e, 32'shd134cf80, 
               32'shd135e1d9, 32'shd136f43a, 32'shd13806a2, 32'shd1391911, 32'shd13a2b87, 32'shd13b3e04, 32'shd13c5089, 32'shd13d6315, 
               32'shd13e75a8, 32'shd13f8842, 32'shd1409ae3, 32'shd141ad8c, 32'shd142c03c, 32'shd143d2f3, 32'shd144e5b1, 32'shd145f877, 
               32'shd1470b44, 32'shd1481e17, 32'shd14930f3, 32'shd14a43d5, 32'shd14b56be, 32'shd14c69af, 32'shd14d7ca7, 32'shd14e8fa6, 
               32'shd14fa2ad, 32'shd150b5ba, 32'shd151c8cf, 32'shd152dbeb, 32'shd153ef0e, 32'shd1550238, 32'shd156156a, 32'shd15728a2, 
               32'shd1583be2, 32'shd1594f29, 32'shd15a6278, 32'shd15b75cd, 32'shd15c892a, 32'shd15d9c8e, 32'shd15eaff9, 32'shd15fc36b, 
               32'shd160d6e5, 32'shd161ea65, 32'shd162fded, 32'shd164117c, 32'shd1652512, 32'shd16638b0, 32'shd1674c54, 32'shd1686000, 
               32'shd16973b3, 32'shd16a876d, 32'shd16b9b2f, 32'shd16caef7, 32'shd16dc2c7, 32'shd16ed69e, 32'shd16fea7c, 32'shd170fe61, 
               32'shd172124d, 32'shd1732641, 32'shd1743a3c, 32'shd1754e3e, 32'shd1766247, 32'shd1777657, 32'shd1788a6f, 32'shd1799e8d, 
               32'shd17ab2b3, 32'shd17bc6e0, 32'shd17cdb14, 32'shd17def50, 32'shd17f0392, 32'shd18017dc, 32'shd1812c2d, 32'shd1824085, 
               32'shd18354e4, 32'shd184694a, 32'shd1857db8, 32'shd186922d, 32'shd187a6a8, 32'shd188bb2b, 32'shd189cfb6, 32'shd18ae447, 
               32'shd18bf8e0, 32'shd18d0d7f, 32'shd18e2226, 32'shd18f36d4, 32'shd1904b89, 32'shd1916046, 32'shd1927509, 32'shd19389d4, 
               32'shd1949ea6, 32'shd195b37f, 32'shd196c85f, 32'shd197dd46, 32'shd198f235, 32'shd19a072a, 32'shd19b1c27, 32'shd19c312b, 
               32'shd19d4636, 32'shd19e5b48, 32'shd19f7062, 32'shd1a08582, 32'shd1a19aaa, 32'shd1a2afd9, 32'shd1a3c50f, 32'shd1a4da4c, 
               32'shd1a5ef90, 32'shd1a704dc, 32'shd1a81a2e, 32'shd1a92f88, 32'shd1aa44e9, 32'shd1ab5a51, 32'shd1ac6fc0, 32'shd1ad8536, 
               32'shd1ae9ab4, 32'shd1afb038, 32'shd1b0c5c4, 32'shd1b1db57, 32'shd1b2f0f1, 32'shd1b40692, 32'shd1b51c3a, 32'shd1b631ea, 
               32'shd1b747a0, 32'shd1b85d5e, 32'shd1b97323, 32'shd1ba88ef, 32'shd1bb9ec2, 32'shd1bcb49c, 32'shd1bdca7e, 32'shd1bee066, 
               32'shd1bff656, 32'shd1c10c4d, 32'shd1c2224b, 32'shd1c33850, 32'shd1c44e5c, 32'shd1c5646f, 32'shd1c67a8a, 32'shd1c790ab, 
               32'shd1c8a6d4, 32'shd1c9bd04, 32'shd1cad33b, 32'shd1cbe979, 32'shd1ccffbe, 32'shd1ce160a, 32'shd1cf2c5e, 32'shd1d042b8, 
               32'shd1d1591a, 32'shd1d26f83, 32'shd1d385f3, 32'shd1d49c6a, 32'shd1d5b2e8, 32'shd1d6c96d, 32'shd1d7dffa, 32'shd1d8f68d, 
               32'shd1da0d28, 32'shd1db23ca, 32'shd1dc3a73, 32'shd1dd5123, 32'shd1de67da, 32'shd1df7e98, 32'shd1e0955d, 32'shd1e1ac2a, 
               32'shd1e2c2fd, 32'shd1e3d9d8, 32'shd1e4f0ba, 32'shd1e607a3, 32'shd1e71e93, 32'shd1e8358a, 32'shd1e94c88, 32'shd1ea638d, 
               32'shd1eb7a9a, 32'shd1ec91ad, 32'shd1eda8c8, 32'shd1eebfea, 32'shd1efd713, 32'shd1f0ee43, 32'shd1f2057a, 32'shd1f31cb8, 
               32'shd1f433fd, 32'shd1f54b49, 32'shd1f6629d, 32'shd1f779f8, 32'shd1f89159, 32'shd1f9a8c2, 32'shd1fac032, 32'shd1fbd7a9, 
               32'shd1fcef27, 32'shd1fe06ac, 32'shd1ff1e38, 32'shd20035cc, 32'shd2014d66, 32'shd2026508, 32'shd2037cb0, 32'shd2049460, 
               32'shd205ac17, 32'shd206c3d5, 32'shd207db9a, 32'shd208f366, 32'shd20a0b39, 32'shd20b2313, 32'shd20c3af4, 32'shd20d52dd, 
               32'shd20e6acc, 32'shd20f82c3, 32'shd2109ac1, 32'shd211b2c5, 32'shd212cad1, 32'shd213e2e4, 32'shd214fafe, 32'shd216131f, 
               32'shd2172b48, 32'shd2184377, 32'shd2195bad, 32'shd21a73eb, 32'shd21b8c2f, 32'shd21ca47b, 32'shd21dbccd, 32'shd21ed527, 
               32'shd21fed88, 32'shd22105f0, 32'shd2221e5f, 32'shd22336d5, 32'shd2244f52, 32'shd22567d6, 32'shd2268061, 32'shd22798f3, 
               32'shd228b18d, 32'shd229ca2d, 32'shd22ae2d5, 32'shd22bfb83, 32'shd22d1439, 32'shd22e2cf6, 32'shd22f45b9, 32'shd2305e84, 
               32'shd2317756, 32'shd232902f, 32'shd233a90f, 32'shd234c1f6, 32'shd235dae4, 32'shd236f3da, 32'shd2380cd6, 32'shd23925d9, 
               32'shd23a3ee4, 32'shd23b57f5, 32'shd23c710e, 32'shd23d8a2d, 32'shd23ea354, 32'shd23fbc82, 32'shd240d5b6, 32'shd241eef2, 
               32'shd2430835, 32'shd244217f, 32'shd2453ad0, 32'shd2465428, 32'shd2476d87, 32'shd24886ed, 32'shd249a05a, 32'shd24ab9ce, 
               32'shd24bd34a, 32'shd24ceccc, 32'shd24e0655, 32'shd24f1fe6, 32'shd250397d, 32'shd251531c, 32'shd2526cc1, 32'shd253866e, 
               32'shd254a021, 32'shd255b9dc, 32'shd256d39e, 32'shd257ed67, 32'shd2590736, 32'shd25a210d, 32'shd25b3aeb, 32'shd25c54d0, 
               32'shd25d6ebc, 32'shd25e88af, 32'shd25fa2a9, 32'shd260bcaa, 32'shd261d6b2, 32'shd262f0c1, 32'shd2640ad7, 32'shd26524f5, 
               32'shd2663f19, 32'shd2675944, 32'shd2687376, 32'shd2698db0, 32'shd26aa7f0, 32'shd26bc237, 32'shd26cdc86, 32'shd26df6db, 
               32'shd26f1138, 32'shd2702b9b, 32'shd2714606, 32'shd2726077, 32'shd2737af0, 32'shd2749570, 32'shd275aff6, 32'shd276ca84, 
               32'shd277e518, 32'shd278ffb4, 32'shd27a1a57, 32'shd27b3501, 32'shd27c4fb1, 32'shd27d6a69, 32'shd27e8528, 32'shd27f9fee, 
               32'shd280babb, 32'shd281d58e, 32'shd282f069, 32'shd2840b4b, 32'shd2852634, 32'shd2864124, 32'shd2875c1b, 32'shd2887719, 
               32'shd289921e, 32'shd28aad2a, 32'shd28bc83d, 32'shd28ce357, 32'shd28dfe77, 32'shd28f199f, 32'shd29034ce, 32'shd2915004, 
               32'shd2926b41, 32'shd2938685, 32'shd294a1d0, 32'shd295bd23, 32'shd296d87c, 32'shd297f3dc, 32'shd2990f43, 32'shd29a2ab1, 
               32'shd29b4626, 32'shd29c61a2, 32'shd29d7d25, 32'shd29e98af, 32'shd29fb440, 32'shd2a0cfd8, 32'shd2a1eb77, 32'shd2a3071d, 
               32'shd2a422ca, 32'shd2a53e7e, 32'shd2a65a39, 32'shd2a775fb, 32'shd2a891c4, 32'shd2a9ad94, 32'shd2aac96b, 32'shd2abe549, 
               32'shd2ad012e, 32'shd2ae1d1a, 32'shd2af390d, 32'shd2b05506, 32'shd2b17107, 32'shd2b28d0f, 32'shd2b3a91e, 32'shd2b4c534, 
               32'shd2b5e151, 32'shd2b6fd75, 32'shd2b8199f, 32'shd2b935d1, 32'shd2ba520a, 32'shd2bb6e4a, 32'shd2bc8a91, 32'shd2bda6de, 
               32'shd2bec333, 32'shd2bfdf8f, 32'shd2c0fbf1, 32'shd2c2185b, 32'shd2c334cc, 32'shd2c45143, 32'shd2c56dc2, 32'shd2c68a47, 
               32'shd2c7a6d4, 32'shd2c8c367, 32'shd2c9e002, 32'shd2cafca3, 32'shd2cc194c, 32'shd2cd35fb, 32'shd2ce52b1, 32'shd2cf6f6f, 
               32'shd2d08c33, 32'shd2d1a8fe, 32'shd2d2c5d0, 32'shd2d3e2aa, 32'shd2d4ff8a, 32'shd2d61c71, 32'shd2d7395f, 32'shd2d85654, 
               32'shd2d97350, 32'shd2da9053, 32'shd2dbad5d, 32'shd2dcca6e, 32'shd2dde786, 32'shd2df04a5, 32'shd2e021ca, 32'shd2e13ef7, 
               32'shd2e25c2b, 32'shd2e37965, 32'shd2e496a7, 32'shd2e5b3f0, 32'shd2e6d13f, 32'shd2e7ee96, 32'shd2e90bf3, 32'shd2ea2957, 
               32'shd2eb46c3, 32'shd2ec6435, 32'shd2ed81ae, 32'shd2ee9f2e, 32'shd2efbcb6, 32'shd2f0da44, 32'shd2f1f7d9, 32'shd2f31575, 
               32'shd2f43318, 32'shd2f550c2, 32'shd2f66e72, 32'shd2f78c2a, 32'shd2f8a9e9, 32'shd2f9c7ae, 32'shd2fae57b, 32'shd2fc034f, 
               32'shd2fd2129, 32'shd2fe3f0b, 32'shd2ff5cf3, 32'shd3007ae2, 32'shd30198d8, 32'shd302b6d6, 32'shd303d4da, 32'shd304f2e5, 
               32'shd30610f7, 32'shd3072f10, 32'shd3084d30, 32'shd3096b56, 32'shd30a8984, 32'shd30ba7b9, 32'shd30cc5f4, 32'shd30de437, 
               32'shd30f0280, 32'shd31020d1, 32'shd3113f28, 32'shd3125d86, 32'shd3137bec, 32'shd3149a58, 32'shd315b8cb, 32'shd316d745, 
               32'shd317f5c6, 32'shd319144e, 32'shd31a32dc, 32'shd31b5172, 32'shd31c700f, 32'shd31d8eb2, 32'shd31ead5c, 32'shd31fcc0e, 
               32'shd320eac6, 32'shd3220985, 32'shd323284b, 32'shd3244718, 32'shd32565ec, 32'shd32684c7, 32'shd327a3a9, 32'shd328c292, 
               32'shd329e181, 32'shd32b0078, 32'shd32c1f75, 32'shd32d3e7a, 32'shd32e5d85, 32'shd32f7c97, 32'shd3309bb0, 32'shd331bad0, 
               32'shd332d9f7, 32'shd333f925, 32'shd335185a, 32'shd3363795, 32'shd33756d8, 32'shd3387621, 32'shd3399572, 32'shd33ab4c9, 
               32'shd33bd427, 32'shd33cf38c, 32'shd33e12f8, 32'shd33f326b, 32'shd34051e5, 32'shd3417165, 32'shd34290ed, 32'shd343b07b, 
               32'shd344d011, 32'shd345efad, 32'shd3470f50, 32'shd3482efa, 32'shd3494eab, 32'shd34a6e63, 32'shd34b8e22, 32'shd34cade8, 
               32'shd34dcdb4, 32'shd34eed88, 32'shd3500d62, 32'shd3512d43, 32'shd3524d2b, 32'shd3536d1a, 32'shd3548d10, 32'shd355ad0d, 
               32'shd356cd11, 32'shd357ed1b, 32'shd3590d2c, 32'shd35a2d45, 32'shd35b4d64, 32'shd35c6d8a, 32'shd35d8db7, 32'shd35eadeb, 
               32'shd35fce26, 32'shd360ee67, 32'shd3620eb0, 32'shd3632eff, 32'shd3644f55, 32'shd3656fb3, 32'shd3669017, 32'shd367b082, 
               32'shd368d0f3, 32'shd369f16c, 32'shd36b11eb, 32'shd36c3272, 32'shd36d52ff, 32'shd36e7393, 32'shd36f942e, 32'shd370b4d0, 
               32'shd371d579, 32'shd372f629, 32'shd37416df, 32'shd375379d, 32'shd3765861, 32'shd377792c, 32'shd37899fe, 32'shd379bad7, 
               32'shd37adbb6, 32'shd37bfc9d, 32'shd37d1d8a, 32'shd37e3e7f, 32'shd37f5f7a, 32'shd380807c, 32'shd381a185, 32'shd382c295, 
               32'shd383e3ab, 32'shd38504c9, 32'shd38625ed, 32'shd3874718, 32'shd388684a, 32'shd3898983, 32'shd38aaac3, 32'shd38bcc0a, 
               32'shd38ced57, 32'shd38e0eac, 32'shd38f3007, 32'shd3905169, 32'shd39172d2, 32'shd3929441, 32'shd393b5b8, 32'shd394d735, 
               32'shd395f8ba, 32'shd3971a45, 32'shd3983bd7, 32'shd3995d70, 32'shd39a7f0f, 32'shd39ba0b6, 32'shd39cc263, 32'shd39de418, 
               32'shd39f05d3, 32'shd3a02795, 32'shd3a1495d, 32'shd3a26b2d, 32'shd3a38d03, 32'shd3a4aee1, 32'shd3a5d0c5, 32'shd3a6f2b0, 
               32'shd3a814a2, 32'shd3a9369a, 32'shd3aa589a, 32'shd3ab7aa0, 32'shd3ac9cad, 32'shd3adbec1, 32'shd3aee0dc, 32'shd3b002fe, 
               32'shd3b12526, 32'shd3b24756, 32'shd3b3698c, 32'shd3b48bc9, 32'shd3b5ae0d, 32'shd3b6d057, 32'shd3b7f2a9, 32'shd3b91501, 
               32'shd3ba3760, 32'shd3bb59c6, 32'shd3bc7c33, 32'shd3bd9ea7, 32'shd3bec121, 32'shd3bfe3a2, 32'shd3c1062a, 32'shd3c228b9, 
               32'shd3c34b4f, 32'shd3c46dec, 32'shd3c5908f, 32'shd3c6b339, 32'shd3c7d5ea, 32'shd3c8f8a2, 32'shd3ca1b61, 32'shd3cb3e26, 
               32'shd3cc60f2, 32'shd3cd83c6, 32'shd3cea69f, 32'shd3cfc980, 32'shd3d0ec68, 32'shd3d20f56, 32'shd3d3324b, 32'shd3d45547, 
               32'shd3d5784a, 32'shd3d69b54, 32'shd3d7be64, 32'shd3d8e17b, 32'shd3da049a, 32'shd3db27be, 32'shd3dc4aea, 32'shd3dd6e1c, 
               32'shd3de9156, 32'shd3dfb496, 32'shd3e0d7dd, 32'shd3e1fb2a, 32'shd3e31e7f, 32'shd3e441da, 32'shd3e5653c, 32'shd3e688a5, 
               32'shd3e7ac15, 32'shd3e8cf8b, 32'shd3e9f309, 32'shd3eb168d, 32'shd3ec3a18, 32'shd3ed5da9, 32'shd3ee8142, 32'shd3efa4e1, 
               32'shd3f0c887, 32'shd3f1ec34, 32'shd3f30fe8, 32'shd3f433a2, 32'shd3f55764, 32'shd3f67b2c, 32'shd3f79efa, 32'shd3f8c2d0, 
               32'shd3f9e6ad, 32'shd3fb0a90, 32'shd3fc2e7a, 32'shd3fd526a, 32'shd3fe7662, 32'shd3ff9a60, 32'shd400be66, 32'shd401e271, 
               32'shd4030684, 32'shd4042a9e, 32'shd4054ebe, 32'shd40672e5, 32'shd4079713, 32'shd408bb48, 32'shd409df83, 32'shd40b03c5, 
               32'shd40c280e, 32'shd40d4c5e, 32'shd40e70b4, 32'shd40f9512, 32'shd410b976, 32'shd411dde1, 32'shd4130252, 32'shd41426cb, 
               32'shd4154b4a, 32'shd4166fd0, 32'shd417945c, 32'shd418b8f0, 32'shd419dd8a, 32'shd41b022b, 32'shd41c26d3, 32'shd41d4b81, 
               32'shd41e7037, 32'shd41f94f3, 32'shd420b9b6, 32'shd421de7f, 32'shd4230350, 32'shd4242827, 32'shd4254d05, 32'shd42671ea, 
               32'shd42796d5, 32'shd428bbc7, 32'shd429e0c0, 32'shd42b05c0, 32'shd42c2ac6, 32'shd42d4fd4, 32'shd42e74e8, 32'shd42f9a02, 
               32'shd430bf24, 32'shd431e44c, 32'shd433097b, 32'shd4342eb1, 32'shd43553ee, 32'shd4367931, 32'shd4379e7b, 32'shd438c3cc, 
               32'shd439e923, 32'shd43b0e81, 32'shd43c33e7, 32'shd43d5952, 32'shd43e7ec5, 32'shd43fa43e, 32'shd440c9be, 32'shd441ef45, 
               32'shd44314d3, 32'shd4443a67, 32'shd4456002, 32'shd44685a4, 32'shd447ab4c, 32'shd448d0fb, 32'shd449f6b1, 32'shd44b1c6e, 
               32'shd44c4232, 32'shd44d67fc, 32'shd44e8dcd, 32'shd44fb3a4, 32'shd450d983, 32'shd451ff68, 32'shd4532554, 32'shd4544b46, 
               32'shd4557140, 32'shd4569740, 32'shd457bd47, 32'shd458e354, 32'shd45a0969, 32'shd45b2f84, 32'shd45c55a5, 32'shd45d7bce, 
               32'shd45ea1fd, 32'shd45fc833, 32'shd460ee70, 32'shd46214b3, 32'shd4633afd, 32'shd464614e, 32'shd46587a6, 32'shd466ae04, 
               32'shd467d469, 32'shd468fad5, 32'shd46a2147, 32'shd46b47c0, 32'shd46c6e40, 32'shd46d94c7, 32'shd46ebb54, 32'shd46fe1e8, 
               32'shd4710883, 32'shd4722f25, 32'shd47355cd, 32'shd4747c7c, 32'shd475a332, 32'shd476c9ee, 32'shd477f0b1, 32'shd479177b, 
               32'shd47a3e4b, 32'shd47b6523, 32'shd47c8c00, 32'shd47db2e5, 32'shd47ed9d0, 32'shd48000c2, 32'shd48127bb, 32'shd4824ebb, 
               32'shd48375c1, 32'shd4849cce, 32'shd485c3e1, 32'shd486eafc, 32'shd488121d, 32'shd4893944, 32'shd48a6073, 32'shd48b87a8, 
               32'shd48caee4, 32'shd48dd626, 32'shd48efd6f, 32'shd49024bf, 32'shd4914c16, 32'shd4927373, 32'shd4939ad7, 32'shd494c242, 
               32'shd495e9b3, 32'shd497112b, 32'shd49838aa, 32'shd4996030, 32'shd49a87bc, 32'shd49baf4f, 32'shd49cd6e8, 32'shd49dfe89, 
               32'shd49f2630, 32'shd4a04ddd, 32'shd4a17591, 32'shd4a29d4c, 32'shd4a3c50e, 32'shd4a4ecd7, 32'shd4a614a6, 32'shd4a73c7b, 
               32'shd4a86458, 32'shd4a98c3b, 32'shd4aab425, 32'shd4abdc15, 32'shd4ad040c, 32'shd4ae2c0a, 32'shd4af540f, 32'shd4b07c1a, 
               32'shd4b1a42c, 32'shd4b2cc44, 32'shd4b3f464, 32'shd4b51c8a, 32'shd4b644b6, 32'shd4b76ce9, 32'shd4b89523, 32'shd4b9bd64, 
               32'shd4bae5ab, 32'shd4bc0df9, 32'shd4bd364e, 32'shd4be5ea9, 32'shd4bf870b, 32'shd4c0af74, 32'shd4c1d7e3, 32'shd4c30059, 
               32'shd4c428d6, 32'shd4c55159, 32'shd4c679e3, 32'shd4c7a274, 32'shd4c8cb0b, 32'shd4c9f3a9, 32'shd4cb1c4e, 32'shd4cc44f9, 
               32'shd4cd6dab, 32'shd4ce9664, 32'shd4cfbf23, 32'shd4d0e7e9, 32'shd4d210b5, 32'shd4d33989, 32'shd4d46263, 32'shd4d58b43, 
               32'shd4d6b42b, 32'shd4d7dd18, 32'shd4d9060d, 32'shd4da2f08, 32'shd4db580a, 32'shd4dc8113, 32'shd4ddaa22, 32'shd4ded338, 
               32'shd4dffc54, 32'shd4e12577, 32'shd4e24ea1, 32'shd4e377d1, 32'shd4e4a108, 32'shd4e5ca46, 32'shd4e6f38b, 32'shd4e81cd6, 
               32'shd4e94627, 32'shd4ea6f80, 32'shd4eb98de, 32'shd4ecc244, 32'shd4edebb0, 32'shd4ef1523, 32'shd4f03e9d, 32'shd4f1681d, 
               32'shd4f291a4, 32'shd4f3bb31, 32'shd4f4e4c5, 32'shd4f60e60, 32'shd4f73801, 32'shd4f861a9, 32'shd4f98b58, 32'shd4fab50d, 
               32'shd4fbdec9, 32'shd4fd088c, 32'shd4fe3255, 32'shd4ff5c24, 32'shd50085fb, 32'shd501afd8, 32'shd502d9bc, 32'shd50403a6, 
               32'shd5052d97, 32'shd506578e, 32'shd507818d, 32'shd508ab91, 32'shd509d59d, 32'shd50affaf, 32'shd50c29c8, 32'shd50d53e7, 
               32'shd50e7e0d, 32'shd50fa83a, 32'shd510d26d, 32'shd511fca7, 32'shd51326e7, 32'shd514512e, 32'shd5157b7c, 32'shd516a5d0, 
               32'shd517d02b, 32'shd518fa8c, 32'shd51a24f5, 32'shd51b4f63, 32'shd51c79d9, 32'shd51da455, 32'shd51eced7, 32'shd51ff960, 
               32'shd52123f0, 32'shd5224e87, 32'shd5237924, 32'shd524a3c7, 32'shd525ce72, 32'shd526f923, 32'shd52823da, 32'shd5294e98, 
               32'shd52a795d, 32'shd52ba428, 32'shd52ccefa, 32'shd52df9d3, 32'shd52f24b2, 32'shd5304f97, 32'shd5317a84, 32'shd532a577, 
               32'shd533d070, 32'shd534fb70, 32'shd5362677, 32'shd5375184, 32'shd5387c98, 32'shd539a7b3, 32'shd53ad2d4, 32'shd53bfdfb, 
               32'shd53d292a, 32'shd53e545f, 32'shd53f7f9a, 32'shd540aadc, 32'shd541d625, 32'shd5430174, 32'shd5442cca, 32'shd5455826, 
               32'shd5468389, 32'shd547aef3, 32'shd548da63, 32'shd54a05da, 32'shd54b3157, 32'shd54c5cdb, 32'shd54d8866, 32'shd54eb3f7, 
               32'shd54fdf8f, 32'shd5510b2d, 32'shd55236d2, 32'shd553627d, 32'shd5548e30, 32'shd555b9e8, 32'shd556e5a7, 32'shd558116d, 
               32'shd5593d3a, 32'shd55a690c, 32'shd55b94e6, 32'shd55cc0c6, 32'shd55decad, 32'shd55f189a, 32'shd560448e, 32'shd5617088, 
               32'shd5629c89, 32'shd563c891, 32'shd564f49f, 32'shd56620b3, 32'shd5674ccf, 32'shd56878f1, 32'shd569a519, 32'shd56ad148, 
               32'shd56bfd7d, 32'shd56d29b9, 32'shd56e55fc, 32'shd56f8245, 32'shd570ae95, 32'shd571daeb, 32'shd5730748, 32'shd57433ac, 
               32'shd5756016, 32'shd5768c86, 32'shd577b8fe, 32'shd578e57b, 32'shd57a1200, 32'shd57b3e8a, 32'shd57c6b1c, 32'shd57d97b4, 
               32'shd57ec452, 32'shd57ff0f7, 32'shd5811da3, 32'shd5824a55, 32'shd583770e, 32'shd584a3cd, 32'shd585d093, 32'shd586fd5f, 
               32'shd5882a32, 32'shd589570b, 32'shd58a83eb, 32'shd58bb0d2, 32'shd58cddbf, 32'shd58e0ab3, 32'shd58f37ad, 32'shd59064ae, 
               32'shd59191b5, 32'shd592bec3, 32'shd593ebd7, 32'shd59518f2, 32'shd5964614, 32'shd597733c, 32'shd598a06a, 32'shd599cd9f, 
               32'shd59afadb, 32'shd59c281d, 32'shd59d5566, 32'shd59e82b5, 32'shd59fb00b, 32'shd5a0dd67, 32'shd5a20aca, 32'shd5a33833, 
               32'shd5a465a3, 32'shd5a59319, 32'shd5a6c096, 32'shd5a7ee1a, 32'shd5a91ba4, 32'shd5aa4934, 32'shd5ab76cb, 32'shd5aca469, 
               32'shd5add20d, 32'shd5aeffb8, 32'shd5b02d69, 32'shd5b15b21, 32'shd5b288df, 32'shd5b3b6a4, 32'shd5b4e46f, 32'shd5b61241, 
               32'shd5b74019, 32'shd5b86df8, 32'shd5b99bdd, 32'shd5bac9c9, 32'shd5bbf7bc, 32'shd5bd25b4, 32'shd5be53b4, 32'shd5bf81ba, 
               32'shd5c0afc6, 32'shd5c1ddd9, 32'shd5c30bf3, 32'shd5c43a13, 32'shd5c56839, 32'shd5c69666, 32'shd5c7c49a, 32'shd5c8f2d4, 
               32'shd5ca2115, 32'shd5cb4f5c, 32'shd5cc7da9, 32'shd5cdabfd, 32'shd5ceda58, 32'shd5d008b9, 32'shd5d13721, 32'shd5d2658f, 
               32'shd5d39403, 32'shd5d4c27e, 32'shd5d5f100, 32'shd5d71f88, 32'shd5d84e17, 32'shd5d97cac, 32'shd5daab48, 32'shd5dbd9ea, 
               32'shd5dd0892, 32'shd5de3742, 32'shd5df65f7, 32'shd5e094b3, 32'shd5e1c376, 32'shd5e2f23f, 32'shd5e4210f, 32'shd5e54fe5, 
               32'shd5e67ec1, 32'shd5e7ada4, 32'shd5e8dc8e, 32'shd5ea0b7e, 32'shd5eb3a75, 32'shd5ec6972, 32'shd5ed9875, 32'shd5eec77f, 
               32'shd5eff690, 32'shd5f125a7, 32'shd5f254c4, 32'shd5f383e8, 32'shd5f4b313, 32'shd5f5e244, 32'shd5f7117b, 32'shd5f840b9, 
               32'shd5f96ffd, 32'shd5fa9f48, 32'shd5fbce9a, 32'shd5fcfdf1, 32'shd5fe2d50, 32'shd5ff5cb4, 32'shd6008c20, 32'shd601bb91, 
               32'shd602eb0a, 32'shd6041a88, 32'shd6054a0d, 32'shd6067999, 32'shd607a92b, 32'shd608d8c4, 32'shd60a0863, 32'shd60b3808, 
               32'shd60c67b4, 32'shd60d9767, 32'shd60ec720, 32'shd60ff6df, 32'shd61126a5, 32'shd6125671, 32'shd6138644, 32'shd614b61d, 
               32'shd615e5fd, 32'shd61715e3, 32'shd61845d0, 32'shd61975c3, 32'shd61aa5bd, 32'shd61bd5bd, 32'shd61d05c3, 32'shd61e35d0, 
               32'shd61f65e4, 32'shd62095fe, 32'shd621c61e, 32'shd622f645, 32'shd6242672, 32'shd62556a6, 32'shd62686e0, 32'shd627b720, 
               32'shd628e767, 32'shd62a17b5, 32'shd62b4809, 32'shd62c7863, 32'shd62da8c4, 32'shd62ed92c, 32'shd6300999, 32'shd6313a0e, 
               32'shd6326a88, 32'shd6339b09, 32'shd634cb91, 32'shd635fc1f, 32'shd6372cb3, 32'shd6385d4e, 32'shd6398df0, 32'shd63abe97, 
               32'shd63bef46, 32'shd63d1ffa, 32'shd63e50b5, 32'shd63f8177, 32'shd640b23f, 32'shd641e30d, 32'shd64313e2, 32'shd64444bd, 
               32'shd645759f, 32'shd646a687, 32'shd647d776, 32'shd649086b, 32'shd64a3966, 32'shd64b6a68, 32'shd64c9b71, 32'shd64dcc7f, 
               32'shd64efd94, 32'shd6502eb0, 32'shd6515fd2, 32'shd65290fb, 32'shd653c229, 32'shd654f35f, 32'shd656249b, 32'shd65755dd, 
               32'shd6588725, 32'shd659b874, 32'shd65ae9ca, 32'shd65c1b26, 32'shd65d4c88, 32'shd65e7df1, 32'shd65faf60, 32'shd660e0d5, 
               32'shd6621251, 32'shd66343d4, 32'shd664755c, 32'shd665a6ec, 32'shd666d881, 32'shd6680a1d, 32'shd6693bc0, 32'shd66a6d69, 
               32'shd66b9f18, 32'shd66cd0ce, 32'shd66e028a, 32'shd66f344c, 32'shd6706615, 32'shd67197e5, 32'shd672c9ba, 32'shd673fb97, 
               32'shd6752d79, 32'shd6765f62, 32'shd6779151, 32'shd678c347, 32'shd679f543, 32'shd67b2746, 32'shd67c594f, 32'shd67d8b5e, 
               32'shd67ebd74, 32'shd67fef90, 32'shd68121b3, 32'shd68253dc, 32'shd683860b, 32'shd684b841, 32'shd685ea7d, 32'shd6871cc0, 
               32'shd6884f09, 32'shd6898158, 32'shd68ab3ae, 32'shd68be60a, 32'shd68d186d, 32'shd68e4ad6, 32'shd68f7d45, 32'shd690afbb, 
               32'shd691e237, 32'shd69314b9, 32'shd6944742, 32'shd69579d2, 32'shd696ac67, 32'shd697df03, 32'shd69911a6, 32'shd69a444f, 
               32'shd69b76fe, 32'shd69ca9b3, 32'shd69ddc6f, 32'shd69f0f32, 32'shd6a041fa, 32'shd6a174ca, 32'shd6a2a79f, 32'shd6a3da7b, 
               32'shd6a50d5d, 32'shd6a64046, 32'shd6a77335, 32'shd6a8a62a, 32'shd6a9d926, 32'shd6ab0c28, 32'shd6ac3f31, 32'shd6ad7240, 
               32'shd6aea555, 32'shd6afd870, 32'shd6b10b92, 32'shd6b23ebb, 32'shd6b371ea, 32'shd6b4a51f, 32'shd6b5d85a, 32'shd6b70b9c, 
               32'shd6b83ee4, 32'shd6b97233, 32'shd6baa588, 32'shd6bbd8e3, 32'shd6bd0c45, 32'shd6be3fad, 32'shd6bf731b, 32'shd6c0a690, 
               32'shd6c1da0b, 32'shd6c30d8c, 32'shd6c44114, 32'shd6c574a2, 32'shd6c6a837, 32'shd6c7dbd2, 32'shd6c90f73, 32'shd6ca431b, 
               32'shd6cb76c9, 32'shd6ccaa7d, 32'shd6cdde38, 32'shd6cf11f9, 32'shd6d045c0, 32'shd6d1798e, 32'shd6d2ad62, 32'shd6d3e13d, 
               32'shd6d5151d, 32'shd6d64904, 32'shd6d77cf2, 32'shd6d8b0e6, 32'shd6d9e4e0, 32'shd6db18e0, 32'shd6dc4ce7, 32'shd6dd80f5, 
               32'shd6deb508, 32'shd6dfe922, 32'shd6e11d42, 32'shd6e25169, 32'shd6e38596, 32'shd6e4b9c9, 32'shd6e5ee03, 32'shd6e72243, 
               32'shd6e85689, 32'shd6e98ad6, 32'shd6eabf28, 32'shd6ebf382, 32'shd6ed27e1, 32'shd6ee5c47, 32'shd6ef90b4, 32'shd6f0c526, 
               32'shd6f1f99f, 32'shd6f32e1f, 32'shd6f462a4, 32'shd6f59730, 32'shd6f6cbc2, 32'shd6f8005b, 32'shd6f934fa, 32'shd6fa699f, 
               32'shd6fb9e4b, 32'shd6fcd2fd, 32'shd6fe07b5, 32'shd6ff3c73, 32'shd7007138, 32'shd701a604, 32'shd702dad5, 32'shd7040fad, 
               32'shd705448b, 32'shd7067970, 32'shd707ae5a, 32'shd708e34c, 32'shd70a1843, 32'shd70b4d41, 32'shd70c8245, 32'shd70db74f, 
               32'shd70eec60, 32'shd7102177, 32'shd7115694, 32'shd7128bb8, 32'shd713c0e2, 32'shd714f612, 32'shd7162b49, 32'shd7176086, 
               32'shd71895c9, 32'shd719cb12, 32'shd71b0062, 32'shd71c35b8, 32'shd71d6b15, 32'shd71ea077, 32'shd71fd5e0, 32'shd7210b50, 
               32'shd72240c5, 32'shd7237641, 32'shd724abc4, 32'shd725e14c, 32'shd72716db, 32'shd7284c70, 32'shd729820c, 32'shd72ab7ad, 
               32'shd72bed55, 32'shd72d2304, 32'shd72e58b8, 32'shd72f8e73, 32'shd730c434, 32'shd731f9fc, 32'shd7332fca, 32'shd734659e, 
               32'shd7359b78, 32'shd736d159, 32'shd7380740, 32'shd7393d2d, 32'shd73a7321, 32'shd73ba91a, 32'shd73cdf1b, 32'shd73e1521, 
               32'shd73f4b2e, 32'shd7408141, 32'shd741b75a, 32'shd742ed79, 32'shd744239f, 32'shd74559cb, 32'shd7468ffe, 32'shd747c636, 
               32'shd748fc75, 32'shd74a32bb, 32'shd74b6906, 32'shd74c9f58, 32'shd74dd5b0, 32'shd74f0c0e, 32'shd7504273, 32'shd75178de, 
               32'shd752af4f, 32'shd753e5c6, 32'shd7551c44, 32'shd75652c8, 32'shd7578952, 32'shd758bfe3, 32'shd759f679, 32'shd75b2d17, 
               32'shd75c63ba, 32'shd75d9a63, 32'shd75ed113, 32'shd76007c9, 32'shd7613e86, 32'shd7627548, 32'shd763ac11, 32'shd764e2e0, 
               32'shd76619b6, 32'shd7675092, 32'shd7688774, 32'shd769be5c, 32'shd76af54a, 32'shd76c2c3f, 32'shd76d633a, 32'shd76e9a3b, 
               32'shd76fd143, 32'shd7710850, 32'shd7723f64, 32'shd773767f, 32'shd774ad9f, 32'shd775e4c6, 32'shd7771bf3, 32'shd7785326, 
               32'shd7798a60, 32'shd77ac1a0, 32'shd77bf8e6, 32'shd77d3032, 32'shd77e6784, 32'shd77f9edd, 32'shd780d63c, 32'shd7820da1, 
               32'shd783450d, 32'shd7847c7f, 32'shd785b3f7, 32'shd786eb75, 32'shd78822f9, 32'shd7895a84, 32'shd78a9215, 32'shd78bc9ac, 
               32'shd78d014a, 32'shd78e38ed, 32'shd78f7097, 32'shd790a847, 32'shd791dffe, 32'shd79317ba, 32'shd7944f7d, 32'shd7958746, 
               32'shd796bf16, 32'shd797f6eb, 32'shd7992ec7, 32'shd79a66a9, 32'shd79b9e91, 32'shd79cd680, 32'shd79e0e74, 32'shd79f466f, 
               32'shd7a07e70, 32'shd7a1b678, 32'shd7a2ee85, 32'shd7a42699, 32'shd7a55eb3, 32'shd7a696d3, 32'shd7a7cefa, 32'shd7a90727, 
               32'shd7aa3f5a, 32'shd7ab7793, 32'shd7acafd2, 32'shd7ade818, 32'shd7af2063, 32'shd7b058b6, 32'shd7b1910e, 32'shd7b2c96c, 
               32'shd7b401d1, 32'shd7b53a3c, 32'shd7b672ad, 32'shd7b7ab24, 32'shd7b8e3a2, 32'shd7ba1c25, 32'shd7bb54af, 32'shd7bc8d40, 
               32'shd7bdc5d6, 32'shd7befe72, 32'shd7c03715, 32'shd7c16fbe, 32'shd7c2a86d, 32'shd7c3e123, 32'shd7c519de, 32'shd7c652a0, 
               32'shd7c78b68, 32'shd7c8c436, 32'shd7c9fd0b, 32'shd7cb35e6, 32'shd7cc6ec6, 32'shd7cda7ad, 32'shd7cee09b, 32'shd7d0198e, 
               32'shd7d15288, 32'shd7d28b87, 32'shd7d3c48d, 32'shd7d4fd9a, 32'shd7d636ac, 32'shd7d76fc5, 32'shd7d8a8e3, 32'shd7d9e208, 
               32'shd7db1b34, 32'shd7dc5465, 32'shd7dd8d9c, 32'shd7dec6da, 32'shd7e0001e, 32'shd7e13968, 32'shd7e272b8, 32'shd7e3ac0f, 
               32'shd7e4e56c, 32'shd7e61ece, 32'shd7e75838, 32'shd7e891a7, 32'shd7e9cb1c, 32'shd7eb0498, 32'shd7ec3e1a, 32'shd7ed77a1, 
               32'shd7eeb130, 32'shd7efeac4, 32'shd7f1245e, 32'shd7f25dff, 32'shd7f397a6, 32'shd7f4d153, 32'shd7f60b06, 32'shd7f744bf, 
               32'shd7f87e7f, 32'shd7f9b845, 32'shd7faf211, 32'shd7fc2be3, 32'shd7fd65bb, 32'shd7fe9f99, 32'shd7ffd97e, 32'shd8011369, 
               32'shd8024d59, 32'shd8038751, 32'shd804c14e, 32'shd805fb51, 32'shd807355b, 32'shd8086f6a, 32'shd809a980, 32'shd80ae39c, 
               32'shd80c1dbf, 32'shd80d57e7, 32'shd80e9216, 32'shd80fcc4a, 32'shd8110685, 32'shd81240c6, 32'shd8137b0d, 32'shd814b55b, 
               32'shd815efae, 32'shd8172a08, 32'shd8186468, 32'shd8199ecd, 32'shd81ad93a, 32'shd81c13ac, 32'shd81d4e24, 32'shd81e88a3, 
               32'shd81fc328, 32'shd820fdb2, 32'shd8223843, 32'shd82372db, 32'shd824ad78, 32'shd825e81b, 32'shd82722c5, 32'shd8285d75, 
               32'shd829982b, 32'shd82ad2e7, 32'shd82c0da9, 32'shd82d4871, 32'shd82e833f, 32'shd82fbe14, 32'shd830f8ef, 32'shd83233d0, 
               32'shd8336eb7, 32'shd834a9a4, 32'shd835e497, 32'shd8371f91, 32'shd8385a90, 32'shd8399596, 32'shd83ad0a2, 32'shd83c0bb4, 
               32'shd83d46cc, 32'shd83e81ea, 32'shd83fbd0e, 32'shd840f839, 32'shd8423369, 32'shd8436ea0, 32'shd844a9dd, 32'shd845e520, 
               32'shd8472069, 32'shd8485bb8, 32'shd849970e, 32'shd84ad269, 32'shd84c0dcb, 32'shd84d4933, 32'shd84e84a0, 32'shd84fc014, 
               32'shd850fb8e, 32'shd852370f, 32'shd8537295, 32'shd854ae21, 32'shd855e9b4, 32'shd857254d, 32'shd85860ec, 32'shd8599c91, 
               32'shd85ad83c, 32'shd85c13ed, 32'shd85d4fa4, 32'shd85e8b61, 32'shd85fc725, 32'shd86102ee, 32'shd8623ebe, 32'shd8637a94, 
               32'shd864b670, 32'shd865f252, 32'shd8672e3a, 32'shd8686a28, 32'shd869a61d, 32'shd86ae217, 32'shd86c1e18, 32'shd86d5a1e, 
               32'shd86e962b, 32'shd86fd23e, 32'shd8710e57, 32'shd8724a76, 32'shd873869b, 32'shd874c2c7, 32'shd875fef8, 32'shd8773b2f, 
               32'shd878776d, 32'shd879b3b1, 32'shd87aeffa, 32'shd87c2c4a, 32'shd87d68a0, 32'shd87ea4fc, 32'shd87fe15e, 32'shd8811dc7, 
               32'shd8825a35, 32'shd88396a9, 32'shd884d324, 32'shd8860fa4, 32'shd8874c2b, 32'shd88888b8, 32'shd889c54b, 32'shd88b01e4, 
               32'shd88c3e83, 32'shd88d7b28, 32'shd88eb7d3, 32'shd88ff484, 32'shd891313b, 32'shd8926df9, 32'shd893aabc, 32'shd894e786, 
               32'shd8962456, 32'shd897612b, 32'shd8989e07, 32'shd899dae9, 32'shd89b17d1, 32'shd89c54bf, 32'shd89d91b3, 32'shd89ecead, 
               32'shd8a00bae, 32'shd8a148b4, 32'shd8a285c0, 32'shd8a3c2d3, 32'shd8a4ffec, 32'shd8a63d0a, 32'shd8a77a2f, 32'shd8a8b75a, 
               32'shd8a9f48a, 32'shd8ab31c1, 32'shd8ac6efe, 32'shd8adac41, 32'shd8aee98a, 32'shd8b026da, 32'shd8b1642f, 32'shd8b2a18a, 
               32'shd8b3deeb, 32'shd8b51c53, 32'shd8b659c0, 32'shd8b79734, 32'shd8b8d4ad, 32'shd8ba122d, 32'shd8bb4fb3, 32'shd8bc8d3e, 
               32'shd8bdcad0, 32'shd8bf0868, 32'shd8c04606, 32'shd8c183aa, 32'shd8c2c154, 32'shd8c3ff04, 32'shd8c53cba, 32'shd8c67a76, 
               32'shd8c7b838, 32'shd8c8f601, 32'shd8ca33cf, 32'shd8cb71a3, 32'shd8ccaf7e, 32'shd8cded5e, 32'shd8cf2b45, 32'shd8d06931, 
               32'shd8d1a724, 32'shd8d2e51c, 32'shd8d4231b, 32'shd8d56120, 32'shd8d69f2a, 32'shd8d7dd3b, 32'shd8d91b52, 32'shd8da596f, 
               32'shd8db9792, 32'shd8dcd5bb, 32'shd8de13ea, 32'shd8df521f, 32'shd8e0905a, 32'shd8e1ce9b, 32'shd8e30ce2, 32'shd8e44b2f, 
               32'shd8e58982, 32'shd8e6c7db, 32'shd8e8063a, 32'shd8e944a0, 32'shd8ea830b, 32'shd8ebc17c, 32'shd8ecfff4, 32'shd8ee3e71, 
               32'shd8ef7cf4, 32'shd8f0bb7e, 32'shd8f1fa0d, 32'shd8f338a3, 32'shd8f4773e, 32'shd8f5b5df, 32'shd8f6f487, 32'shd8f83335, 
               32'shd8f971e8, 32'shd8fab0a2, 32'shd8fbef61, 32'shd8fd2e27, 32'shd8fe6cf2, 32'shd8ffabc4, 32'shd900ea9c, 32'shd9022979, 
               32'shd903685d, 32'shd904a747, 32'shd905e636, 32'shd907252c, 32'shd9086428, 32'shd909a32a, 32'shd90ae231, 32'shd90c213f, 
               32'shd90d6053, 32'shd90e9f6d, 32'shd90fde8c, 32'shd9111db2, 32'shd9125cde, 32'shd9139c10, 32'shd914db47, 32'shd9161a85, 
               32'shd91759c9, 32'shd9189913, 32'shd919d863, 32'shd91b17b8, 32'shd91c5714, 32'shd91d9676, 32'shd91ed5de, 32'shd920154b, 
               32'shd92154bf, 32'shd9229439, 32'shd923d3b9, 32'shd925133e, 32'shd92652ca, 32'shd927925c, 32'shd928d1f4, 32'shd92a1191, 
               32'shd92b5135, 32'shd92c90df, 32'shd92dd08e, 32'shd92f1044, 32'shd9305000, 32'shd9318fc1, 32'shd932cf89, 32'shd9340f56, 
               32'shd9354f2a, 32'shd9368f04, 32'shd937cee3, 32'shd9390ec9, 32'shd93a4eb4, 32'shd93b8ea6, 32'shd93cce9d, 32'shd93e0e9b, 
               32'shd93f4e9e, 32'shd9408ea7, 32'shd941ceb7, 32'shd9430ecc, 32'shd9444ee7, 32'shd9458f09, 32'shd946cf30, 32'shd9480f5d, 
               32'shd9494f90, 32'shd94a8fca, 32'shd94bd009, 32'shd94d104e, 32'shd94e5099, 32'shd94f90ea, 32'shd950d141, 32'shd952119e, 
               32'shd9535201, 32'shd954926a, 32'shd955d2d9, 32'shd957134d, 32'shd95853c8, 32'shd9599449, 32'shd95ad4d0, 32'shd95c155c, 
               32'shd95d55ef, 32'shd95e9688, 32'shd95fd726, 32'shd96117cb, 32'shd9625875, 32'shd9639926, 32'shd964d9dc, 32'shd9661a98, 
               32'shd9675b5a, 32'shd9689c23, 32'shd969dcf1, 32'shd96b1dc5, 32'shd96c5e9f, 32'shd96d9f7f, 32'shd96ee065, 32'shd9702151, 
               32'shd9716243, 32'shd972a33b, 32'shd973e438, 32'shd975253c, 32'shd9766646, 32'shd977a755, 32'shd978e86b, 32'shd97a2986, 
               32'shd97b6aa8, 32'shd97cabcf, 32'shd97decfd, 32'shd97f2e30, 32'shd9806f69, 32'shd981b0a8, 32'shd982f1ed, 32'shd9843338, 
               32'shd9857489, 32'shd986b5e0, 32'shd987f73d, 32'shd989389f, 32'shd98a7a08, 32'shd98bbb77, 32'shd98cfceb, 32'shd98e3e66, 
               32'shd98f7fe6, 32'shd990c16c, 32'shd99202f8, 32'shd993448b, 32'shd9948623, 32'shd995c7c1, 32'shd9970965, 32'shd9984b0e, 
               32'shd9998cbe, 32'shd99ace74, 32'shd99c102f, 32'shd99d51f1, 32'shd99e93b8, 32'shd99fd586, 32'shd9a11759, 32'shd9a25932, 
               32'shd9a39b11, 32'shd9a4dcf6, 32'shd9a61ee1, 32'shd9a760d2, 32'shd9a8a2c9, 32'shd9a9e4c6, 32'shd9ab26c8, 32'shd9ac68d1, 
               32'shd9adaadf, 32'shd9aeecf4, 32'shd9b02f0e, 32'shd9b1712e, 32'shd9b2b354, 32'shd9b3f580, 32'shd9b537b2, 32'shd9b679ea, 
               32'shd9b7bc27, 32'shd9b8fe6b, 32'shd9ba40b5, 32'shd9bb8304, 32'shd9bcc559, 32'shd9be07b4, 32'shd9bf4a15, 32'shd9c08c7c, 
               32'shd9c1cee9, 32'shd9c3115c, 32'shd9c453d5, 32'shd9c59653, 32'shd9c6d8d8, 32'shd9c81b62, 32'shd9c95df3, 32'shd9caa089, 
               32'shd9cbe325, 32'shd9cd25c7, 32'shd9ce686e, 32'shd9cfab1c, 32'shd9d0edd0, 32'shd9d23089, 32'shd9d37349, 32'shd9d4b60e, 
               32'shd9d5f8d9, 32'shd9d73baa, 32'shd9d87e81, 32'shd9d9c15e, 32'shd9db0441, 32'shd9dc4729, 32'shd9dd8a18, 32'shd9decd0c, 
               32'shd9e01006, 32'shd9e15306, 32'shd9e2960c, 32'shd9e3d918, 32'shd9e51c2a, 32'shd9e65f42, 32'shd9e7a25f, 32'shd9e8e582, 
               32'shd9ea28ac, 32'shd9eb6bdb, 32'shd9ecaf10, 32'shd9edf24b, 32'shd9ef358b, 32'shd9f078d2, 32'shd9f1bc1e, 32'shd9f2ff71, 
               32'shd9f442c9, 32'shd9f58627, 32'shd9f6c98b, 32'shd9f80cf5, 32'shd9f95064, 32'shd9fa93da, 32'shd9fbd755, 32'shd9fd1ad6, 
               32'shd9fe5e5e, 32'shd9ffa1eb, 32'shda00e57d, 32'shda022916, 32'shda036cb5, 32'shda04b059, 32'shda05f403, 32'shda0737b3, 
               32'shda087b69, 32'shda09bf25, 32'shda0b02e7, 32'shda0c46af, 32'shda0d8a7c, 32'shda0ece4f, 32'shda101228, 32'shda115607, 
               32'shda1299ec, 32'shda13ddd7, 32'shda1521c7, 32'shda1665be, 32'shda17a9ba, 32'shda18edbc, 32'shda1a31c4, 32'shda1b75d1, 
               32'shda1cb9e5, 32'shda1dfdfe, 32'shda1f421e, 32'shda208643, 32'shda21ca6e, 32'shda230e9e, 32'shda2452d5, 32'shda259711, 
               32'shda26db54, 32'shda281f9c, 32'shda2963ea, 32'shda2aa83e, 32'shda2bec97, 32'shda2d30f7, 32'shda2e755c, 32'shda2fb9c7, 
               32'shda30fe38, 32'shda3242af, 32'shda33872c, 32'shda34cbae, 32'shda361036, 32'shda3754c4, 32'shda389958, 32'shda39ddf2, 
               32'shda3b2292, 32'shda3c6737, 32'shda3dabe2, 32'shda3ef093, 32'shda40354a, 32'shda417a07, 32'shda42beca, 32'shda440392, 
               32'shda454860, 32'shda468d34, 32'shda47d20e, 32'shda4916ed, 32'shda4a5bd3, 32'shda4ba0be, 32'shda4ce5af, 32'shda4e2aa6, 
               32'shda4f6fa3, 32'shda50b4a5, 32'shda51f9ae, 32'shda533ebc, 32'shda5483d0, 32'shda55c8e9, 32'shda570e09, 32'shda58532e, 
               32'shda599859, 32'shda5add8a, 32'shda5c22c1, 32'shda5d67fe, 32'shda5ead40, 32'shda5ff288, 32'shda6137d6, 32'shda627d2a, 
               32'shda63c284, 32'shda6507e3, 32'shda664d48, 32'shda6792b3, 32'shda68d824, 32'shda6a1d9b, 32'shda6b6317, 32'shda6ca899, 
               32'shda6dee21, 32'shda6f33af, 32'shda707942, 32'shda71bedc, 32'shda73047b, 32'shda744a20, 32'shda758fcb, 32'shda76d57b, 
               32'shda781b31, 32'shda7960ed, 32'shda7aa6af, 32'shda7bec77, 32'shda7d3244, 32'shda7e7818, 32'shda7fbdf1, 32'shda8103cf, 
               32'shda8249b4, 32'shda838f9e, 32'shda84d58f, 32'shda861b84, 32'shda876180, 32'shda88a782, 32'shda89ed89, 32'shda8b3396, 
               32'shda8c79a9, 32'shda8dbfc1, 32'shda8f05e0, 32'shda904c04, 32'shda91922e, 32'shda92d85d, 32'shda941e93, 32'shda9564ce, 
               32'shda96ab0f, 32'shda97f156, 32'shda9937a2, 32'shda9a7df5, 32'shda9bc44d, 32'shda9d0aab, 32'shda9e510e, 32'shda9f9778, 
               32'shdaa0dde7, 32'shdaa2245c, 32'shdaa36ad6, 32'shdaa4b157, 32'shdaa5f7dd, 32'shdaa73e69, 32'shdaa884fa, 32'shdaa9cb92, 
               32'shdaab122f, 32'shdaac58d2, 32'shdaad9f7b, 32'shdaaee629, 32'shdab02cdd, 32'shdab17397, 32'shdab2ba57, 32'shdab4011d, 
               32'shdab547e8, 32'shdab68eb9, 32'shdab7d590, 32'shdab91c6c, 32'shdaba634e, 32'shdabbaa36, 32'shdabcf124, 32'shdabe3818, 
               32'shdabf7f11, 32'shdac0c610, 32'shdac20d15, 32'shdac3541f, 32'shdac49b2f, 32'shdac5e245, 32'shdac72961, 32'shdac87082, 
               32'shdac9b7a9, 32'shdacafed6, 32'shdacc4609, 32'shdacd8d41, 32'shdaced47f, 32'shdad01bc3, 32'shdad1630d, 32'shdad2aa5c, 
               32'shdad3f1b1, 32'shdad5390c, 32'shdad6806d, 32'shdad7c7d3, 32'shdad90f3f, 32'shdada56b0, 32'shdadb9e28, 32'shdadce5a5, 
               32'shdade2d28, 32'shdadf74b1, 32'shdae0bc3f, 32'shdae203d3, 32'shdae34b6d, 32'shdae4930c, 32'shdae5dab2, 32'shdae7225c, 
               32'shdae86a0d, 32'shdae9b1c4, 32'shdaeaf980, 32'shdaec4141, 32'shdaed8909, 32'shdaeed0d6, 32'shdaf018a9, 32'shdaf16082, 
               32'shdaf2a860, 32'shdaf3f045, 32'shdaf5382e, 32'shdaf6801e, 32'shdaf7c813, 32'shdaf9100e, 32'shdafa580f, 32'shdafba015, 
               32'shdafce821, 32'shdafe3033, 32'shdaff784b, 32'shdb00c068, 32'shdb02088b, 32'shdb0350b4, 32'shdb0498e2, 32'shdb05e116, 
               32'shdb072950, 32'shdb08718f, 32'shdb09b9d4, 32'shdb0b021f, 32'shdb0c4a70, 32'shdb0d92c6, 32'shdb0edb22, 32'shdb102383, 
               32'shdb116beb, 32'shdb12b458, 32'shdb13fccb, 32'shdb154543, 32'shdb168dc1, 32'shdb17d645, 32'shdb191ece, 32'shdb1a675e, 
               32'shdb1baff2, 32'shdb1cf88d, 32'shdb1e412d, 32'shdb1f89d3, 32'shdb20d27f, 32'shdb221b30, 32'shdb2363e7, 32'shdb24aca4, 
               32'shdb25f566, 32'shdb273e2e, 32'shdb2886fc, 32'shdb29cfcf, 32'shdb2b18a9, 32'shdb2c6187, 32'shdb2daa6c, 32'shdb2ef356, 
               32'shdb303c46, 32'shdb31853b, 32'shdb32ce36, 32'shdb341737, 32'shdb35603e, 32'shdb36a94a, 32'shdb37f25c, 32'shdb393b73, 
               32'shdb3a8491, 32'shdb3bcdb3, 32'shdb3d16dc, 32'shdb3e600a, 32'shdb3fa93e, 32'shdb40f278, 32'shdb423bb7, 32'shdb4384fc, 
               32'shdb44ce46, 32'shdb461797, 32'shdb4760ec, 32'shdb48aa48, 32'shdb49f3a9, 32'shdb4b3d10, 32'shdb4c867d, 32'shdb4dcfef, 
               32'shdb4f1967, 32'shdb5062e4, 32'shdb51ac67, 32'shdb52f5f0, 32'shdb543f7e, 32'shdb558913, 32'shdb56d2ac, 32'shdb581c4c, 
               32'shdb5965f1, 32'shdb5aaf9c, 32'shdb5bf94c, 32'shdb5d4302, 32'shdb5e8cbe, 32'shdb5fd67f, 32'shdb612046, 32'shdb626a13, 
               32'shdb63b3e5, 32'shdb64fdbd, 32'shdb66479b, 32'shdb67917e, 32'shdb68db67, 32'shdb6a2555, 32'shdb6b6f49, 32'shdb6cb943, 
               32'shdb6e0342, 32'shdb6f4d48, 32'shdb709752, 32'shdb71e163, 32'shdb732b79, 32'shdb747594, 32'shdb75bfb5, 32'shdb7709dc, 
               32'shdb785409, 32'shdb799e3b, 32'shdb7ae873, 32'shdb7c32b0, 32'shdb7d7cf3, 32'shdb7ec73c, 32'shdb80118a, 32'shdb815bde, 
               32'shdb82a638, 32'shdb83f097, 32'shdb853afc, 32'shdb868566, 32'shdb87cfd6, 32'shdb891a4c, 32'shdb8a64c7, 32'shdb8baf48, 
               32'shdb8cf9cf, 32'shdb8e445b, 32'shdb8f8eed, 32'shdb90d984, 32'shdb922421, 32'shdb936ec4, 32'shdb94b96c, 32'shdb96041a, 
               32'shdb974ece, 32'shdb989987, 32'shdb99e445, 32'shdb9b2f0a, 32'shdb9c79d4, 32'shdb9dc4a3, 32'shdb9f0f78, 32'shdba05a53, 
               32'shdba1a534, 32'shdba2f01a, 32'shdba43b05, 32'shdba585f7, 32'shdba6d0ed, 32'shdba81bea, 32'shdba966ec, 32'shdbaab1f3, 
               32'shdbabfd01, 32'shdbad4814, 32'shdbae932c, 32'shdbafde4a, 32'shdbb1296e, 32'shdbb27497, 32'shdbb3bfc6, 32'shdbb50afa, 
               32'shdbb65634, 32'shdbb7a174, 32'shdbb8ecb9, 32'shdbba3804, 32'shdbbb8354, 32'shdbbcceaa, 32'shdbbe1a06, 32'shdbbf6567, 
               32'shdbc0b0ce, 32'shdbc1fc3a, 32'shdbc347ac, 32'shdbc49324, 32'shdbc5dea1, 32'shdbc72a24, 32'shdbc875ac, 32'shdbc9c13a, 
               32'shdbcb0cce, 32'shdbcc5867, 32'shdbcda405, 32'shdbceefaa, 32'shdbd03b53, 32'shdbd18703, 32'shdbd2d2b8, 32'shdbd41e72, 
               32'shdbd56a32, 32'shdbd6b5f8, 32'shdbd801c3, 32'shdbd94d94, 32'shdbda996b, 32'shdbdbe547, 32'shdbdd3128, 32'shdbde7d10, 
               32'shdbdfc8fc, 32'shdbe114ef, 32'shdbe260e6, 32'shdbe3ace4, 32'shdbe4f8e7, 32'shdbe644ef, 32'shdbe790fe, 32'shdbe8dd11, 
               32'shdbea292b, 32'shdbeb7549, 32'shdbecc16e, 32'shdbee0d98, 32'shdbef59c7, 32'shdbf0a5fc, 32'shdbf1f237, 32'shdbf33e77, 
               32'shdbf48abd, 32'shdbf5d708, 32'shdbf72359, 32'shdbf86fb0, 32'shdbf9bc0c, 32'shdbfb086d, 32'shdbfc54d4, 32'shdbfda141, 
               32'shdbfeedb3, 32'shdc003a2b, 32'shdc0186a8, 32'shdc02d32b, 32'shdc041fb4, 32'shdc056c42, 32'shdc06b8d5, 32'shdc08056e, 
               32'shdc09520d, 32'shdc0a9eb1, 32'shdc0beb5b, 32'shdc0d380a, 32'shdc0e84bf, 32'shdc0fd179, 32'shdc111e39, 32'shdc126afe, 
               32'shdc13b7c9, 32'shdc15049a, 32'shdc165170, 32'shdc179e4c, 32'shdc18eb2d, 32'shdc1a3813, 32'shdc1b8500, 32'shdc1cd1f1, 
               32'shdc1e1ee9, 32'shdc1f6be5, 32'shdc20b8e8, 32'shdc2205f0, 32'shdc2352fd, 32'shdc24a010, 32'shdc25ed28, 32'shdc273a46, 
               32'shdc28876a, 32'shdc29d493, 32'shdc2b21c1, 32'shdc2c6ef5, 32'shdc2dbc2f, 32'shdc2f096e, 32'shdc3056b3, 32'shdc31a3fd, 
               32'shdc32f14d, 32'shdc343ea2, 32'shdc358bfd, 32'shdc36d95d, 32'shdc3826c3, 32'shdc39742e, 32'shdc3ac19f, 32'shdc3c0f15, 
               32'shdc3d5c91, 32'shdc3eaa12, 32'shdc3ff799, 32'shdc414526, 32'shdc4292b8, 32'shdc43e04f, 32'shdc452dec, 32'shdc467b8e, 
               32'shdc47c936, 32'shdc4916e4, 32'shdc4a6497, 32'shdc4bb24f, 32'shdc4d000d, 32'shdc4e4dd1, 32'shdc4f9b9a, 32'shdc50e968, 
               32'shdc52373c, 32'shdc538516, 32'shdc54d2f5, 32'shdc5620d9, 32'shdc576ec3, 32'shdc58bcb3, 32'shdc5a0aa8, 32'shdc5b58a2, 
               32'shdc5ca6a2, 32'shdc5df4a7, 32'shdc5f42b2, 32'shdc6090c3, 32'shdc61ded9, 32'shdc632cf4, 32'shdc647b15, 32'shdc65c93c, 
               32'shdc671768, 32'shdc686599, 32'shdc69b3d0, 32'shdc6b020c, 32'shdc6c504e, 32'shdc6d9e96, 32'shdc6eece2, 32'shdc703b35, 
               32'shdc71898d, 32'shdc72d7ea, 32'shdc74264d, 32'shdc7574b5, 32'shdc76c323, 32'shdc781196, 32'shdc79600f, 32'shdc7aae8d, 
               32'shdc7bfd11, 32'shdc7d4b9a, 32'shdc7e9a28, 32'shdc7fe8bc, 32'shdc813756, 32'shdc8285f5, 32'shdc83d49a, 32'shdc852344, 
               32'shdc8671f3, 32'shdc87c0a8, 32'shdc890f62, 32'shdc8a5e22, 32'shdc8bace8, 32'shdc8cfbb2, 32'shdc8e4a83, 32'shdc8f9958, 
               32'shdc90e834, 32'shdc923714, 32'shdc9385fa, 32'shdc94d4e6, 32'shdc9623d7, 32'shdc9772ce, 32'shdc98c1ca, 32'shdc9a10cb, 
               32'shdc9b5fd2, 32'shdc9caede, 32'shdc9dfdf0, 32'shdc9f4d07, 32'shdca09c24, 32'shdca1eb46, 32'shdca33a6e, 32'shdca4899b, 
               32'shdca5d8cd, 32'shdca72805, 32'shdca87743, 32'shdca9c686, 32'shdcab15ce, 32'shdcac651c, 32'shdcadb46f, 32'shdcaf03c8, 
               32'shdcb05326, 32'shdcb1a28a, 32'shdcb2f1f3, 32'shdcb44161, 32'shdcb590d5, 32'shdcb6e04e, 32'shdcb82fcd, 32'shdcb97f51, 
               32'shdcbacedb, 32'shdcbc1e6a, 32'shdcbd6dff, 32'shdcbebd99, 32'shdcc00d38, 32'shdcc15cdd, 32'shdcc2ac87, 32'shdcc3fc37, 
               32'shdcc54bec, 32'shdcc69ba7, 32'shdcc7eb67, 32'shdcc93b2c, 32'shdcca8af7, 32'shdccbdac7, 32'shdccd2a9d, 32'shdcce7a78, 
               32'shdccfca59, 32'shdcd11a3f, 32'shdcd26a2a, 32'shdcd3ba1b, 32'shdcd50a12, 32'shdcd65a0d, 32'shdcd7aa0e, 32'shdcd8fa15, 
               32'shdcda4a21, 32'shdcdb9a32, 32'shdcdcea49, 32'shdcde3a66, 32'shdcdf8a87, 32'shdce0daae, 32'shdce22adb, 32'shdce37b0d, 
               32'shdce4cb44, 32'shdce61b81, 32'shdce76bc3, 32'shdce8bc0b, 32'shdcea0c58, 32'shdceb5caa, 32'shdcecad02, 32'shdcedfd5f, 
               32'shdcef4dc2, 32'shdcf09e2a, 32'shdcf1ee97, 32'shdcf33f0a, 32'shdcf48f82, 32'shdcf5e000, 32'shdcf73083, 32'shdcf8810b, 
               32'shdcf9d199, 32'shdcfb222c, 32'shdcfc72c5, 32'shdcfdc363, 32'shdcff1407, 32'shdd0064af, 32'shdd01b55e, 32'shdd030611, 
               32'shdd0456ca, 32'shdd05a789, 32'shdd06f84d, 32'shdd084916, 32'shdd0999e4, 32'shdd0aeab9, 32'shdd0c3b92, 32'shdd0d8c71, 
               32'shdd0edd55, 32'shdd102e3e, 32'shdd117f2d, 32'shdd12d022, 32'shdd14211b, 32'shdd15721b, 32'shdd16c31f, 32'shdd181429, 
               32'shdd196538, 32'shdd1ab64d, 32'shdd1c0767, 32'shdd1d5886, 32'shdd1ea9ab, 32'shdd1ffad5, 32'shdd214c05, 32'shdd229d3a, 
               32'shdd23ee74, 32'shdd253fb4, 32'shdd2690f9, 32'shdd27e243, 32'shdd293393, 32'shdd2a84e8, 32'shdd2bd643, 32'shdd2d27a3, 
               32'shdd2e7908, 32'shdd2fca73, 32'shdd311be3, 32'shdd326d58, 32'shdd33bed3, 32'shdd351053, 32'shdd3661d8, 32'shdd37b363, 
               32'shdd3904f4, 32'shdd3a5689, 32'shdd3ba824, 32'shdd3cf9c4, 32'shdd3e4b6a, 32'shdd3f9d15, 32'shdd40eec5, 32'shdd42407b, 
               32'shdd439236, 32'shdd44e3f7, 32'shdd4635bd, 32'shdd478788, 32'shdd48d958, 32'shdd4a2b2e, 32'shdd4b7d09, 32'shdd4cceea, 
               32'shdd4e20d0, 32'shdd4f72bb, 32'shdd50c4ac, 32'shdd5216a2, 32'shdd53689d, 32'shdd54ba9e, 32'shdd560ca4, 32'shdd575eaf, 
               32'shdd58b0c0, 32'shdd5a02d6, 32'shdd5b54f1, 32'shdd5ca712, 32'shdd5df938, 32'shdd5f4b64, 32'shdd609d94, 32'shdd61efcb, 
               32'shdd634206, 32'shdd649447, 32'shdd65e68d, 32'shdd6738d8, 32'shdd688b29, 32'shdd69dd7f, 32'shdd6b2fdb, 32'shdd6c823b, 
               32'shdd6dd4a2, 32'shdd6f270d, 32'shdd70797e, 32'shdd71cbf4, 32'shdd731e6f, 32'shdd7470f0, 32'shdd75c376, 32'shdd771602, 
               32'shdd786892, 32'shdd79bb29, 32'shdd7b0dc4, 32'shdd7c6065, 32'shdd7db30b, 32'shdd7f05b6, 32'shdd805867, 32'shdd81ab1d, 
               32'shdd82fdd8, 32'shdd845099, 32'shdd85a35f, 32'shdd86f62a, 32'shdd8848fb, 32'shdd899bd1, 32'shdd8aeeac, 32'shdd8c418c, 
               32'shdd8d9472, 32'shdd8ee75d, 32'shdd903a4e, 32'shdd918d44, 32'shdd92e03f, 32'shdd94333f, 32'shdd958645, 32'shdd96d950, 
               32'shdd982c60, 32'shdd997f76, 32'shdd9ad291, 32'shdd9c25b1, 32'shdd9d78d7, 32'shdd9ecc01, 32'shdda01f32, 32'shdda17267, 
               32'shdda2c5a2, 32'shdda418e2, 32'shdda56c27, 32'shdda6bf72, 32'shdda812c2, 32'shdda96617, 32'shddaab972, 32'shddac0cd1, 
               32'shddad6036, 32'shddaeb3a1, 32'shddb00711, 32'shddb15a86, 32'shddb2ae00, 32'shddb4017f, 32'shddb55504, 32'shddb6a88f, 
               32'shddb7fc1e, 32'shddb94fb3, 32'shddbaa34d, 32'shddbbf6ec, 32'shddbd4a91, 32'shddbe9e3a, 32'shddbff1ea, 32'shddc1459e, 
               32'shddc29958, 32'shddc3ed17, 32'shddc540db, 32'shddc694a5, 32'shddc7e873, 32'shddc93c48, 32'shddca9021, 32'shddcbe400, 
               32'shddcd37e4, 32'shddce8bcd, 32'shddcfdfbb, 32'shddd133af, 32'shddd287a8, 32'shddd3dba6, 32'shddd52faa, 32'shddd683b3, 
               32'shddd7d7c1, 32'shddd92bd4, 32'shddda7fed, 32'shdddbd40b, 32'shdddd282e, 32'shddde7c56, 32'shdddfd084, 32'shdde124b7, 
               32'shdde278ef, 32'shdde3cd2d, 32'shdde5216f, 32'shdde675b7, 32'shdde7ca05, 32'shdde91e57, 32'shddea72af, 32'shddebc70c, 
               32'shdded1b6e, 32'shddee6fd6, 32'shddefc443, 32'shddf118b5, 32'shddf26d2c, 32'shddf3c1a9, 32'shddf5162a, 32'shddf66ab1, 
               32'shddf7bf3e, 32'shddf913cf, 32'shddfa6866, 32'shddfbbd02, 32'shddfd11a3, 32'shddfe664a, 32'shddffbaf6, 32'shde010fa7, 
               32'shde02645d, 32'shde03b919, 32'shde050dd9, 32'shde06629f, 32'shde07b76b, 32'shde090c3b, 32'shde0a6111, 32'shde0bb5ec, 
               32'shde0d0acc, 32'shde0e5fb1, 32'shde0fb49c, 32'shde11098c, 32'shde125e81, 32'shde13b37b, 32'shde15087b, 32'shde165d80, 
               32'shde17b28a, 32'shde190799, 32'shde1a5cad, 32'shde1bb1c7, 32'shde1d06e6, 32'shde1e5c0a, 32'shde1fb134, 32'shde210662, 
               32'shde225b96, 32'shde23b0cf, 32'shde25060e, 32'shde265b51, 32'shde27b09a, 32'shde2905e8, 32'shde2a5b3b, 32'shde2bb093, 
               32'shde2d05f1, 32'shde2e5b54, 32'shde2fb0bc, 32'shde310629, 32'shde325b9b, 32'shde33b113, 32'shde350690, 32'shde365c12, 
               32'shde37b199, 32'shde390726, 32'shde3a5cb8, 32'shde3bb24f, 32'shde3d07eb, 32'shde3e5d8c, 32'shde3fb333, 32'shde4108de, 
               32'shde425e8f, 32'shde43b446, 32'shde450a01, 32'shde465fc2, 32'shde47b587, 32'shde490b52, 32'shde4a6122, 32'shde4bb6f8, 
               32'shde4d0cd2, 32'shde4e62b2, 32'shde4fb897, 32'shde510e81, 32'shde526471, 32'shde53ba65, 32'shde55105f, 32'shde56665e, 
               32'shde57bc62, 32'shde59126b, 32'shde5a687a, 32'shde5bbe8d, 32'shde5d14a6, 32'shde5e6ac4, 32'shde5fc0e8, 32'shde611710, 
               32'shde626d3e, 32'shde63c371, 32'shde6519a9, 32'shde666fe6, 32'shde67c628, 32'shde691c70, 32'shde6a72bc, 32'shde6bc90e, 
               32'shde6d1f65, 32'shde6e75c2, 32'shde6fcc23, 32'shde71228a, 32'shde7278f5, 32'shde73cf66, 32'shde7525dc, 32'shde767c58, 
               32'shde77d2d8, 32'shde79295e, 32'shde7a7fe9, 32'shde7bd679, 32'shde7d2d0e, 32'shde7e83a8, 32'shde7fda48, 32'shde8130ec, 
               32'shde828796, 32'shde83de45, 32'shde8534f9, 32'shde868bb2, 32'shde87e271, 32'shde893935, 32'shde8a8ffd, 32'shde8be6cb, 
               32'shde8d3d9e, 32'shde8e9477, 32'shde8feb54, 32'shde914237, 32'shde92991e, 32'shde93f00b, 32'shde9546fd, 32'shde969df5, 
               32'shde97f4f1, 32'shde994bf2, 32'shde9aa2f9, 32'shde9bfa05, 32'shde9d5116, 32'shde9ea82c, 32'shde9fff47, 32'shdea15668, 
               32'shdea2ad8d, 32'shdea404b8, 32'shdea55be8, 32'shdea6b31d, 32'shdea80a57, 32'shdea96196, 32'shdeaab8da, 32'shdeac1024, 
               32'shdead6773, 32'shdeaebec6, 32'shdeb0161f, 32'shdeb16d7d, 32'shdeb2c4e1, 32'shdeb41c49, 32'shdeb573b7, 32'shdeb6cb29, 
               32'shdeb822a1, 32'shdeb97a1e, 32'shdebad1a0, 32'shdebc2927, 32'shdebd80b3, 32'shdebed845, 32'shdec02fdb, 32'shdec18777, 
               32'shdec2df18, 32'shdec436be, 32'shdec58e69, 32'shdec6e619, 32'shdec83dce, 32'shdec99589, 32'shdecaed48, 32'shdecc450d, 
               32'shdecd9cd7, 32'shdecef4a6, 32'shded04c7a, 32'shded1a453, 32'shded2fc31, 32'shded45414, 32'shded5abfd, 32'shded703eb, 
               32'shded85bdd, 32'shded9b3d5, 32'shdedb0bd2, 32'shdedc63d4, 32'shdeddbbdb, 32'shdedf13e8, 32'shdee06bf9, 32'shdee1c40f, 
               32'shdee31c2b, 32'shdee4744c, 32'shdee5cc72, 32'shdee7249c, 32'shdee87ccc, 32'shdee9d502, 32'shdeeb2d3c, 32'shdeec857b, 
               32'shdeedddc0, 32'shdeef3609, 32'shdef08e58, 32'shdef1e6ab, 32'shdef33f04, 32'shdef49762, 32'shdef5efc5, 32'shdef7482d, 
               32'shdef8a09b, 32'shdef9f90d, 32'shdefb5184, 32'shdefcaa01, 32'shdefe0282, 32'shdeff5b09, 32'shdf00b395, 32'shdf020c26, 
               32'shdf0364bc, 32'shdf04bd57, 32'shdf0615f7, 32'shdf076e9c, 32'shdf08c746, 32'shdf0a1ff5, 32'shdf0b78aa, 32'shdf0cd163, 
               32'shdf0e2a22, 32'shdf0f82e6, 32'shdf10dbaf, 32'shdf12347c, 32'shdf138d4f, 32'shdf14e627, 32'shdf163f04, 32'shdf1797e7, 
               32'shdf18f0ce, 32'shdf1a49ba, 32'shdf1ba2ab, 32'shdf1cfba2, 32'shdf1e549d, 32'shdf1fad9e, 32'shdf2106a4, 32'shdf225fae, 
               32'shdf23b8be, 32'shdf2511d3, 32'shdf266aed, 32'shdf27c40c, 32'shdf291d30, 32'shdf2a7659, 32'shdf2bcf87, 32'shdf2d28bb, 
               32'shdf2e81f3, 32'shdf2fdb30, 32'shdf313473, 32'shdf328dba, 32'shdf33e707, 32'shdf354058, 32'shdf3699af, 32'shdf37f30b, 
               32'shdf394c6b, 32'shdf3aa5d1, 32'shdf3bff3c, 32'shdf3d58ac, 32'shdf3eb221, 32'shdf400b9b, 32'shdf41651a, 32'shdf42be9e, 
               32'shdf441828, 32'shdf4571b6, 32'shdf46cb49, 32'shdf4824e1, 32'shdf497e7f, 32'shdf4ad821, 32'shdf4c31c9, 32'shdf4d8b75, 
               32'shdf4ee527, 32'shdf503edd, 32'shdf519899, 32'shdf52f25a, 32'shdf544c1f, 32'shdf55a5ea, 32'shdf56ffba, 32'shdf58598f, 
               32'shdf59b369, 32'shdf5b0d48, 32'shdf5c672b, 32'shdf5dc114, 32'shdf5f1b02, 32'shdf6074f5, 32'shdf61ceee, 32'shdf6328eb, 
               32'shdf6482ed, 32'shdf65dcf4, 32'shdf673700, 32'shdf689111, 32'shdf69eb27, 32'shdf6b4543, 32'shdf6c9f63, 32'shdf6df988, 
               32'shdf6f53b3, 32'shdf70ade2, 32'shdf720816, 32'shdf736250, 32'shdf74bc8e, 32'shdf7616d2, 32'shdf77711a, 32'shdf78cb67, 
               32'shdf7a25ba, 32'shdf7b8011, 32'shdf7cda6e, 32'shdf7e34cf, 32'shdf7f8f36, 32'shdf80e9a2, 32'shdf824412, 32'shdf839e88, 
               32'shdf84f902, 32'shdf865382, 32'shdf87ae06, 32'shdf890890, 32'shdf8a631f, 32'shdf8bbdb2, 32'shdf8d184b, 32'shdf8e72e8, 
               32'shdf8fcd8b, 32'shdf912833, 32'shdf9282df, 32'shdf93dd91, 32'shdf953848, 32'shdf969303, 32'shdf97edc4, 32'shdf99488a, 
               32'shdf9aa354, 32'shdf9bfe24, 32'shdf9d58f8, 32'shdf9eb3d2, 32'shdfa00eb1, 32'shdfa16994, 32'shdfa2c47d, 32'shdfa41f6a, 
               32'shdfa57a5d, 32'shdfa6d554, 32'shdfa83051, 32'shdfa98b53, 32'shdfaae659, 32'shdfac4165, 32'shdfad9c75, 32'shdfaef78b, 
               32'shdfb052a5, 32'shdfb1adc4, 32'shdfb308e9, 32'shdfb46412, 32'shdfb5bf41, 32'shdfb71a74, 32'shdfb875ac, 32'shdfb9d0ea, 
               32'shdfbb2c2c, 32'shdfbc8773, 32'shdfbde2bf, 32'shdfbf3e11, 32'shdfc09967, 32'shdfc1f4c2, 32'shdfc35022, 32'shdfc4ab87, 
               32'shdfc606f1, 32'shdfc76260, 32'shdfc8bdd4, 32'shdfca194d, 32'shdfcb74cb, 32'shdfccd04e, 32'shdfce2bd6, 32'shdfcf8763, 
               32'shdfd0e2f5, 32'shdfd23e8c, 32'shdfd39a27, 32'shdfd4f5c8, 32'shdfd6516e, 32'shdfd7ad18, 32'shdfd908c8, 32'shdfda647d, 
               32'shdfdbc036, 32'shdfdd1bf5, 32'shdfde77b8, 32'shdfdfd380, 32'shdfe12f4e, 32'shdfe28b20, 32'shdfe3e6f7, 32'shdfe542d3, 
               32'shdfe69eb4, 32'shdfe7fa9b, 32'shdfe95686, 32'shdfeab276, 32'shdfec0e6a, 32'shdfed6a64, 32'shdfeec663, 32'shdff02267, 
               32'shdff17e70, 32'shdff2da7d, 32'shdff43690, 32'shdff592a7, 32'shdff6eec4, 32'shdff84ae5, 32'shdff9a70c, 32'shdffb0337, 
               32'shdffc5f67, 32'shdffdbb9c, 32'shdfff17d7, 32'she0007416, 32'she001d05a, 32'she0032ca2, 32'she00488f0, 32'she005e543, 
               32'she007419b, 32'she0089df7, 32'she009fa59, 32'she00b56bf, 32'she00cb32b, 32'she00e0f9b, 32'she00f6c11, 32'she010c88b, 
               32'she012250a, 32'she013818e, 32'she014de17, 32'she0163aa5, 32'she0179738, 32'she018f3cf, 32'she01a506c, 32'she01bad0e, 
               32'she01d09b4, 32'she01e6660, 32'she01fc310, 32'she0211fc5, 32'she0227c7f, 32'she023d93e, 32'she0253602, 32'she02692cb, 
               32'she027ef99, 32'she0294c6c, 32'she02aa943, 32'she02c0620, 32'she02d6301, 32'she02ebfe8, 32'she0301cd3, 32'she03179c3, 
               32'she032d6b8, 32'she03433b2, 32'she03590b1, 32'she036edb5, 32'she0384abe, 32'she039a7cb, 32'she03b04de, 32'she03c61f5, 
               32'she03dbf11, 32'she03f1c33, 32'she0407959, 32'she041d684, 32'she04333b3, 32'she04490e8, 32'she045ee22, 32'she0474b60, 
               32'she048a8a4, 32'she04a05ec, 32'she04b6339, 32'she04cc08c, 32'she04e1de3, 32'she04f7b3e, 32'she050d89f, 32'she0523605, 
               32'she053936f, 32'she054f0df, 32'she0564e53, 32'she057abcc, 32'she059094a, 32'she05a66cd, 32'she05bc455, 32'she05d21e2, 
               32'she05e7f74, 32'she05fdd0a, 32'she0613aa5, 32'she0629846, 32'she063f5eb, 32'she0655395, 32'she066b144, 32'she0680ef7, 
               32'she0696cb0, 32'she06aca6d, 32'she06c2830, 32'she06d85f7, 32'she06ee3c3, 32'she0704194, 32'she0719f6a, 32'she072fd44, 
               32'she0745b24, 32'she075b908, 32'she07716f2, 32'she07874e0, 32'she079d2d3, 32'she07b30cb, 32'she07c8ec7, 32'she07decc9, 
               32'she07f4acf, 32'she080a8db, 32'she08206eb, 32'she0836500, 32'she084c31a, 32'she0862139, 32'she0877f5c, 32'she088dd85, 
               32'she08a3bb2, 32'she08b99e4, 32'she08cf81b, 32'she08e5657, 32'she08fb497, 32'she09112dd, 32'she0927127, 32'she093cf77, 
               32'she0952dcb, 32'she0968c24, 32'she097ea81, 32'she09948e4, 32'she09aa74b, 32'she09c05b8, 32'she09d6429, 32'she09ec29f, 
               32'she0a0211a, 32'she0a17f99, 32'she0a2de1e, 32'she0a43ca7, 32'she0a59b35, 32'she0a6f9c8, 32'she0a85860, 32'she0a9b6fd, 
               32'she0ab159e, 32'she0ac7445, 32'she0add2f0, 32'she0af31a0, 32'she0b09055, 32'she0b1ef0e, 32'she0b34dcd, 32'she0b4ac90, 
               32'she0b60b58, 32'she0b76a25, 32'she0b8c8f7, 32'she0ba27cd, 32'she0bb86a9, 32'she0bce589, 32'she0be446e, 32'she0bfa358, 
               32'she0c10247, 32'she0c2613a, 32'she0c3c033, 32'she0c51f30, 32'she0c67e32, 32'she0c7dd39, 32'she0c93c44, 32'she0ca9b55, 
               32'she0cbfa6a, 32'she0cd5984, 32'she0ceb8a3, 32'she0d017c6, 32'she0d176ef, 32'she0d2d61c, 32'she0d4354e, 32'she0d59485, 
               32'she0d6f3c1, 32'she0d85301, 32'she0d9b247, 32'she0db1191, 32'she0dc70e0, 32'she0ddd033, 32'she0df2f8c, 32'she0e08ee9, 
               32'she0e1ee4b, 32'she0e34db2, 32'she0e4ad1e, 32'she0e60c8e, 32'she0e76c04, 32'she0e8cb7e, 32'she0ea2afd, 32'she0eb8a80, 
               32'she0ecea09, 32'she0ee4996, 32'she0efa928, 32'she0f108bf, 32'she0f2685b, 32'she0f3c7fb, 32'she0f527a0, 32'she0f6874a, 
               32'she0f7e6f9, 32'she0f946ad, 32'she0faa665, 32'she0fc0622, 32'she0fd65e4, 32'she0fec5ab, 32'she1002577, 32'she1018547, 
               32'she102e51c, 32'she10444f6, 32'she105a4d4, 32'she10704b8, 32'she10864a0, 32'she109c48d, 32'she10b247f, 32'she10c8475, 
               32'she10de470, 32'she10f4470, 32'she110a475, 32'she112047f, 32'she113648d, 32'she114c4a0, 32'she11624b8, 32'she11784d5, 
               32'she118e4f6, 32'she11a451c, 32'she11ba547, 32'she11d0577, 32'she11e65ac, 32'she11fc5e5, 32'she1212623, 32'she1228666, 
               32'she123e6ad, 32'she12546f9, 32'she126a74a, 32'she12807a0, 32'she12967fb, 32'she12ac85a, 32'she12c28be, 32'she12d8927, 
               32'she12ee995, 32'she1304a07, 32'she131aa7e, 32'she1330afa, 32'she1346b7a, 32'she135cc00, 32'she1372c8a, 32'she1388d19, 
               32'she139edac, 32'she13b4e44, 32'she13caee1, 32'she13e0f83, 32'she13f702a, 32'she140d0d5, 32'she1423185, 32'she143923a, 
               32'she144f2f3, 32'she14653b2, 32'she147b475, 32'she149153c, 32'she14a7609, 32'she14bd6da, 32'she14d37b0, 32'she14e988b, 
               32'she14ff96a, 32'she1515a4e, 32'she152bb37, 32'she1541c25, 32'she1557d17, 32'she156de0e, 32'she1583f0a, 32'she159a00a, 
               32'she15b0110, 32'she15c621a, 32'she15dc328, 32'she15f243c, 32'she1608554, 32'she161e671, 32'she1634792, 32'she164a8b8, 
               32'she16609e3, 32'she1676b13, 32'she168cc48, 32'she16a2d81, 32'she16b8ebf, 32'she16cf001, 32'she16e5149, 32'she16fb295, 
               32'she17113e5, 32'she172753b, 32'she173d695, 32'she17537f4, 32'she1769958, 32'she177fac0, 32'she1795c2d, 32'she17abd9f, 
               32'she17c1f15, 32'she17d8090, 32'she17ee210, 32'she1804395, 32'she181a51e, 32'she18306ac, 32'she184683e, 32'she185c9d6, 
               32'she1872b72, 32'she1888d13, 32'she189eeb8, 32'she18b5062, 32'she18cb211, 32'she18e13c4, 32'she18f757d, 32'she190d73a, 
               32'she19238fb, 32'she1939ac2, 32'she194fc8d, 32'she1965e5c, 32'she197c031, 32'she199220a, 32'she19a83e7, 32'she19be5ca, 
               32'she19d47b1, 32'she19ea99d, 32'she1a00b8d, 32'she1a16d83, 32'she1a2cf7c, 32'she1a4317b, 32'she1a5937e, 32'she1a6f586, 
               32'she1a85793, 32'she1a9b9a4, 32'she1ab1bba, 32'she1ac7dd5, 32'she1addff4, 32'she1af4218, 32'she1b0a441, 32'she1b2066e, 
               32'she1b368a0, 32'she1b4cad7, 32'she1b62d12, 32'she1b78f52, 32'she1b8f197, 32'she1ba53e0, 32'she1bbb62e, 32'she1bd1881, 
               32'she1be7ad8, 32'she1bfdd34, 32'she1c13f95, 32'she1c2a1fa, 32'she1c40464, 32'she1c566d3, 32'she1c6c946, 32'she1c82bbe, 
               32'she1c98e3b, 32'she1caf0bc, 32'she1cc5342, 32'she1cdb5cd, 32'she1cf185c, 32'she1d07af0, 32'she1d1dd89, 32'she1d34026, 
               32'she1d4a2c8, 32'she1d6056f, 32'she1d7681a, 32'she1d8caca, 32'she1da2d7e, 32'she1db9037, 32'she1dcf2f5, 32'she1de55b8, 
               32'she1dfb87f, 32'she1e11b4b, 32'she1e27e1b, 32'she1e3e0f0, 32'she1e543ca, 32'she1e6a6a8, 32'she1e8098b, 32'she1e96c73, 
               32'she1eacf5f, 32'she1ec3250, 32'she1ed9545, 32'she1eef83f, 32'she1f05b3e, 32'she1f1be42, 32'she1f3214a, 32'she1f48457, 
               32'she1f5e768, 32'she1f74a7e, 32'she1f8ad98, 32'she1fa10b8, 32'she1fb73dc, 32'she1fcd704, 32'she1fe3a31, 32'she1ff9d63, 
               32'she2010099, 32'she20263d4, 32'she203c714, 32'she2052a58, 32'she2068da1, 32'she207f0ef, 32'she2095441, 32'she20ab798, 
               32'she20c1af3, 32'she20d7e53, 32'she20ee1b7, 32'she2104521, 32'she211a88f, 32'she2130c01, 32'she2146f78, 32'she215d2f4, 
               32'she2173674, 32'she21899f9, 32'she219fd82, 32'she21b6111, 32'she21cc4a3, 32'she21e283b, 32'she21f8bd7, 32'she220ef77, 
               32'she222531c, 32'she223b6c6, 32'she2251a75, 32'she2267e28, 32'she227e1df, 32'she229459b, 32'she22aa95c, 32'she22c0d21, 
               32'she22d70eb, 32'she22ed4ba, 32'she230388d, 32'she2319c65, 32'she2330041, 32'she2346422, 32'she235c808, 32'she2372bf2, 
               32'she2388fe1, 32'she239f3d4, 32'she23b57cc, 32'she23cbbc9, 32'she23e1fca, 32'she23f83d0, 32'she240e7da, 32'she2424be9, 
               32'she243affc, 32'she2451414, 32'she2467831, 32'she247dc52, 32'she2494078, 32'she24aa4a2, 32'she24c08d1, 32'she24d6d05, 
               32'she24ed13d, 32'she250357a, 32'she25199bb, 32'she252fe01, 32'she254624b, 32'she255c69b, 32'she2572aee, 32'she2588f46, 
               32'she259f3a3, 32'she25b5804, 32'she25cbc6a, 32'she25e20d5, 32'she25f8544, 32'she260e9b7, 32'she2624e2f, 32'she263b2ac, 
               32'she265172e, 32'she2667bb3, 32'she267e03e, 32'she26944cd, 32'she26aa960, 32'she26c0df9, 32'she26d7295, 32'she26ed736, 
               32'she2703bdc, 32'she271a087, 32'she2730536, 32'she27469e9, 32'she275cea1, 32'she277335e, 32'she278981f, 32'she279fce4, 
               32'she27b61af, 32'she27cc67d, 32'she27e2b51, 32'she27f9029, 32'she280f505, 32'she28259e6, 32'she283becc, 32'she28523b6, 
               32'she28688a4, 32'she287ed98, 32'she289528f, 32'she28ab78c, 32'she28c1c8c, 32'she28d8192, 32'she28ee69c, 32'she2904baa, 
               32'she291b0bd, 32'she29315d5, 32'she2947af1, 32'she295e011, 32'she2974536, 32'she298aa60, 32'she29a0f8e, 32'she29b74c1, 
               32'she29cd9f8, 32'she29e3f34, 32'she29fa474, 32'she2a109b9, 32'she2a26f03, 32'she2a3d451, 32'she2a539a3, 32'she2a69efa, 
               32'she2a80456, 32'she2a969b6, 32'she2aacf1a, 32'she2ac3483, 32'she2ad99f1, 32'she2aeff63, 32'she2b064da, 32'she2b1ca55, 
               32'she2b32fd4, 32'she2b49559, 32'she2b5fae1, 32'she2b7606e, 32'she2b8c600, 32'she2ba2b96, 32'she2bb9131, 32'she2bcf6d1, 
               32'she2be5c74, 32'she2bfc21d, 32'she2c127c9, 32'she2c28d7b, 32'she2c3f331, 32'she2c558eb, 32'she2c6beaa, 32'she2c8246d, 
               32'she2c98a35, 32'she2caf001, 32'she2cc55d2, 32'she2cdbba8, 32'she2cf2182, 32'she2d08760, 32'she2d1ed43, 32'she2d3532a, 
               32'she2d4b916, 32'she2d61f07, 32'she2d784fb, 32'she2d8eaf5, 32'she2da50f3, 32'she2dbb6f5, 32'she2dd1cfc, 32'she2de8307, 
               32'she2dfe917, 32'she2e14f2b, 32'she2e2b544, 32'she2e41b62, 32'she2e58183, 32'she2e6e7aa, 32'she2e84dd4, 32'she2e9b404, 
               32'she2eb1a37, 32'she2ec8070, 32'she2ede6ac, 32'she2ef4cee, 32'she2f0b333, 32'she2f2197e, 32'she2f37fcc, 32'she2f4e61f, 
               32'she2f64c77, 32'she2f7b2d3, 32'she2f91934, 32'she2fa7f99, 32'she2fbe602, 32'she2fd4c70, 32'she2feb2e3, 32'she300195a, 
               32'she3017fd5, 32'she302e655, 32'she3044cd9, 32'she305b362, 32'she30719ef, 32'she3088081, 32'she309e717, 32'she30b4db2, 
               32'she30cb451, 32'she30e1af5, 32'she30f819d, 32'she310e849, 32'she3124efa, 32'she313b5b0, 32'she3151c6a, 32'she3168328, 
               32'she317e9eb, 32'she31950b2, 32'she31ab77e, 32'she31c1e4e, 32'she31d8523, 32'she31eebfc, 32'she32052da, 32'she321b9bc, 
               32'she32320a2, 32'she324878d, 32'she325ee7d, 32'she3275570, 32'she328bc69, 32'she32a2365, 32'she32b8a67, 32'she32cf16c, 
               32'she32e5876, 32'she32fbf85, 32'she3312698, 32'she3328daf, 32'she333f4cb, 32'she3355beb, 32'she336c310, 32'she3382a39, 
               32'she3399167, 32'she33af899, 32'she33c5fcf, 32'she33dc70a, 32'she33f2e4a, 32'she340958d, 32'she341fcd6, 32'she3436422, 
               32'she344cb73, 32'she34632c9, 32'she3479a23, 32'she3490181, 32'she34a68e4, 32'she34bd04b, 32'she34d37b7, 32'she34e9f27, 
               32'she350069b, 32'she3516e14, 32'she352d592, 32'she3543d13, 32'she355a49a, 32'she3570c24, 32'she35873b3, 32'she359db47, 
               32'she35b42df, 32'she35caa7b, 32'she35e121c, 32'she35f79c1, 32'she360e16a, 32'she3624918, 32'she363b0cb, 32'she3651881, 
               32'she366803c, 32'she367e7fc, 32'she3694fc0, 32'she36ab788, 32'she36c1f55, 32'she36d8727, 32'she36eeefc, 32'she37056d6, 
               32'she371beb5, 32'she3732697, 32'she3748e7f, 32'she375f66a, 32'she3775e5a, 32'she378c64f, 32'she37a2e48, 32'she37b9645, 
               32'she37cfe47, 32'she37e664d, 32'she37fce57, 32'she3813666, 32'she3829e79, 32'she3840691, 32'she3856ead, 32'she386d6cd, 
               32'she3883ef2, 32'she389a71b, 32'she38b0f49, 32'she38c777b, 32'she38ddfb1, 32'she38f47ec, 32'she390b02b, 32'she392186f, 
               32'she39380b6, 32'she394e903, 32'she3965153, 32'she397b9a8, 32'she3992202, 32'she39a8a60, 32'she39bf2c2, 32'she39d5b28, 
               32'she39ec393, 32'she3a02c03, 32'she3a19476, 32'she3a2fcee, 32'she3a4656b, 32'she3a5cdec, 32'she3a73671, 32'she3a89efa, 
               32'she3aa0788, 32'she3ab701b, 32'she3acd8b1, 32'she3ae414c, 32'she3afa9ec, 32'she3b1128f, 32'she3b27b38, 32'she3b3e3e4, 
               32'she3b54c95, 32'she3b6b54a, 32'she3b81e04, 32'she3b986c2, 32'she3baef84, 32'she3bc584b, 32'she3bdc116, 32'she3bf29e5, 
               32'she3c092b9, 32'she3c1fb91, 32'she3c3646d, 32'she3c4cd4e, 32'she3c63633, 32'she3c79f1d, 32'she3c9080b, 32'she3ca70fd, 
               32'she3cbd9f4, 32'she3cd42ee, 32'she3ceabee, 32'she3d014f1, 32'she3d17df9, 32'she3d2e706, 32'she3d45016, 32'she3d5b92b, 
               32'she3d72245, 32'she3d88b62, 32'she3d9f484, 32'she3db5dab, 32'she3dcc6d5, 32'she3de3004, 32'she3df9938, 32'she3e1026f, 
               32'she3e26bac, 32'she3e3d4ec, 32'she3e53e31, 32'she3e6a77a, 32'she3e810c7, 32'she3e97a19, 32'she3eae36f, 32'she3ec4cc9, 
               32'she3edb628, 32'she3ef1f8b, 32'she3f088f2, 32'she3f1f25e, 32'she3f35bce, 32'she3f4c542, 32'she3f62ebb, 32'she3f79838, 
               32'she3f901ba, 32'she3fa6b3f, 32'she3fbd4c9, 32'she3fd3e57, 32'she3fea7ea, 32'she4001181, 32'she4017b1c, 32'she402e4bc, 
               32'she4044e60, 32'she405b808, 32'she40721b4, 32'she4088b65, 32'she409f51a, 32'she40b5ed4, 32'she40cc891, 32'she40e3254, 
               32'she40f9c1a, 32'she41105e5, 32'she4126fb4, 32'she413d987, 32'she415435f, 32'she416ad3a, 32'she418171b, 32'she41980ff, 
               32'she41aeae8, 32'she41c54d5, 32'she41dbec7, 32'she41f28bc, 32'she42092b6, 32'she421fcb5, 32'she42366b7, 32'she424d0be, 
               32'she4263ac9, 32'she427a4d9, 32'she4290eed, 32'she42a7905, 32'she42be321, 32'she42d4d42, 32'she42eb767, 32'she4302190, 
               32'she4318bbe, 32'she432f5ef, 32'she4346026, 32'she435ca60, 32'she437349f, 32'she4389ee2, 32'she43a0929, 32'she43b7374, 
               32'she43cddc4, 32'she43e4818, 32'she43fb271, 32'she4411ccd, 32'she442872e, 32'she443f194, 32'she4455bfd, 32'she446c66b, 
               32'she44830dd, 32'she4499b53, 32'she44b05ce, 32'she44c704d, 32'she44ddad0, 32'she44f4557, 32'she450afe3, 32'she4521a73, 
               32'she4538507, 32'she454efa0, 32'she4565a3c, 32'she457c4de, 32'she4592f83, 32'she45a9a2c, 32'she45c04da, 32'she45d6f8c, 
               32'she45eda43, 32'she46044fd, 32'she461afbc, 32'she4631a7f, 32'she4648547, 32'she465f012, 32'she4675ae2, 32'she468c5b6, 
               32'she46a308f, 32'she46b9b6b, 32'she46d064c, 32'she46e7131, 32'she46fdc1b, 32'she4714709, 32'she472b1fa, 32'she4741cf1, 
               32'she47587eb, 32'she476f2ea, 32'she4785ded, 32'she479c8f4, 32'she47b33ff, 32'she47c9f0f, 32'she47e0a23, 32'she47f753b, 
               32'she480e057, 32'she4824b78, 32'she483b69d, 32'she48521c6, 32'she4868cf3, 32'she487f825, 32'she489635a, 32'she48ace94, 
               32'she48c39d3, 32'she48da515, 32'she48f105c, 32'she4907ba7, 32'she491e6f6, 32'she4935249, 32'she494bda1, 32'she49628fd, 
               32'she497945d, 32'she498ffc1, 32'she49a6b2a, 32'she49bd697, 32'she49d4208, 32'she49ead7d, 32'she4a018f7, 32'she4a18474, 
               32'she4a2eff6, 32'she4a45b7c, 32'she4a5c707, 32'she4a73295, 32'she4a89e28, 32'she4aa09bf, 32'she4ab755a, 32'she4ace0fa, 
               32'she4ae4c9d, 32'she4afb845, 32'she4b123f1, 32'she4b28fa1, 32'she4b3fb56, 32'she4b5670f, 32'she4b6d2cb, 32'she4b83e8d, 
               32'she4b9aa52, 32'she4bb161b, 32'she4bc81e9, 32'she4bdedbb, 32'she4bf5991, 32'she4c0c56b, 32'she4c2314a, 32'she4c39d2d, 
               32'she4c50914, 32'she4c674ff, 32'she4c7e0ee, 32'she4c94ce2, 32'she4cab8d9, 32'she4cc24d5, 32'she4cd90d5, 32'she4cefcda, 
               32'she4d068e2, 32'she4d1d4ef, 32'she4d34100, 32'she4d4ad15, 32'she4d6192e, 32'she4d7854c, 32'she4d8f16d, 32'she4da5d93, 
               32'she4dbc9bd, 32'she4dd35eb, 32'she4dea21e, 32'she4e00e54, 32'she4e17a8f, 32'she4e2e6ce, 32'she4e45311, 32'she4e5bf59, 
               32'she4e72ba4, 32'she4e897f4, 32'she4ea0448, 32'she4eb70a0, 32'she4ecdcfc, 32'she4ee495c, 32'she4efb5c1, 32'she4f12229, 
               32'she4f28e96, 32'she4f3fb07, 32'she4f5677d, 32'she4f6d3f6, 32'she4f84074, 32'she4f9acf5, 32'she4fb197b, 32'she4fc8605, 
               32'she4fdf294, 32'she4ff5f26, 32'she500cbbc, 32'she5023857, 32'she503a4f6, 32'she5051199, 32'she5067e40, 32'she507eaec, 
               32'she509579b, 32'she50ac44f, 32'she50c3107, 32'she50d9dc3, 32'she50f0a83, 32'she5107747, 32'she511e410, 32'she51350dc, 
               32'she514bdad, 32'she5162a82, 32'she517975b, 32'she5190438, 32'she51a711a, 32'she51bddff, 32'she51d4ae9, 32'she51eb7d7, 
               32'she52024c9, 32'she52191bf, 32'she522feb9, 32'she5246bb8, 32'she525d8ba, 32'she52745c1, 32'she528b2cc, 32'she52a1fdb, 
               32'she52b8cee, 32'she52cfa05, 32'she52e6720, 32'she52fd440, 32'she5314163, 32'she532ae8b, 32'she5341bb7, 32'she53588e7, 
               32'she536f61b, 32'she5386354, 32'she539d090, 32'she53b3dd1, 32'she53cab15, 32'she53e185e, 32'she53f85ab, 32'she540f2fc, 
               32'she5426051, 32'she543cdab, 32'she5453b08, 32'she546a86a, 32'she54815cf, 32'she5498339, 32'she54af0a7, 32'she54c5e19, 
               32'she54dcb8f, 32'she54f3909, 32'she550a688, 32'she552140a, 32'she5538191, 32'she554ef1c, 32'she5565cab, 32'she557ca3e, 
               32'she55937d5, 32'she55aa570, 32'she55c130f, 32'she55d80b2, 32'she55eee5a, 32'she5605c06, 32'she561c9b5, 32'she5633769, 
               32'she564a521, 32'she56612dd, 32'she567809d, 32'she568ee61, 32'she56a5c2a, 32'she56bc9f6, 32'she56d37c7, 32'she56ea59b, 
               32'she5701374, 32'she5718151, 32'she572ef32, 32'she5745d17, 32'she575cb00, 32'she57738ed, 32'she578a6de, 32'she57a14d4, 
               32'she57b82cd, 32'she57cf0cb, 32'she57e5ecc, 32'she57fccd2, 32'she5813adc, 32'she582a8ea, 32'she58416fc, 32'she5858512, 
               32'she586f32c, 32'she588614a, 32'she589cf6d, 32'she58b3d93, 32'she58cabbe, 32'she58e19ec, 32'she58f881f, 32'she590f656, 
               32'she5926490, 32'she593d2cf, 32'she5954112, 32'she596af59, 32'she5981da4, 32'she5998bf3, 32'she59afa47, 32'she59c689e, 
               32'she59dd6f9, 32'she59f4559, 32'she5a0b3bc, 32'she5a22224, 32'she5a39090, 32'she5a4feff, 32'she5a66d73, 32'she5a7dbeb, 
               32'she5a94a67, 32'she5aab8e7, 32'she5ac276b, 32'she5ad95f3, 32'she5af047f, 32'she5b0730f, 32'she5b1e1a3, 32'she5b3503c, 
               32'she5b4bed8, 32'she5b62d79, 32'she5b79c1d, 32'she5b90ac6, 32'she5ba7972, 32'she5bbe823, 32'she5bd56d7, 32'she5bec590, 
               32'she5c0344d, 32'she5c1a30e, 32'she5c311d3, 32'she5c4809c, 32'she5c5ef69, 32'she5c75e3a, 32'she5c8cd0f, 32'she5ca3be8, 
               32'she5cbaac5, 32'she5cd19a6, 32'she5ce888b, 32'she5cff775, 32'she5d16662, 32'she5d2d553, 32'she5d44449, 32'she5d5b342, 
               32'she5d72240, 32'she5d89141, 32'she5da0047, 32'she5db6f50, 32'she5dcde5e, 32'she5de4d6f, 32'she5dfbc85, 32'she5e12b9f, 
               32'she5e29abc, 32'she5e409de, 32'she5e57904, 32'she5e6e82e, 32'she5e8575b, 32'she5e9c68d, 32'she5eb35c3, 32'she5eca4fd, 
               32'she5ee143b, 32'she5ef837d, 32'she5f0f2c3, 32'she5f2620d, 32'she5f3d15b, 32'she5f540ad, 32'she5f6b003, 32'she5f81f5d, 
               32'she5f98ebb, 32'she5fafe1d, 32'she5fc6d83, 32'she5fddced, 32'she5ff4c5b, 32'she600bbcd, 32'she6022b43, 32'she6039abd, 
               32'she6050a3b, 32'she60679bd, 32'she607e944, 32'she60958ce, 32'she60ac85c, 32'she60c37ee, 32'she60da784, 32'she60f171e, 
               32'she61086bc, 32'she611f65e, 32'she6136605, 32'she614d5af, 32'she616455d, 32'she617b50f, 32'she61924c5, 32'she61a947f, 
               32'she61c043d, 32'she61d73ff, 32'she61ee3c6, 32'she6205390, 32'she621c35e, 32'she6233330, 32'she624a306, 32'she62612e0, 
               32'she62782be, 32'she628f2a0, 32'she62a6286, 32'she62bd270, 32'she62d425e, 32'she62eb250, 32'she6302246, 32'she6319240, 
               32'she633023e, 32'she6347240, 32'she635e245, 32'she637524f, 32'she638c25d, 32'she63a326f, 32'she63ba285, 32'she63d129e, 
               32'she63e82bc, 32'she63ff2de, 32'she6416303, 32'she642d32d, 32'she644435a, 32'she645b38c, 32'she64723c2, 32'she64893fb, 
               32'she64a0438, 32'she64b747a, 32'she64ce4bf, 32'she64e5509, 32'she64fc556, 32'she65135a7, 32'she652a5fc, 32'she6541656, 
               32'she65586b3, 32'she656f714, 32'she6586779, 32'she659d7e2, 32'she65b484f, 32'she65cb8c0, 32'she65e2935, 32'she65f99ae, 
               32'she6610a2a, 32'she6627aab, 32'she663eb30, 32'she6655bb8, 32'she666cc45, 32'she6683cd5, 32'she669ad6a, 32'she66b1e02, 
               32'she66c8e9f, 32'she66dff3f, 32'she66f6fe3, 32'she670e08c, 32'she6725138, 32'she673c1e8, 32'she675329c, 32'she676a354, 
               32'she6781410, 32'she67984cf, 32'she67af593, 32'she67c665b, 32'she67dd727, 32'she67f47f6, 32'she680b8ca, 32'she68229a1, 
               32'she6839a7c, 32'she6850b5c, 32'she6867c3f, 32'she687ed26, 32'she6895e11, 32'she68acf00, 32'she68c3ff3, 32'she68db0ea, 
               32'she68f21e5, 32'she69092e4, 32'she69203e6, 32'she69374ed, 32'she694e5f7, 32'she6965706, 32'she697c818, 32'she699392e, 
               32'she69aaa48, 32'she69c1b66, 32'she69d8c88, 32'she69efdae, 32'she6a06ed8, 32'she6a1e006, 32'she6a35137, 32'she6a4c26d, 
               32'she6a633a6, 32'she6a7a4e4, 32'she6a91625, 32'she6aa876a, 32'she6abf8b3, 32'she6ad6a00, 32'she6aedb51, 32'she6b04ca6, 
               32'she6b1bdff, 32'she6b32f5b, 32'she6b4a0bc, 32'she6b61220, 32'she6b78389, 32'she6b8f4f5, 32'she6ba6665, 32'she6bbd7d9, 
               32'she6bd4951, 32'she6bebacd, 32'she6c02c4c, 32'she6c19dd0, 32'she6c30f57, 32'she6c480e3, 32'she6c5f272, 32'she6c76405, 
               32'she6c8d59c, 32'she6ca4737, 32'she6cbb8d6, 32'she6cd2a79, 32'she6ce9c1f, 32'she6d00dca, 32'she6d17f78, 32'she6d2f12a, 
               32'she6d462e1, 32'she6d5d49b, 32'she6d74658, 32'she6d8b81a, 32'she6da29e0, 32'she6db9ba9, 32'she6dd0d77, 32'she6de7f48, 
               32'she6dff11d, 32'she6e162f6, 32'she6e2d4d3, 32'she6e446b4, 32'she6e5b899, 32'she6e72a81, 32'she6e89c6d, 32'she6ea0e5e, 
               32'she6eb8052, 32'she6ecf24a, 32'she6ee6446, 32'she6efd645, 32'she6f14849, 32'she6f2ba51, 32'she6f42c5c, 32'she6f59e6b, 
               32'she6f7107e, 32'she6f88295, 32'she6f9f4b0, 32'she6fb66ce, 32'she6fcd8f1, 32'she6fe4b17, 32'she6ffbd41, 32'she7012f6f, 
               32'she702a1a1, 32'she70413d7, 32'she7058611, 32'she706f84e, 32'she7086a8f, 32'she709dcd5, 32'she70b4f1e, 32'she70cc16b, 
               32'she70e33bb, 32'she70fa610, 32'she7111868, 32'she7128ac4, 32'she713fd25, 32'she7156f89, 32'she716e1f0, 32'she718545c, 
               32'she719c6cb, 32'she71b393f, 32'she71cabb6, 32'she71e1e31, 32'she71f90b0, 32'she7210332, 32'she72275b9, 32'she723e843, 
               32'she7255ad1, 32'she726cd63, 32'she7283ff9, 32'she729b293, 32'she72b2530, 32'she72c97d1, 32'she72e0a77, 32'she72f7d20, 
               32'she730efcc, 32'she732627d, 32'she733d531, 32'she73547ea, 32'she736baa6, 32'she7382d66, 32'she739a029, 32'she73b12f1, 
               32'she73c85bc, 32'she73df88c, 32'she73f6b5f, 32'she740de35, 32'she7425110, 32'she743c3ef, 32'she74536d1, 32'she746a9b7, 
               32'she7481ca1, 32'she7498f8f, 32'she74b0280, 32'she74c7575, 32'she74de86f, 32'she74f5b6b, 32'she750ce6c, 32'she7524171, 
               32'she753b479, 32'she7552785, 32'she7569a95, 32'she7580da9, 32'she75980c1, 32'she75af3dc, 32'she75c66fb, 32'she75dda1e, 
               32'she75f4d45, 32'she760c070, 32'she762339e, 32'she763a6d0, 32'she7651a06, 32'she7668d40, 32'she768007e, 32'she76973bf, 
               32'she76ae704, 32'she76c5a4d, 32'she76dcd9a, 32'she76f40ea, 32'she770b43e, 32'she7722797, 32'she7739af2, 32'she7750e52, 
               32'she77681b6, 32'she777f51d, 32'she7796888, 32'she77adbf7, 32'she77c4f69, 32'she77dc2e0, 32'she77f365a, 32'she780a9d8, 
               32'she7821d59, 32'she78390df, 32'she7850468, 32'she78677f5, 32'she787eb86, 32'she7895f1a, 32'she78ad2b3, 32'she78c464f, 
               32'she78db9ef, 32'she78f2d92, 32'she790a13a, 32'she79214e5, 32'she7938894, 32'she794fc47, 32'she7966ffd, 32'she797e3b8, 
               32'she7995776, 32'she79acb37, 32'she79c3efd, 32'she79db2c6, 32'she79f2693, 32'she7a09a64, 32'she7a20e39, 32'she7a38211, 
               32'she7a4f5ed, 32'she7a669cd, 32'she7a7ddb1, 32'she7a95198, 32'she7aac583, 32'she7ac3972, 32'she7adad65, 32'she7af215b, 
               32'she7b09555, 32'she7b20953, 32'she7b37d55, 32'she7b4f15a, 32'she7b66563, 32'she7b7d970, 32'she7b94d80, 32'she7bac195, 
               32'she7bc35ad, 32'she7bda9c9, 32'she7bf1de8, 32'she7c0920c, 32'she7c20633, 32'she7c37a5e, 32'she7c4ee8c, 32'she7c662be, 
               32'she7c7d6f4, 32'she7c94b2e, 32'she7cabf6c, 32'she7cc33ad, 32'she7cda7f2, 32'she7cf1c3a, 32'she7d09087, 32'she7d204d7, 
               32'she7d3792b, 32'she7d4ed82, 32'she7d661de, 32'she7d7d63d, 32'she7d94a9f, 32'she7dabf06, 32'she7dc3370, 32'she7dda7de, 
               32'she7df1c50, 32'she7e090c5, 32'she7e2053e, 32'she7e379bb, 32'she7e4ee3c, 32'she7e662c0, 32'she7e7d748, 32'she7e94bd3, 
               32'she7eac063, 32'she7ec34f6, 32'she7eda98d, 32'she7ef1e27, 32'she7f092c6, 32'she7f20768, 32'she7f37c0d, 32'she7f4f0b7, 
               32'she7f66564, 32'she7f7da14, 32'she7f94ec9, 32'she7fac381, 32'she7fc383d, 32'she7fdacfd, 32'she7ff21c0, 32'she8009687, 
               32'she8020b52, 32'she8038020, 32'she804f4f2, 32'she80669c8, 32'she807dea2, 32'she809537f, 32'she80ac860, 32'she80c3d44, 
               32'she80db22d, 32'she80f2719, 32'she8109c08, 32'she81210fc, 32'she81385f3, 32'she814faed, 32'she8166fec, 32'she817e4ee, 
               32'she81959f4, 32'she81acefd, 32'she81c440a, 32'she81db91b, 32'she81f2e30, 32'she820a348, 32'she8221864, 32'she8238d84, 
               32'she82502a7, 32'she82677ce, 32'she827ecf8, 32'she8296227, 32'she82ad759, 32'she82c4c8e, 32'she82dc1c8, 32'she82f3705, 
               32'she830ac45, 32'she832218a, 32'she83396d2, 32'she8350c1d, 32'she836816d, 32'she837f6c0, 32'she8396c16, 32'she83ae171, 
               32'she83c56cf, 32'she83dcc31, 32'she83f4196, 32'she840b6ff, 32'she8422c6c, 32'she843a1dc, 32'she8451750, 32'she8468cc8, 
               32'she8480243, 32'she84977c2, 32'she84aed45, 32'she84c62cb, 32'she84dd855, 32'she84f4de2, 32'she850c374, 32'she8523909, 
               32'she853aea1, 32'she855243d, 32'she85699dd, 32'she8580f81, 32'she8598528, 32'she85afad3, 32'she85c7081, 32'she85de633, 
               32'she85f5be9, 32'she860d1a2, 32'she862475f, 32'she863bd20, 32'she86532e4, 32'she866a8ac, 32'she8681e78, 32'she8699447, 
               32'she86b0a1a, 32'she86c7ff0, 32'she86df5cb, 32'she86f6ba8, 32'she870e18a, 32'she872576f, 32'she873cd57, 32'she8754344, 
               32'she876b934, 32'she8782f27, 32'she879a51e, 32'she87b1b19, 32'she87c9118, 32'she87e071a, 32'she87f7d1f, 32'she880f329, 
               32'she8826936, 32'she883df46, 32'she885555a, 32'she886cb72, 32'she888418e, 32'she889b7ad, 32'she88b2dcf, 32'she88ca3f6, 
               32'she88e1a20, 32'she88f904d, 32'she891067e, 32'she8927cb3, 32'she893f2eb, 32'she8956927, 32'she896df67, 32'she89855aa, 
               32'she899cbf1, 32'she89b423b, 32'she89cb889, 32'she89e2edb, 32'she89fa530, 32'she8a11b89, 32'she8a291e5, 32'she8a40845, 
               32'she8a57ea9, 32'she8a6f510, 32'she8a86b7b, 32'she8a9e1ea, 32'she8ab585c, 32'she8acced1, 32'she8ae454b, 32'she8afbbc7, 
               32'she8b13248, 32'she8b2a8cc, 32'she8b41f53, 32'she8b595df, 32'she8b70c6d, 32'she8b88300, 32'she8b9f996, 32'she8bb702f, 
               32'she8bce6cd, 32'she8be5d6d, 32'she8bfd412, 32'she8c14aba, 32'she8c2c165, 32'she8c43814, 32'she8c5aec7, 32'she8c7257d, 
               32'she8c89c37, 32'she8ca12f4, 32'she8cb89b5, 32'she8cd007a, 32'she8ce7742, 32'she8cfee0e, 32'she8d164dd, 32'she8d2dbb0, 
               32'she8d45286, 32'she8d5c960, 32'she8d7403e, 32'she8d8b71f, 32'she8da2e04, 32'she8dba4ec, 32'she8dd1bd8, 32'she8de92c7, 
               32'she8e009ba, 32'she8e180b1, 32'she8e2f7ab, 32'she8e46ea9, 32'she8e5e5aa, 32'she8e75caf, 32'she8e8d3b7, 32'she8ea4ac3, 
               32'she8ebc1d3, 32'she8ed38e6, 32'she8eeaffd, 32'she8f02717, 32'she8f19e34, 32'she8f31556, 32'she8f48c7b, 32'she8f603a3, 
               32'she8f77acf, 32'she8f8f1ff, 32'she8fa6932, 32'she8fbe068, 32'she8fd57a2, 32'she8fecee0, 32'she9004621, 32'she901bd66, 
               32'she90334af, 32'she904abfa, 32'she906234a, 32'she9079a9d, 32'she90911f3, 32'she90a894d, 32'she90c00ab, 32'she90d780c, 
               32'she90eef71, 32'she91066d9, 32'she911de45, 32'she91355b4, 32'she914cd27, 32'she916449d, 32'she917bc17, 32'she9193395, 
               32'she91aab16, 32'she91c229a, 32'she91d9a22, 32'she91f11ae, 32'she920893d, 32'she92200cf, 32'she9237866, 32'she924efff, 
               32'she926679c, 32'she927df3d, 32'she92956e1, 32'she92ace89, 32'she92c4634, 32'she92dbde3, 32'she92f3596, 32'she930ad4b, 
               32'she9322505, 32'she9339cc2, 32'she9351482, 32'she9368c46, 32'she938040d, 32'she9397bd8, 32'she93af3a7, 32'she93c6b79, 
               32'she93de34e, 32'she93f5b27, 32'she940d304, 32'she9424ae4, 32'she943c2c7, 32'she9453aae, 32'she946b299, 32'she9482a87, 
               32'she949a278, 32'she94b1a6d, 32'she94c9266, 32'she94e0a62, 32'she94f8261, 32'she950fa64, 32'she952726b, 32'she953ea75, 
               32'she9556282, 32'she956da93, 32'she95852a8, 32'she959cac0, 32'she95b42db, 32'she95cbafa, 32'she95e331d, 32'she95fab43, 
               32'she961236c, 32'she9629b99, 32'she96413c9, 32'she9658bfd, 32'she9670435, 32'she9687c70, 32'she969f4ae, 32'she96b6cf0, 
               32'she96ce535, 32'she96e5d7e, 32'she96fd5ca, 32'she9714e1a, 32'she972c66d, 32'she9743ec4, 32'she975b71e, 32'she9772f7c, 
               32'she978a7dd, 32'she97a2042, 32'she97b98aa, 32'she97d1115, 32'she97e8984, 32'she98001f7, 32'she9817a6d, 32'she982f2e6, 
               32'she9846b63, 32'she985e3e4, 32'she9875c68, 32'she988d4ef, 32'she98a4d7a, 32'she98bc608, 32'she98d3e9a, 32'she98eb72f, 
               32'she9902fc7, 32'she991a864, 32'she9932103, 32'she99499a6, 32'she996124d, 32'she9978af7, 32'she99903a4, 32'she99a7c55, 
               32'she99bf509, 32'she99d6dc1, 32'she99ee67c, 32'she9a05f3b, 32'she9a1d7fd, 32'she9a350c2, 32'she9a4c98b, 32'she9a64258, 
               32'she9a7bb28, 32'she9a933fb, 32'she9aaacd2, 32'she9ac25ac, 32'she9ad9e8a, 32'she9af176b, 32'she9b0904f, 32'she9b20937, 
               32'she9b38223, 32'she9b4fb12, 32'she9b67404, 32'she9b7ecfa, 32'she9b965f3, 32'she9badeef, 32'she9bc57f0, 32'she9bdd0f3, 
               32'she9bf49fa, 32'she9c0c304, 32'she9c23c12, 32'she9c3b523, 32'she9c52e38, 32'she9c6a750, 32'she9c8206b, 32'she9c9998a, 
               32'she9cb12ad, 32'she9cc8bd3, 32'she9ce04fc, 32'she9cf7e28, 32'she9d0f758, 32'she9d2708c, 32'she9d3e9c3, 32'she9d562fd, 
               32'she9d6dc3b, 32'she9d8557c, 32'she9d9cec0, 32'she9db4808, 32'she9dcc154, 32'she9de3aa3, 32'she9dfb3f5, 32'she9e12d4a, 
               32'she9e2a6a3, 32'she9e42000, 32'she9e59960, 32'she9e712c3, 32'she9e88c2a, 32'she9ea0594, 32'she9eb7f01, 32'she9ecf872, 
               32'she9ee71e6, 32'she9efeb5e, 32'she9f164d9, 32'she9f2de58, 32'she9f457da, 32'she9f5d15f, 32'she9f74ae8, 32'she9f8c474, 
               32'she9fa3e03, 32'she9fbb796, 32'she9fd312c, 32'she9feaac6, 32'shea002463, 32'shea019e04, 32'shea0317a7, 32'shea04914f, 
               32'shea060af9, 32'shea0784a7, 32'shea08fe59, 32'shea0a780e, 32'shea0bf1c6, 32'shea0d6b81, 32'shea0ee540, 32'shea105f03, 
               32'shea11d8c8, 32'shea135291, 32'shea14cc5e, 32'shea16462e, 32'shea17c001, 32'shea1939d8, 32'shea1ab3b2, 32'shea1c2d8f, 
               32'shea1da770, 32'shea1f2154, 32'shea209b3b, 32'shea221526, 32'shea238f15, 32'shea250906, 32'shea2682fb, 32'shea27fcf4, 
               32'shea2976ef, 32'shea2af0ee, 32'shea2c6af1, 32'shea2de4f7, 32'shea2f5f00, 32'shea30d90c, 32'shea32531c, 32'shea33cd30, 
               32'shea354746, 32'shea36c160, 32'shea383b7e, 32'shea39b59e, 32'shea3b2fc2, 32'shea3ca9ea, 32'shea3e2415, 32'shea3f9e43, 
               32'shea411874, 32'shea4292a9, 32'shea440ce1, 32'shea45871d, 32'shea47015c, 32'shea487b9e, 32'shea49f5e4, 32'shea4b702d, 
               32'shea4cea79, 32'shea4e64c9, 32'shea4fdf1c, 32'shea515972, 32'shea52d3cc, 32'shea544e29, 32'shea55c889, 32'shea5742ed, 
               32'shea58bd54, 32'shea5a37be, 32'shea5bb22c, 32'shea5d2c9d, 32'shea5ea712, 32'shea602189, 32'shea619c04, 32'shea631683, 
               32'shea649105, 32'shea660b8a, 32'shea678612, 32'shea69009e, 32'shea6a7b2d, 32'shea6bf5bf, 32'shea6d7055, 32'shea6eeaee, 
               32'shea70658a, 32'shea71e02a, 32'shea735acd, 32'shea74d573, 32'shea76501d, 32'shea77caca, 32'shea79457a, 32'shea7ac02e, 
               32'shea7c3ae5, 32'shea7db59f, 32'shea7f305d, 32'shea80ab1e, 32'shea8225e2, 32'shea83a0a9, 32'shea851b74, 32'shea869642, 
               32'shea881114, 32'shea898be9, 32'shea8b06c1, 32'shea8c819c, 32'shea8dfc7b, 32'shea8f775d, 32'shea90f242, 32'shea926d2b, 
               32'shea93e817, 32'shea956306, 32'shea96ddf9, 32'shea9858ee, 32'shea99d3e8, 32'shea9b4ee4, 32'shea9cc9e4, 32'shea9e44e7, 
               32'shea9fbfed, 32'sheaa13af7, 32'sheaa2b604, 32'sheaa43114, 32'sheaa5ac27, 32'sheaa7273e, 32'sheaa8a258, 32'sheaaa1d76, 
               32'sheaab9896, 32'sheaad13ba, 32'sheaae8ee2, 32'sheab00a0c, 32'sheab1853a, 32'sheab3006b, 32'sheab47b9f, 32'sheab5f6d7, 
               32'sheab77212, 32'sheab8ed50, 32'sheaba6892, 32'sheabbe3d7, 32'sheabd5f1f, 32'sheabeda6a, 32'sheac055b9, 32'sheac1d10b, 
               32'sheac34c60, 32'sheac4c7b8, 32'sheac64314, 32'sheac7be73, 32'sheac939d5, 32'sheacab53b, 32'sheacc30a4, 32'sheacdac10, 
               32'sheacf277f, 32'shead0a2f2, 32'shead21e68, 32'shead399e1, 32'shead5155d, 32'shead690dd, 32'shead80c60, 32'shead987e6, 
               32'sheadb0370, 32'sheadc7efd, 32'sheaddfa8d, 32'sheadf7620, 32'sheae0f1b6, 32'sheae26d50, 32'sheae3e8ed, 32'sheae5648e, 
               32'sheae6e031, 32'sheae85bd8, 32'sheae9d782, 32'sheaeb532f, 32'sheaeccee0, 32'sheaee4a94, 32'sheaefc64b, 32'sheaf14205, 
               32'sheaf2bdc3, 32'sheaf43983, 32'sheaf5b547, 32'sheaf7310f, 32'sheaf8acd9, 32'sheafa28a7, 32'sheafba478, 32'sheafd204c, 
               32'sheafe9c24, 32'sheb0017ff, 32'sheb0193dd, 32'sheb030fbe, 32'sheb048ba2, 32'sheb06078a, 32'sheb078375, 32'sheb08ff63, 
               32'sheb0a7b54, 32'sheb0bf749, 32'sheb0d7341, 32'sheb0eef3c, 32'sheb106b3a, 32'sheb11e73c, 32'sheb136341, 32'sheb14df49, 
               32'sheb165b54, 32'sheb17d762, 32'sheb195374, 32'sheb1acf89, 32'sheb1c4ba1, 32'sheb1dc7bc, 32'sheb1f43db, 32'sheb20bffd, 
               32'sheb223c22, 32'sheb23b84a, 32'sheb253475, 32'sheb26b0a4, 32'sheb282cd6, 32'sheb29a90b, 32'sheb2b2543, 32'sheb2ca17f, 
               32'sheb2e1dbe, 32'sheb2f99ff, 32'sheb311645, 32'sheb32928d, 32'sheb340ed9, 32'sheb358b27, 32'sheb370779, 32'sheb3883ce, 
               32'sheb3a0027, 32'sheb3b7c82, 32'sheb3cf8e1, 32'sheb3e7543, 32'sheb3ff1a8, 32'sheb416e11, 32'sheb42ea7c, 32'sheb4466eb, 
               32'sheb45e35d, 32'sheb475fd2, 32'sheb48dc4b, 32'sheb4a58c6, 32'sheb4bd545, 32'sheb4d51c7, 32'sheb4ece4c, 32'sheb504ad4, 
               32'sheb51c760, 32'sheb5343ef, 32'sheb54c081, 32'sheb563d16, 32'sheb57b9ae, 32'sheb593649, 32'sheb5ab2e8, 32'sheb5c2f8a, 
               32'sheb5dac2f, 32'sheb5f28d7, 32'sheb60a582, 32'sheb622231, 32'sheb639ee3, 32'sheb651b98, 32'sheb669850, 32'sheb68150b, 
               32'sheb6991ca, 32'sheb6b0e8b, 32'sheb6c8b50, 32'sheb6e0818, 32'sheb6f84e3, 32'sheb7101b1, 32'sheb727e83, 32'sheb73fb57, 
               32'sheb75782f, 32'sheb76f50a, 32'sheb7871e8, 32'sheb79eeca, 32'sheb7b6bae, 32'sheb7ce896, 32'sheb7e6581, 32'sheb7fe26f, 
               32'sheb815f60, 32'sheb82dc54, 32'sheb84594c, 32'sheb85d646, 32'sheb875344, 32'sheb88d045, 32'sheb8a4d49, 32'sheb8bca50, 
               32'sheb8d475b, 32'sheb8ec468, 32'sheb904179, 32'sheb91be8d, 32'sheb933ba4, 32'sheb94b8be, 32'sheb9635db, 32'sheb97b2fc, 
               32'sheb99301f, 32'sheb9aad46, 32'sheb9c2a70, 32'sheb9da79d, 32'sheb9f24cd, 32'sheba0a200, 32'sheba21f37, 32'sheba39c71, 
               32'sheba519ad, 32'sheba696ed, 32'sheba81430, 32'sheba99176, 32'shebab0ec0, 32'shebac8c0c, 32'shebae095c, 32'shebaf86ae, 
               32'shebb10404, 32'shebb2815d, 32'shebb3feb9, 32'shebb57c18, 32'shebb6f97b, 32'shebb876e0, 32'shebb9f449, 32'shebbb71b5, 
               32'shebbcef23, 32'shebbe6c95, 32'shebbfea0b, 32'shebc16783, 32'shebc2e4fe, 32'shebc4627d, 32'shebc5dffe, 32'shebc75d83, 
               32'shebc8db0b, 32'shebca5896, 32'shebcbd624, 32'shebcd53b5, 32'shebced149, 32'shebd04ee1, 32'shebd1cc7b, 32'shebd34a19, 
               32'shebd4c7ba, 32'shebd6455d, 32'shebd7c304, 32'shebd940ae, 32'shebdabe5c, 32'shebdc3c0c, 32'shebddb9bf, 32'shebdf3776, 
               32'shebe0b52f, 32'shebe232ec, 32'shebe3b0ac, 32'shebe52e6f, 32'shebe6ac35, 32'shebe829fe, 32'shebe9a7ca, 32'shebeb259a, 
               32'shebeca36c, 32'shebee2141, 32'shebef9f1a, 32'shebf11cf6, 32'shebf29ad4, 32'shebf418b6, 32'shebf5969b, 32'shebf71483, 
               32'shebf8926f, 32'shebfa105d, 32'shebfb8e4e, 32'shebfd0c42, 32'shebfe8a3a, 32'shec000835, 32'shec018632, 32'shec030433, 
               32'shec048237, 32'shec06003e, 32'shec077e48, 32'shec08fc55, 32'shec0a7a65, 32'shec0bf878, 32'shec0d768e, 32'shec0ef4a8, 
               32'shec1072c4, 32'shec11f0e4, 32'shec136f06, 32'shec14ed2c, 32'shec166b55, 32'shec17e981, 32'shec1967b0, 32'shec1ae5e2, 
               32'shec1c6417, 32'shec1de24f, 32'shec1f608a, 32'shec20dec8, 32'shec225d09, 32'shec23db4e, 32'shec255995, 32'shec26d7e0, 
               32'shec28562d, 32'shec29d47e, 32'shec2b52d1, 32'shec2cd128, 32'shec2e4f82, 32'shec2fcddf, 32'shec314c3f, 32'shec32caa2, 
               32'shec344908, 32'shec35c771, 32'shec3745dd, 32'shec38c44c, 32'shec3a42be, 32'shec3bc133, 32'shec3d3fac, 32'shec3ebe27, 
               32'shec403ca5, 32'shec41bb27, 32'shec4339ab, 32'shec44b833, 32'shec4636bd, 32'shec47b54b, 32'shec4933dc, 32'shec4ab26f, 
               32'shec4c3106, 32'shec4dafa0, 32'shec4f2e3d, 32'shec50acdc, 32'shec522b7f, 32'shec53aa25, 32'shec5528ce, 32'shec56a77a, 
               32'shec582629, 32'shec59a4db, 32'shec5b2390, 32'shec5ca248, 32'shec5e2103, 32'shec5f9fc2, 32'shec611e83, 32'shec629d47, 
               32'shec641c0e, 32'shec659ad9, 32'shec6719a6, 32'shec689876, 32'shec6a1749, 32'shec6b9620, 32'shec6d14f9, 32'shec6e93d6, 
               32'shec7012b5, 32'shec719197, 32'shec73107d, 32'shec748f65, 32'shec760e51, 32'shec778d3f, 32'shec790c31, 32'shec7a8b25, 
               32'shec7c0a1d, 32'shec7d8917, 32'shec7f0815, 32'shec808715, 32'shec820619, 32'shec83851f, 32'shec850429, 32'shec868335, 
               32'shec880245, 32'shec898158, 32'shec8b006d, 32'shec8c7f86, 32'shec8dfea1, 32'shec8f7dc0, 32'shec90fce1, 32'shec927c06, 
               32'shec93fb2e, 32'shec957a58, 32'shec96f986, 32'shec9878b6, 32'shec99f7ea, 32'shec9b7720, 32'shec9cf65a, 32'shec9e7596, 
               32'shec9ff4d6, 32'sheca17418, 32'sheca2f35e, 32'sheca472a6, 32'sheca5f1f2, 32'sheca77140, 32'sheca8f091, 32'shecaa6fe6, 
               32'shecabef3d, 32'shecad6e97, 32'shecaeedf5, 32'shecb06d55, 32'shecb1ecb8, 32'shecb36c1f, 32'shecb4eb88, 32'shecb66af4, 
               32'shecb7ea63, 32'shecb969d5, 32'shecbae94b, 32'shecbc68c3, 32'shecbde83e, 32'shecbf67bc, 32'shecc0e73d, 32'shecc266c1, 
               32'shecc3e648, 32'shecc565d2, 32'shecc6e55f, 32'shecc864ee, 32'shecc9e481, 32'sheccb6417, 32'sheccce3b0, 32'shecce634b, 
               32'sheccfe2ea, 32'shecd1628c, 32'shecd2e230, 32'shecd461d8, 32'shecd5e182, 32'shecd76130, 32'shecd8e0e0, 32'shecda6093, 
               32'shecdbe04a, 32'shecdd6003, 32'shecdedfbf, 32'shece05f7e, 32'shece1df40, 32'shece35f06, 32'shece4dece, 32'shece65e98, 
               32'shece7de66, 32'shece95e37, 32'sheceade0b, 32'shecec5de2, 32'shecedddbb, 32'shecef5d98, 32'shecf0dd78, 32'shecf25d5a, 
               32'shecf3dd3f, 32'shecf55d28, 32'shecf6dd13, 32'shecf85d01, 32'shecf9dcf3, 32'shecfb5ce7, 32'shecfcdcde, 32'shecfe5cd8, 
               32'shecffdcd4, 32'shed015cd4, 32'shed02dcd7, 32'shed045cdd, 32'shed05dce5, 32'shed075cf1, 32'shed08dcff, 32'shed0a5d11, 
               32'shed0bdd25, 32'shed0d5d3c, 32'shed0edd56, 32'shed105d74, 32'shed11dd94, 32'shed135db6, 32'shed14dddc, 32'shed165e05, 
               32'shed17de31, 32'shed195e5f, 32'shed1ade91, 32'shed1c5ec5, 32'shed1ddefd, 32'shed1f5f37, 32'shed20df74, 32'shed225fb4, 
               32'shed23dff7, 32'shed25603d, 32'shed26e086, 32'shed2860d1, 32'shed29e120, 32'shed2b6171, 32'shed2ce1c6, 32'shed2e621d, 
               32'shed2fe277, 32'shed3162d4, 32'shed32e334, 32'shed346397, 32'shed35e3fd, 32'shed376466, 32'shed38e4d2, 32'shed3a6540, 
               32'shed3be5b1, 32'shed3d6626, 32'shed3ee69d, 32'shed406717, 32'shed41e794, 32'shed436814, 32'shed44e897, 32'shed46691c, 
               32'shed47e9a5, 32'shed496a30, 32'shed4aeabe, 32'shed4c6b50, 32'shed4debe4, 32'shed4f6c7b, 32'shed50ed14, 32'shed526db1, 
               32'shed53ee51, 32'shed556ef3, 32'shed56ef99, 32'shed587041, 32'shed59f0ec, 32'shed5b719a, 32'shed5cf24b, 32'shed5e72fe, 
               32'shed5ff3b5, 32'shed61746f, 32'shed62f52b, 32'shed6475ea, 32'shed65f6ac, 32'shed677771, 32'shed68f839, 32'shed6a7904, 
               32'shed6bf9d1, 32'shed6d7aa2, 32'shed6efb75, 32'shed707c4b, 32'shed71fd24, 32'shed737e00, 32'shed74fedf, 32'shed767fc0, 
               32'shed7800a5, 32'shed79818c, 32'shed7b0276, 32'shed7c8363, 32'shed7e0453, 32'shed7f8546, 32'shed81063b, 32'shed828734, 
               32'shed84082f, 32'shed85892d, 32'shed870a2e, 32'shed888b32, 32'shed8a0c39, 32'shed8b8d42, 32'shed8d0e4f, 32'shed8e8f5e, 
               32'shed901070, 32'shed919185, 32'shed93129d, 32'shed9493b7, 32'shed9614d5, 32'shed9795f5, 32'shed991718, 32'shed9a983e, 
               32'shed9c1967, 32'shed9d9a92, 32'shed9f1bc1, 32'sheda09cf2, 32'sheda21e26, 32'sheda39f5d, 32'sheda52097, 32'sheda6a1d4, 
               32'sheda82313, 32'sheda9a455, 32'shedab259a, 32'shedaca6e2, 32'shedae282d, 32'shedafa97b, 32'shedb12acb, 32'shedb2ac1e, 
               32'shedb42d74, 32'shedb5aecd, 32'shedb73029, 32'shedb8b187, 32'shedba32e9, 32'shedbbb44d, 32'shedbd35b4, 32'shedbeb71e, 
               32'shedc0388a, 32'shedc1b9fa, 32'shedc33b6c, 32'shedc4bce1, 32'shedc63e59, 32'shedc7bfd3, 32'shedc94151, 32'shedcac2d1, 
               32'shedcc4454, 32'shedcdc5da, 32'shedcf4763, 32'shedd0c8ee, 32'shedd24a7d, 32'shedd3cc0e, 32'shedd54da2, 32'shedd6cf38, 
               32'shedd850d2, 32'shedd9d26e, 32'sheddb540d, 32'sheddcd5af, 32'shedde5754, 32'sheddfd8fb, 32'shede15aa6, 32'shede2dc53, 
               32'shede45e03, 32'shede5dfb5, 32'shede7616b, 32'shede8e323, 32'shedea64de, 32'shedebe69c, 32'sheded685d, 32'shedeeea20, 
               32'shedf06be6, 32'shedf1edaf, 32'shedf36f7b, 32'shedf4f14a, 32'shedf6731b, 32'shedf7f4ef, 32'shedf976c6, 32'shedfaf8a0, 
               32'shedfc7a7c, 32'shedfdfc5b, 32'shedff7e3d, 32'shee010022, 32'shee02820a, 32'shee0403f4, 32'shee0585e1, 32'shee0707d1, 
               32'shee0889c4, 32'shee0a0bb9, 32'shee0b8db1, 32'shee0d0fac, 32'shee0e91aa, 32'shee1013ab, 32'shee1195ae, 32'shee1317b4, 
               32'shee1499bd, 32'shee161bc8, 32'shee179dd7, 32'shee191fe8, 32'shee1aa1fc, 32'shee1c2412, 32'shee1da62c, 32'shee1f2848, 
               32'shee20aa67, 32'shee222c88, 32'shee23aead, 32'shee2530d4, 32'shee26b2fe, 32'shee28352a, 32'shee29b75a, 32'shee2b398c, 
               32'shee2cbbc1, 32'shee2e3df8, 32'shee2fc033, 32'shee314270, 32'shee32c4b0, 32'shee3446f2, 32'shee35c938, 32'shee374b80, 
               32'shee38cdcb, 32'shee3a5018, 32'shee3bd269, 32'shee3d54bc, 32'shee3ed712, 32'shee40596a, 32'shee41dbc6, 32'shee435e24, 
               32'shee44e084, 32'shee4662e8, 32'shee47e54e, 32'shee4967b7, 32'shee4aea23, 32'shee4c6c91, 32'shee4def02, 32'shee4f7176, 
               32'shee50f3ed, 32'shee527666, 32'shee53f8e2, 32'shee557b61, 32'shee56fde3, 32'shee588067, 32'shee5a02ee, 32'shee5b8578, 
               32'shee5d0804, 32'shee5e8a93, 32'shee600d25, 32'shee618fba, 32'shee631251, 32'shee6494eb, 32'shee661788, 32'shee679a27, 
               32'shee691cc9, 32'shee6a9f6e, 32'shee6c2216, 32'shee6da4c0, 32'shee6f276d, 32'shee70aa1d, 32'shee722ccf, 32'shee73af84, 
               32'shee75323c, 32'shee76b4f7, 32'shee7837b4, 32'shee79ba74, 32'shee7b3d36, 32'shee7cbffc, 32'shee7e42c4, 32'shee7fc58f, 
               32'shee81485c, 32'shee82cb2c, 32'shee844dff, 32'shee85d0d4, 32'shee8753ad, 32'shee88d688, 32'shee8a5965, 32'shee8bdc46, 
               32'shee8d5f29, 32'shee8ee20e, 32'shee9064f7, 32'shee91e7e2, 32'shee936acf, 32'shee94edc0, 32'shee9670b3, 32'shee97f3a9, 
               32'shee9976a1, 32'shee9af99d, 32'shee9c7c9a, 32'shee9dff9b, 32'shee9f829e, 32'sheea105a4, 32'sheea288ad, 32'sheea40bb8, 
               32'sheea58ec6, 32'sheea711d6, 32'sheea894ea, 32'sheeaa1800, 32'sheeab9b18, 32'sheead1e34, 32'sheeaea152, 32'sheeb02472, 
               32'sheeb1a796, 32'sheeb32abc, 32'sheeb4ade4, 32'sheeb63110, 32'sheeb7b43e, 32'sheeb9376e, 32'sheebabaa2, 32'sheebc3dd8, 
               32'sheebdc110, 32'sheebf444c, 32'sheec0c78a, 32'sheec24aca, 32'sheec3ce0d, 32'sheec55153, 32'sheec6d49c, 32'sheec857e7, 
               32'sheec9db35, 32'sheecb5e86, 32'sheecce1d9, 32'sheece652f, 32'sheecfe887, 32'sheed16be3, 32'sheed2ef40, 32'sheed472a1, 
               32'sheed5f604, 32'sheed7796a, 32'sheed8fcd2, 32'sheeda803d, 32'sheedc03ab, 32'sheedd871b, 32'sheedf0a8e, 32'sheee08e04, 
               32'sheee2117c, 32'sheee394f7, 32'sheee51875, 32'sheee69bf5, 32'sheee81f78, 32'sheee9a2fd, 32'sheeeb2685, 32'sheeecaa10, 
               32'sheeee2d9d, 32'sheeefb12d, 32'sheef134c0, 32'sheef2b855, 32'sheef43bed, 32'sheef5bf88, 32'sheef74325, 32'sheef8c6c5, 
               32'sheefa4a67, 32'sheefbce0c, 32'sheefd51b4, 32'sheefed55e, 32'shef00590b, 32'shef01dcba, 32'shef03606c, 32'shef04e421, 
               32'shef0667d9, 32'shef07eb93, 32'shef096f4f, 32'shef0af30e, 32'shef0c76d0, 32'shef0dfa95, 32'shef0f7e5c, 32'shef110225, 
               32'shef1285f2, 32'shef1409c1, 32'shef158d92, 32'shef171166, 32'shef18953d, 32'shef1a1916, 32'shef1b9cf2, 32'shef1d20d1, 
               32'shef1ea4b2, 32'shef202896, 32'shef21ac7c, 32'shef233065, 32'shef24b451, 32'shef26383f, 32'shef27bc2f, 32'shef294023, 
               32'shef2ac419, 32'shef2c4811, 32'shef2dcc0c, 32'shef2f500a, 32'shef30d40a, 32'shef32580d, 32'shef33dc13, 32'shef35601b, 
               32'shef36e426, 32'shef386833, 32'shef39ec43, 32'shef3b7055, 32'shef3cf46a, 32'shef3e7882, 32'shef3ffc9c, 32'shef4180b9, 
               32'shef4304d8, 32'shef4488fa, 32'shef460d1f, 32'shef479146, 32'shef491570, 32'shef4a999c, 32'shef4c1dcb, 32'shef4da1fc, 
               32'shef4f2630, 32'shef50aa67, 32'shef522ea0, 32'shef53b2dc, 32'shef55371a, 32'shef56bb5b, 32'shef583f9e, 32'shef59c3e4, 
               32'shef5b482d, 32'shef5ccc78, 32'shef5e50c6, 32'shef5fd516, 32'shef615969, 32'shef62ddbe, 32'shef646216, 32'shef65e670, 
               32'shef676ace, 32'shef68ef2d, 32'shef6a738f, 32'shef6bf7f4, 32'shef6d7c5b, 32'shef6f00c5, 32'shef708532, 32'shef7209a1, 
               32'shef738e12, 32'shef751286, 32'shef7696fd, 32'shef781b76, 32'shef799ff2, 32'shef7b2470, 32'shef7ca8f1, 32'shef7e2d74, 
               32'shef7fb1fa, 32'shef813683, 32'shef82bb0e, 32'shef843f9b, 32'shef85c42b, 32'shef8748be, 32'shef88cd53, 32'shef8a51eb, 
               32'shef8bd685, 32'shef8d5b22, 32'shef8edfc1, 32'shef906463, 32'shef91e907, 32'shef936dae, 32'shef94f258, 32'shef967704, 
               32'shef97fbb2, 32'shef998063, 32'shef9b0517, 32'shef9c89cd, 32'shef9e0e85, 32'shef9f9341, 32'shefa117fe, 32'shefa29cbe, 
               32'shefa42181, 32'shefa5a646, 32'shefa72b0e, 32'shefa8afd9, 32'shefaa34a5, 32'shefabb975, 32'shefad3e47, 32'shefaec31b, 
               32'shefb047f2, 32'shefb1cccb, 32'shefb351a7, 32'shefb4d686, 32'shefb65b66, 32'shefb7e04a, 32'shefb96530, 32'shefbaea18, 
               32'shefbc6f03, 32'shefbdf3f1, 32'shefbf78e1, 32'shefc0fdd3, 32'shefc282c8, 32'shefc407c0, 32'shefc58cba, 32'shefc711b6, 
               32'shefc896b5, 32'shefca1bb7, 32'shefcba0bb, 32'shefcd25c1, 32'shefceaacb, 32'shefd02fd6, 32'shefd1b4e4, 32'shefd339f5, 
               32'shefd4bf08, 32'shefd6441d, 32'shefd7c935, 32'shefd94e50, 32'shefdad36c, 32'shefdc588c, 32'shefddddae, 32'shefdf62d2, 
               32'shefe0e7f9, 32'shefe26d23, 32'shefe3f24f, 32'shefe5777d, 32'shefe6fcae, 32'shefe881e1, 32'shefea0717, 32'shefeb8c4f, 
               32'shefed118a, 32'shefee96c7, 32'sheff01c07, 32'sheff1a149, 32'sheff3268e, 32'sheff4abd5, 32'sheff6311f, 32'sheff7b66b, 
               32'sheff93bba, 32'sheffac10b, 32'sheffc465e, 32'sheffdcbb4, 32'shefff510d, 32'shf000d668, 32'shf0025bc5, 32'shf003e125, 
               32'shf0056687, 32'shf006ebec, 32'shf0087153, 32'shf009f6bd, 32'shf00b7c29, 32'shf00d0198, 32'shf00e8709, 32'shf0100c7d, 
               32'shf01191f3, 32'shf013176b, 32'shf0149ce6, 32'shf0162263, 32'shf017a7e3, 32'shf0192d66, 32'shf01ab2ea, 32'shf01c3871, 
               32'shf01dbdfb, 32'shf01f4387, 32'shf020c916, 32'shf0224ea7, 32'shf023d43a, 32'shf02559d0, 32'shf026df68, 32'shf0286503, 
               32'shf029eaa1, 32'shf02b7040, 32'shf02cf5e2, 32'shf02e7b87, 32'shf030012e, 32'shf03186d7, 32'shf0330c83, 32'shf0349231, 
               32'shf03617e2, 32'shf0379d95, 32'shf039234b, 32'shf03aa903, 32'shf03c2ebd, 32'shf03db47a, 32'shf03f3a3a, 32'shf040bffb, 
               32'shf04245c0, 32'shf043cb86, 32'shf045514f, 32'shf046d71b, 32'shf0485ce9, 32'shf049e2b9, 32'shf04b688c, 32'shf04cee61, 
               32'shf04e7438, 32'shf04ffa12, 32'shf0517fef, 32'shf05305ce, 32'shf0548baf, 32'shf0561193, 32'shf0579779, 32'shf0591d61, 
               32'shf05aa34c, 32'shf05c293a, 32'shf05daf29, 32'shf05f351b, 32'shf060bb10, 32'shf0624107, 32'shf063c700, 32'shf0654cfc, 
               32'shf066d2fa, 32'shf06858fb, 32'shf069defe, 32'shf06b6503, 32'shf06ceb0b, 32'shf06e7115, 32'shf06ff722, 32'shf0717d31, 
               32'shf0730342, 32'shf0748956, 32'shf0760f6c, 32'shf0779585, 32'shf0791ba0, 32'shf07aa1bd, 32'shf07c27dd, 32'shf07dadff, 
               32'shf07f3424, 32'shf080ba4b, 32'shf0824074, 32'shf083c6a0, 32'shf0854cce, 32'shf086d2ff, 32'shf0885932, 32'shf089df67, 
               32'shf08b659f, 32'shf08cebd9, 32'shf08e7215, 32'shf08ff854, 32'shf0917e95, 32'shf09304d9, 32'shf0948b1f, 32'shf0961167, 
               32'shf09797b2, 32'shf0991dff, 32'shf09aa44e, 32'shf09c2aa0, 32'shf09db0f4, 32'shf09f374b, 32'shf0a0bda4, 32'shf0a243ff, 
               32'shf0a3ca5d, 32'shf0a550bd, 32'shf0a6d71f, 32'shf0a85d84, 32'shf0a9e3eb, 32'shf0ab6a55, 32'shf0acf0c1, 32'shf0ae772f, 
               32'shf0affda0, 32'shf0b18413, 32'shf0b30a88, 32'shf0b49100, 32'shf0b6177a, 32'shf0b79df6, 32'shf0b92475, 32'shf0baaaf6, 
               32'shf0bc317a, 32'shf0bdb7ff, 32'shf0bf3e88, 32'shf0c0c512, 32'shf0c24b9f, 32'shf0c3d22e, 32'shf0c558c0, 32'shf0c6df54, 
               32'shf0c865ea, 32'shf0c9ec83, 32'shf0cb731e, 32'shf0ccf9bb, 32'shf0ce805b, 32'shf0d006fd, 32'shf0d18da1, 32'shf0d31448, 
               32'shf0d49af1, 32'shf0d6219c, 32'shf0d7a84a, 32'shf0d92efa, 32'shf0dab5ad, 32'shf0dc3c61, 32'shf0ddc318, 32'shf0df49d2, 
               32'shf0e0d08d, 32'shf0e2574c, 32'shf0e3de0c, 32'shf0e564cf, 32'shf0e6eb94, 32'shf0e8725b, 32'shf0e9f925, 32'shf0eb7ff1, 
               32'shf0ed06bf, 32'shf0ee8d90, 32'shf0f01463, 32'shf0f19b38, 32'shf0f32210, 32'shf0f4a8ea, 32'shf0f62fc6, 32'shf0f7b6a5, 
               32'shf0f93d86, 32'shf0fac469, 32'shf0fc4b4f, 32'shf0fdd236, 32'shf0ff5921, 32'shf100e00d, 32'shf10266fc, 32'shf103eded, 
               32'shf10574e0, 32'shf106fbd6, 32'shf10882ce, 32'shf10a09c9, 32'shf10b90c5, 32'shf10d17c4, 32'shf10e9ec6, 32'shf11025c9, 
               32'shf111accf, 32'shf11333d7, 32'shf114bae2, 32'shf11641ef, 32'shf117c8fe, 32'shf119500f, 32'shf11ad723, 32'shf11c5e39, 
               32'shf11de551, 32'shf11f6c6c, 32'shf120f389, 32'shf1227aa8, 32'shf12401c9, 32'shf12588ed, 32'shf1271013, 32'shf128973b, 
               32'shf12a1e66, 32'shf12ba593, 32'shf12d2cc2, 32'shf12eb3f4, 32'shf1303b27, 32'shf131c25d, 32'shf1334996, 32'shf134d0d0, 
               32'shf136580d, 32'shf137df4d, 32'shf139668e, 32'shf13aedd2, 32'shf13c7518, 32'shf13dfc60, 32'shf13f83ab, 32'shf1410af8, 
               32'shf1429247, 32'shf1441998, 32'shf145a0ec, 32'shf1472842, 32'shf148af9a, 32'shf14a36f4, 32'shf14bbe51, 32'shf14d45b0, 
               32'shf14ecd11, 32'shf1505475, 32'shf151dbdb, 32'shf1536343, 32'shf154eaad, 32'shf156721a, 32'shf157f989, 32'shf15980fa, 
               32'shf15b086d, 32'shf15c8fe3, 32'shf15e175b, 32'shf15f9ed5, 32'shf1612651, 32'shf162add0, 32'shf1643551, 32'shf165bcd4, 
               32'shf1674459, 32'shf168cbe1, 32'shf16a536b, 32'shf16bdaf7, 32'shf16d6286, 32'shf16eea16, 32'shf17071a9, 32'shf171f93e, 
               32'shf17380d6, 32'shf175086f, 32'shf176900b, 32'shf17817a9, 32'shf1799f4a, 32'shf17b26ec, 32'shf17cae91, 32'shf17e3638, 
               32'shf17fbde2, 32'shf181458d, 32'shf182cd3b, 32'shf18454eb, 32'shf185dc9d, 32'shf1876452, 32'shf188ec09, 32'shf18a73c2, 
               32'shf18bfb7d, 32'shf18d833a, 32'shf18f0afa, 32'shf19092bc, 32'shf1921a80, 32'shf193a246, 32'shf1952a0f, 32'shf196b1d9, 
               32'shf19839a6, 32'shf199c176, 32'shf19b4947, 32'shf19cd11b, 32'shf19e58f1, 32'shf19fe0c9, 32'shf1a168a3, 32'shf1a2f080, 
               32'shf1a4785e, 32'shf1a6003f, 32'shf1a78822, 32'shf1a91008, 32'shf1aa97ef, 32'shf1ac1fd9, 32'shf1ada7c5, 32'shf1af2fb3, 
               32'shf1b0b7a4, 32'shf1b23f97, 32'shf1b3c78b, 32'shf1b54f82, 32'shf1b6d77c, 32'shf1b85f77, 32'shf1b9e775, 32'shf1bb6f75, 
               32'shf1bcf777, 32'shf1be7f7b, 32'shf1c00781, 32'shf1c18f8a, 32'shf1c31795, 32'shf1c49fa2, 32'shf1c627b1, 32'shf1c7afc3, 
               32'shf1c937d6, 32'shf1cabfec, 32'shf1cc4804, 32'shf1cdd01e, 32'shf1cf583b, 32'shf1d0e059, 32'shf1d2687a, 32'shf1d3f09d, 
               32'shf1d578c2, 32'shf1d700ea, 32'shf1d88913, 32'shf1da113f, 32'shf1db996d, 32'shf1dd219d, 32'shf1dea9cf, 32'shf1e03203, 
               32'shf1e1ba3a, 32'shf1e34273, 32'shf1e4caae, 32'shf1e652eb, 32'shf1e7db2a, 32'shf1e9636b, 32'shf1eaebaf, 32'shf1ec73f5, 
               32'shf1edfc3d, 32'shf1ef8487, 32'shf1f10cd3, 32'shf1f29522, 32'shf1f41d72, 32'shf1f5a5c5, 32'shf1f72e1a, 32'shf1f8b671, 
               32'shf1fa3ecb, 32'shf1fbc726, 32'shf1fd4f84, 32'shf1fed7e4, 32'shf2006046, 32'shf201e8aa, 32'shf2037110, 32'shf204f978, 
               32'shf20681e3, 32'shf2080a50, 32'shf20992bf, 32'shf20b1b30, 32'shf20ca3a3, 32'shf20e2c18, 32'shf20fb490, 32'shf2113d09, 
               32'shf212c585, 32'shf2144e03, 32'shf215d683, 32'shf2175f06, 32'shf218e78a, 32'shf21a7010, 32'shf21bf899, 32'shf21d8124, 
               32'shf21f09b1, 32'shf2209240, 32'shf2221ad1, 32'shf223a365, 32'shf2252bfa, 32'shf226b492, 32'shf2283d2c, 32'shf229c5c7, 
               32'shf22b4e66, 32'shf22cd706, 32'shf22e5fa8, 32'shf22fe84c, 32'shf23170f3, 32'shf232f99c, 32'shf2348247, 32'shf2360af4, 
               32'shf23793a3, 32'shf2391c54, 32'shf23aa507, 32'shf23c2dbd, 32'shf23db674, 32'shf23f3f2e, 32'shf240c7ea, 32'shf24250a8, 
               32'shf243d968, 32'shf245622a, 32'shf246eaee, 32'shf24873b5, 32'shf249fc7d, 32'shf24b8548, 32'shf24d0e15, 32'shf24e96e4, 
               32'shf2501fb5, 32'shf251a888, 32'shf253315d, 32'shf254ba34, 32'shf256430e, 32'shf257cbe9, 32'shf25954c7, 32'shf25adda7, 
               32'shf25c6688, 32'shf25def6c, 32'shf25f7852, 32'shf261013b, 32'shf2628a25, 32'shf2641311, 32'shf2659c00, 32'shf26724f0, 
               32'shf268ade3, 32'shf26a36d8, 32'shf26bbfce, 32'shf26d48c7, 32'shf26ed1c2, 32'shf2705abf, 32'shf271e3bf, 32'shf2736cc0, 
               32'shf274f5c3, 32'shf2767ec9, 32'shf27807d0, 32'shf27990da, 32'shf27b19e6, 32'shf27ca2f4, 32'shf27e2c04, 32'shf27fb516, 
               32'shf2813e2a, 32'shf282c740, 32'shf2845058, 32'shf285d972, 32'shf287628f, 32'shf288ebad, 32'shf28a74ce, 32'shf28bfdf0, 
               32'shf28d8715, 32'shf28f103c, 32'shf2909965, 32'shf2922290, 32'shf293abbd, 32'shf29534ec, 32'shf296be1d, 32'shf2984750, 
               32'shf299d085, 32'shf29b59bc, 32'shf29ce2f6, 32'shf29e6c31, 32'shf29ff56f, 32'shf2a17eae, 32'shf2a307f0, 32'shf2a49134, 
               32'shf2a61a7a, 32'shf2a7a3c1, 32'shf2a92d0b, 32'shf2aab657, 32'shf2ac3fa5, 32'shf2adc8f5, 32'shf2af5247, 32'shf2b0db9b, 
               32'shf2b264f2, 32'shf2b3ee4a, 32'shf2b577a4, 32'shf2b70101, 32'shf2b88a5f, 32'shf2ba13c0, 32'shf2bb9d22, 32'shf2bd2687, 
               32'shf2beafed, 32'shf2c03956, 32'shf2c1c2c0, 32'shf2c34c2d, 32'shf2c4d59c, 32'shf2c65f0d, 32'shf2c7e880, 32'shf2c971f5, 
               32'shf2cafb6b, 32'shf2cc84e4, 32'shf2ce0e5f, 32'shf2cf97dc, 32'shf2d1215b, 32'shf2d2aadd, 32'shf2d43460, 32'shf2d5bde5, 
               32'shf2d7476c, 32'shf2d8d0f5, 32'shf2da5a81, 32'shf2dbe40e, 32'shf2dd6d9d, 32'shf2def72e, 32'shf2e080c2, 32'shf2e20a57, 
               32'shf2e393ef, 32'shf2e51d88, 32'shf2e6a723, 32'shf2e830c1, 32'shf2e9ba60, 32'shf2eb4402, 32'shf2eccda5, 32'shf2ee574b, 
               32'shf2efe0f2, 32'shf2f16a9c, 32'shf2f2f448, 32'shf2f47df5, 32'shf2f607a5, 32'shf2f79156, 32'shf2f91b0a, 32'shf2faa4c0, 
               32'shf2fc2e77, 32'shf2fdb831, 32'shf2ff41ed, 32'shf300cbaa, 32'shf302556a, 32'shf303df2c, 32'shf30568ef, 32'shf306f2b5, 
               32'shf3087c7d, 32'shf30a0646, 32'shf30b9012, 32'shf30d19e0, 32'shf30ea3af, 32'shf3102d81, 32'shf311b755, 32'shf313412a, 
               32'shf314cb02, 32'shf31654db, 32'shf317deb7, 32'shf3196895, 32'shf31af274, 32'shf31c7c56, 32'shf31e0639, 32'shf31f901f, 
               32'shf3211a07, 32'shf322a3f0, 32'shf3242ddc, 32'shf325b7c9, 32'shf32741b9, 32'shf328cbaa, 32'shf32a559e, 32'shf32bdf93, 
               32'shf32d698a, 32'shf32ef384, 32'shf3307d7f, 32'shf332077c, 32'shf333917c, 32'shf3351b7d, 32'shf336a580, 32'shf3382f86, 
               32'shf339b98d, 32'shf33b4396, 32'shf33ccda1, 32'shf33e57ae, 32'shf33fe1bd, 32'shf3416bce, 32'shf342f5e1, 32'shf3447ff6, 
               32'shf3460a0d, 32'shf3479426, 32'shf3491e41, 32'shf34aa85e, 32'shf34c327c, 32'shf34dbc9d, 32'shf34f46c0, 32'shf350d0e5, 
               32'shf3525b0b, 32'shf353e534, 32'shf3556f5e, 32'shf356f98b, 32'shf35883b9, 32'shf35a0de9, 32'shf35b981c, 32'shf35d2250, 
               32'shf35eac86, 32'shf36036be, 32'shf361c0f9, 32'shf3634b35, 32'shf364d573, 32'shf3665fb3, 32'shf367e9f4, 32'shf3697438, 
               32'shf36afe7e, 32'shf36c88c6, 32'shf36e130f, 32'shf36f9d5b, 32'shf37127a9, 32'shf372b1f8, 32'shf3743c49, 32'shf375c69d, 
               32'shf37750f2, 32'shf378db49, 32'shf37a65a2, 32'shf37beffe, 32'shf37d7a5b, 32'shf37f04b9, 32'shf3808f1a, 32'shf382197d, 
               32'shf383a3e2, 32'shf3852e48, 32'shf386b8b1, 32'shf388431b, 32'shf389cd88, 32'shf38b57f6, 32'shf38ce266, 32'shf38e6cd9, 
               32'shf38ff74d, 32'shf39181c3, 32'shf3930c3b, 32'shf39496b4, 32'shf3962130, 32'shf397abae, 32'shf399362d, 32'shf39ac0af, 
               32'shf39c4b32, 32'shf39dd5b8, 32'shf39f603f, 32'shf3a0eac8, 32'shf3a27553, 32'shf3a3ffe0, 32'shf3a58a6f, 32'shf3a71500, 
               32'shf3a89f92, 32'shf3aa2a27, 32'shf3abb4bd, 32'shf3ad3f56, 32'shf3aec9f0, 32'shf3b0548c, 32'shf3b1df2a, 32'shf3b369ca, 
               32'shf3b4f46c, 32'shf3b67f10, 32'shf3b809b6, 32'shf3b9945d, 32'shf3bb1f07, 32'shf3bca9b2, 32'shf3be345f, 32'shf3bfbf0e, 
               32'shf3c149bf, 32'shf3c2d472, 32'shf3c45f27, 32'shf3c5e9de, 32'shf3c77496, 32'shf3c8ff51, 32'shf3ca8a0d, 32'shf3cc14cb, 
               32'shf3cd9f8b, 32'shf3cf2a4d, 32'shf3d0b511, 32'shf3d23fd7, 32'shf3d3ca9e, 32'shf3d55568, 32'shf3d6e033, 32'shf3d86b00, 
               32'shf3d9f5cf, 32'shf3db80a0, 32'shf3dd0b73, 32'shf3de9648, 32'shf3e0211f, 32'shf3e1abf7, 32'shf3e336d1, 32'shf3e4c1ae, 
               32'shf3e64c8c, 32'shf3e7d76c, 32'shf3e9624d, 32'shf3eaed31, 32'shf3ec7817, 32'shf3ee02fe, 32'shf3ef8de7, 32'shf3f118d2, 
               32'shf3f2a3bf, 32'shf3f42eae, 32'shf3f5b99f, 32'shf3f74491, 32'shf3f8cf86, 32'shf3fa5a7c, 32'shf3fbe574, 32'shf3fd706e, 
               32'shf3fefb6a, 32'shf4008668, 32'shf4021167, 32'shf4039c68, 32'shf405276c, 32'shf406b271, 32'shf4083d78, 32'shf409c880, 
               32'shf40b538b, 32'shf40cde97, 32'shf40e69a6, 32'shf40ff4b6, 32'shf4117fc8, 32'shf4130adc, 32'shf41495f1, 32'shf4162109, 
               32'shf417ac22, 32'shf419373d, 32'shf41ac25a, 32'shf41c4d79, 32'shf41dd89a, 32'shf41f63bc, 32'shf420eee1, 32'shf4227a07, 
               32'shf424052f, 32'shf4259058, 32'shf4271b84, 32'shf428a6b2, 32'shf42a31e1, 32'shf42bbd12, 32'shf42d4845, 32'shf42ed37a, 
               32'shf4305eb0, 32'shf431e9e9, 32'shf4337523, 32'shf435005f, 32'shf4368b9d, 32'shf43816dd, 32'shf439a21e, 32'shf43b2d61, 
               32'shf43cb8a7, 32'shf43e43ed, 32'shf43fcf36, 32'shf4415a81, 32'shf442e5cd, 32'shf444711b, 32'shf445fc6b, 32'shf44787bd, 
               32'shf4491311, 32'shf44a9e66, 32'shf44c29be, 32'shf44db517, 32'shf44f4071, 32'shf450cbce, 32'shf452572c, 32'shf453e28d, 
               32'shf4556def, 32'shf456f953, 32'shf45884b8, 32'shf45a1020, 32'shf45b9b89, 32'shf45d26f4, 32'shf45eb261, 32'shf4603dcf, 
               32'shf461c940, 32'shf46354b2, 32'shf464e026, 32'shf4666b9c, 32'shf467f713, 32'shf469828d, 32'shf46b0e08, 32'shf46c9985, 
               32'shf46e2504, 32'shf46fb084, 32'shf4713c06, 32'shf472c78a, 32'shf4745310, 32'shf475de98, 32'shf4776a21, 32'shf478f5ad, 
               32'shf47a8139, 32'shf47c0cc8, 32'shf47d9859, 32'shf47f23eb, 32'shf480af7f, 32'shf4823b15, 32'shf483c6ad, 32'shf4855246, 
               32'shf486dde1, 32'shf488697e, 32'shf489f51d, 32'shf48b80bd, 32'shf48d0c5f, 32'shf48e9803, 32'shf49023a9, 32'shf491af51, 
               32'shf4933afa, 32'shf494c6a5, 32'shf4965252, 32'shf497de00, 32'shf49969b1, 32'shf49af563, 32'shf49c8117, 32'shf49e0ccc, 
               32'shf49f9884, 32'shf4a1243d, 32'shf4a2aff8, 32'shf4a43bb4, 32'shf4a5c773, 32'shf4a75333, 32'shf4a8def5, 32'shf4aa6ab8, 
               32'shf4abf67e, 32'shf4ad8245, 32'shf4af0e0d, 32'shf4b099d8, 32'shf4b225a4, 32'shf4b3b173, 32'shf4b53d42, 32'shf4b6c914, 
               32'shf4b854e7, 32'shf4b9e0bc, 32'shf4bb6c93, 32'shf4bcf86c, 32'shf4be8446, 32'shf4c01022, 32'shf4c19c00, 32'shf4c327df, 
               32'shf4c4b3c0, 32'shf4c63fa3, 32'shf4c7cb88, 32'shf4c9576e, 32'shf4cae356, 32'shf4cc6f40, 32'shf4cdfb2c, 32'shf4cf8719, 
               32'shf4d11308, 32'shf4d29ef9, 32'shf4d42aeb, 32'shf4d5b6e0, 32'shf4d742d6, 32'shf4d8cecd, 32'shf4da5ac7, 32'shf4dbe6c2, 
               32'shf4dd72be, 32'shf4defebd, 32'shf4e08abd, 32'shf4e216bf, 32'shf4e3a2c3, 32'shf4e52ec8, 32'shf4e6bacf, 32'shf4e846d8, 
               32'shf4e9d2e3, 32'shf4eb5eef, 32'shf4eceafd, 32'shf4ee770c, 32'shf4f0031e, 32'shf4f18f31, 32'shf4f31b46, 32'shf4f4a75c, 
               32'shf4f63374, 32'shf4f7bf8e, 32'shf4f94baa, 32'shf4fad7c7, 32'shf4fc63e6, 32'shf4fdf007, 32'shf4ff7c29, 32'shf501084d, 
               32'shf5029473, 32'shf504209a, 32'shf505acc3, 32'shf50738ee, 32'shf508c51b, 32'shf50a5149, 32'shf50bdd79, 32'shf50d69aa, 
               32'shf50ef5de, 32'shf5108213, 32'shf5120e49, 32'shf5139a82, 32'shf51526bc, 32'shf516b2f7, 32'shf5183f35, 32'shf519cb74, 
               32'shf51b57b5, 32'shf51ce3f7, 32'shf51e703b, 32'shf51ffc81, 32'shf52188c9, 32'shf5231512, 32'shf524a15d, 32'shf5262da9, 
               32'shf527b9f7, 32'shf5294647, 32'shf52ad299, 32'shf52c5eec, 32'shf52deb41, 32'shf52f7797, 32'shf53103ef, 32'shf5329049, 
               32'shf5341ca5, 32'shf535a902, 32'shf5373561, 32'shf538c1c1, 32'shf53a4e24, 32'shf53bda87, 32'shf53d66ed, 32'shf53ef354, 
               32'shf5407fbd, 32'shf5420c27, 32'shf5439893, 32'shf5452501, 32'shf546b171, 32'shf5483de2, 32'shf549ca55, 32'shf54b56c9, 
               32'shf54ce33f, 32'shf54e6fb7, 32'shf54ffc30, 32'shf55188ab, 32'shf5531528, 32'shf554a1a6, 32'shf5562e26, 32'shf557baa8, 
               32'shf559472b, 32'shf55ad3b0, 32'shf55c6036, 32'shf55decbe, 32'shf55f7948, 32'shf56105d4, 32'shf5629261, 32'shf5641eef, 
               32'shf565ab80, 32'shf5673812, 32'shf568c4a5, 32'shf56a513b, 32'shf56bddd1, 32'shf56d6a6a, 32'shf56ef704, 32'shf57083a0, 
               32'shf572103d, 32'shf5739cdc, 32'shf575297d, 32'shf576b61f, 32'shf57842c3, 32'shf579cf69, 32'shf57b5c10, 32'shf57ce8b9, 
               32'shf57e7563, 32'shf580020f, 32'shf5818ebd, 32'shf5831b6c, 32'shf584a81d, 32'shf58634cf, 32'shf587c183, 32'shf5894e39, 
               32'shf58adaf0, 32'shf58c67a9, 32'shf58df464, 32'shf58f8120, 32'shf5910dde, 32'shf5929a9d, 32'shf594275e, 32'shf595b421, 
               32'shf59740e5, 32'shf598cdab, 32'shf59a5a72, 32'shf59be73b, 32'shf59d7406, 32'shf59f00d2, 32'shf5a08da0, 32'shf5a21a6f, 
               32'shf5a3a740, 32'shf5a53413, 32'shf5a6c0e7, 32'shf5a84dbd, 32'shf5a9da94, 32'shf5ab676d, 32'shf5acf448, 32'shf5ae8124, 
               32'shf5b00e02, 32'shf5b19ae1, 32'shf5b327c2, 32'shf5b4b4a5, 32'shf5b64189, 32'shf5b7ce6f, 32'shf5b95b56, 32'shf5bae83f, 
               32'shf5bc7529, 32'shf5be0215, 32'shf5bf8f03, 32'shf5c11bf2, 32'shf5c2a8e3, 32'shf5c435d5, 32'shf5c5c2c9, 32'shf5c74fbf, 
               32'shf5c8dcb6, 32'shf5ca69af, 32'shf5cbf6a9, 32'shf5cd83a5, 32'shf5cf10a2, 32'shf5d09da1, 32'shf5d22aa2, 32'shf5d3b7a4, 
               32'shf5d544a7, 32'shf5d6d1ad, 32'shf5d85eb3, 32'shf5d9ebbc, 32'shf5db78c6, 32'shf5dd05d1, 32'shf5de92de, 32'shf5e01fed, 
               32'shf5e1acfd, 32'shf5e33a0f, 32'shf5e4c722, 32'shf5e65437, 32'shf5e7e14e, 32'shf5e96e66, 32'shf5eafb7f, 32'shf5ec889a, 
               32'shf5ee15b7, 32'shf5efa2d5, 32'shf5f12ff5, 32'shf5f2bd16, 32'shf5f44a39, 32'shf5f5d75e, 32'shf5f76484, 32'shf5f8f1ab, 
               32'shf5fa7ed4, 32'shf5fc0bff, 32'shf5fd992b, 32'shf5ff2659, 32'shf600b388, 32'shf60240b9, 32'shf603cdeb, 32'shf6055b1f, 
               32'shf606e854, 32'shf608758b, 32'shf60a02c3, 32'shf60b8ffd, 32'shf60d1d39, 32'shf60eaa76, 32'shf61037b5, 32'shf611c4f5, 
               32'shf6135237, 32'shf614df7a, 32'shf6166cbe, 32'shf617fa05, 32'shf619874c, 32'shf61b1496, 32'shf61ca1e1, 32'shf61e2f2d, 
               32'shf61fbc7b, 32'shf62149ca, 32'shf622d71b, 32'shf624646e, 32'shf625f1c2, 32'shf6277f17, 32'shf6290c6e, 32'shf62a99c7, 
               32'shf62c2721, 32'shf62db47c, 32'shf62f41d9, 32'shf630cf38, 32'shf6325c98, 32'shf633e9fa, 32'shf635775d, 32'shf63704c1, 
               32'shf6389228, 32'shf63a1f8f, 32'shf63bacf8, 32'shf63d3a63, 32'shf63ec7cf, 32'shf640553d, 32'shf641e2ac, 32'shf643701d, 
               32'shf644fd8f, 32'shf6468b03, 32'shf6481878, 32'shf649a5ef, 32'shf64b3367, 32'shf64cc0e0, 32'shf64e4e5c, 32'shf64fdbd8, 
               32'shf6516956, 32'shf652f6d6, 32'shf6548457, 32'shf65611da, 32'shf6579f5e, 32'shf6592ce4, 32'shf65aba6b, 32'shf65c47f3, 
               32'shf65dd57d, 32'shf65f6309, 32'shf660f096, 32'shf6627e24, 32'shf6640bb4, 32'shf6659946, 32'shf66726d9, 32'shf668b46d, 
               32'shf66a4203, 32'shf66bcf9b, 32'shf66d5d34, 32'shf66eeace, 32'shf670786a, 32'shf6720607, 32'shf67393a6, 32'shf6752146, 
               32'shf676aee8, 32'shf6783c8b, 32'shf679ca30, 32'shf67b57d6, 32'shf67ce57e, 32'shf67e7327, 32'shf68000d1, 32'shf6818e7d, 
               32'shf6831c2b, 32'shf684a9da, 32'shf686378a, 32'shf687c53c, 32'shf68952ef, 32'shf68ae0a4, 32'shf68c6e5a, 32'shf68dfc12, 
               32'shf68f89cb, 32'shf6911786, 32'shf692a542, 32'shf69432ff, 32'shf695c0be, 32'shf6974e7f, 32'shf698dc41, 32'shf69a6a04, 
               32'shf69bf7c9, 32'shf69d858f, 32'shf69f1357, 32'shf6a0a120, 32'shf6a22eea, 32'shf6a3bcb6, 32'shf6a54a84, 32'shf6a6d853, 
               32'shf6a86623, 32'shf6a9f3f5, 32'shf6ab81c8, 32'shf6ad0f9d, 32'shf6ae9d73, 32'shf6b02b4a, 32'shf6b1b923, 32'shf6b346fe, 
               32'shf6b4d4d9, 32'shf6b662b7, 32'shf6b7f095, 32'shf6b97e76, 32'shf6bb0c57, 32'shf6bc9a3a, 32'shf6be281e, 32'shf6bfb604, 
               32'shf6c143ec, 32'shf6c2d1d4, 32'shf6c45fbe, 32'shf6c5edaa, 32'shf6c77b97, 32'shf6c90985, 32'shf6ca9775, 32'shf6cc2566, 
               32'shf6cdb359, 32'shf6cf414d, 32'shf6d0cf43, 32'shf6d25d39, 32'shf6d3eb32, 32'shf6d5792c, 32'shf6d70727, 32'shf6d89523, 
               32'shf6da2321, 32'shf6dbb121, 32'shf6dd3f21, 32'shf6decd24, 32'shf6e05b27, 32'shf6e1e92c, 32'shf6e37733, 32'shf6e5053a, 
               32'shf6e69344, 32'shf6e8214e, 32'shf6e9af5a, 32'shf6eb3d68, 32'shf6eccb77, 32'shf6ee5987, 32'shf6efe798, 32'shf6f175ac, 
               32'shf6f303c0, 32'shf6f491d6, 32'shf6f61fed, 32'shf6f7ae06, 32'shf6f93c20, 32'shf6faca3b, 32'shf6fc5858, 32'shf6fde676, 
               32'shf6ff7496, 32'shf70102b6, 32'shf70290d9, 32'shf7041efd, 32'shf705ad22, 32'shf7073b48, 32'shf708c970, 32'shf70a5799, 
               32'shf70be5c4, 32'shf70d73f0, 32'shf70f021d, 32'shf710904c, 32'shf7121e7c, 32'shf713acae, 32'shf7153ae1, 32'shf716c915, 
               32'shf718574b, 32'shf719e582, 32'shf71b73ba, 32'shf71d01f4, 32'shf71e902f, 32'shf7201e6c, 32'shf721acaa, 32'shf7233ae9, 
               32'shf724c92a, 32'shf726576c, 32'shf727e5af, 32'shf72973f4, 32'shf72b023a, 32'shf72c9081, 32'shf72e1eca, 32'shf72fad14, 
               32'shf7313b60, 32'shf732c9ad, 32'shf73457fb, 32'shf735e64a, 32'shf737749b, 32'shf73902ee, 32'shf73a9141, 32'shf73c1f96, 
               32'shf73daded, 32'shf73f3c44, 32'shf740ca9d, 32'shf74258f8, 32'shf743e754, 32'shf74575b1, 32'shf747040f, 32'shf748926f, 
               32'shf74a20d0, 32'shf74baf33, 32'shf74d3d96, 32'shf74ecbfc, 32'shf7505a62, 32'shf751e8ca, 32'shf7537733, 32'shf755059e, 
               32'shf756940a, 32'shf7582277, 32'shf759b0e5, 32'shf75b3f55, 32'shf75ccdc6, 32'shf75e5c39, 32'shf75feaad, 32'shf7617922, 
               32'shf7630799, 32'shf7649610, 32'shf766248a, 32'shf767b304, 32'shf7694180, 32'shf76acffd, 32'shf76c5e7c, 32'shf76decfb, 
               32'shf76f7b7d, 32'shf77109ff, 32'shf7729883, 32'shf7742708, 32'shf775b58e, 32'shf7774416, 32'shf778d29f, 32'shf77a6129, 
               32'shf77befb5, 32'shf77d7e42, 32'shf77f0cd0, 32'shf7809b60, 32'shf78229f1, 32'shf783b883, 32'shf7854717, 32'shf786d5ab, 
               32'shf7886442, 32'shf789f2d9, 32'shf78b8172, 32'shf78d100c, 32'shf78e9ea7, 32'shf7902d44, 32'shf791bbe2, 32'shf7934a81, 
               32'shf794d922, 32'shf79667c4, 32'shf797f667, 32'shf799850b, 32'shf79b13b1, 32'shf79ca258, 32'shf79e3100, 32'shf79fbfaa, 
               32'shf7a14e55, 32'shf7a2dd01, 32'shf7a46baf, 32'shf7a5fa5d, 32'shf7a7890d, 32'shf7a917bf, 32'shf7aaa671, 32'shf7ac3525, 
               32'shf7adc3db, 32'shf7af5291, 32'shf7b0e149, 32'shf7b27002, 32'shf7b3febc, 32'shf7b58d78, 32'shf7b71c35, 32'shf7b8aaf3, 
               32'shf7ba39b3, 32'shf7bbc873, 32'shf7bd5735, 32'shf7bee5f9, 32'shf7c074bd, 32'shf7c20383, 32'shf7c3924a, 32'shf7c52112, 
               32'shf7c6afdc, 32'shf7c83ea7, 32'shf7c9cd73, 32'shf7cb5c41, 32'shf7cceb0f, 32'shf7ce79df, 32'shf7d008b1, 32'shf7d19783, 
               32'shf7d32657, 32'shf7d4b52c, 32'shf7d64402, 32'shf7d7d2da, 32'shf7d961b3, 32'shf7daf08d, 32'shf7dc7f68, 32'shf7de0e44, 
               32'shf7df9d22, 32'shf7e12c01, 32'shf7e2bae2, 32'shf7e449c3, 32'shf7e5d8a6, 32'shf7e7678a, 32'shf7e8f670, 32'shf7ea8556, 
               32'shf7ec143e, 32'shf7eda327, 32'shf7ef3211, 32'shf7f0c0fd, 32'shf7f24fea, 32'shf7f3ded8, 32'shf7f56dc7, 32'shf7f6fcb8, 
               32'shf7f88ba9, 32'shf7fa1a9c, 32'shf7fba991, 32'shf7fd3886, 32'shf7fec77d, 32'shf8005675, 32'shf801e56e, 32'shf8037468, 
               32'shf8050364, 32'shf8069261, 32'shf808215f, 32'shf809b05e, 32'shf80b3f5f, 32'shf80cce61, 32'shf80e5d64, 32'shf80fec68, 
               32'shf8117b6d, 32'shf8130a74, 32'shf814997c, 32'shf8162885, 32'shf817b78f, 32'shf819469b, 32'shf81ad5a8, 32'shf81c64b6, 
               32'shf81df3c5, 32'shf81f82d5, 32'shf82111e7, 32'shf822a0fa, 32'shf824300e, 32'shf825bf23, 32'shf8274e3a, 32'shf828dd51, 
               32'shf82a6c6a, 32'shf82bfb84, 32'shf82d8aa0, 32'shf82f19bc, 32'shf830a8da, 32'shf83237f9, 32'shf833c719, 32'shf835563b, 
               32'shf836e55d, 32'shf8387481, 32'shf83a03a6, 32'shf83b92cc, 32'shf83d21f3, 32'shf83eb11c, 32'shf8404046, 32'shf841cf71, 
               32'shf8435e9d, 32'shf844edca, 32'shf8467cf9, 32'shf8480c28, 32'shf8499b59, 32'shf84b2a8b, 32'shf84cb9bf, 32'shf84e48f3, 
               32'shf84fd829, 32'shf8516760, 32'shf852f698, 32'shf85485d1, 32'shf856150b, 32'shf857a447, 32'shf8593383, 32'shf85ac2c1, 
               32'shf85c5201, 32'shf85de141, 32'shf85f7082, 32'shf860ffc5, 32'shf8628f09, 32'shf8641e4e, 32'shf865ad94, 32'shf8673cdb, 
               32'shf868cc24, 32'shf86a5b6d, 32'shf86beab8, 32'shf86d7a04, 32'shf86f0952, 32'shf87098a0, 32'shf87227ef, 32'shf873b740, 
               32'shf8754692, 32'shf876d5e5, 32'shf8786539, 32'shf879f48e, 32'shf87b83e5, 32'shf87d133d, 32'shf87ea295, 32'shf88031ef, 
               32'shf881c14b, 32'shf88350a7, 32'shf884e004, 32'shf8866f63, 32'shf887fec3, 32'shf8898e23, 32'shf88b1d86, 32'shf88cace9, 
               32'shf88e3c4d, 32'shf88fcbb3, 32'shf8915b19, 32'shf892ea81, 32'shf89479ea, 32'shf8960954, 32'shf89798bf, 32'shf899282c, 
               32'shf89ab799, 32'shf89c4708, 32'shf89dd678, 32'shf89f65e8, 32'shf8a0f55b, 32'shf8a284ce, 32'shf8a41442, 32'shf8a5a3b8, 
               32'shf8a7332e, 32'shf8a8c2a6, 32'shf8aa521f, 32'shf8abe199, 32'shf8ad7114, 32'shf8af0090, 32'shf8b0900d, 32'shf8b21f8c, 
               32'shf8b3af0c, 32'shf8b53e8c, 32'shf8b6ce0e, 32'shf8b85d91, 32'shf8b9ed15, 32'shf8bb7c9b, 32'shf8bd0c21, 32'shf8be9ba9, 
               32'shf8c02b31, 32'shf8c1babb, 32'shf8c34a46, 32'shf8c4d9d2, 32'shf8c6695f, 32'shf8c7f8ed, 32'shf8c9887c, 32'shf8cb180d, 
               32'shf8cca79e, 32'shf8ce3731, 32'shf8cfc6c5, 32'shf8d1565a, 32'shf8d2e5f0, 32'shf8d47587, 32'shf8d6051f, 32'shf8d794b8, 
               32'shf8d92452, 32'shf8dab3ee, 32'shf8dc438b, 32'shf8ddd328, 32'shf8df62c7, 32'shf8e0f267, 32'shf8e28208, 32'shf8e411aa, 
               32'shf8e5a14d, 32'shf8e730f2, 32'shf8e8c097, 32'shf8ea503d, 32'shf8ebdfe5, 32'shf8ed6f8e, 32'shf8eeff37, 32'shf8f08ee2, 
               32'shf8f21e8e, 32'shf8f3ae3b, 32'shf8f53de9, 32'shf8f6cd98, 32'shf8f85d49, 32'shf8f9ecfa, 32'shf8fb7cac, 32'shf8fd0c60, 
               32'shf8fe9c15, 32'shf9002bca, 32'shf901bb81, 32'shf9034b39, 32'shf904daf2, 32'shf9066aac, 32'shf907fa67, 32'shf9098a23, 
               32'shf90b19e0, 32'shf90ca99e, 32'shf90e395e, 32'shf90fc91e, 32'shf91158e0, 32'shf912e8a2, 32'shf9147866, 32'shf916082b, 
               32'shf91797f0, 32'shf91927b7, 32'shf91ab77f, 32'shf91c4748, 32'shf91dd712, 32'shf91f66dd, 32'shf920f6a9, 32'shf9228677, 
               32'shf9241645, 32'shf925a614, 32'shf92735e5, 32'shf928c5b6, 32'shf92a5589, 32'shf92be55c, 32'shf92d7531, 32'shf92f0506, 
               32'shf93094dd, 32'shf93224b5, 32'shf933b48e, 32'shf9354468, 32'shf936d442, 32'shf938641e, 32'shf939f3fb, 32'shf93b83d9, 
               32'shf93d13b8, 32'shf93ea399, 32'shf940337a, 32'shf941c35c, 32'shf943533f, 32'shf944e323, 32'shf9467309, 32'shf94802ef, 
               32'shf94992d7, 32'shf94b22bf, 32'shf94cb2a8, 32'shf94e4293, 32'shf94fd27f, 32'shf951626b, 32'shf952f259, 32'shf9548247, 
               32'shf9561237, 32'shf957a228, 32'shf9593219, 32'shf95ac20c, 32'shf95c5200, 32'shf95de1f5, 32'shf95f71ea, 32'shf96101e1, 
               32'shf96291d9, 32'shf96421d2, 32'shf965b1cc, 32'shf96741c7, 32'shf968d1c3, 32'shf96a61c0, 32'shf96bf1be, 32'shf96d81bc, 
               32'shf96f11bc, 32'shf970a1bd, 32'shf97231bf, 32'shf973c1c2, 32'shf97551c6, 32'shf976e1cc, 32'shf97871d2, 32'shf97a01d9, 
               32'shf97b91e1, 32'shf97d21ea, 32'shf97eb1f4, 32'shf98041ff, 32'shf981d20b, 32'shf9836218, 32'shf984f226, 32'shf9868235, 
               32'shf9881245, 32'shf989a256, 32'shf98b3268, 32'shf98cc27b, 32'shf98e528f, 32'shf98fe2a5, 32'shf99172bb, 32'shf99302d2, 
               32'shf99492ea, 32'shf9962303, 32'shf997b31d, 32'shf9994338, 32'shf99ad354, 32'shf99c6371, 32'shf99df38e, 32'shf99f83ad, 
               32'shf9a113cd, 32'shf9a2a3ee, 32'shf9a43410, 32'shf9a5c433, 32'shf9a75457, 32'shf9a8e47c, 32'shf9aa74a1, 32'shf9ac04c8, 
               32'shf9ad94f0, 32'shf9af2519, 32'shf9b0b542, 32'shf9b2456d, 32'shf9b3d599, 32'shf9b565c5, 32'shf9b6f5f3, 32'shf9b88621, 
               32'shf9ba1651, 32'shf9bba681, 32'shf9bd36b3, 32'shf9bec6e5, 32'shf9c05719, 32'shf9c1e74d, 32'shf9c37782, 32'shf9c507b9, 
               32'shf9c697f0, 32'shf9c82828, 32'shf9c9b861, 32'shf9cb489b, 32'shf9ccd8d6, 32'shf9ce6912, 32'shf9cff94f, 32'shf9d1898d, 
               32'shf9d319cc, 32'shf9d4aa0c, 32'shf9d63a4d, 32'shf9d7ca8f, 32'shf9d95ad1, 32'shf9daeb15, 32'shf9dc7b5a, 32'shf9de0b9f, 
               32'shf9df9be6, 32'shf9e12c2d, 32'shf9e2bc75, 32'shf9e44cbf, 32'shf9e5dd09, 32'shf9e76d54, 32'shf9e8fda0, 32'shf9ea8ded, 
               32'shf9ec1e3b, 32'shf9edae8a, 32'shf9ef3eda, 32'shf9f0cf2b, 32'shf9f25f7d, 32'shf9f3efcf, 32'shf9f58023, 32'shf9f71078, 
               32'shf9f8a0cd, 32'shf9fa3123, 32'shf9fbc17b, 32'shf9fd51d3, 32'shf9fee22c, 32'shfa007286, 32'shfa0202e1, 32'shfa03933d, 
               32'shfa05239a, 32'shfa06b3f8, 32'shfa084457, 32'shfa09d4b7, 32'shfa0b6517, 32'shfa0cf579, 32'shfa0e85db, 32'shfa10163e, 
               32'shfa11a6a3, 32'shfa133708, 32'shfa14c76e, 32'shfa1657d5, 32'shfa17e83d, 32'shfa1978a6, 32'shfa1b090f, 32'shfa1c997a, 
               32'shfa1e29e5, 32'shfa1fba52, 32'shfa214abf, 32'shfa22db2d, 32'shfa246b9d, 32'shfa25fc0d, 32'shfa278c7e, 32'shfa291cf0, 
               32'shfa2aad62, 32'shfa2c3dd6, 32'shfa2dce4b, 32'shfa2f5ec0, 32'shfa30ef36, 32'shfa327fae, 32'shfa341026, 32'shfa35a09f, 
               32'shfa373119, 32'shfa38c194, 32'shfa3a520f, 32'shfa3be28c, 32'shfa3d7309, 32'shfa3f0388, 32'shfa409407, 32'shfa422487, 
               32'shfa43b508, 32'shfa45458a, 32'shfa46d60d, 32'shfa486691, 32'shfa49f715, 32'shfa4b879b, 32'shfa4d1821, 32'shfa4ea8a8, 
               32'shfa503930, 32'shfa51c9b9, 32'shfa535a43, 32'shfa54eace, 32'shfa567b5a, 32'shfa580be6, 32'shfa599c73, 32'shfa5b2d02, 
               32'shfa5cbd91, 32'shfa5e4e21, 32'shfa5fdeb1, 32'shfa616f43, 32'shfa62ffd6, 32'shfa649069, 32'shfa6620fd, 32'shfa67b193, 
               32'shfa694229, 32'shfa6ad2bf, 32'shfa6c6357, 32'shfa6df3f0, 32'shfa6f8489, 32'shfa711524, 32'shfa72a5bf, 32'shfa74365b, 
               32'shfa75c6f8, 32'shfa775795, 32'shfa78e834, 32'shfa7a78d3, 32'shfa7c0974, 32'shfa7d9a15, 32'shfa7f2ab7, 32'shfa80bb5a, 
               32'shfa824bfd, 32'shfa83dca2, 32'shfa856d47, 32'shfa86fded, 32'shfa888e95, 32'shfa8a1f3c, 32'shfa8bafe5, 32'shfa8d408f, 
               32'shfa8ed139, 32'shfa9061e5, 32'shfa91f291, 32'shfa93833e, 32'shfa9513eb, 32'shfa96a49a, 32'shfa98354a, 32'shfa99c5fa, 
               32'shfa9b56ab, 32'shfa9ce75d, 32'shfa9e7810, 32'shfaa008c3, 32'shfaa19978, 32'shfaa32a2d, 32'shfaa4bae3, 32'shfaa64b9a, 
               32'shfaa7dc52, 32'shfaa96d0a, 32'shfaaafdc4, 32'shfaac8e7e, 32'shfaae1f39, 32'shfaafaff5, 32'shfab140b2, 32'shfab2d16f, 
               32'shfab4622d, 32'shfab5f2ed, 32'shfab783ad, 32'shfab9146d, 32'shfabaa52f, 32'shfabc35f1, 32'shfabdc6b4, 32'shfabf5778, 
               32'shfac0e83d, 32'shfac27903, 32'shfac409c9, 32'shfac59a91, 32'shfac72b59, 32'shfac8bc22, 32'shfaca4ceb, 32'shfacbddb6, 
               32'shfacd6e81, 32'shfaceff4d, 32'shfad0901a, 32'shfad220e8, 32'shfad3b1b6, 32'shfad54285, 32'shfad6d355, 32'shfad86426, 
               32'shfad9f4f8, 32'shfadb85ca, 32'shfadd169e, 32'shfadea772, 32'shfae03847, 32'shfae1c91c, 32'shfae359f3, 32'shfae4eaca, 
               32'shfae67ba2, 32'shfae80c7a, 32'shfae99d54, 32'shfaeb2e2e, 32'shfaecbf0a, 32'shfaee4fe5, 32'shfaefe0c2, 32'shfaf171a0, 
               32'shfaf3027e, 32'shfaf4935d, 32'shfaf6243d, 32'shfaf7b51d, 32'shfaf945ff, 32'shfafad6e1, 32'shfafc67c4, 32'shfafdf8a7, 
               32'shfaff898c, 32'shfb011a71, 32'shfb02ab57, 32'shfb043c3e, 32'shfb05cd25, 32'shfb075e0e, 32'shfb08eef7, 32'shfb0a7fe1, 
               32'shfb0c10cb, 32'shfb0da1b6, 32'shfb0f32a3, 32'shfb10c38f, 32'shfb12547d, 32'shfb13e56c, 32'shfb15765b, 32'shfb17074b, 
               32'shfb18983b, 32'shfb1a292d, 32'shfb1bba1f, 32'shfb1d4b12, 32'shfb1edc06, 32'shfb206cfa, 32'shfb21fdef, 32'shfb238ee5, 
               32'shfb251fdc, 32'shfb26b0d3, 32'shfb2841cc, 32'shfb29d2c5, 32'shfb2b63be, 32'shfb2cf4b9, 32'shfb2e85b4, 32'shfb3016b0, 
               32'shfb31a7ac, 32'shfb3338aa, 32'shfb34c9a8, 32'shfb365aa7, 32'shfb37eba7, 32'shfb397ca7, 32'shfb3b0da8, 32'shfb3c9eaa, 
               32'shfb3e2fac, 32'shfb3fc0b0, 32'shfb4151b4, 32'shfb42e2b9, 32'shfb4473be, 32'shfb4604c4, 32'shfb4795cb, 32'shfb4926d3, 
               32'shfb4ab7db, 32'shfb4c48e4, 32'shfb4dd9ee, 32'shfb4f6af9, 32'shfb50fc04, 32'shfb528d10, 32'shfb541e1d, 32'shfb55af2a, 
               32'shfb574039, 32'shfb58d148, 32'shfb5a6257, 32'shfb5bf368, 32'shfb5d8479, 32'shfb5f158a, 32'shfb60a69d, 32'shfb6237b0, 
               32'shfb63c8c4, 32'shfb6559d9, 32'shfb66eaee, 32'shfb687c04, 32'shfb6a0d1b, 32'shfb6b9e32, 32'shfb6d2f4a, 32'shfb6ec063, 
               32'shfb70517d, 32'shfb71e297, 32'shfb7373b2, 32'shfb7504ce, 32'shfb7695ea, 32'shfb782707, 32'shfb79b825, 32'shfb7b4944, 
               32'shfb7cda63, 32'shfb7e6b83, 32'shfb7ffca3, 32'shfb818dc4, 32'shfb831ee6, 32'shfb84b009, 32'shfb86412c, 32'shfb87d250, 
               32'shfb896375, 32'shfb8af49b, 32'shfb8c85c1, 32'shfb8e16e7, 32'shfb8fa80f, 32'shfb913937, 32'shfb92ca60, 32'shfb945b89, 
               32'shfb95ecb4, 32'shfb977ddf, 32'shfb990f0a, 32'shfb9aa036, 32'shfb9c3163, 32'shfb9dc291, 32'shfb9f53bf, 32'shfba0e4ee, 
               32'shfba2761e, 32'shfba4074e, 32'shfba5987f, 32'shfba729b1, 32'shfba8bae3, 32'shfbaa4c16, 32'shfbabdd49, 32'shfbad6e7e, 
               32'shfbaeffb3, 32'shfbb090e8, 32'shfbb2221f, 32'shfbb3b356, 32'shfbb5448d, 32'shfbb6d5c6, 32'shfbb866ff, 32'shfbb9f838, 
               32'shfbbb8973, 32'shfbbd1aad, 32'shfbbeabe9, 32'shfbc03d25, 32'shfbc1ce62, 32'shfbc35fa0, 32'shfbc4f0de, 32'shfbc6821d, 
               32'shfbc8135c, 32'shfbc9a49d, 32'shfbcb35dd, 32'shfbccc71f, 32'shfbce5861, 32'shfbcfe9a4, 32'shfbd17ae7, 32'shfbd30c2b, 
               32'shfbd49d70, 32'shfbd62eb5, 32'shfbd7bffb, 32'shfbd95142, 32'shfbdae289, 32'shfbdc73d1, 32'shfbde0519, 32'shfbdf9663, 
               32'shfbe127ac, 32'shfbe2b8f7, 32'shfbe44a42, 32'shfbe5db8e, 32'shfbe76cda, 32'shfbe8fe27, 32'shfbea8f75, 32'shfbec20c3, 
               32'shfbedb212, 32'shfbef4361, 32'shfbf0d4b1, 32'shfbf26602, 32'shfbf3f753, 32'shfbf588a5, 32'shfbf719f8, 32'shfbf8ab4b, 
               32'shfbfa3c9f, 32'shfbfbcdf4, 32'shfbfd5f49, 32'shfbfef09f, 32'shfc0081f5, 32'shfc02134c, 32'shfc03a4a3, 32'shfc0535fc, 
               32'shfc06c754, 32'shfc0858ae, 32'shfc09ea08, 32'shfc0b7b62, 32'shfc0d0cbe, 32'shfc0e9e1a, 32'shfc102f76, 32'shfc11c0d3, 
               32'shfc135231, 32'shfc14e38f, 32'shfc1674ee, 32'shfc18064d, 32'shfc1997ae, 32'shfc1b290e, 32'shfc1cba6f, 32'shfc1e4bd1, 
               32'shfc1fdd34, 32'shfc216e97, 32'shfc22fffb, 32'shfc24915f, 32'shfc2622c4, 32'shfc27b429, 32'shfc29458f, 32'shfc2ad6f6, 
               32'shfc2c685d, 32'shfc2df9c5, 32'shfc2f8b2e, 32'shfc311c97, 32'shfc32ae00, 32'shfc343f6a, 32'shfc35d0d5, 32'shfc376240, 
               32'shfc38f3ac, 32'shfc3a8519, 32'shfc3c1686, 32'shfc3da7f4, 32'shfc3f3962, 32'shfc40cad1, 32'shfc425c40, 32'shfc43edb0, 
               32'shfc457f21, 32'shfc471092, 32'shfc48a204, 32'shfc4a3376, 32'shfc4bc4e9, 32'shfc4d565c, 32'shfc4ee7d0, 32'shfc507945, 
               32'shfc520aba, 32'shfc539c30, 32'shfc552da6, 32'shfc56bf1d, 32'shfc585094, 32'shfc59e20c, 32'shfc5b7385, 32'shfc5d04fe, 
               32'shfc5e9678, 32'shfc6027f2, 32'shfc61b96d, 32'shfc634ae8, 32'shfc64dc64, 32'shfc666de0, 32'shfc67ff5d, 32'shfc6990db, 
               32'shfc6b2259, 32'shfc6cb3d8, 32'shfc6e4557, 32'shfc6fd6d7, 32'shfc716857, 32'shfc72f9d8, 32'shfc748b59, 32'shfc761cdb, 
               32'shfc77ae5e, 32'shfc793fe1, 32'shfc7ad164, 32'shfc7c62e8, 32'shfc7df46d, 32'shfc7f85f2, 32'shfc811778, 32'shfc82a8fe, 
               32'shfc843a85, 32'shfc85cc0d, 32'shfc875d95, 32'shfc88ef1d, 32'shfc8a80a6, 32'shfc8c122f, 32'shfc8da3ba, 32'shfc8f3544, 
               32'shfc90c6cf, 32'shfc92585b, 32'shfc93e9e7, 32'shfc957b74, 32'shfc970d01, 32'shfc989e8f, 32'shfc9a301d, 32'shfc9bc1ac, 
               32'shfc9d533b, 32'shfc9ee4cb, 32'shfca0765b, 32'shfca207ec, 32'shfca3997e, 32'shfca52b0f, 32'shfca6bca2, 32'shfca84e35, 
               32'shfca9dfc8, 32'shfcab715c, 32'shfcad02f1, 32'shfcae9486, 32'shfcb0261b, 32'shfcb1b7b1, 32'shfcb34948, 32'shfcb4dadf, 
               32'shfcb66c77, 32'shfcb7fe0f, 32'shfcb98fa7, 32'shfcbb2140, 32'shfcbcb2da, 32'shfcbe4474, 32'shfcbfd60e, 32'shfcc167aa, 
               32'shfcc2f945, 32'shfcc48ae1, 32'shfcc61c7e, 32'shfcc7ae1b, 32'shfcc93fb9, 32'shfccad157, 32'shfccc62f5, 32'shfccdf494, 
               32'shfccf8634, 32'shfcd117d4, 32'shfcd2a974, 32'shfcd43b15, 32'shfcd5ccb7, 32'shfcd75e59, 32'shfcd8effb, 32'shfcda819e, 
               32'shfcdc1342, 32'shfcdda4e6, 32'shfcdf368a, 32'shfce0c82f, 32'shfce259d5, 32'shfce3eb7a, 32'shfce57d21, 32'shfce70ec8, 
               32'shfce8a06f, 32'shfcea3217, 32'shfcebc3bf, 32'shfced5568, 32'shfceee711, 32'shfcf078bb, 32'shfcf20a65, 32'shfcf39c0f, 
               32'shfcf52dbb, 32'shfcf6bf66, 32'shfcf85112, 32'shfcf9e2bf, 32'shfcfb746c, 32'shfcfd0619, 32'shfcfe97c7, 32'shfd002975, 
               32'shfd01bb24, 32'shfd034cd3, 32'shfd04de83, 32'shfd067033, 32'shfd0801e4, 32'shfd099395, 32'shfd0b2547, 32'shfd0cb6f9, 
               32'shfd0e48ab, 32'shfd0fda5e, 32'shfd116c12, 32'shfd12fdc6, 32'shfd148f7a, 32'shfd16212f, 32'shfd17b2e4, 32'shfd194499, 
               32'shfd1ad650, 32'shfd1c6806, 32'shfd1df9bd, 32'shfd1f8b74, 32'shfd211d2c, 32'shfd22aee5, 32'shfd24409d, 32'shfd25d257, 
               32'shfd276410, 32'shfd28f5ca, 32'shfd2a8785, 32'shfd2c1940, 32'shfd2daafb, 32'shfd2f3cb7, 32'shfd30ce73, 32'shfd326030, 
               32'shfd33f1ed, 32'shfd3583ab, 32'shfd371569, 32'shfd38a727, 32'shfd3a38e6, 32'shfd3bcaa5, 32'shfd3d5c65, 32'shfd3eee25, 
               32'shfd407fe6, 32'shfd4211a7, 32'shfd43a368, 32'shfd45352a, 32'shfd46c6ec, 32'shfd4858af, 32'shfd49ea72, 32'shfd4b7c35, 
               32'shfd4d0df9, 32'shfd4e9fbe, 32'shfd503182, 32'shfd51c348, 32'shfd53550d, 32'shfd54e6d3, 32'shfd56789a, 32'shfd580a60, 
               32'shfd599c28, 32'shfd5b2def, 32'shfd5cbfb7, 32'shfd5e5180, 32'shfd5fe348, 32'shfd617512, 32'shfd6306db, 32'shfd6498a5, 
               32'shfd662a70, 32'shfd67bc3b, 32'shfd694e06, 32'shfd6adfd2, 32'shfd6c719e, 32'shfd6e036a, 32'shfd6f9537, 32'shfd712704, 
               32'shfd72b8d2, 32'shfd744aa0, 32'shfd75dc6e, 32'shfd776e3d, 32'shfd79000d, 32'shfd7a91dc, 32'shfd7c23ac, 32'shfd7db57c, 
               32'shfd7f474d, 32'shfd80d91e, 32'shfd826af0, 32'shfd83fcc2, 32'shfd858e94, 32'shfd872067, 32'shfd88b23a, 32'shfd8a440d, 
               32'shfd8bd5e1, 32'shfd8d67b5, 32'shfd8ef98a, 32'shfd908b5f, 32'shfd921d34, 32'shfd93af0a, 32'shfd9540e0, 32'shfd96d2b7, 
               32'shfd98648d, 32'shfd99f665, 32'shfd9b883c, 32'shfd9d1a14, 32'shfd9eabec, 32'shfda03dc5, 32'shfda1cf9e, 32'shfda36178, 
               32'shfda4f351, 32'shfda6852b, 32'shfda81706, 32'shfda9a8e1, 32'shfdab3abc, 32'shfdaccc98, 32'shfdae5e74, 32'shfdaff050, 
               32'shfdb1822c, 32'shfdb31409, 32'shfdb4a5e7, 32'shfdb637c5, 32'shfdb7c9a3, 32'shfdb95b81, 32'shfdbaed60, 32'shfdbc7f3f, 
               32'shfdbe111e, 32'shfdbfa2fe, 32'shfdc134de, 32'shfdc2c6bf, 32'shfdc458a0, 32'shfdc5ea81, 32'shfdc77c62, 32'shfdc90e44, 
               32'shfdcaa027, 32'shfdcc3209, 32'shfdcdc3ec, 32'shfdcf55cf, 32'shfdd0e7b3, 32'shfdd27997, 32'shfdd40b7b, 32'shfdd59d60, 
               32'shfdd72f45, 32'shfdd8c12a, 32'shfdda530f, 32'shfddbe4f5, 32'shfddd76dc, 32'shfddf08c2, 32'shfde09aa9, 32'shfde22c90, 
               32'shfde3be78, 32'shfde55060, 32'shfde6e248, 32'shfde87431, 32'shfdea0619, 32'shfdeb9803, 32'shfded29ec, 32'shfdeebbd6, 
               32'shfdf04dc0, 32'shfdf1dfab, 32'shfdf37195, 32'shfdf50380, 32'shfdf6956c, 32'shfdf82758, 32'shfdf9b944, 32'shfdfb4b30, 
               32'shfdfcdd1d, 32'shfdfe6f0a, 32'shfe0000f7, 32'shfe0192e4, 32'shfe0324d2, 32'shfe04b6c0, 32'shfe0648af, 32'shfe07da9e, 
               32'shfe096c8d, 32'shfe0afe7c, 32'shfe0c906c, 32'shfe0e225c, 32'shfe0fb44c, 32'shfe11463d, 32'shfe12d82e, 32'shfe146a1f, 
               32'shfe15fc11, 32'shfe178e02, 32'shfe191ff5, 32'shfe1ab1e7, 32'shfe1c43da, 32'shfe1dd5cd, 32'shfe1f67c0, 32'shfe20f9b3, 
               32'shfe228ba7, 32'shfe241d9b, 32'shfe25af90, 32'shfe274184, 32'shfe28d379, 32'shfe2a656f, 32'shfe2bf764, 32'shfe2d895a, 
               32'shfe2f1b50, 32'shfe30ad47, 32'shfe323f3d, 32'shfe33d134, 32'shfe35632c, 32'shfe36f523, 32'shfe38871b, 32'shfe3a1913, 
               32'shfe3bab0b, 32'shfe3d3d04, 32'shfe3ecefd, 32'shfe4060f6, 32'shfe41f2ef, 32'shfe4384e9, 32'shfe4516e3, 32'shfe46a8dd, 
               32'shfe483ad8, 32'shfe49ccd2, 32'shfe4b5ecd, 32'shfe4cf0c9, 32'shfe4e82c4, 32'shfe5014c0, 32'shfe51a6bc, 32'shfe5338b8, 
               32'shfe54cab5, 32'shfe565cb2, 32'shfe57eeaf, 32'shfe5980ac, 32'shfe5b12aa, 32'shfe5ca4a8, 32'shfe5e36a6, 32'shfe5fc8a4, 
               32'shfe615aa3, 32'shfe62eca2, 32'shfe647ea1, 32'shfe6610a0, 32'shfe67a2a0, 32'shfe6934a0, 32'shfe6ac6a0, 32'shfe6c58a0, 
               32'shfe6deaa1, 32'shfe6f7ca1, 32'shfe710ea2, 32'shfe72a0a4, 32'shfe7432a5, 32'shfe75c4a7, 32'shfe7756a9, 32'shfe78e8ab, 
               32'shfe7a7aae, 32'shfe7c0cb1, 32'shfe7d9eb4, 32'shfe7f30b7, 32'shfe80c2ba, 32'shfe8254be, 32'shfe83e6c2, 32'shfe8578c6, 
               32'shfe870aca, 32'shfe889ccf, 32'shfe8a2ed4, 32'shfe8bc0d9, 32'shfe8d52de, 32'shfe8ee4e3, 32'shfe9076e9, 32'shfe9208ef, 
               32'shfe939af5, 32'shfe952cfb, 32'shfe96bf02, 32'shfe985109, 32'shfe99e310, 32'shfe9b7517, 32'shfe9d071e, 32'shfe9e9926, 
               32'shfea02b2e, 32'shfea1bd36, 32'shfea34f3e, 32'shfea4e147, 32'shfea6734f, 32'shfea80558, 32'shfea99761, 32'shfeab296b, 
               32'shfeacbb74, 32'shfeae4d7e, 32'shfeafdf88, 32'shfeb17192, 32'shfeb3039d, 32'shfeb495a7, 32'shfeb627b2, 32'shfeb7b9bd, 
               32'shfeb94bc8, 32'shfebaddd3, 32'shfebc6fdf, 32'shfebe01ea, 32'shfebf93f6, 32'shfec12603, 32'shfec2b80f, 32'shfec44a1b, 
               32'shfec5dc28, 32'shfec76e35, 32'shfec90042, 32'shfeca924f, 32'shfecc245d, 32'shfecdb66a, 32'shfecf4878, 32'shfed0da86, 
               32'shfed26c94, 32'shfed3fea3, 32'shfed590b1, 32'shfed722c0, 32'shfed8b4cf, 32'shfeda46de, 32'shfedbd8ed, 32'shfedd6afd, 
               32'shfedefd0c, 32'shfee08f1c, 32'shfee2212c, 32'shfee3b33c, 32'shfee5454c, 32'shfee6d75d, 32'shfee8696d, 32'shfee9fb7e, 
               32'shfeeb8d8f, 32'shfeed1fa0, 32'shfeeeb1b2, 32'shfef043c3, 32'shfef1d5d5, 32'shfef367e6, 32'shfef4f9f8, 32'shfef68c0b, 
               32'shfef81e1d, 32'shfef9b02f, 32'shfefb4242, 32'shfefcd455, 32'shfefe6668, 32'shfefff87b, 32'shff018a8e, 32'shff031ca1, 
               32'shff04aeb5, 32'shff0640c8, 32'shff07d2dc, 32'shff0964f0, 32'shff0af704, 32'shff0c8919, 32'shff0e1b2d, 32'shff0fad41, 
               32'shff113f56, 32'shff12d16b, 32'shff146380, 32'shff15f595, 32'shff1787aa, 32'shff1919c0, 32'shff1aabd5, 32'shff1c3deb, 
               32'shff1dd001, 32'shff1f6217, 32'shff20f42d, 32'shff228643, 32'shff24185a, 32'shff25aa70, 32'shff273c87, 32'shff28ce9e, 
               32'shff2a60b4, 32'shff2bf2cb, 32'shff2d84e3, 32'shff2f16fa, 32'shff30a911, 32'shff323b29, 32'shff33cd40, 32'shff355f58, 
               32'shff36f170, 32'shff388388, 32'shff3a15a0, 32'shff3ba7b9, 32'shff3d39d1, 32'shff3ecbe9, 32'shff405e02, 32'shff41f01b, 
               32'shff438234, 32'shff45144c, 32'shff46a666, 32'shff48387f, 32'shff49ca98, 32'shff4b5cb1, 32'shff4ceecb, 32'shff4e80e5, 
               32'shff5012fe, 32'shff51a518, 32'shff533732, 32'shff54c94c, 32'shff565b66, 32'shff57ed80, 32'shff597f9b, 32'shff5b11b5, 
               32'shff5ca3d0, 32'shff5e35ea, 32'shff5fc805, 32'shff615a20, 32'shff62ec3b, 32'shff647e56, 32'shff661071, 32'shff67a28c, 
               32'shff6934a8, 32'shff6ac6c3, 32'shff6c58de, 32'shff6deafa, 32'shff6f7d16, 32'shff710f31, 32'shff72a14d, 32'shff743369, 
               32'shff75c585, 32'shff7757a1, 32'shff78e9bd, 32'shff7a7bda, 32'shff7c0df6, 32'shff7da012, 32'shff7f322f, 32'shff80c44b, 
               32'shff825668, 32'shff83e885, 32'shff857aa2, 32'shff870cbe, 32'shff889edb, 32'shff8a30f8, 32'shff8bc316, 32'shff8d5533, 
               32'shff8ee750, 32'shff90796d, 32'shff920b8b, 32'shff939da8, 32'shff952fc5, 32'shff96c1e3, 32'shff985401, 32'shff99e61e, 
               32'shff9b783c, 32'shff9d0a5a, 32'shff9e9c78, 32'shffa02e96, 32'shffa1c0b4, 32'shffa352d2, 32'shffa4e4f0, 32'shffa6770e, 
               32'shffa8092c, 32'shffa99b4a, 32'shffab2d69, 32'shffacbf87, 32'shffae51a5, 32'shffafe3c4, 32'shffb175e2, 32'shffb30801, 
               32'shffb49a1f, 32'shffb62c3e, 32'shffb7be5d, 32'shffb9507c, 32'shffbae29a, 32'shffbc74b9, 32'shffbe06d8, 32'shffbf98f7, 
               32'shffc12b16, 32'shffc2bd35, 32'shffc44f54, 32'shffc5e173, 32'shffc77392, 32'shffc905b1, 32'shffca97d0, 32'shffcc29ef, 
               32'shffcdbc0f, 32'shffcf4e2e, 32'shffd0e04d, 32'shffd2726c, 32'shffd4048c, 32'shffd596ab, 32'shffd728ca, 32'shffd8baea, 
               32'shffda4d09, 32'shffdbdf29, 32'shffdd7148, 32'shffdf0368, 32'shffe09587, 32'shffe227a7, 32'shffe3b9c6, 32'shffe54be6, 
               32'shffe6de05, 32'shffe87025, 32'shffea0245, 32'shffeb9464, 32'shffed2684, 32'shffeeb8a3, 32'shfff04ac3, 32'shfff1dce3, 
               32'shfff36f02, 32'shfff50122, 32'shfff69342, 32'shfff82561, 32'shfff9b781, 32'shfffb49a1, 32'shfffcdbc1, 32'shfffe6de0
            };

            reg signed [31:0] W_Re_reg, W_Im_reg;
            always_ff @(posedge clk) begin
               W_Re_reg <= W_Re_table[k];
               W_Im_reg <= W_Im_table[k];
            end

            round32 #(.WIDTH(W_WIDTH)) round_re(W_Re_reg, W_Re);
            round32 #(.WIDTH(W_WIDTH)) round_im(W_Im_reg, W_Im);
         end
   endgenerate
endmodule :W_int32

`endif
