$dumpfile("dump.vcd");
$dumpvars;
