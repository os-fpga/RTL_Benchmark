----------------------------------------------------------------------------------
-- Company: Bluechip Technology
-- Engineer: Istvan Nagy, buenos@freemail.hu
-- 
-- Create Date:    15:58:13 05/30/2010
-- Design Name: 
-- Module Name:    op2p Port 
-- Project Name: 
-- Target Devices: Xilinx Spartan-6 LXT XC6SLX45T (for a 1.5GGbit/s 1x2 CAT-6-UTP), or other.
--   An optimal device for backplane applications could be the Xilinx Kintex XC7K355T-2FFG901 
--   (10.3Gbit/s 4x4, for 6U VPX), or a Kintex XC7K160T-2FFG676 (10.3Gbit/s 4x1, for 3U VPX).
-- Tool versions: ISE DS 12.1 M.53d
--
-- Dependencies: 
--  This design includes the aurora interface core which was generated by the Xilinx 
--  CoreGenerator. All the VHD files were copied here, including the ones from the 
--  "Reference Design" folder. This file is the top level source of the module, 
--  and is not generated by CoreGen. Search for all VHD files in all subfolders, then copy all.
--  2 files had to be modified (the ones from the example design folder): 
--     aurora_8b10b_v5_1_reset_logic.vhd
--     aurora_8b10b_v5_1_example_des_modified.vhd 
--  The last one has its filename and module name also modified, not only the internal logic.
--  If we use different Refclk/Linerate/widths/device-type, then we have to regenerate the
--  the Aurora core, and re-modify the files.
--  See the details at the bottom of this file in comment.
--
-- Revision 1.0 - Proof of concept
-- Additional Comments: 
--
-- Description: Open Peer to Peer Interface, Wishbone to Aurora Bridge (OP2P).
--   This is only one port. In a plug-in board or blade server we would need an FPGA
--   as the backplane bridge. The OP2P interface is optimized for mesh backplane
--   topologies. The backplane bridge needs a separate port for each backplane link.
--   There has to be a higher level scheduler logic or a soft processor to implement it.
--   To support bigger than purtnum^2 elements in a mesh, the bridge has to implement
--   packet forwarding. This way not every node will be directly conencted to every other.
--   It may be obvious that the forwarding involves 2 ports and some interaction from a DMA
--   or processor. The backplane bridge would normally consist of 4 OP2P ports, a host 
--   interface (PCIe), a local memory buffer interface (1 DRAM chip on-board, or BRAM on-chip)
--   and a local-host (soft proc or statemachine-type DMA logic)
--
-- Electrical Interface:
-- The data line rate is set to 1.5Gbps / diffpair, with 2 lanes in each direction, so
-- this gives a total of 6Gbps bandwidth. The reference clock is expected to be 75MHz LVDS
-- differential, but if we want to regenerate the core for a different linerate then we 
-- need to change the ref lock frequency. The reference clock must come from an on-board 
-- external clock generator, the Spartan6's internal clock networks dont meet the GTP's 
-- jitter specs. The external clock chip frequency can be controlled through the PR0,PR1,
-- OD0, OD1, OD2 pins.
--
-- Limitations:
-- This code is a proof of concept only. The data bandwidth is limited, since the on-chip
-- data buses/processing is 32-bit. The Spartan-6 (-2 speed grade) device is able to run
-- the interface with an around 100MHz on-chip parallel bus, but since the valid PLL settings
-- don't allow for parallel bus speed in this range, the on-chip logic runs on 75MHz with
-- serial line rate of 1.5Gbps. On a newer 7-series FPGA (Kintex, Virtex), it would run faster.
-- To utilize the 10.3Gbps speed on a 4x4 lane 6U-VPX backplane application, we would need
-- around 1.03GT/sec on-chip parallel buses with long burst support. At the moment the core
-- has 32-bit buses (FIFOs, Wishbone-bus to DRAM) and no burst support on the Wishbone side.
-- If we change the design to have 128bit on-chip parallel buses, then it would need a 250MHz
-- parallel-bus-clock speed, which might work on a Virtex-7 or Kintex-7 device. This would
-- mean a 4GBytes/s/port/direction data bandwidth (32GB/s/card total) on each backplane port 
-- (6U VPX at 10.3Gbps). On ISE-12.1 for Series-6 FPGAs, 128bit bus is only available for min x4.
-- A 3U VPX system at 10.3Gbps line-rate would have 1GBytes/sec/dir data bandwidth on each port,
-- which could still be achieved with a 32-bit on-chip bus at 250MHz. At 10.3Gbps (6U VPX), x4 
-- link width (instead of x1) would not provide additional bandwidth when using 32-bit parallel 
-- bus at 250MHz. 250MHz is around at the device limit with this core for Xilinx series-6/7.
-- A 64-bit 66MHz Compact-PCI interface only has a 0.528GBytes/sec aggregate bandwidth used 
-- by all cards and directions together.
-- The serial and the Wishbone transactions overlap to save time (latency), but transferring the
-- same amount of data on the Wishbone bus takes 3-10-times more time than it is on the serial
-- side. Currently at every 3-10 clock cycles there is a new Wishbone transaction when processing
-- a single OP2P packet. A long burst support would mean one WB transfer at every clock cycle.
--
-- Protocol: 
-- The lower layers are based on the Xilinx Aurora protocol, and generated by the Xilinx 
-- Coregenerator tool and instantiated in this file. The higher layers are implemented in 
-- this file.
-- All transactions are peer to peer, non-transparent, and implementing buffer-copy from 
-- devive/address to device/address.
-- Transmit can be initiated by localhost (it writes into local memory, then sets a registerbit 
-- accessed through the op2p_config_wb bus) or by arrived read request packet from remote device.
-- What happens during transmit: The IP reads the data from the local buffer, and sends it to the 
-- specified destination (target), then generates an interrupt. Receive: when receiving a packet, 
-- the aurora IP writes it into the memory (address is specified in the packet), then generates
-- an interrupt to the local host. So, all transfers happen directly between the memory and the 
-- aurora link, the host can not write the data into the aurora IP.
--
-- Packet format: Header + payload data. Max 2kBytes in one packet. If the request is targeting
--  a larger than 2kBytes memory area, then the scheduler has to divide the data into 2kB packets.
--  Header: 
--    1st DW: source ID (16bit 31:16), destination ID (16bit 15:0)
--    2nd DW: destination address (32bit)
--    3rd DW: source address (32bit)
--    4th DW: byte count(16bit: 1-64k 31:16), packet-type (4bit 15:12), status (4bit 11:8), 
--            first byte enable (4bit 7:4), RFU (4bit 3:0)
--       Packet type: 0000=wr_req, 0001=rd_request, 0010=rd_completion, 1010=retransmit_req, 
--							 others: RFU
--       Status: 0000=succesful_transaction, 0001=no_further_hop, 0010=unknown_error
--
-- Addressing: device identification is based on ID. Every packet copies a specified amount
--  of data from source_address in source device to destination_address in destination device (wr) or 
--  requests a read in the opposite way. The Aurora bridge normally has its own 4G or less address
--  space, which is a DRAM chip connected to the bridge (FPGA), typically 64MBytes. Every board 
--  has its own 0...MAX address space, which is indepenent from the other board's address spaces.
--  The local host is a processor, which can be the board's main x86/PPC/MIPS processor or a dedicated 
--  small processor inside or attached-to the aurora bridge (FPGA).
--  The completion swaps the source/destination ID/address fields!
-- ID: 10-bit chassys address and 6-bit slot address. The slot address can be figured out from 
--  the backplane's geographical addressing pins. The chassys address have to be specified by the 
--  user in a software or stored on the backplane in an EEPROM. The ID is programmed into the 
--  aurora interface registers after powerup by the local host. There is no plug and play device
--  discovery by hardware, although software can initiate discovery by pinging all possible device 
--  numbers in the chassys or in the server room. 
--  ID=0 means that the destination of the transaction is the device immediately found at the other end 
--  of the physical link, which also means that chassys addresses start from 1 till 1023, slot 
--  addresses from 0 till 63. ID0 can be used for discovery in backplanes, or for communication
--  in pint-to-point logical/physical connections in dedicated cable-links (system with 2 devices only).
-- Discovery: in the backplane, the port/link connectionsa re known based on the geographical 
--  addressing and the fixed topology. Only slot-0 has access to other chassys. At powerup, every 
--  slot pings the other slots to see if they are there, by a dummy 1-byte read.
-- Multi-hop transactions (FORWARDING) in multi-mesh topologies: if a device receives a packet which does 
--  not match its ID, then it has to store the packet in local DRAM, and the localhost has to retransmit in 
--  the appropriate port (another aurora block), based on the discovery or map. Packets to other chassys 
--  have to go through slot-0. When a port forwards a packet, the host writes the original source ID into
--  the source ID fifo, not the local ID. Sending forwarding (posted-write or read-request) request packets
--  is done like sending normal request through the same command FIFOs, with source-ID/=local_id written
--  into the FIFO. Receiving a forwarding (not matching ID) packet: store the whole packet in DRAM at an
--  automatically allocated location. The host can see in the siso_status_reg if there is anything, and read
--  the latest packet's address from the op2p_forwreq_pointer_reg FIFO. Later when the local host processor 
--  initiates a re-transmit, it should tell the port logic to free-up the memory buffer portion used by the 
--  packet. This is done by using the op2p_forw_freeupaddr_reg command FIFO. The buffer in use starts at a 
--  pre-programmed point set by op2p_forwarding_bufferbase_reg. The buffer can have max 512 entries, each 
--  2kByte (to accomodate a 1kBytes data + 4*32bit header), 1MByte total.
--  If a device is the actual destination for a forwarding packet, then it will see it as a notmal packet,
--  since the destination ID will match its local_id, and it will act as it would to a normal request packet.
--  
--
-- Software requirements:
--  Each board's local host processor has to have a complete map of the system. This can come from a discovery
--  protocol (not detailed here) or from a user manual entry (non plug and play, requires an administrator to
--  maintain the system, instead of "end users" like in case of commercial products). This map tells which port 
--  we find the node that we want to talk to, and which port we send the forwarding packets to. The local host
--  interaction to the system can be done two ways: a) simple system where one processor handles all transactions
--  at a register-level, b) a local DMA controller or soft processor inside the FPGA handles all packets at the 
--  register level but the local host processor only handles the user data and port mapping. In a possible
--  discovery protocol we do iterations, where node requests information from their neighbours in every iteration.
--  The data requested/provided contains data gathered in the previous iterations. In the first iteration we detect
--  only the direct neighbours (link partners) and their slot/chassys addresses. The number of iterations needed
--  equal to the number of hops needed plus one. In a room of four 8-slot chassys we need 4 iterations. Handling
--  this should be done by a software layer.
--
--  Registers (op2p_config_wb bus):
--   WRITE REQ (local host writes): source address (local), destination address, source ID, destination ID, 
--    byte-count.
--   WRITE_COMPLETION (this IP writes it): source address (remote), destination address (local), source ID, destination ID 
--    (check for match or forwarding), byte-count.
--   READ REQ (local host writes): source address (local), destination address, source ID (set up once), destination ID, 
--    byte-count.
--   READ completion status: completed_localaddress
--   Forwarding REQUEST received: buffer start address pointer and buffer size (local host writes it, not a FIFO), Packet 
--     pointer (FIFO, the aurora IP writes it). The complete packet with header is stored in memory. the packet size is in the header
--     Forwarding buffer freeup: free up buffer area already forwarded. address and size.
--   Control registers: FIFO status for every FIFO.
--   All of these registers are FIFOs, one transaction involves reading or writing 5 FIFOs (a COMMAND). Source ID is local ID 
--    for most of the transactions, except for the forwarded packets. 
--   Initiate outgoing transactions: Write all resuired registers in a set (wr, rdreq). Where more than one FIFO has to be 
--    written, the last written one will initiate the OP2P transaction. (all regs in a set must be written once).
--   If a read request arrives, the core will send the completion back with data, and will mark the source ID from the localid_reg,
--    that has to be written after system initialization once.
--   Link health: The host software should read the op2p_link_status_reg before initiating any op2p transactions, because if the 
--    link is not alive and trying to send packets then (due to broken connection or unpowered link partner) the system might hang.
--    The logic will not initiate any transactions if the link is not alive, this can cause command buffer overflow.
--
--	  Register Addresses (BYTE ADDRESSES):
--	  -------------------
--		--00h - op2p_fifostatus_reg		
--			Tells the status flags of the command FIFOs	
--		--04h - op2p_wr_sourceaddress_reg			(write command)
--		--08h - op2p_wr_destinationaddress_reg		(write command)
--		--0Ch - op2p_wr_sourceid_reg					(write command) 
--		--10h - op2p_wr_destinationid_reg			(write command)
--		--14h - op2p_wr_bytecount_reg					(write command)
--		--18h - op2p_rdreq_localaddress_reg			 (read request command)
--		--1Ch - op2p_rdreq_destinationaddress_reg	 (read request command)
--		--20h - op2p_rdreq_sourceid_reg				 (read request command)
--		--24h - op2p_rdreq_destinationid_reg		 (read request command)
--		--28h - op2p_rdreq_bytecount_reg				 (read request command)
--		--2Ch - op2p_rdcompl_localaddress_reg
--			If a read is completed, this FIFO will show the address where the data has been stored.
--			This can be used to poll the status of the read operation.
--		--30h - op2p_forwarding_bufferbase_reg		(forwarding buffer setup)
--			At startup write here the base address of the 1MBytes forwarding buffer in the DRAM buffer
--		--38h - op2p_forw_freeupaddr_reg			(forw buf runtime management)
--			After retransmitting a forwarding packet, the local host proc/DMA should write the
--			value from the op2p_forwreq_pointer_reg back into this FIFO to free-up the bufefr entry.
--		--40h - op2p_forwreq_pointer_reg			(forw buf runtime management)
--			If a packed arrived without ID-match, then it got stored in the local DRAM buffer
--			for retransmitting. The starting addresses are stored in this FIFO for the cpu to read.
--		--44h - op2p_arrivedwrite_address_reg
--			If a write has arrived, this FIFO will show the address where the data has been stored.
--			This can be used to to see if anyoone wrote data to us.
--		--48h - op2p_localid_reg
--			The local ID of this device. written by local host. Receiving completion 
--			or addressed (dest ID/=0) packet without setting this is not poosible. Set after startup.
--		--4Ch - op2p_link_status_reg
--			Tells if the link is alive, and also which lanes
--		--50h - op2p_port_reset_reg
--			We can initiate a soft reset to this OP2P port by register write
--		--54h - link_error_count_reg
--			This counts errors found in incoming packets. Counts forever from reset
--			8b10b encoding-based "non-existing-code" and disparity errors get detected.
--
--   Register bits:
--     op2p_link_status_reg: 
--        bit-0=CHANNEL_UP, 
--        bit-n:1=LANE_UP(0:n), 
--			 other bits are zero
--        bit-29: fc_haltlinkpartner   
--        bit-30: fc_halted_bylinkpartner   
--        bit-31: HARD_ERROR (needs port-reset)
--     op2p_fifostatus_reg
--			(0) <=  op2p_forwreq_pointer_regempty;       --empty
--			(1) <=  op2p_rdcompl_localaddress_regempty;
--			(2) <=  op2p_arrivedwrite_address_regempty; 
--			(3) <=  op2p_wr_sourceaddress_regfull;       --full
--			(4) <=  op2p_wr_destinationaddress_regfull;
--			(5) <=  op2p_wr_sourceid_regfull;
--			(6) <=  op2p_wr_destinationid_regfull;
--			(7) <=  op2p_wr_bytecount_regfull;
--			(8) <=  op2p_rdreq_localaddress_regfull;
--			(9) <=  op2p_rdreq_destinationaddress_regfull;
--			(10) <=  op2p_rdreq_sourceid_regfull;
--			(11) <=  op2p_rdreq_destinationid_regfull;
--			(12) <=  op2p_rdreq_bytecount_regfull;
--			(13) <=  op2p_forw_freeupaddr_regfull;
--			(14) <=  RFU
--			(31 downto 15) <=  (OTHERS => '0');
--		op2p_port_reset_reg
--			bit-0: set 1 to hold reset, set 0 to release from reset. After startup the port is not in reset.
--		Address registers:
--			all 32 bits are used. 4GB address space in the local DRAM buffer. (not x86 host memory space address)
--		ID registers: 
--			bit [15:0] are used for the 16-bit IDs.
--		Byte count registers
--			The number of bytes to be transferred. This must be 32bit aligned, 2 LSBs will be ignored.
--
--  Interrupts to local host:
--   - read completion (fifo was written)
--   - forwarding request
--   - write arrived
--   if any of the readable FIFOs is not empty, the interrupt stays asserted.
--
--  Trigger for (DRAM) WB transfer:
--   From Local-Host (op2p_config_wb bus, command registers filled) or request or response packet from
--   remote device.
--
--  Clocking architecture:
--   Every chip has its own reference clock, to refclk is wired between boards, only the data is 
--   connected. 
--   Clock Compensation: The Aurora 8B/10B protocol specifies a clock compensation mechanism 
--   that allows up to +/- 100 ppm difference between reference clocks on each side of the link.
--   This is a part of the Coregen-Aurora IP and it automatically inserts CC messages into 
--   the communication channel, using up around 1-2% of the data bandwidth.
--   Refclk: From external pin, on-board (on the PCB) 75MHz low jitter clock generator/pll/oscillator.
--   For the prototype board, a Texas Instruments CDCM61001 was used.
--   The reference clock source must be at least +/-50ppm accurate.
--   The DRAM/buffer interface is in the same clock domain as the rest of the OP2P/Aurora logic,
--   while the host interface is separate and isolated by command FIFOs.
--
-- Device Type Migration:
--  This core should work on any Xilinx Series-5/6/7 FPGAs, but at now it runs on XC6SLX45T.
--  For a new device (not an XC6SLX45T) we have to regenerate the Coregenerator cores,
--  replace all BUFIO2/MGT/BUFG/BRAM (and other) to the chosen device's appropriate resources,
--  in both the VHDL and the UCF sources. Also in the UCF the BUFIO2 and MGT placements 
--  will have to be re-specified with the appropriate resources/locations. The coregenerator
--  will have to be set up to generate cores with the same parameters and ports as they are
--  used here (to be useable as a drop-in replacement). Some resources are instantiated as
--  part of the Coregen cores, so they will be chosen by Coregen appropriately, we just need
--  to adjust their LOC placement constraints in the UCF file.
--
-- Coregenerator parameters:
--  Aurora8b10b: Name=aurora_8b10b_v5_1, Lanes=2, LaneWidth=2 (bytes on parallel bus from one lane), 
--               LineRate=1.5, GT_REFCLK=75MHz. These first few parameters have to be set accordingly, 
--               to achieve a 32bit databus (lanes x LaneW =4), valid PLL settings (from datasheet: 
--               a valid SerialRate-parallelclock-REFCLK combination), STA result on the parallel bus  
--               clock (check max possible CLK speed in STA report).
--               DataFlowMode=Duplex, Interface=Framing, FlowControl=CompletionNFC, GTP-LOC:X1Y0-GT0=1/GT1=2,
--               Clock source=GTPD1. The LOC has to work with the board schematics and other cores (PCIe).
--               See the instructions about source modifications at the bottom of this file (in comment).
--  Blockram: Name=blk_mem_gen_v4_1, Type=SimpleDpRAM, WriteEn=off, Algor=MinArea, 
--            WriteWidth=32, WriteDepth=512, Ena=AlwaysEnabled, ReadWidth=32, RegisterPorttB=off
--            LoadInitFile=off, Fill=off, UseRSTB=off.
--  FIFOs:  Name=fifo_generator_v6_1, R/W-ClockDomains=IndependentClocks/DistrRAM, ReadMode=StandardFIFO,
--          WriteWidth=32, WriteDepth=16, AlmostFull/Empty=off, WriteACK=off, WrOverflow=on, RdValid=off, 
--          RdEnderflow=on, ResetPin=on, EnableResSync=on, FullFlagResVal=0, UseDoutReset=on, DoutResVal=0,
--          ProgrammableFlags(full/emp)=No, DataCount=AllOff, 
--
---------------------------------------------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity op2p is
    Port ( --FPGA PINS (EXTERNAL):
           GTPD1_P  : in std_logic; --aurora GTP refclk P
           GTPD1_N  : in std_logic; --aurora GTP refclk N
           op2p_RXP  : in std_logic_vector(0 to 1);
           op2p_RXN  : in std_logic_vector(0 to 1);
           op2p_TXP  : out std_logic_vector(0 to 1);
           op2p_TXN  : out std_logic_vector(0 to 1);
			  --INTERNAL PORTS:
			  --DATA BUS (wishbone, to local DRAM): this IP is master on this
			  op2p_memory_wb_data_o : out std_logic_vector(31 downto 0); 
			  op2p_memory_wb_data_i : in std_logic_vector(31 downto 0);
			  op2p_memory_wb_addr_o : out std_logic_vector(25 downto 0);
			  op2p_memory_wb_cyc_o : out std_logic;
			  op2p_memory_wb_stb_o : out std_logic;
			  op2p_memory_wb_wr_o : out std_logic;
			  op2p_memory_wb_ack_i : in std_logic;
			  op2p_memory_wb_clk_o : out std_logic; 
			  op2p_memory_wb_sel_o : out std_logic_vector(3 downto 0);
			  --instruction registers wb-bus : this IP is slave on this
			  op2p_config_wb_data_o : in std_logic_vector(31 downto 0); 
			  op2p_config_wb_data_i : out std_logic_vector(31 downto 0);
			  op2p_config_wb_addr_i : in std_logic_vector(6 downto 0);
			  op2p_config_wb_cyc_i : in std_logic;
			  op2p_config_wb_stb_i : in std_logic;
			  op2p_config_wb_wr_i : in std_logic;
			  op2p_config_wb_ack_o : out std_logic;
			  op2p_config_wb_clk_i : in std_logic; 	
			  op2p_config_wb_sel_o :  in std_logic_vector(3 downto 0);
			  --system signals			  
			  op2p_reset : in std_logic;
			  x25m_clk : in std_logic;
			  CHANNEL_UP_copy : out std_logic;
			  --reference clock setting:
			  op2p_refclkset_od0 : out std_logic;
			  op2p_refclkset_od1 : out std_logic;
			  op2p_refclkset_od2 : out std_logic;
			  op2p_refclkset_pr0 : out std_logic;
			  op2p_refclkset_pr1 : out std_logic;
			  --interrupt out:	
			  op2p_irq : out  STD_LOGIC
			 );
end op2p;

-- ----- ARCHITECTURE START -------------------------------------------------------------------
architecture Behavioral of op2p is

-----------------------------------------------------------------------------------------------
   -- Internal Signals ------------------------------------------------------------------------
	--SIGNAL dummy : std_logic_vector(15 downto 0);	
  SIGNAL  RESET     : std_logic;
  SIGNAL  HARD_ERROR        : std_logic;
  SIGNAL  SOFT_ERROR        : std_logic;
  SIGNAL  FRAME_ERROR       : std_logic;
  SIGNAL  ERR_COUNT         : std_logic_vector(0 to 7);
  SIGNAL  LANE_UP           : std_logic_vector(0 to 1);
  SIGNAL  CHANNEL_UP        : std_logic;
  SIGNAL  INIT_CLK          :  std_logic;
  SIGNAL  GT_RESET_IN       :  std_logic;
  SIGNAL  TX_D    :  std_logic_vector(0 to 31); 
  SIGNAL  TX_REM          :  std_logic_vector(0 to 1);     
  SIGNAL  TX_SOF_N        :  std_logic;
  SIGNAL  TX_EOF_N        :  std_logic;
  SIGNAL  TX_SRC_RDY_N    :  std_logic;
  SIGNAL  TX_DST_RDY_N    :   std_logic;  
  SIGNAL  NFC_REQ_N       :  std_logic;
  SIGNAL  NFC_NB          :  std_logic_vector(0 to 3);     
  SIGNAL  NFC_ACK_N       :   std_logic;  
  SIGNAL  RX_D    :  std_logic_vector(0 to 31); 
  SIGNAL  RX_REM          :  std_logic_vector(0 to 1);     
  SIGNAL  RX_SOF_N        :  std_logic;
  SIGNAL  RX_EOF_N        :  std_logic;
  SIGNAL  RX_SRC_RDY_N    :  std_logic; 
  SIGNAL  RX_SNF          :  std_logic;
  SIGNAL  RX_FC_NB        :  std_logic_vector(0 to 3);  

  --received packet properties -not fifo
  SIGNAL op2p_wr_sourceaddress  : std_logic_vector(31 downto 0);
  SIGNAL op2p_wr_destinationaddress_reg : std_logic_vector(31 downto 0);
  SIGNAL op2p_wr_sourceid_reg  : std_logic_vector(31 downto 0);
  SIGNAL op2p_wr_destinationid_reg  : std_logic_vector(31 downto 0);
  --SIGNAL op2p_wr_destinationid_reg : std_logic_vector(31 downto 0);
  SIGNAL op2p_wr_bytecount_reg  : std_logic_vector(31 downto 0);
  SIGNAL op2p_wr_sourceaddressrd_en : std_logic;
  SIGNAL op2p_wr_sourceaddressdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_wr_sourceaddressempty : std_logic;
  
  --FIFO signals to the wb-slave interface:
  SIGNAL op2p_wr_sourceaddress_regrd_en : std_logic;
  SIGNAL op2p_wr_destinationaddress_regrd_en : std_logic;
  SIGNAL op2p_wr_sourceid_regrd_en : std_logic;
  SIGNAL op2p_wr_destinationid_regrd_en : std_logic;
  SIGNAL op2p_wr_bytecount_regrd_en : std_logic;
  SIGNAL op2p_rdreq_localaddress_regrd_en : std_logic;
  SIGNAL op2p_rdreq_destinationaddress_regrd_en : std_logic;
  SIGNAL op2p_rdreq_sourceid_regrd_en : std_logic;
  SIGNAL op2p_rdreq_destinationid_regrd_en : std_logic;
  SIGNAL op2p_rdreq_bytecount_regrd_en : std_logic;
  SIGNAL op2p_forw_freeupaddr_regrd_en : std_logic;
  SIGNAL op2p_forw_freeupsize_regrd_en : std_logic;
  SIGNAL op2p_forwreq_pointer_regdin : std_logic_vector(31 downto 0);
  SIGNAL op2p_forwreq_pointer_regwr_en : std_logic;
  SIGNAL op2p_rdcompl_localaddress_regdin : std_logic_vector(31 downto 0);
  SIGNAL op2p_rdcompl_localaddress_regwr_en : std_logic;
  SIGNAL op2p_arrivedwrite_address_regdin : std_logic_vector(31 downto 0);
  SIGNAL op2p_arrivedwrite_address_regwr_en : std_logic;          
  --SIGNAL op2p_config_wb_data_i : std_logic_vector(31 downto 0);
  --SIGNAL op2p_config_wb_ack_o : std_logic;
  SIGNAL op2p_irq_not_used : std_logic;
  SIGNAL op2p_wr_sourceaddress_regdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_wr_sourceaddress_regempty : std_logic;
  SIGNAL op2p_wr_destinationaddress_regdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_wr_destinationaddress_regempty : std_logic;
  SIGNAL op2p_wr_sourceid_regdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_wr_sourceid_regempty : std_logic;
  SIGNAL op2p_wr_destinationid_regdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_wr_destinationid_regempty : std_logic;
  SIGNAL op2p_wr_bytecount_regdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_wr_bytecount_regempty : std_logic;
  SIGNAL op2p_rdreq_localaddress_regdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_rdreq_localaddress_regempty : std_logic;
  SIGNAL op2p_rdreq_destinationaddress_regdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_rdreq_destinationaddress_regempty : std_logic;
  SIGNAL op2p_rdreq_sourceid_regdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_rdreq_sourceid_regempty : std_logic;
  SIGNAL op2p_rdreq_destinationid_regdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_rdreq_destinationid_regempty : std_logic;
  SIGNAL op2p_rdreq_bytecount_regdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_rdreq_bytecount_regempty : std_logic;
  SIGNAL op2p_forw_freeupaddr_regdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_forw_freeupaddr_regempty : std_logic;
  SIGNAL op2p_forw_freeupsize_regdout : std_logic_vector(31 downto 0);
  SIGNAL op2p_forw_freeupsize_regempty : std_logic;
  SIGNAL op2p_forwarding_bufferbase_reg : std_logic_vector(31 downto 0);
  SIGNAL op2p_forwarding_bufsize_reg : std_logic_vector(31 downto 0);
  SIGNAL op2p_forwreq_pointer_regfull : std_logic;
  SIGNAL op2p_rdcompl_localaddress_regfull : std_logic;
  SIGNAL op2p_arrivedwrite_address_regfull : std_logic;
  SIGNAL op2p_local_id : std_logic_vector(15 downto 0);

  SIGNAL bram_rxpacket_we  : std_logic_vector(0 downto 0);
  SIGNAL bram_rxpacket_writeaddress : std_logic_vector(8 downto 0);
  SIGNAL bram_rxpacket_writedata : std_logic_vector(31 downto 0);
  SIGNAL bram_rxpacket_readaddress : std_logic_vector(8 downto 0);
  SIGNAL bram_rxpacket_readdata : std_logic_vector(31 downto 0);
  SIGNAL bram_txpacket_we : std_logic_vector(0 downto 0);
  SIGNAL bram_txpacket_writeaddress : std_logic_vector(8 downto 0);
  SIGNAL bram_txpacket_writedata : std_logic_vector(31 downto 0);
  SIGNAL bram_txpacket_readaddress : std_logic_vector(8 downto 0);
  SIGNAL bram_txpacket_readdata : std_logic_vector(31 downto 0);
  
  SIGNAL packetstm_counter : std_logic_vector(7 downto 0);
  SIGNAL fbm_nextraddress_req : std_logic;
  SIGNAL fbm_nextraddress : std_logic_vector(31 downto 0);
  
  SIGNAL destination_address : std_logic_vector(31 downto 0);
  SIGNAL source_id : std_logic_vector(15 downto 0);
  SIGNAL destination_id : std_logic_vector(15 downto 0);
  SIGNAL source_address : std_logic_vector(31 downto 0);
  SIGNAL byte_count  : std_logic_vector(31 downto 0);

	--
  SIGNAL forw_packetaddr_allocated : std_logic;
  --SIGNAL fbm_nextraddress : std_logic_vector(31 downto 0);
  --SIGNAL fbm_nextraddress_req : std_logic_vector(31 downto 0);

  SIGNAL forwbuf_descriptor_ddword0 : std_logic_vector(63 downto 0);
  SIGNAL forwbuf_descriptor_ddword1 : std_logic_vector(63 downto 0);
  SIGNAL forwbuf_descriptor_ddword2 : std_logic_vector(63 downto 0);
  SIGNAL forwbuf_descriptor_ddword3 : std_logic_vector(63 downto 0);
  SIGNAL forwbuf_descriptor_ddword4 : std_logic_vector(63 downto 0);
  SIGNAL forwbuf_descriptor_ddword5 : std_logic_vector(63 downto 0);
  SIGNAL forwbuf_descriptor_ddword6 : std_logic_vector(63 downto 0);
  SIGNAL forwbuf_descriptor_ddword7 : std_logic_vector(63 downto 0);

  SIGNAL forwbuf_descriptor_byte0 : std_logic_vector(7 downto 0);
  SIGNAL forwbuf_descriptor_byte1 : std_logic_vector(7 downto 0);
  SIGNAL forwbuf_descriptor_byte2 : std_logic_vector(7 downto 0);
  SIGNAL forwbuf_descriptor_byte3 : std_logic_vector(7 downto 0);
  SIGNAL forwbuf_descriptor_byte4 : std_logic_vector(7 downto 0);
  SIGNAL forwbuf_descriptor_byte5 : std_logic_vector(7 downto 0);
  SIGNAL forwbuf_descriptor_byte6 : std_logic_vector(7 downto 0);
  SIGNAL forwbuf_descriptor_byte7 : std_logic_vector(7 downto 0);

  SIGNAL forwbuf_descriptor_bit0 : std_logic;
  SIGNAL forwbuf_descriptor_bit1  : std_logic;
  SIGNAL forwbuf_descriptor_bit2  : std_logic;
  SIGNAL forwbuf_descriptor_bit3 : std_logic;
  SIGNAL forwbuf_descriptor_bit4 : std_logic;
  SIGNAL forwbuf_descriptor_bit5 : std_logic;
  SIGNAL forwbuf_descriptor_bit6 : std_logic;
  SIGNAL forwbuf_descriptor_bit7 : std_logic;
  SIGNAL forwbuff_position_byteoffset : std_logic_vector(19 downto 0);
  SIGNAL forwbuff_position_bitoffset : std_logic_vector(5 downto 0);
  --SIGNAL forwbuff_position_byteoffset : std_logic_vector(18 downto 0);
  SIGNAL forwbuff_position : std_logic_vector(8 downto 0);

  --SIGNAL forwbuff_position_byteoffset : std_logic_vector(18 downto 0);
  --SIGNAL forwbuff_position_bitoffset : std_logic_vector(5 downto 0);
  SIGNAL free_this_location  : std_logic_vector(31 downto 0); --(18 downto 0);
  SIGNAL which_64bit_isit_tofreeup  : std_logic_vector(2 downto 0);
  SIGNAL which_bit_isit_tofreeup : std_logic_vector(5 downto 0);
  SIGNAL fbm_state : std_logic_vector(7 downto 0);
  
  SIGNAL user_clk_i : std_logic;
  
  SIGNAL wb0_state : std_logic_vector(7 downto 0);
  SIGNAL wb_transaction_complete : std_logic;
  SIGNAL op2p_wb_addr_o_feed : std_logic_vector(31 downto 0);
  SIGNAL op2p_wb_sel_o_feed : std_logic_vector(3 downto 0);
  SIGNAL op2p_wb_data_o_feed : std_logic_vector(31 downto 0);
  SIGNAL start_write_wb0 : std_logic;
  SIGNAL op2p_memory_wb_data_i_latched : std_logic_vector(31 downto 0);
  SIGNAL start_read_wb0 : std_logic;
  SIGNAL rx_fc_nb_latched : std_logic_vector(3 downto 0);
  SIGNAL epif_tx_state : std_logic_vector(7 downto 0);
  SIGNAL pcie_packet_tx_complete : std_logic;
  SIGNAL txtrn_counter : std_logic_vector(7 downto 0);
  SIGNAL packet_state : std_logic_vector(7 downto 0);
  SIGNAL op2p_there_is_a_new_packet_to_transmit : std_logic;
  SIGNAL packet_payloadsize_dwords : std_logic_vector(31 downto 0);
  SIGNAL packet_payloadsize_dwords_p4 : std_logic_vector(31 downto 0);
  SIGNAL op2p_just_received_a_new_packet : std_logic;
  SIGNAL epif_rx_state : std_logic_vector(7 downto 0);
  SIGNAL rx_dst_rdy_n : std_logic;
  SIGNAL trn_rx_counter : std_logic_vector(7 downto 0);
  SIGNAL rxpacket_decodedaddress : std_logic_vector(31 downto 0);
  SIGNAL rxpacket_firstdw_be : std_logic_vector(3 downto 0);
  SIGNAL rxpacket_lastdw_be : std_logic_vector(3 downto 0);
  SIGNAL rxpacket_requesterid : std_logic_vector(15 downto 0);
  SIGNAL packet_state_copy : std_logic_vector(7 downto 0);
  SIGNAL bram_rxpacket_firstdata_address : std_logic_vector(31 downto 0);
  SIGNAL rxpacket_header_dw1 : std_logic_vector(31 downto 0);
  SIGNAL rxpacket_header_dw2 : std_logic_vector(31 downto 0);
  SIGNAL rxpacket_header_dw3 : std_logic_vector(31 downto 0);
  SIGNAL rxpacket_header_dw4 : std_logic_vector(31 downto 0);
  SIGNAL packet_datacount : std_logic_vector(15 downto 0);
  SIGNAL rxpacket_type : std_logic_vector(3 downto 0);
  SIGNAL rxpacket_status : std_logic_vector(3 downto 0);
  SIGNAL rxpacket_sourceid : std_logic_vector(15 downto 0);
  SIGNAL rxpacket_destinationid : std_logic_vector(15 downto 0);
  SIGNAL rxpacket_destinationaddress : std_logic_vector(31 downto 0);
  SIGNAL rxpacket_sourceaddress : std_logic_vector(31 downto 0);
  SIGNAL bit10 : std_logic_vector(1 downto 0);
  SIGNAL op2p_mem_wb_data_i_latched : std_logic_vector(31 downto 0);
  SIGNAL op2p_packet_tx_complete : std_logic;
  --SIGNAL op2p_rdreq_destinationid_regdout : std_logic_vector(31 downto 0);
  SIGNAL trn_reset_n : std_logic;
  SIGNAL cfg_completer_id : std_logic_vector(15 downto 0);
  SIGNAL op2p_forw_freeupaddr_regrd_en_copy : std_logic;
  SIGNAL forwbus_64bit : std_logic_vector(63 downto 0);
  SIGNAL which_64bit_isit : std_logic_vector(2 downto 0);
  SIGNAL forwbus_8bit : std_logic_vector(7 downto 0);
  SIGNAL which_8bit_isit : std_logic_vector(2 downto 0);
  SIGNAL which_bit_isit : std_logic_vector(2 downto 0);
  SIGNAL packetstm_isin_idle : std_logic;
  SIGNAL op2p_wr_anybuffers_empty : std_logic;
  SIGNAL op2p_rdreq_anybuffers_empty : std_logic;
  SIGNAL idmatch : std_logic;

  SIGNAL op2p_local_id_reclocked : std_logic_vector(15 downto 0);
  SIGNAL op2p_local_id_reclocked2 : std_logic_vector(15 downto 0);
  SIGNAL op2p_link_status_reg : std_logic_vector(31 downto 0);
  SIGNAL change_flag_packetstm :  std_logic;
  SIGNAL bram_txpacket_readdata_inrtm : std_logic_vector(31 downto 0);
  SIGNAL txstm_reenable_fc  :  std_logic;
  SIGNAL op2p_reset2  :  std_logic;
  SIGNAL op2p_soft_reset  :  std_logic;
  SIGNAL txstm_haltdata_fc1  :  std_logic;
  SIGNAL txstm_haltdata_fc2  :  std_logic;
  SIGNAL op2p_event_pulse  :  std_logic;
  SIGNAL op2p_forwreq_pointer_regempty2  :  std_logic;
  SIGNAL link_error_count_reg : std_logic_vector(31 downto 0);
  SIGNAL link_errcnt_latchedinidle : std_logic_vector(31 downto 0);
  SIGNAL fc_haltlinkpartner   :  std_logic;
  SIGNAL fc_halted_bylinkpartner   :  std_logic;
  SIGNAL it_is_a_retransmit  :  std_logic;
  SIGNAL op2p_event_pulse_xl  :  std_logic;
  SIGNAL op2p_event_pulse_xl_counter : std_logic_vector(3 downto 0);
  SIGNAL rx_detected :  std_logic;
  SIGNAL rx_detect_ff_clear :  std_logic;




  
-----------------------------------------------------------------------------------------------
	-- COMPONENT DECLARATIONS (introducing the IPs) --------------------------------------------
	
	component aurora_exmpl_des_modified
	port
	 (
    -- User I/O
            RESET             : in std_logic;
            HARD_ERROR        : out std_logic;
            SOFT_ERROR        : out std_logic;
            FRAME_ERROR       : out std_logic;
            ERR_COUNT         : out std_logic_vector(0 to 7);
            LANE_UP           : out std_logic_vector(0 to 1);
            CHANNEL_UP        : out std_logic;
            INIT_CLK          : in  std_logic;
            GT_RESET_IN       : in  std_logic;
	-- Clocks
           GTPD1_P   : in  std_logic;
           GTPD1_N   : in  std_logic;
			  user_clk_i : out std_logic;
			  x25m_clkin  : in  std_logic;
	--from the Frame Generator in the original reference design: (gtp-tx)
        -- User Interface
        TX_D            : in  std_logic_vector(0 to 31); 
        TX_REM          : in  std_logic_vector(0 to 1);     
        TX_SOF_N        : in  std_logic;
        TX_EOF_N        : in  std_logic;
        TX_SRC_RDY_N    : in  std_logic;
        TX_DST_RDY_N    : out   std_logic;  
        -- NFC Interface
        NFC_REQ_N       : in  std_logic;
        NFC_NB          : in  std_logic_vector(0 to 3);     
        NFC_ACK_N       : out   std_logic;  
	--from the Frame Check module in the original reference design: (gtp-rx)
        -- User Interface
        RX_D            : out  std_logic_vector(0 to 31); 
        RX_REM          : out  std_logic_vector(0 to 1);     
        RX_SOF_N        : out  std_logic;
        RX_EOF_N        : out  std_logic;
        RX_SRC_RDY_N    : out  std_logic; 
        -- NFC Interface
        RX_SNF          : out  std_logic;
        RX_FC_NB        : out  std_logic_vector(0 to 3);   
   -- Gbit I/O
            RXP               : in std_logic_vector(0 to 1);
            RXN               : in std_logic_vector(0 to 1);
            TXP               : out std_logic_vector(0 to 1);
            TXN               : out std_logic_vector(0 to 1)
	 );
	end component;

	COMPONENT op2p_host_wb_if
	PORT(
		op2p_config_wb_data_o : IN std_logic_vector(31 downto 0);
		op2p_config_wb_addr_i : IN std_logic_vector(6 downto 0);
		op2p_config_wb_cyc_i : IN std_logic;
		op2p_config_wb_stb_i : IN std_logic;
		op2p_config_wb_wr_i : IN std_logic;
		op2p_config_wb_clk_i : IN std_logic;
		op2p_config_wb_sel_o : IN std_logic_vector(3 downto 0);
		op2p_reset : IN std_logic;
		x25m_clk : IN std_logic;
		user_clk_i : in std_logic;
		op2p_wr_sourceaddress_regrd_en : IN std_logic;
		op2p_wr_destinationaddress_regrd_en : IN std_logic;
		op2p_wr_sourceid_regrd_en : IN std_logic;
		op2p_wr_destinationid_regrd_en : IN std_logic;
		op2p_wr_bytecount_regrd_en : IN std_logic;
		op2p_rdreq_localaddress_regrd_en : IN std_logic;
		op2p_rdreq_destinationaddress_regrd_en : IN std_logic;
		op2p_rdreq_sourceid_regrd_en : IN std_logic;
		op2p_rdreq_destinationid_regrd_en : IN std_logic;
		op2p_rdreq_bytecount_regrd_en : IN std_logic;
		op2p_forw_freeupaddr_regrd_en : IN std_logic;
		op2p_forw_freeupsize_regrd_en : IN std_logic;
		op2p_forwreq_pointer_regdin : IN std_logic_vector(31 downto 0);
		op2p_forwreq_pointer_regwr_en : IN std_logic;
		op2p_rdcompl_localaddress_regdin : IN std_logic_vector(31 downto 0);
		op2p_rdcompl_localaddress_regwr_en : IN std_logic;
		op2p_arrivedwrite_address_regdin : IN std_logic_vector(31 downto 0);
		op2p_arrivedwrite_address_regwr_en : IN std_logic;          
		op2p_config_wb_data_i : OUT std_logic_vector(31 downto 0);
		op2p_config_wb_ack_o : OUT std_logic;
		op2p_irq : OUT std_logic;
		op2p_wr_sourceaddress_regdout : OUT std_logic_vector(31 downto 0);
		op2p_wr_sourceaddress_regempty : OUT std_logic;
		op2p_wr_destinationaddress_regdout : OUT std_logic_vector(31 downto 0);
		op2p_wr_destinationaddress_regempty : OUT std_logic;
		op2p_wr_sourceid_regdout : OUT std_logic_vector(31 downto 0);
		op2p_wr_sourceid_regempty : OUT std_logic;
		op2p_wr_destinationid_regdout : OUT std_logic_vector(31 downto 0);
		op2p_wr_destinationid_regempty : OUT std_logic;
		op2p_wr_bytecount_regdout : OUT std_logic_vector(31 downto 0);
		op2p_wr_bytecount_regempty : OUT std_logic;
		op2p_rdreq_localaddress_regdout : OUT std_logic_vector(31 downto 0);
		op2p_rdreq_localaddress_regempty : OUT std_logic;
		op2p_rdreq_destinationaddress_regdout : OUT std_logic_vector(31 downto 0);
		op2p_rdreq_destinationaddress_regempty : OUT std_logic;
		op2p_rdreq_sourceid_regdout : OUT std_logic_vector(31 downto 0);
		op2p_rdreq_sourceid_regempty : OUT std_logic;
		op2p_rdreq_destinationid_regdout : OUT std_logic_vector(31 downto 0);
		op2p_rdreq_destinationid_regempty : OUT std_logic;
		op2p_rdreq_bytecount_regdout : OUT std_logic_vector(31 downto 0);
		op2p_rdreq_bytecount_regempty : OUT std_logic;
		op2p_local_id : out  std_logic_vector(15 downto 0); 
		op2p_forw_freeupaddr_regdout : OUT std_logic_vector(31 downto 0);
		op2p_forw_freeupaddr_regempty : OUT std_logic;
		op2p_forw_freeupsize_regdout : OUT std_logic_vector(31 downto 0);
		op2p_forw_freeupsize_regempty : OUT std_logic;
		op2p_forwarding_bufferbase_reg : OUT std_logic_vector(31 downto 0);
		op2p_forwarding_bufsize_reg : OUT std_logic_vector(31 downto 0);
		op2p_forwreq_pointer_regfull : OUT std_logic;
		op2p_rdcompl_localaddress_regfull : OUT std_logic;
		op2p_link_status_reg : IN std_logic_vector(31 downto 0);
		op2p_soft_reset  : OUT std_logic;
		op2p_forwreq_pointer_regempty2  : OUT std_logic;
		link_error_count_reg  : IN std_logic_vector(31 downto 0);
		op2p_arrivedwrite_address_regfull : OUT std_logic
		);
	END COMPONENT;

	COMPONENT blk_mem_gen_v4_1
	PORT(
		clka : IN std_logic;
		wea : IN std_logic_vector(0 to 0);
		addra : IN std_logic_vector(8 downto 0);
		dina : IN std_logic_vector(31 downto 0);
		clkb : IN std_logic;
		addrb : IN std_logic_vector(8 downto 0);          
		doutb : OUT std_logic_vector(31 downto 0)
		);
	END COMPONENT;




-- ------- SYNTHESIS ATTRIBUTES: --------------------------------------------------
--attribute keep_hierarchy : string; 
--attribute keep_hierarchy of op2p: entity is "yes"; 
 -- KEEP HIERARCHY
 -- attribute keep : string; 
 -- attribute keep of clock_signal_name: signal is "true"; 
 attribute keep : string; 
 --attribute keep of op2p_memory_wb_clk_o: signal is "true";
 attribute keep of user_clk_i: signal is "true"; 


-----------------------------------------------------------------------------------------------
-- --------ARCHITECTURE BODY BEGINS -----------------------------------------------------------
begin



-----------------------------------------------------------------------------------------------
	-- COMPONENT INSTALLATIONS (connecting the IPs to local signals) ---------------------------
	Inst_aurora_exmpl_des_modified : aurora_exmpl_des_modified
	  port map
		(
		--  User I/O      
		 RESET   =>  op2p_reset2  ,   -- : in std_logic;     
		 HARD_ERROR   =>  HARD_ERROR  ,   -- : out std_logic;     
		 SOFT_ERROR   =>  SOFT_ERROR  ,   -- : out std_logic;     
		 FRAME_ERROR   =>  FRAME_ERROR  ,   -- : out std_logic;     
		 ERR_COUNT   =>  ERR_COUNT  ,   -- : out std_logic_vector(0 to 7);   
		 LANE_UP   =>  LANE_UP  ,   -- : out std_logic_vector(0 to 1);   
		 CHANNEL_UP   =>  CHANNEL_UP  ,   -- : out std_logic;     
		 INIT_CLK   =>  INIT_CLK  ,   -- : in std_logic;     
		 GT_RESET_IN   =>  GT_RESET_IN  ,   -- : in std_logic;     
		 -- Clocks       
		 GTPD1_P   =>  GTPD1_P  ,   -- : in std_logic;     
		 GTPD1_N   =>  GTPD1_N  ,   -- : in std_logic;
		 user_clk_i => user_clk_i,
		 x25m_clkin  => x25m_clk,
		-- the Frame Generator in the original reference design:
		 -- User Interface      
		 TX_D   =>  TX_D  ,   -- : out std_logic_vector(0 to 31);   
		 TX_REM   =>  TX_REM  ,   -- : out std_logic_vector(0 to 1);    
		 TX_SOF_N   =>  TX_SOF_N  ,   -- : out std_logic;      
		 TX_EOF_N   =>  TX_EOF_N  ,   -- : out std_logic;      
		 TX_SRC_RDY_N   =>  TX_SRC_RDY_N  ,   -- : out std_logic;      
		 TX_DST_RDY_N   =>  TX_DST_RDY_N  ,   -- : in std_logic;      
		 -- NFC Interface       
		 NFC_REQ_N   =>  NFC_REQ_N  ,   -- : out std_logic;      
		 NFC_NB   =>  NFC_NB  ,   -- : out std_logic_vector(0 to 3);    
		 NFC_ACK_N   =>  NFC_ACK_N  ,   -- : in std_logic;        
		-- the Frame Check module in the original reference design:
		 -- User Interface       
		 RX_D   =>  RX_D  ,   -- : in std_logic_vector(0 to 31);    
		 RX_REM   =>  RX_REM  ,   -- : in std_logic_vector(0 to 1);
		 RX_SOF_N   =>  RX_SOF_N  ,   -- : in std_logic;  
		 RX_EOF_N   =>  RX_EOF_N  ,   -- : in std_logic;  
		 RX_SRC_RDY_N   =>  RX_SRC_RDY_N  ,   -- : in std_logic;  
		 -- NFC Interface   
		 RX_SNF   =>  RX_SNF  ,   -- : in std_logic;  
		 RX_FC_NB   =>  RX_FC_NB  ,   -- : in std_logic_vector(0 to 3); 
		-- V5 I/O   
		 RXP   =>  op2p_RXP  ,   -- : in std_logic_vector(0 to 1);
		 RXN   =>  op2p_RXN  ,   -- : in std_logic_vector(0 to 1);
		 TXP   =>  op2p_TXP  ,   -- : out std_logic_vector(0 to 1);
		 TXN   =>  op2p_TXN     -- : out std_logic_vector(0 to 1)
		 ); 


	--the wishbone slave interface with its FIFOs.
	Inst_op2p_host_wb_if: op2p_host_wb_if PORT MAP(
	 op2p_config_wb_data_o => op2p_config_wb_data_o ,
	 op2p_config_wb_data_i => op2p_config_wb_data_i ,
	 op2p_config_wb_addr_i => op2p_config_wb_addr_i ,
	 op2p_config_wb_cyc_i => op2p_config_wb_cyc_i ,
	 op2p_config_wb_stb_i => op2p_config_wb_stb_i ,
	 op2p_config_wb_wr_i => op2p_config_wb_wr_i ,
	 op2p_config_wb_ack_o => op2p_config_wb_ack_o ,
	 op2p_config_wb_clk_i => op2p_config_wb_clk_i ,
	 op2p_config_wb_sel_o => op2p_config_wb_sel_o ,
	 op2p_reset => op2p_reset ,
	 x25m_clk => x25m_clk ,
	 user_clk_i => user_clk_i,
	 op2p_irq => op2p_irq_not_used ,
	 op2p_wr_sourceaddress_regrd_en => op2p_wr_sourceaddress_regrd_en ,
	 op2p_wr_sourceaddress_regdout => op2p_wr_sourceaddress_regdout ,
	 op2p_wr_sourceaddress_regempty => op2p_wr_sourceaddress_regempty ,
	 op2p_wr_destinationaddress_regrd_en => op2p_wr_destinationaddress_regrd_en ,
	 op2p_wr_destinationaddress_regdout => op2p_wr_destinationaddress_regdout ,
	 op2p_wr_destinationaddress_regempty => op2p_wr_destinationaddress_regempty ,
	 op2p_wr_sourceid_regrd_en => op2p_wr_sourceid_regrd_en ,
	 op2p_wr_sourceid_regdout => op2p_wr_sourceid_regdout ,
	 op2p_wr_sourceid_regempty => op2p_wr_sourceid_regempty ,
	 op2p_wr_destinationid_regrd_en => op2p_wr_destinationid_regrd_en ,
	 op2p_wr_destinationid_regdout => op2p_wr_destinationid_regdout ,
	 op2p_wr_destinationid_regempty => op2p_wr_destinationid_regempty ,
	 op2p_wr_bytecount_regrd_en => op2p_wr_bytecount_regrd_en ,
	 op2p_wr_bytecount_regdout => op2p_wr_bytecount_regdout ,
	 op2p_wr_bytecount_regempty => op2p_wr_bytecount_regempty ,
	 op2p_rdreq_localaddress_regrd_en => op2p_rdreq_localaddress_regrd_en ,
	 op2p_rdreq_localaddress_regdout => op2p_rdreq_localaddress_regdout ,
	 op2p_rdreq_localaddress_regempty => op2p_rdreq_localaddress_regempty ,
	 op2p_rdreq_destinationaddress_regrd_en => op2p_rdreq_destinationaddress_regrd_en ,
	 op2p_rdreq_destinationaddress_regdout => op2p_rdreq_destinationaddress_regdout ,
	 op2p_rdreq_destinationaddress_regempty => op2p_rdreq_destinationaddress_regempty ,
	 op2p_rdreq_sourceid_regrd_en => op2p_rdreq_sourceid_regrd_en ,
	 op2p_rdreq_sourceid_regdout => op2p_rdreq_sourceid_regdout ,
	 op2p_rdreq_sourceid_regempty => op2p_rdreq_sourceid_regempty ,
	 op2p_rdreq_destinationid_regrd_en => op2p_rdreq_destinationid_regrd_en ,
	 op2p_rdreq_destinationid_regdout => op2p_rdreq_destinationid_regdout ,
	 op2p_rdreq_destinationid_regempty => op2p_rdreq_destinationid_regempty ,
	 op2p_rdreq_bytecount_regrd_en => op2p_rdreq_bytecount_regrd_en ,
	 op2p_rdreq_bytecount_regdout => op2p_rdreq_bytecount_regdout ,
	 op2p_rdreq_bytecount_regempty => op2p_rdreq_bytecount_regempty ,
	 op2p_local_id => op2p_local_id,
	 op2p_forw_freeupaddr_regrd_en => op2p_forw_freeupaddr_regrd_en ,
	 op2p_forw_freeupaddr_regdout => op2p_forw_freeupaddr_regdout ,
	 op2p_forw_freeupaddr_regempty => op2p_forw_freeupaddr_regempty ,
	 op2p_forw_freeupsize_regrd_en => op2p_forw_freeupsize_regrd_en ,
	 op2p_forw_freeupsize_regdout => op2p_forw_freeupsize_regdout ,
	 op2p_forw_freeupsize_regempty => op2p_forw_freeupsize_regempty ,
	 op2p_forwarding_bufferbase_reg => op2p_forwarding_bufferbase_reg ,
	 op2p_forwarding_bufsize_reg => op2p_forwarding_bufsize_reg ,
	 op2p_forwreq_pointer_regdin => op2p_forwreq_pointer_regdin ,
	 op2p_forwreq_pointer_regwr_en => op2p_forwreq_pointer_regwr_en ,
	 op2p_forwreq_pointer_regfull => op2p_forwreq_pointer_regfull ,
	 op2p_rdcompl_localaddress_regdin => op2p_rdcompl_localaddress_regdin ,
	 op2p_rdcompl_localaddress_regwr_en => op2p_rdcompl_localaddress_regwr_en ,
	 op2p_rdcompl_localaddress_regfull => op2p_rdcompl_localaddress_regfull ,
	 op2p_arrivedwrite_address_regdin => op2p_arrivedwrite_address_regdin ,
	 op2p_arrivedwrite_address_regwr_en => op2p_arrivedwrite_address_regwr_en ,
	 op2p_link_status_reg => op2p_link_status_reg ,
	 op2p_soft_reset  => op2p_soft_reset,
	 op2p_forwreq_pointer_regempty2  => op2p_forwreq_pointer_regempty2,
	 link_error_count_reg => link_error_count_reg,
	 op2p_arrivedwrite_address_regfull => op2p_arrivedwrite_address_regfull 
	);

	--block ram for RX packet:
	Inst_bram_rxpacket: blk_mem_gen_v4_1 PORT MAP(
		clka => user_clk_i,
		wea => bram_rxpacket_we,
		addra => bram_rxpacket_writeaddress(8 downto 0),
		dina => bram_rxpacket_writedata,
		clkb => user_clk_i,
		addrb => bram_rxpacket_readaddress(8 downto 0),
		doutb => bram_rxpacket_readdata
	);

	--block ram for TX packet:
	Inst_bram_txpacket: blk_mem_gen_v4_1 PORT MAP(
		clka => user_clk_i,
		wea => bram_txpacket_we,
		addra => bram_txpacket_writeaddress(8 downto 0),
		dina => bram_txpacket_writedata,
		clkb => user_clk_i,
		addrb => bram_txpacket_readaddress(8 downto 0),
		doutb => bram_txpacket_readdata
	); 
				
				
				
-----------------------------------------------------------------------------------------------
	-- MAIN LOGIC: -----------------------------------------------------------------------------



	--controlled reset:
	--from 2 sources: HW reset from host (PCIe) and from a soft port reset register
	op2p_reset2 <= op2p_reset or op2p_soft_reset;
	
	
	--INTERRUPT TO HOST:
	--Active high
	--This gets asserted if any data arrived, if outgoing write has finished, if  forwarding buffer has something in it.
	op2p_irq <= op2p_event_pulse_xl;
	--op2p_irq <= op2p_event_pulse or (not op2p_forwreq_pointer_regempty2); --event pulse gets asserted even when a fw packet is stored.
	--the fifo status register tells if there is a pointer in the forw_req FIFO.
	--or use it from the wb slave state machine:
	--op2p_irq <= op2p_irq_not_used;
	--Generate a longer/detectable pulse, since it will cross clock domains
	process (trn_reset_n, user_clk_i) 
	begin
	if (trn_reset_n='0') then 
		op2p_event_pulse_xl <= '0';
		op2p_event_pulse_xl_counter <= (OTHERS => '0');
	else
		if (user_clk_i'event and user_clk_i = '1') then
			if (op2p_event_pulse='1') then
			  op2p_event_pulse_xl <= '1';
			  op2p_event_pulse_xl_counter <= (OTHERS => '0');
			elsif (op2p_event_pulse_xl_counter="1000") then
			  op2p_event_pulse_xl <= '0';
			  --counter stays at value
			else
			  op2p_event_pulse_xl_counter <= op2p_event_pulse_xl_counter +1;
			end if;
		end if;        
	end if;
	end process;


	--LINK STATUS connections:
	--THIS HAS TO BE MODIFIED BASED ON THE NUMBER OF LANES USED
	op2p_link_status_reg(0) <= CHANNEL_UP;
	op2p_link_status_reg(2 downto 1) <= LANE_UP (0 to 1); --LANE_UP : out std_logic_vector(0 to 1)
	op2p_link_status_reg(28 downto 3)  <= (OTHERS => '0');
	op2p_link_status_reg(29) <= fc_haltlinkpartner;
	op2p_link_status_reg(30) <= fc_halted_bylinkpartner;
	op2p_link_status_reg(31) <= HARD_ERROR;
	CHANNEL_UP_copy <= CHANNEL_UP;


	--aurora interface FIX conenctions:
	RESET <= op2p_reset;
	trn_reset_n <= not op2p_reset2;
	INIT_CLK <= x25m_clk; --Debounce the GT_RESET_IN signal using the INIT_CLK
	GT_RESET_IN <= op2p_reset2;
	op2p_memory_wb_clk_o <=  user_clk_i;
	
	
	--Set reference clock to be 75MHz (generated from 25MHz source driven by the FPGA):
	--On-board CDCM61001 clock chip setting:
			  op2p_refclkset_od0  <= '1';
			  op2p_refclkset_od1  <= '1';
			  op2p_refclkset_od2  <= '1';
			  op2p_refclkset_pr0  <= '0';
			  op2p_refclkset_pr1  <= '0';


	--check if a new command has arrived.
	--Do this by checking the empty flags of the FIFOs.
	--Wait until all necessary FIFOs are filled up, before initiating an OP2P transaction.
	process (trn_reset_n, user_clk_i) 
	begin
	if (trn_reset_n='0') then 
			op2p_wr_anybuffers_empty <= '1';
			op2p_rdreq_anybuffers_empty <= '1';
	else
		if (user_clk_i'event and user_clk_i = '1') then
			--wr:
			op2p_wr_anybuffers_empty <=  op2p_wr_sourceaddress_regempty 
					or op2p_wr_destinationaddress_regempty 
					or op2p_wr_sourceid_regempty 
					or op2p_wr_destinationid_regempty 
					or op2p_wr_bytecount_regempty ;
			--rd:
			op2p_rdreq_anybuffers_empty <=  op2p_rdreq_localaddress_regempty
					or op2p_rdreq_destinationaddress_regempty 
					or op2p_rdreq_sourceid_regempty 
					or op2p_rdreq_destinationid_regempty 
					or op2p_rdreq_bytecount_regempty ;		
		end if;        
	end if;
	end process;


	--CHECK FOR IDMATCH.
	process (trn_reset_n, user_clk_i, packet_state) 
	begin
	if (trn_reset_n='0') then 
		idmatch <= '0';
		op2p_local_id_reclocked <= (OTHERS => '0');
		op2p_local_id_reclocked2 <= (OTHERS => '0');
	else
		if (user_clk_i'event and user_clk_i = '1') then
			op2p_local_id_reclocked <= op2p_local_id;
			op2p_local_id_reclocked2 <= op2p_local_id_reclocked;
			if (packet_state = "00000001") then
				if ((rxpacket_destinationid (15 downto 0) = op2p_local_id_reclocked2(15 downto 0))
						or (rxpacket_destinationid (15 downto 0) = "0000000000000000")) then
					idmatch <= '1';
				else
					idmatch <= '0';
				end if;
			end if;  
		end if;        
	end if;
	end process;
  
  
	--Count link errors: (max 4 billion)
	process (trn_reset_n, user_clk_i) 
	begin
	if (trn_reset_n='0') then 
		link_error_count_reg <= (OTHERS => '0');
	else
		if (user_clk_i'event and user_clk_i = '1') then
			if (SOFT_ERROR='1' or FRAME_ERROR='1') then
			  link_error_count_reg <= link_error_count_reg +1;
			end if;
		end if;        
	end if;
	end process;


	--RX detection flip-flop
	process (trn_reset_n, user_clk_i)
	begin
	if (trn_reset_n='0') then 
		rx_detected <= '0';
	else
		if (user_clk_i'event and user_clk_i = '1') then
			if (op2p_just_received_a_new_packet ='1') then
			  rx_detected <= '1';
			elsif (rx_detect_ff_clear ='1') then
			  rx_detected <= '0';
			end if;
		end if;        
	end if;
	end process;





	-- -----------------------------------------------------------------------------
	-- WISBONE Master INTERFACE ----------------------------------------------------
	--This is for accessing the local memory.

    --main state machine: set states, capture inputs, set addr/data outputs
	 --minimum 2 clock cycles / transaction. writes are posted, reads have wait states.
    process (op2p_reset2, user_clk_i, wb0_state, start_read_wb0, start_write_wb0,
				op2p_wb_addr_o_feed, op2p_wb_data_o_feed, op2p_wb_sel_o_feed) 
    begin
    if (op2p_reset2='1') then 
       wb0_state <= "00000000";
       wb_transaction_complete <= '0';
		 op2p_memory_wb_addr_o <= "00000000000000000000000000";
		 op2p_memory_wb_sel_o <= "0000";
		 op2p_memory_wb_data_o <= "00000000000000000000000000000000";
		 op2p_mem_wb_data_i_latched <= (OTHERS => '0');
		 
    else
      if (user_clk_i'event and user_clk_i = '1') then
                case ( wb0_state ) is

                --********** IDLE STATE  **********
                when "00000000" =>   --state 0        
                    wb_transaction_complete <='0';
                    op2p_memory_wb_addr_o <= op2p_wb_addr_o_feed (25 downto 0);
                    op2p_memory_wb_sel_o <= op2p_wb_sel_o_feed;
                    op2p_memory_wb_data_o <= op2p_wb_data_o_feed;
						  if (start_read_wb0 ='1') then --go to read
						    wb0_state <= "00000001";
						  elsif (start_write_wb0 ='1') then --go to write
						    wb0_state <= "00000010";
						  end if;

                --********** READ STATE ********** 
					 --set the outputs, 
					 --if ACK asserted, sample the data input
					 --The hold requirements are oversatisfyed by going back to idle, 
					 --and by the fact that the slave uses the cyc/stb/wr strobes synchronously.
                when "00000001" =>   --state 1
                    if (op2p_memory_wb_ack_i='1') then
						    op2p_mem_wb_data_i_latched <= op2p_memory_wb_data_i; --sample the incoming data
							 wb_transaction_complete <='1'; --signalling ready, but only for one clock cycle
							 wb0_state <= "00000000"; --go to state 0
						  else
						  	 wb_transaction_complete <='0';
						  end if;	   		  

                --********** WRITE STATE **********     
					 --if ACK asserted, go back to idle
					 --The hold requirements are oversatisfyed by waiting for ACK to remove write data					 
                when "00000010" =>   --state 2
                    if (op2p_memory_wb_ack_i='1') then
							 wb0_state <= "00000000"; --go to state 0
							 wb_transaction_complete <='1';
						  else
						     wb_transaction_complete <='0';
						  end if;
						  
                when others => --error
                      wb0_state <= "00000000"; --go to state 0
                end case;     
       end if;        
    end if;
    end process;
    --sync control on wb-control signals:
    process (op2p_reset2, wb0_state) 
    begin
    if (op2p_reset2='1') then 
		op2p_memory_wb_cyc_o  <= '0';
		op2p_memory_wb_stb_o  <= '0';
		op2p_memory_wb_wr_o  <= '0';
    else
      if (wb0_state = "00000000") then --idle
			op2p_memory_wb_cyc_o  <= '0';
			op2p_memory_wb_stb_o  <= '0';
			op2p_memory_wb_wr_o  <= '0';
      elsif (wb0_state = "00000001") then --read 
			op2p_memory_wb_cyc_o  <= '1';
			op2p_memory_wb_stb_o  <= '1';
			op2p_memory_wb_wr_o  <= '0';
      elsif (wb0_state = "00000010") then --write 
			op2p_memory_wb_cyc_o  <= '1';
			op2p_memory_wb_stb_o  <= '1';
			op2p_memory_wb_wr_o  <= '1';
		else
			op2p_memory_wb_cyc_o  <= '0';
			op2p_memory_wb_stb_o  <= '0';
			op2p_memory_wb_wr_o  <= '0';
		end if;
    end if;
    end process;







	-- -----------------------------------------------------------------------------------
	-- INTERFACE TO THE aurora-IP --------------------------------------------------------
	
	--what to do with these?
        --TX_REM          : in  std_logic_vector(0 to 1); 
		  --Specifies the number of valid bytes in the last data beat;
		  --valid only while TX_EOF_N is asserted. REM bus widths
		  --are given by [0:r(n)], where r(n) = ceiling [{log2(n)}-1].
		  --The TX_REM bus is used to indicate the number of valid bytes in the final word of the frame.
		  TX_REM <= "11"; --always all 4 bytes of a dword valid.
		  
        --RX_REM          : out  std_logic_vector(0 to 1); 
		  --Specifies the number of valid bytes in the last data beat;
		  --valid only when RX_EOF_N is asserted. REM bus widths
		  --are given by [0:r(n)], where r(n) = ceiling [{log2(n)}-1].
		  --dont conenct.

	--FLOW CONTROL ---------------------------------------
	--Flow control logic is built into the TX statemachine.
	--The Aurora 8B/10B protocol includes native flow control (NFC) to allow receivers to
	--control the rate at which data is sent to them by specifying a number of idle data beats that
	--must be placed into the data stream. The data flow can even be turned off completely by
	--requesting that the transmitter temporarily send only idles (XOFF).
	--To send an NFC message to a channel partner, the user application asserts NFC_REQ_N
	--and writes an NFC code to NFC_NB. The NFC code indicates the minimum number of idle
	--cycles the channel partner should insert in its TX data stream. The user application must
	--hold NFC_REQ_N and NFC_NB until NFC_ACK_N is asserted on a positive USER_CLK
	--edge, indicating the Aurora 8B/10B core will transmit the NFC message.
	--Aurora 8B/10B cores cannot transmit data while sending NFC messages.
	--
	 --In this code, we only support NFC_NB=1111=wait or 0000=ready
	 --only allow packets to arrive when the packet buffer is not in use by the scheduler. 
	 
	 --latch the latest flow control state. 0000=ready, 1111=wait, others not supported (assumes wait)
	 process ( op2p_reset2, user_clk_i, RX_FC_NB)
    begin
       if (op2p_reset2='1') then
         RX_FC_NB_latched <= "0000";
			fc_halted_bylinkpartner <= '0';
       elsif (user_clk_i'event and user_clk_i='1') then
         if (RX_SNF='1') then
			  RX_FC_NB_latched <= RX_FC_NB;
			  if (RX_FC_NB="1111") then
			     fc_halted_bylinkpartner <= '1';
			  else
			     fc_halted_bylinkpartner <= '0';
			  end if;
			end if;
       end if;
    end process;	


	-- TX: INTERFACE TO THE aurora-IP: TRANSMIT  PACKETS:-----
    process (op2p_reset2, user_clk_i, epif_tx_state, bram_txpacket_readdata, bram_txpacket_readaddress, txstm_reenable_fc,
				op2p_there_is_a_new_packet_to_transmit, packet_payloadsize_dwords, txtrn_counter, packetstm_isin_idle,
				NFC_ACK_N, RX_SNF, RX_FC_NB, op2p_forwreq_pointer_regfull, bram_txpacket_readdata_inrtm) 
    begin
    if (op2p_reset2='1') then 
      epif_tx_state <= "00000000";
      TX_SRC_RDY_N <='1';
		TX_SOF_N <= '1';
		TX_EOF_N <= '1';
		TX_D <= (OTHERS => '0');
		op2p_packet_tx_complete <= '0';
		txtrn_counter <= "00000001";
		bram_txpacket_readaddress <= (OTHERS => '0');
		NFC_REQ_N <= '1'; --flow control wait request off
		NFC_NB <= "0000";
		fc_haltlinkpartner <= '0';
    else
      if (user_clk_i'event and user_clk_i = '1') then
                bram_txpacket_readdata_inrtm <= bram_txpacket_readdata; --break timing path
					 case ( epif_tx_state ) is

                --********** idle STATE  **********
                when "00000000" =>   --state 0        
                    --if there is a new packet assembled and the EP is ready,  
						  --start the tx-trn bus transaction.
						  if (op2p_there_is_a_new_packet_to_transmit='1' --scheduler ordered a transmit
								and TX_DST_RDY_N='0'							--aurora ip ready
								and fc_halted_bylinkpartner = '0') then    --other end did not request a wait
						    epif_tx_state <= "00000001"; --next state 1
						  elsif (txstm_reenable_fc = '1') then --main scheduler finished last transaction
						  --elsif ((txstm_reenable_fc = '1') and (op2p_forwreq_pointer_regfull='0')) then
						    epif_tx_state <= "00000101"; --re-enable flow control, to allow packets to arrive here.
						  elsif (op2p_forwreq_pointer_regfull='1' --dont send more forwarding or any packet
									or txstm_haltdata_fc2 = '1' --main sch initiated some transaction. single pulse
									or txstm_haltdata_fc1 = '1') then --RXSTM finished filling up buffer. single pulse
									--or packet_state="00000001" --the local scheduler is processing the last received packed data
									--or packet_state="00000010" 
									--or packet_state="00000110" 
									--or packet_state="00000111" 
									--or packet_state="00001000") then --scheduler's read state 
						    epif_tx_state <= "00000100"; --flow control wait request  STATE
						  end if;
                    TX_SRC_RDY_N <='1';
						  TX_SOF_N <= '1';
						  TX_EOF_N <= '1';
						  TX_D <= (OTHERS => '0');
						  op2p_packet_tx_complete <= '0';
						  txtrn_counter <= "00000001";
						  bram_txpacket_readaddress <= (OTHERS => '0');
						  NFC_REQ_N <= '1'; --flow control wait request off

                --********** ready-wait STATE  **********
                when "00000001" =>   --state 1        
                    --if there is a new TLP assembled and the EP is ready, 
						  --start the tx-trn bus transaction.
						  if (TX_DST_RDY_N='0') then
						    epif_tx_state <= "00000010"; --next state
							 bram_txpacket_readaddress <= bram_txpacket_readaddress +1;
						  else
						    bram_txpacket_readaddress <= (OTHERS => '0');
						  end if;
                    TX_SRC_RDY_N <='1';
						  TX_SOF_N <= '1';
						  TX_EOF_N <= '1';
						  TX_D <= (OTHERS => '0');
						  op2p_packet_tx_complete <= '0';
						  txtrn_counter <= "00000001";
						  
						  
                --********** transfer STATE **********     				 
                when "00000010" =>   --state 2
                    TX_SRC_RDY_N <='0';
						  --Lounch data, and turn it around as well:
						  TX_D (0) <= bram_txpacket_readdata_inrtm(31);
						  TX_D (1) <= bram_txpacket_readdata_inrtm(30);
						  TX_D (2) <= bram_txpacket_readdata_inrtm(29);
						  TX_D (3) <= bram_txpacket_readdata_inrtm(28);
						  TX_D (4) <= bram_txpacket_readdata_inrtm(27);
						  TX_D (5) <= bram_txpacket_readdata_inrtm(26);
						  TX_D (6) <= bram_txpacket_readdata_inrtm(25);
						  TX_D (7) <= bram_txpacket_readdata_inrtm(24);
						  TX_D (8) <= bram_txpacket_readdata_inrtm(23);
						  TX_D (9) <= bram_txpacket_readdata_inrtm(22);
						  TX_D (10) <= bram_txpacket_readdata_inrtm(21);
						  TX_D (11) <= bram_txpacket_readdata_inrtm(20);
						  TX_D (12) <= bram_txpacket_readdata_inrtm(19);
						  TX_D (13) <= bram_txpacket_readdata_inrtm(18);
						  TX_D (14) <= bram_txpacket_readdata_inrtm(17);
						  TX_D (15) <= bram_txpacket_readdata_inrtm(16);
						  TX_D (16) <= bram_txpacket_readdata_inrtm(15);
						  TX_D (17) <= bram_txpacket_readdata_inrtm(14);
						  TX_D (18) <= bram_txpacket_readdata_inrtm(13);
						  TX_D (19) <= bram_txpacket_readdata_inrtm(12);
						  TX_D (20) <= bram_txpacket_readdata_inrtm(11);
						  TX_D (21) <= bram_txpacket_readdata_inrtm(10);
						  TX_D (22) <= bram_txpacket_readdata_inrtm(9);
						  TX_D (23) <= bram_txpacket_readdata_inrtm(8);
						  TX_D (24) <= bram_txpacket_readdata_inrtm(7);
						  TX_D (25) <= bram_txpacket_readdata_inrtm(6);
						  TX_D (26) <= bram_txpacket_readdata_inrtm(5);
						  TX_D (27) <= bram_txpacket_readdata_inrtm(4);
						  TX_D (28) <= bram_txpacket_readdata_inrtm(3);
						  TX_D (29) <= bram_txpacket_readdata_inrtm(2);
						  TX_D (30) <= bram_txpacket_readdata_inrtm(1);
						  TX_D (31) <= bram_txpacket_readdata_inrtm(0);
						  if (TX_DST_RDY_N='0') then 
						    txtrn_counter <= txtrn_counter +1;
							 bram_txpacket_readaddress <= bram_txpacket_readaddress +1;
						  end if;
						  if (txtrn_counter = "00000010") then
						    TX_SOF_N <= '0'; --start
						  else
						    TX_SOF_N <= '1';
						  end if;
						  --test number of dwords:
						  if (txtrn_counter = packet_payloadsize_dwords +5) then -- "+4" is the header and "+1" is for the delay
						  --this is the last dword, next clk is next state
							 epif_tx_state <= "01100100"; --back to idle, since finished, after an intermediate wait state
						    TX_EOF_N <= '0'; --end
						    op2p_packet_tx_complete <= '1'; --assert for 1 clk
						  else
						    TX_EOF_N <= '1'; --not end yet
						    op2p_packet_tx_complete <= '0'; --not complete yet
						  end if;

                --********** wait STATE **********
					 --wait one clock cycle before going back to idle
                when "01100100" =>   --state x
						  epif_tx_state <= "00000000";
                    TX_SRC_RDY_N <='1';
						  TX_SOF_N <= '1';
						  TX_EOF_N <= '1';
						  TX_D <= (OTHERS => '0');
						  op2p_packet_tx_complete <= '0';
						  txtrn_counter <= "00000001";
						  bram_txpacket_readaddress <= (OTHERS => '0');
						  NFC_REQ_N <= '1'; --flow control wait request off

                --********** flow control wait request STATE **********
					 --ask the link partner to wait
                when "00000100" =>   --state 4
                    NFC_NB <= "1111"; --pause: do not send me more data for now
						  fc_haltlinkpartner <= '1'; --registerbit, telling that we have halted the link partner
						  if ( NFC_ACK_N='0') then
						    NFC_REQ_N <= '1'; --flow control wait request off
							 epif_tx_state <= "00000000"; --back to idle
 						  else
						    NFC_REQ_N <= '0'; --flow control wait request on
						  end if;

                --********** flow control re-enable STATE ********** 
					 --Re-enable (for the link-partner) the transmission , if the scheduler 
					 --is in idle, or at least not currently using the RX_packet packet buffer.
                when "00000101" =>   --state 5
                    NFC_NB <= "0000"; --enable data flow
						  fc_haltlinkpartner <= '0';  --registerbit, telling that we have reenabled the link partner
							  if ( NFC_ACK_N='0') then
								 NFC_REQ_N <= '1'; --flow control wait request off
								 epif_tx_state <= "00000000"; --back to idle
							  else
								 NFC_REQ_N <= '0'; --flow control wait request on
							  end if;


                when others => --error
                    epif_tx_state <= "00000000"; --back to idle
                    TX_SRC_RDY_N <='1';
						  TX_SOF_N <= '1';
						  TX_EOF_N <= '1';
						  TX_D <= (OTHERS => '0');
						  op2p_packet_tx_complete <= '0';
						  txtrn_counter <= "00000001";
						  
                end case;     
       end if;        
    end if;
    end process;
	 



	-- RX: INTERFACE TO THE aurora-IP: GET the received packet PACKETS:- ----
    process (op2p_reset2, user_clk_i, epif_rx_state, packet_state, trn_rx_counter,
				bram_rxpacket_writeaddress, packetstm_isin_idle) 
    begin
    if (op2p_reset2='1') then 
       bram_rxpacket_writedata <= (OTHERS => '0');
		 bram_rxpacket_we <=  "0"; 
		 op2p_just_received_a_new_packet <= '0'; 
		 epif_rx_state	<= "00000000"; 
		 RX_Dst_rdy_n <= '1';
		 trn_rx_counter <= (OTHERS => '0');
		 bram_rxpacket_writeaddress <=  (OTHERS => '0');
		 txstm_haltdata_fc1 <= '0'; --data can come in 
    else
      if (user_clk_i'event and user_clk_i = '1') then

                case ( epif_rx_state ) is

                --********** idle STATE  **********
                when "00000000" =>   --state 0
						  op2p_just_received_a_new_packet <= '0';
						  bram_rxpacket_writedata  <= RX_D;
						  txstm_haltdata_fc1 <= '0'; --reset this signal
						  if (RX_SRC_RDY_N='0' and RX_SOF_N='0' and packetstm_isin_idle = '1' and RX_Dst_rdy_n='0') then 
						    trn_rx_counter <= trn_rx_counter +1;
							 bram_rxpacket_writeaddress <= bram_rxpacket_writeaddress +1;
							 epif_rx_state <= "00000001";
						  else
						    trn_rx_counter <= (OTHERS => '0');
							 bram_rxpacket_writeaddress  <= (OTHERS => '0');
						  end if;
						  --destination ready:
						  if (packetstm_isin_idle = '1')then
							  RX_Dst_rdy_n <= '0';
						  else
							  RX_Dst_rdy_n <= '1';
						  end if;
						  --write into buffer:
						  if (RX_SRC_RDY_N='0' and RX_SOF_N='0' and packetstm_isin_idle = '1') then 
							 bram_rxpacket_we <= "1";
						  else
							 bram_rxpacket_we <= "0";
						  end if;

                --********** read STATE ********** 
                when "00000001" =>   --state 1
						  if (RX_EOF_N ='0') then --last dw
						    epif_rx_state <= "00000010"; --for the next clk cycle
							 RX_Dst_rdy_n <= '1'; --ok, dont send more yet
							 txstm_haltdata_fc1 <= '1'; --dont send more yet
						  end if;
						  if (RX_SRC_RDY_N='0') then --only act if the EP was ready
							  trn_rx_counter <= trn_rx_counter +1;
							  --get the data, and turn it around as well:
							  bram_rxpacket_writedata (0) <= RX_D(31);
							  bram_rxpacket_writedata (1) <= RX_D(30);
							  bram_rxpacket_writedata (2) <= RX_D(29);
							  bram_rxpacket_writedata (3) <= RX_D(28);
							  bram_rxpacket_writedata (4) <= RX_D(27);
							  bram_rxpacket_writedata (5) <= RX_D(26);
							  bram_rxpacket_writedata (6) <= RX_D(25);
							  bram_rxpacket_writedata (7) <= RX_D(24);
							  bram_rxpacket_writedata (8) <= RX_D(23);
							  bram_rxpacket_writedata (9) <= RX_D(22);
							  bram_rxpacket_writedata (10) <= RX_D(21);
							  bram_rxpacket_writedata (11) <= RX_D(20);
							  bram_rxpacket_writedata (12) <= RX_D(19);
							  bram_rxpacket_writedata (13) <= RX_D(18);
							  bram_rxpacket_writedata (14) <= RX_D(17);
							  bram_rxpacket_writedata (15) <= RX_D(16);
							  bram_rxpacket_writedata (16) <= RX_D(15);
							  bram_rxpacket_writedata (17) <= RX_D(14);
							  bram_rxpacket_writedata (18) <= RX_D(13);
							  bram_rxpacket_writedata (19) <= RX_D(12);
							  bram_rxpacket_writedata (20) <= RX_D(11);
							  bram_rxpacket_writedata (21) <= RX_D(10);
							  bram_rxpacket_writedata (22) <= RX_D(9);
							  bram_rxpacket_writedata (23) <= RX_D(8);
							  bram_rxpacket_writedata (24) <= RX_D(7);
							  bram_rxpacket_writedata (25) <= RX_D(6);
							  bram_rxpacket_writedata (26) <= RX_D(5);
							  bram_rxpacket_writedata (27) <= RX_D(4);
							  bram_rxpacket_writedata (28) <= RX_D(3);
							  bram_rxpacket_writedata (29) <= RX_D(2);
							  bram_rxpacket_writedata (30) <= RX_D(1);
							  bram_rxpacket_writedata (31) <= RX_D(0);
							  bram_rxpacket_we <=  "1"; 
							  bram_rxpacket_writeaddress <= bram_rxpacket_writeaddress +1;
						  else
						    bram_rxpacket_we <=  "0"; 
						  end if;
						  if (trn_rx_counter = "00000010") then
						   op2p_just_received_a_new_packet <= '1';--assert for one clk only
						  else
						   op2p_just_received_a_new_packet <= '0';
						  end if;

                --********** finished filling up RX packet STATE **********     				 
                when "00000010" =>   --state 2
                    op2p_just_received_a_new_packet <= '0';--deassert
						  epif_rx_state <= "00000000";
						  trn_rx_counter <= (OTHERS => '0');
						  bram_rxpacket_we <=  "0";
						  bram_rxpacket_writeaddress <=  (OTHERS => '0');
						  
                when others => --error
                      epif_rx_state <= "00000000"; --go to state 0
                end case;     
       end if;        
    end if;
    end process;
	 







	-- -----------------------------------------------------------------------------------
	-- --- MAIN SCHEDULER ----------------------------------------------------------------
	-- --- ALSO PACKET PROCESSING.

	-- Packet format: Header + payload data. Max 2kBytes in one packet. If the request is tergating
	--  a larger than 2kBytes memory area, then the scheduler has to divide the data into 2kB packets.
	--  Header: 
	--    1st DW: source ID (16bit 31:16), destination ID (16bit 15:0)
	--    2nd DW: destination address (32bit)
	--    3rd DW: source address (32bit)
	--    4th DW: byte count(16bit: 1-64k 31:16), packet-type (4bit 15:12), status (4bit 11:8), 
	--            first byte enable (4bit 7:4)
	--       Packet type: 0000=wr_req, 0001=rd_request, 0010=rd_completion, 0011=rd_forwarding request, 
	--          0100=rd_forw_compl, 0101=wr_forwarding, others: RFU
	--       Status: 0000=succesful_transaction, 0001=no_further_hop, 0010=unknown_error
	-- The user must write the local address field last, since that register/FIFO triggers the transfer.


	 --packet-protocol statemachine:
    process (trn_reset_n, user_clk_i, packet_state, 
				op2p_just_received_a_new_packet, packet_datacount, op2p_local_id, RX_FC_NB_latched,
				bram_rxpacket_readdata,  bram_txpacket_writeaddress, bram_rxpacket_readaddress,
				packet_state_copy,  rxpacket_decodedaddress, bram_rxpacket_firstdata_address,
				rxpacket_header_dw1, rxpacket_header_dw2, rxpacket_header_dw3, rxpacket_header_dw4,
				bit10, rxpacket_firstdw_be, wb_transaction_complete, packet_payloadsize_dwords_p4,
				packet_payloadsize_dwords, op2p_mem_wb_data_i_latched, cfg_completer_id,
				rxpacket_requesterid, CHANNEL_UP, change_flag_packetstm) 
    begin
    if (trn_reset_n='0') then 
		start_read_wb0 <= '0';
		start_write_wb0 <= '0';
		op2p_wb_data_o_feed	 <= (others => '0');
		op2p_wb_addr_o_feed <= (others => '0');
		op2p_wb_sel_o_feed  <= (others => '0');
		op2p_there_is_a_new_packet_to_transmit  <= '0';
		rxpacket_decodedaddress<= (others => '0');
		packet_payloadsize_dwords <= (others => '0');
		rxpacket_firstdw_be <= (others => '0');
		rxpacket_lastdw_be <= (others => '0');
		rxpacket_requesterid <= (others => '0');
		packet_state <= (others => '0');
		packet_state_copy  <= (others => '0');
		bram_txpacket_we <= "0";
		bram_txpacket_writeaddress    <= (others => '0');
		bram_txpacket_writedata     <= (others => '0');
		bram_rxpacket_readaddress   <= (others => '0');
		bram_rxpacket_firstdata_address   <= (others => '0');
		rxpacket_header_dw1   <= (others => '0');
		rxpacket_header_dw2   <= (others => '0');
		rxpacket_header_dw3   <= (others => '0');
		rxpacket_header_dw4   <= "00000000000000001111000000000000";
		packetstm_counter <=  (others => '0');
		fbm_nextraddress_req <= '0';
		destination_address <=  (others => '0');
		source_id <=  (others => '0');
		destination_id <=  (others => '0');
		source_address <=  (others => '0');
		byte_count <=  (others => '0');
		packet_datacount <= (others => '0');
		packetstm_isin_idle <= '1';
		op2p_wr_sourceaddress_regrd_en  <=  '0'; 
		op2p_wr_destinationaddress_regrd_en  <=  '0'; 
		op2p_wr_sourceid_regrd_en  <=  '0'; 
		op2p_wr_destinationid_regrd_en  <=  '0';
		op2p_wr_bytecount_regrd_en  <=  '0';
		op2p_rdreq_localaddress_regrd_en  <=  '0'; 
		op2p_rdreq_destinationaddress_regrd_en  <=  '0'; 
		op2p_rdreq_sourceid_regrd_en  <=  '0'; 
		op2p_rdreq_destinationid_regrd_en  <=  '0';
		op2p_rdreq_bytecount_regrd_en  <=  '0';
		change_flag_packetstm <= '0';
		txstm_reenable_fc <= '0';
		txstm_haltdata_fc2 <= '0';
		op2p_event_pulse <= '0';
		op2p_forwreq_pointer_regwr_en  <=  '0';
		op2p_forwreq_pointer_regdin <= (OTHERS => '0');
		link_errcnt_latchedinidle <= (OTHERS => '0');
		it_is_a_retransmit <= '0';
		rx_detect_ff_clear  <= '0';
		
    else
      if (user_clk_i'event and user_clk_i = '1') then
                case ( packet_state ) is

                --********** IDLE STATE  **********
                when "00000000" =>   --state 0   
						  --request from link partner: (write, read req, forw req, forw-compl)					 
						  if ( rx_detected = '1') then
						    packet_state <= "00000001"; --to packet decoding state
							 packetstm_isin_idle <= '0';
						  --request from local host: (write req, read req, forw compl, forw req)
						  elsif (op2p_wr_anybuffers_empty = '0' and CHANNEL_UP='1' and fc_halted_bylinkpartner='0') then
						    packet_state <= "00010000"; --to outgoing write state
							 packetstm_isin_idle <= '0';
							 txstm_haltdata_fc2 <= '1'; --stop data coming in
						  elsif (op2p_rdreq_anybuffers_empty = '0' and CHANNEL_UP='1' and fc_halted_bylinkpartner='0') then
						    packet_state <= "01000000"; --to outgoing RDREQ state
							 packetstm_isin_idle <= '0';
						  else
						    packetstm_isin_idle <= '1';
							 txstm_haltdata_fc2 <= '0'; --let/reenable data coming in
						  end if;
						  --general preparation:				
						  start_write_wb0 <= '0';
						  start_read_wb0 <= '0';
						  packet_state_copy <= packet_state;
							bram_txpacket_we <= "0";
							bram_txpacket_writeaddress   <= (others => '0');
							bram_txpacket_writedata     <= (others => '0');
							bram_rxpacket_readaddress    <= (others => '0');
							packet_datacount <= (others => '0');
							bram_rxpacket_firstdata_address   <= (others => '0');
							packetstm_counter <=  (others => '0');
							rxpacket_header_dw4   <= "00000000000000001111000000000000"; --this is to prevent false decode
							 op2p_wb_data_o_feed	 <= (others => '0');
							op2p_wb_addr_o_feed <= (others => '0');
							op2p_wb_sel_o_feed  <= (others => '0');
							op2p_there_is_a_new_packet_to_transmit  <= '0';
							rxpacket_decodedaddress<= (others => '0');
							--packet_payloadsize_dwords <= (others => '0');
							rxpacket_firstdw_be <= (others => '0');
							rxpacket_lastdw_be <= (others => '0');
							rxpacket_requesterid <= (others => '0');
							rxpacket_header_dw1   <= (others => '0');
							rxpacket_header_dw2   <= (others => '0');
							rxpacket_header_dw3   <= (others => '0');
							fbm_nextraddress_req <= '0';
							destination_address <=  (others => '0');
							source_id <=  (others => '0');
							destination_id <=  (others => '0');
							source_address <=  (others => '0');
							byte_count <=  (others => '0');
							change_flag_packetstm <= '0';
							txstm_reenable_fc <= '0';
							op2p_event_pulse <= '0';
							op2p_forwreq_pointer_regwr_en  <=  '0';
							op2p_forwreq_pointer_regdin <= (OTHERS => '0');
							link_errcnt_latchedinidle <= link_error_count_reg;
							rx_detect_ff_clear <= '0';
							
						  
                --********** packet ARRIVED STATE **********
					 --initiated by link partner
					 --read packet out of EP, decode and decide,
					 --latch address/sel/wr_data
                when "00000001" =>   --state 1
						  packetstm_counter <=  packetstm_counter + 1;
						  packet_state_copy <= packet_state;
						  --set buffer read address:
						  if (packetstm_counter = "00000111") then
						    bram_rxpacket_readaddress <= "000000101"; --point to data
						  elsif (packetstm_counter = "00000110") then
						    bram_rxpacket_readaddress <= "000000101"; --point to data
						  else
						    bram_rxpacket_readaddress <= bram_rxpacket_readaddress + 1;
						  end if;
						  --latch the header:
						  if (packetstm_counter = "000000010") then
						    rxpacket_header_dw1 <= bram_rxpacket_readdata;
							 rx_detect_ff_clear <= '1';
						  elsif (packetstm_counter = "000000011") then
						    rxpacket_header_dw2 <= bram_rxpacket_readdata;
						  elsif (packetstm_counter = "000000100") then
						    rxpacket_header_dw3 <= bram_rxpacket_readdata;
							 rx_detect_ff_clear <= '0';
						  elsif (packetstm_counter = "000000101") then
						    rxpacket_header_dw4 <= bram_rxpacket_readdata;
						  end if;
						  --decode some parameters:
						  --(works at packetstm_counter = "00000110")
						  packet_payloadsize_dwords (7 downto 0) <= rxpacket_header_dw4(25 downto 18); --from bytecount to dword count
						  rxpacket_status <= rxpacket_header_dw4(11 downto 8);
						  rxpacket_firstdw_be <= rxpacket_header_dw4(7 downto 4);
						  rxpacket_requesterid <= rxpacket_header_dw1(31 downto 16); --same as source id, but only for this type of trn
						  rxpacket_sourceid <= rxpacket_header_dw1(31 downto 16);
						  rxpacket_destinationid <= rxpacket_header_dw1(15 downto 0);
						  rxpacket_destinationaddress <= rxpacket_header_dw2(31 downto 0);
						  rxpacket_sourceaddress <= rxpacket_header_dw3(31 downto 0);
						  bram_rxpacket_firstdata_address (8 downto 0)   <= "000000100"; --addr in packet buffer
						  rxpacket_decodedaddress <= rxpacket_destinationaddress;
						  --decide based on header: 
						  -- Packet type: 0000=wr_req, 0001=rd_request, 0010=rd_completion, 0011=forwarding request, 
						  --0100=forw_compl, others: RFU
						  rxpacket_type <= rxpacket_header_dw4(15 downto 12);
						  if (packetstm_counter = "00000111") then --when the parameters are already stored
								--read request arrived. (respond with data)
								if (link_error_count_reg /= link_errcnt_latchedinidle) then 
									--request data retransmit, since error was detected in data stream
									packet_state <= "11110101"; --to retransmit request
								elsif (rxpacket_type="0001" and idmatch='1') then 
									packet_state <= "00000011"; --3
									op2p_wb_addr_o_feed(31 downto 2) <= rxpacket_destinationaddress(31 downto 2);
									op2p_wb_addr_o_feed(1 downto 0) <= bit10(1 downto 0);
									op2p_wb_sel_o_feed  <= rxpacket_firstdw_be;
									bram_txpacket_writeaddress <= "000000011"; --3, point before the first data dw
								--read completion arrived. (put data into memory, same as write arrived state)
								elsif (rxpacket_type="0010" and idmatch='1') then 
									packet_state <= "00000010"; --2
									op2p_wb_addr_o_feed(31 downto 2) <= rxpacket_destinationaddress(31 downto 2);
									op2p_wb_addr_o_feed(1 downto 0) <= bit10(1 downto 0);
									op2p_wb_sel_o_feed  <= rxpacket_firstdw_be;
								--write with data arrived
								elsif (rxpacket_type="0000" and idmatch='1') then 
									packet_state <= "00000010"; --2
									op2p_wb_addr_o_feed(31 downto 2) <= rxpacket_destinationaddress(31 downto 2);
									op2p_wb_addr_o_feed(1 downto 0) <= bit10(1 downto 0);
									op2p_wb_sel_o_feed  <= rxpacket_firstdw_be;
								--rd forwarding request came in (put the whole packet into the memory, except at ID match)
								elsif (rxpacket_type="0001" and idmatch='0') then 
									packet_state <= "01110000";   --state 112
								--rd forwarding completion came in (someone was reading someone, this is the read data)
								elsif (rxpacket_type="0010" and idmatch='0') then 
									packet_state <= "01110000";   --state 112
								--wr forwarding req came in (someone is writing someone with data)
								elsif (rxpacket_type="0000" and idmatch='0') then 
									packet_state <= "01110000";   --state 112
								--Link partner is requesting data retransmit.
								elsif (rxpacket_type="1010") then
								  packet_state <= "11110111";   --state x
								--just wait until this gets a real value
								elsif (rxpacket_type="1111") then 
								 --it also means that the logic will hang here forever if the type=1111.
									packet_state <= "00000001"; --1/decode, stay in this state
								--unsupported request
								else 
								 packet_state <= "00000101";
								 bram_txpacket_writeaddress <= "111111111";
								end if;
						  end if;



                --********** WRITE or other DATA arrived STATE **********
					 --initiated by link partner
					 --This will initiate WB write(s) (1...N DWORD accesses).
					 --This state serves several transaction types:
					 --write arrived, read completion arrived, forwarding packet (req/compl/posted) 
					 --arrived (after pointer manipulation).
                when "00000010" =>   --state 2
						op2p_wb_data_o_feed <= bram_rxpacket_readdata;
						packet_state_copy <= packet_state;
						if (packet_state_copy = packet_state) then 
						  start_write_wb0 <= '0';
						else --generate just one pulse, at the first clk cycle in this state
						  start_write_wb0 <= '1';
						end if;
						if (wb_transaction_complete='1') then  --one DW transfer completed
							if (packet_payloadsize_dwords = packet_datacount + 1)then  --all data completed
							  packet_state <= "00010101"; --to idle (after some detour)
							  if (link_error_count_reg = link_errcnt_latchedinidle ) then
							    txstm_reenable_fc <= '1';
							    op2p_event_pulse <= '1'; --notify host
							  end if;
							else
							  packet_state <= "00010100"; --restart wb transaction with new data
							  bram_rxpacket_readaddress <= bram_rxpacket_readaddress +1;
							  packet_datacount <= packet_datacount +1;
							end if;
						end if;
                --* Write restart state *
                when "00010100" =>   --state 20
 						packet_state <= "00000010";
						packet_state_copy <= packet_state;
						op2p_wb_addr_o_feed(31 downto 2) <= op2p_wb_addr_o_feed(31 downto 2) + 1;
						op2p_wb_addr_o_feed(1 downto 0) <= "00";
						op2p_wb_sel_o_feed <= "1111";
                --* Write finished state *
                when "00010101" =>   --state 21
						packet_state <= "00000000"; --to idle
						if (link_error_count_reg = link_errcnt_latchedinidle ) then
						    --fine, go back to idle
						    packet_state <= "00000000"; --to idle
							 it_is_a_retransmit <= '0'; --next arriving data will be marked as new.
							 -- INFO TO THE LOCAL HOST ABOUT ARRIVED FORWARDING PACKETS 
							 --if the previous wishbone write was a forwarding packet (no ID match), then store pointer
							 if (idmatch='0') then 
								op2p_forwreq_pointer_regwr_en <=  '1';
							 else
								op2p_forwreq_pointer_regwr_en <=  '0';
							 end if;
							 op2p_forwreq_pointer_regdin <= rxpacket_decodedaddress;
						else
						  --request data retransmit, since error was detected in data streem
						  packet_state <= "11110101"; --to retransmit request
						end if;
						packet_state_copy <= packet_state;
						txstm_reenable_fc <= '0';
						op2p_event_pulse <= '0'; 

				 

				 
                --********** READ request arrived STATE **********
					 --requested by link partner
					 --This will initiate WB read(s), then go to completion state to send data to link partner
                when "00000011" =>   --state 3
						op2p_wb_sel_o_feed  <= rxpacket_firstdw_be;
						packet_state_copy <= packet_state;
						it_is_a_retransmit <= '0'; --next arriving packet will be marked as new.
						if (packet_state_copy = packet_state) then 
						  start_read_wb0 <= '0';
						else --generate just one pulse
						  start_read_wb0 <= '1';
						end if;
						if (wb_transaction_complete='1') then 
							bram_txpacket_writedata <= op2p_mem_wb_data_i_latched; --upd val
							bram_txpacket_we <= "1";
							bram_txpacket_writeaddress <= bram_txpacket_writeaddress +1;
							packet_datacount <= packet_datacount +1;
							if (packet_payloadsize_dwords = packet_datacount +1)then 
							  packet_state <= "01111110"; --read completion
							else
							  packet_state <= "00011110"; --one more wb read
							end if;
						else
						  bram_txpacket_we <= "0";
						end if;
                --* read restart STATE  *
                when "00011110" =>   --state 30
						packet_state <= "00000011";
						bram_txpacket_we <= "0";
						packet_state_copy <= packet_state;
						op2p_wb_addr_o_feed(31 downto 2) <= op2p_wb_addr_o_feed(31 downto 2) + 1;
						op2p_wb_addr_o_feed(1 downto 0) <= "00";
						op2p_wb_sel_o_feed <= "1111";
                --intermediate state before completion (to ensure data latch at address-4)
					 when "01111110" =>   --state 126
						packet_state <= "00000100";
						packet_state_copy <= packet_state;
						bram_txpacket_we <= "0";
						bram_txpacket_writeaddress  <=  "111111111";	
						
                --********** READ COMPLETION transmission  STATE **********
					 --requested by link partner (send response with data to link partner)
					 --assemble the tx packet and initiate the transmit
					 --tx packet block ram: bram_txpacket_we, bram_txpacket_writeaddress, bram_txpacket_writedata,
					 --The completion swaps the source/destination ID/address fields!!!!!
                when "00000100" =>   --state 4
                    packet_state_copy <= packet_state;
						  if (bram_txpacket_writeaddress="111111111") then
								bram_txpacket_we <= "1";
								bram_txpacket_writeaddress <= bram_txpacket_writeaddress +1;
								bram_txpacket_writedata (31 downto 16) <= rxpacket_header_dw1(15 downto 0); --source ID** --pre-write header-DW1:
								bram_txpacket_writedata (15 downto 0) <= rxpacket_header_dw1(31 downto 16); --destination ID**
						  elsif (bram_txpacket_writeaddress="000000000") then --pre-write header-DW2:
						    bram_txpacket_we <= "1";
							 bram_txpacket_writeaddress <= bram_txpacket_writeaddress +1;
							  bram_txpacket_writedata (31 downto 0) <= rxpacket_header_dw3; --destination address**
						  elsif (bram_txpacket_writeaddress="000000001") then --pre-write header-DW3:
						    bram_txpacket_we <= "1";
							 bram_txpacket_writeaddress <= bram_txpacket_writeaddress +1;
							  bram_txpacket_writedata (31 downto 0) <= rxpacket_header_dw2;--source address**
						  elsif (bram_txpacket_writeaddress="000000010") then --pre-write header-DW4:
						    bram_txpacket_we <= "1";
							 bram_txpacket_writeaddress <= bram_txpacket_writeaddress +1;
							 --byte count: **
							 --bram_txpacket_writedata (31 downto 16) <= rxpacket_header_dw4 (31 downto 16); 
							 bram_txpacket_writedata (31 downto 26) <= "000000";
							 bram_txpacket_writedata (25 downto 18) <= packet_payloadsize_dwords (7 downto 0);
							 bram_txpacket_writedata (17 downto 16) <= "00";
							  --packet type: Packet type: 0000=wr_req, 0001=rd_request, 0010=rd_completion, 0011=forwarding request, 0100=forw_compl, others: RFU
								  if (rxpacket_type = "0011") then --read forwarding req
									 bram_txpacket_writedata (15 downto 12) <= "0100";
								  else --normal read req
									 bram_txpacket_writedata (15 downto 12) <= "0010";
								  end if;
							  bram_txpacket_writedata (11 downto 8) <= "0000"; --status** : Status: 0000=succesful_transaction, 0001=no_further_hop, 
							    --0010=unknown_error
							  bram_txpacket_writedata (7 downto 4) <= rxpacket_firstdw_be (3 downto 0); --first byte enable**
							  bram_txpacket_writedata (3 downto 0) <= "0000"; --RFU
						  else --data dwords 
						    bram_txpacket_we <= "0";
							 bram_txpacket_writeaddress <=  "111111110";
						  end if;
						  --one pulse to start the ep-if statemachine, upon arriving to this state
							--if (packet_state_copy = packet_state) then 
							--  op2p_there_is_a_new_packet_to_transmit  <= '0';
							--else 
							--  op2p_there_is_a_new_packet_to_transmit  <= '1';
							--end if;
							--back to idle when the ep-if tx is finished: (wait to avoid overwrite)
							if (op2p_packet_tx_complete='1') then 
								packet_state <= "00000000";
								txstm_reenable_fc <= '1';
								op2p_there_is_a_new_packet_to_transmit  <= '0';
							else
							   op2p_there_is_a_new_packet_to_transmit  <= '1';
							end if;



                --********** forwarding PACKET arrived STATE **********
					 --initiated by link partner.
					 --If a packet's destination ID is not a match, then store the packet with header for forwarding.
					 --Allocate memory buffer, then Store the whole packet in DRAM.
					 --if the op2p_forwreq_pointer_reg is full, it automatically requests a FC=halt in the TX state machine.
                when "01110000" =>   --state 112
							packetstm_counter <=  (others => '0');
							packet_state_copy <= packet_state;
							packet_state <= "01110001";
					 when "01110001" =>   --state 113
						  packet_state_copy <= packet_state;
						  bram_rxpacket_readaddress <=  "000000001"; --point to header DW1
						  --this is needed to provide an extra clock for the packet RD data to stabilize before feeding it to WB:
						  if (forw_packetaddr_allocated ='1') then
						    change_flag_packetstm <= '1';
						  end if;
						  if (change_flag_packetstm='1' or it_is_a_retransmit='1') then --now, the mem address should be available, and the BRAM data stable.
						    packetstm_counter <=  (others => '0');
							 rxpacket_decodedaddress <= fbm_nextraddress;
							 if (rxpacket_type="0001" and idmatch='0') then --forwarding read req: no data, just 4DW header
							   packet_payloadsize_dwords <= "00000000000000000000000000000100";
							 else
							   packet_payloadsize_dwords <= packet_payloadsize_dwords_p4; --to copy the header as well
							 end if;
							 fbm_nextraddress_req <= '0';
								op2p_wb_addr_o_feed(31 downto 2) <= fbm_nextraddress(31 downto 2);
								op2p_wb_addr_o_feed(1 downto 0) <= bit10(1 downto 0);
								op2p_wb_sel_o_feed  <= rxpacket_firstdw_be;
								op2p_wb_data_o_feed <= bram_rxpacket_readdata;
								bram_rxpacket_firstdata_address (8 downto 0)   <= "000000001"; --addr in packet buffer
							 packet_state <= "00000010"; --2, go to write state with tricked parameters   ***This state finishes here***
						  elsif (packetstm_counter = "00000010") then --when 2, reset the request pulse
						    fbm_nextraddress_req <= '0';
							 packetstm_counter <=  packetstm_counter; --stop counting
						  else --when counter is 0 or 1, assert request              ***This state starts here***
								if (it_is_a_retransmit='1') then
								  fbm_nextraddress_req <= '0';
								else
								  fbm_nextraddress_req <= '1';
								end if;
							   packetstm_counter <=  packetstm_counter +1;
						  end if;



                --********** UNSUPPORTED REQUEST STATE **********
					 --completion response with status=0010 and no data.
                when "00000101" =>   --state 5
                    packet_state_copy <= packet_state;
						  packet_payloadsize_dwords <=  (OTHERS => '0');
						  bram_txpacket_writeaddress <= bram_txpacket_writeaddress +1;
						  if (bram_txpacket_writeaddress="111111111") then --header 1.dw
						    bram_txpacket_we <= "1";
							  bram_txpacket_writedata (31 downto 16) <= rxpacket_header_dw1(15 downto 0); --source ID**
							  bram_txpacket_writedata (15 downto 0) <= rxpacket_header_dw1(31 downto 16); --destination ID**
						  elsif (bram_txpacket_writeaddress="000000000") then --header 2.dw
						    bram_txpacket_we <= "1";
							  bram_txpacket_writedata (31 downto 0) <= rxpacket_header_dw3; --destination address**
						  elsif (bram_txpacket_writeaddress="000000001") then --header 3.dw
						    bram_txpacket_we <= "1";
							  bram_txpacket_writedata (31 downto 0) <= rxpacket_header_dw2;--source address**
						  elsif (bram_txpacket_writeaddress="000000010") then --header 4.dw
						    bram_txpacket_we <= "1";
						     bram_txpacket_writedata (31 downto 16) <= rxpacket_header_dw4 (31 downto 16); --byte count**
							  --packet type: Packet type: 0000=wr_req, 0001=rd_request, 0010=rd_completion, 0011=forwarding request, 0100=forw_compl, others: RFU
								  if (rxpacket_type = "0011") then --read forwarding req
									 bram_txpacket_writedata (15 downto 12) <= "0100";
								  else --normal read req
									 bram_txpacket_writedata (15 downto 12) <= "0010";
								  end if;
							  bram_txpacket_writedata (11 downto 8) <= "0010"; --status** : Status: 0000=succesful_transaction, 0001=no_further_hop, 
							    --0010=unknown_error
							  bram_txpacket_writedata (7 downto 4) <= rxpacket_header_dw4 (7 downto 4); --first byte enable**
							  bram_txpacket_writedata (3 downto 0) <= "0000"; --RFU
						  else --data dwords 
						    bram_txpacket_we <= "0";
						  end if;
						  --one pulse to start the ep-if statemachine, upon arriving to this state
							--if (packet_state_copy = packet_state) then 
							--  op2p_there_is_a_new_packet_to_transmit  <= '0';
							--else 
							--  op2p_there_is_a_new_packet_to_transmit  <= '1';
							--end if;
							--back to idle when the ep-if tx is finished: (wait to avoid overwrite)
							if (op2p_packet_tx_complete='1') then 
								packet_state <= "00000000";
								txstm_reenable_fc <= '1';
								op2p_there_is_a_new_packet_to_transmit  <= '0';
							else
							   op2p_there_is_a_new_packet_to_transmit  <= '1';								
							end if;



                --********** RETRANSMIT REQUEST STATE **********
					 --error was detected in incoming packet, so request retransmit from link 
					 --partner, with status=0010 and no data.
                when "11110101" =>   --state 245
                    packet_state_copy <= packet_state;
						  packet_payloadsize_dwords <=  (OTHERS => '0');
						  bram_txpacket_writeaddress <= bram_txpacket_writeaddress +1;
						  if (bram_txpacket_writeaddress="111111111") then --header 1.dw
						    bram_txpacket_we <= "1";
							  bram_txpacket_writedata (31 downto 16) <= op2p_local_id_reclocked2(15 downto 0); --source ID**
							  bram_txpacket_writedata (15 downto 0) <= "0000000000000000"; --destination ID (link partner)**
						  elsif (bram_txpacket_writeaddress="000000000") then --header 2.dw
						    bram_txpacket_we <= "1";
							  bram_txpacket_writedata (31 downto 0) <= rxpacket_header_dw3; --destination address**
						  elsif (bram_txpacket_writeaddress="000000001") then --header 3.dw
						    bram_txpacket_we <= "1";
							  bram_txpacket_writedata (31 downto 0) <= rxpacket_header_dw2;--source address**
						  elsif (bram_txpacket_writeaddress="000000010") then --header 4.dw
						    bram_txpacket_we <= "1";
						     bram_txpacket_writedata (31 downto 16) <= rxpacket_header_dw4 (31 downto 16); --byte count**
							  --packet type:  1010=retransmit_req, 
							  bram_txpacket_writedata (15 downto 12) <= "1010";
							  bram_txpacket_writedata (11 downto 8) <= "0010"; --status** : 0010=unknown_error
							  bram_txpacket_writedata (7 downto 4) <= rxpacket_header_dw4 (7 downto 4); --first byte enable**
							  bram_txpacket_writedata (3 downto 0) <= "0000"; --RFU
						  else --data dwords 
						    bram_txpacket_we <= "0";
						  end if;
						  --one pulse to start the ep-if statemachine, upon arriving to this state
							--if (packet_state_copy = packet_state) then 
							--  op2p_there_is_a_new_packet_to_transmit  <= '0';
							--else 
							--  op2p_there_is_a_new_packet_to_transmit  <= '1';
							--end if;
							--back to idle when the ep-if tx is finished: (wait to avoid overwrite)
							if (op2p_packet_tx_complete='1') then 
								packet_state <= "00000000";
								txstm_reenable_fc <= '1';
								it_is_a_retransmit <='1';
								op2p_there_is_a_new_packet_to_transmit  <= '0';
							else
							   op2p_there_is_a_new_packet_to_transmit  <= '1';								
							end if;


                --********** RETRANSMIT STATE **********
					 --send last packet out again, since link partner has requested it.
                when "11110111" =>   --state 247
                    packet_state_copy <= packet_state;
						  --one pulse to start the ep-if statemachine, upon arriving to this state
							--if (packet_state_copy = packet_state) then 
							--  op2p_there_is_a_new_packet_to_transmit  <= '0';
							--else 
							--  op2p_there_is_a_new_packet_to_transmit  <= '1';
							--end if;
							--back to idle when the ep-if tx is finished: (wait to avoid overwrite)
							if (op2p_packet_tx_complete='1') then 
								packet_state <= "00000000";
								txstm_reenable_fc <= '1';
								op2p_there_is_a_new_packet_to_transmit  <= '0';
							else
							   op2p_there_is_a_new_packet_to_transmit  <= '1';								
							end if;						

                --********** Outgoing write STATE **********
                --initiated by local host
                --parameter fetch substate
					 when "00010000" =>   --state x
						packetstm_counter <=  packetstm_counter +1;
						change_flag_packetstm <= '0';
						txstm_haltdata_fc2 <= '0';
						if (packetstm_counter = "00000000") then
							packetstm_counter <=  packetstm_counter +1;
							op2p_wr_sourceaddress_regrd_en  <=  '1'; 
							op2p_wr_destinationaddress_regrd_en  <=  '1'; 
							op2p_wr_sourceid_regrd_en  <=  '1'; 
							op2p_wr_destinationid_regrd_en  <=  '1';
							op2p_wr_bytecount_regrd_en  <=  '1';
						elsif(packetstm_counter = "00000001") then --one more clock until data is stable at the output
						   packetstm_counter <=  packetstm_counter +1;
							op2p_wr_sourceaddress_regrd_en  <=  '0'; 
							op2p_wr_destinationaddress_regrd_en  <=  '0'; 
							op2p_wr_sourceid_regrd_en  <=  '0'; 
							op2p_wr_destinationid_regrd_en  <=  '0';
							op2p_wr_bytecount_regrd_en  <=  '0';
						else --last clock,
							packetstm_counter <=  (OTHERS => '0');
							packet_state <= "00010001"; --to wishbone tr state *****
							source_address <= op2p_wr_sourceaddress_regdout;
							destination_address <= op2p_wr_destinationaddress_regdout;
							source_id <= op2p_wr_sourceid_regdout(15 downto 0);
							destination_id <= op2p_wr_destinationid_regdout(15 downto 0);
							byte_count(31 downto 2) <= op2p_wr_bytecount_regdout(31 downto 2);
							byte_count(1 downto 0) <= "00"; --ignore unaligned data
							packet_payloadsize_dwords(29 downto 0) <= op2p_wr_bytecount_regdout(31 downto 2);
							packet_payloadsize_dwords(31 downto 30) <= "00";
							--prepare wishbone command:
							op2p_wb_addr_o_feed(31 downto 2) <= op2p_wr_sourceaddress_regdout(31 downto 2) ; 
							op2p_wb_addr_o_feed(1 downto 0) <= bit10(1 downto 0);
							op2p_wb_sel_o_feed  <= "1111";
							bram_txpacket_writeaddress <= "000000011"; --start with (before) data field
						end if;
					 --wishbone transactions substate
					 when "00010001" =>   --state x 
						packet_state_copy <= packet_state;
						if (change_flag_packetstm = '1') then 
						  start_read_wb0 <= '0';
						else --generate just one pulse
						  start_read_wb0 <= '1';
						end if;
						if (wb_transaction_complete='1') then
							bram_txpacket_writedata <= op2p_mem_wb_data_i_latched; --upd val
							bram_txpacket_we <= "1";
							packet_datacount <= packet_datacount + 4;
							change_flag_packetstm <= '0';
							bram_txpacket_writeaddress <= bram_txpacket_writeaddress +1;
							if (byte_count = packet_datacount + 4 )then --no more data (pac_dat_c starts at 0, byte_c is min 4)
							  packet_state <= "00010011"; --completion
							else
							  packet_state <= "00010010"; --one more wb read (intermed wait state)
								op2p_wb_addr_o_feed(31 downto 2) <= op2p_wb_addr_o_feed(31 downto 2) + 1; --increm by 4
								op2p_wb_addr_o_feed(1 downto 0) <= "00";
							end if;
						else
						  change_flag_packetstm <= '1';
						  bram_txpacket_we <= "0";
						end if;
                --* intermediate wait STATE  *
                when "00010010" =>   --state 30
						packet_state <= "00010001";
						bram_txpacket_we <= "0";
						change_flag_packetstm <= '0';
					 --packet header assembling substate for outgoing write
					 when "00010011" =>   --state x
                    packet_state_copy <= packet_state;
						  change_flag_packetstm <= '1';
						  if    (change_flag_packetstm='0') then --header 1.dw in next clock cycle
						    bram_txpacket_we <= "1";
							 bram_txpacket_writeaddress <= "000000000"; --set address at dw-zero
							  bram_txpacket_writedata (31 downto 16) <= source_id; --source ID**
							  bram_txpacket_writedata (15 downto 0) <= destination_id; --destination ID**
						  elsif (bram_txpacket_writeaddress="000000000") then --header 2.dw in next clock cycle
						    bram_txpacket_we <= "1";
							 bram_txpacket_writeaddress <= bram_txpacket_writeaddress +1;
							  bram_txpacket_writedata (31 downto 0) <= destination_address; --destination address**
						  elsif (bram_txpacket_writeaddress="000000001") then --header 3.dw in next clock cycle
						    bram_txpacket_we <= "1";
							 bram_txpacket_writeaddress <= bram_txpacket_writeaddress +1;
							  bram_txpacket_writedata (31 downto 0) <= source_address;--source address**
						  elsif (bram_txpacket_writeaddress="000000010") then --header 4.dw in next clock cycle
						    bram_txpacket_we <= "1";
							 bram_txpacket_writeaddress <= bram_txpacket_writeaddress +1;
						     bram_txpacket_writedata (31 downto 16) <= byte_count(15 downto 0); --byte count**
							  bram_txpacket_writedata (15 downto 12) <= "0000"; --packet type** : Packet type: 0000=wr_req, 
							    --0001=rd_request, 0010=rd_completion, 0011=forwarding request, 0100=forw_compl, others: RFU
							  bram_txpacket_writedata (11 downto 8) <= "0000"; --status** : Status: 0000=succesful_transaction, 
							    --0001=no_further_hop, 0010=unknown_error
							  bram_txpacket_writedata (7 downto 4) <= "1111"; --first byte enable**
							  bram_txpacket_writedata (3 downto 0) <= "0000"; --RFU
						  else --data dwords 
						    bram_txpacket_we <= "0";
						  end if;
						  --one pulse to start the ep-if statemachine, upon arriving to this state
							--if (packet_state_copy = packet_state) then 
							--  op2p_there_is_a_new_packet_to_transmit  <= '0';
							--else 
							--  op2p_there_is_a_new_packet_to_transmit  <= '1';
							--end if;
							--back to idle when the ep-if tx is finished: (wait to avoid overwrite)
							if (op2p_packet_tx_complete='1') then 
								packet_state <= "00000000";
								txstm_reenable_fc <= '1';
								op2p_event_pulse <= '1'; --notify host
								op2p_there_is_a_new_packet_to_transmit  <= '0';
							else
							   op2p_there_is_a_new_packet_to_transmit  <= '1';								
							end if;



                --********** Outgoing RD REQ STATE **********
                --initiated by local host
                when "01000000" =>   --state x
						packetstm_counter <=  packetstm_counter +1;
						txstm_haltdata_fc2 <= '0';
						if (packetstm_counter = "00000000") then
							packetstm_counter <=  packetstm_counter +1;
							op2p_rdreq_localaddress_regrd_en  <=  '1'; 
							op2p_rdreq_destinationaddress_regrd_en  <=  '1'; 
							op2p_rdreq_sourceid_regrd_en  <=  '1'; 
							op2p_rdreq_destinationid_regrd_en  <=  '1';
							op2p_rdreq_bytecount_regrd_en  <=  '1';
						elsif(packetstm_counter = "00000001") then --one more clock until data is stable at the output
						   packetstm_counter <=  packetstm_counter +1;
							op2p_rdreq_localaddress_regrd_en  <=  '0'; 
							op2p_rdreq_destinationaddress_regrd_en  <=  '0'; 
							op2p_rdreq_sourceid_regrd_en  <=  '0'; 
							op2p_rdreq_destinationid_regrd_en  <=  '0';
							op2p_rdreq_bytecount_regrd_en  <=  '0';
						else
							packetstm_counter <=  (OTHERS => '0');
							packet_state <= "01000001"; --to next state
							source_address <= op2p_rdreq_localaddress_regdout;
							destination_address <= op2p_rdreq_destinationaddress_regdout;
							source_id <= op2p_rdreq_sourceid_regdout(15 downto 0);
							destination_id <= op2p_rdreq_destinationid_regdout(15 downto 0);
							byte_count(31 downto 2) <= op2p_rdreq_bytecount_regdout(31 downto 2);
							byte_count(1 downto 0) <= "00"; --ignore unaligned data
							 packet_payloadsize_dwords(29 downto 0) <= op2p_rdreq_bytecount_regdout(31 downto 2);
							 packet_payloadsize_dwords(31 downto 30) <= "00";
							 bram_txpacket_writeaddress <= "111111111";
						end if;
					 --packet header assembling substate for outgoing RD REQ 
					 when "01000001" =>   --state x
                    packet_state_copy <= packet_state;
						  bram_txpacket_writeaddress <= bram_txpacket_writeaddress +1;
						  if (bram_txpacket_writeaddress="111111111") then --header 1.dw
						    bram_txpacket_we <= "1";
							  bram_txpacket_writedata (31 downto 16) <= source_id; --source ID**
							  bram_txpacket_writedata (15 downto 0) <= destination_id; --destination ID**
						  elsif (bram_txpacket_writeaddress="000000000") then --header 2.dw
						    bram_txpacket_we <= "1";
							  bram_txpacket_writedata (31 downto 0) <= destination_address; --destination address**
						  elsif (bram_txpacket_writeaddress="000000001") then --header 3.dw
						    bram_txpacket_we <= "1";
							  bram_txpacket_writedata (31 downto 0) <= source_address;--source address** --local address for rd req
						  elsif (bram_txpacket_writeaddress="000000010") then --header 4.dw
						    bram_txpacket_we <= "1";
						     bram_txpacket_writedata (31 downto 16) <= byte_count(15 downto 0); --byte count**
							  bram_txpacket_writedata (15 downto 12) <= "0001"; --packet type** : Packet type: 0000=wr_req, 
							    --0001=rd_request, 0010=rd_completion, 0011=forwarding request, 0100=forw_compl, others: RFU
							  bram_txpacket_writedata (11 downto 8) <= "0000"; --status** : Status: 0000=succesful_transaction, 
							    --0001=no_further_hop, 0010=unknown_error
							  bram_txpacket_writedata (7 downto 4) <= "1111"; --first byte enable**
							  bram_txpacket_writedata (3 downto 0) <= "0000"; --RFU
						  else --data dwords 
						    bram_txpacket_we <= "0";
						  end if;
						  --one pulse to start the ep-if statemachine, upon arriving to this state
							--if (packet_state_copy = packet_state) then 
							--  op2p_there_is_a_new_packet_to_transmit  <= '0';
							--else 
							--  op2p_there_is_a_new_packet_to_transmit  <= '1';
							--end if;
							--back to idle when the ep-if tx is finished: (wait to avoid overwrite)
							if (op2p_packet_tx_complete='1') then 
								packet_state <= "00000000";
								txstm_reenable_fc <= '1';
								op2p_there_is_a_new_packet_to_transmit  <= '0';
							else
							   op2p_there_is_a_new_packet_to_transmit  <= '1';								
							end if;


                when others => --error
                      packet_state <= "00000000"; --go to state 0
                end case;     
					 
       end if;        
    end if;
    end process; --end packet statemachine
	 
	 --speed this up, so do it outside of the synch process:
	 packet_payloadsize_dwords_p4 <= packet_payloadsize_dwords + 4;







	--byte enable encoding to bit1:0
	 process ( trn_reset_n, rxpacket_firstdw_be )
    begin
       if (trn_reset_n = '0') then
           bit10(1 downto 0) <="00";
       else
         if (rxpacket_firstdw_be ="0001") then
			  bit10(1 downto 0) <= "00";
         elsif (rxpacket_firstdw_be ="0010") then
			  bit10(1 downto 0) <= "01";
         elsif (rxpacket_firstdw_be ="0100") then
			  bit10(1 downto 0) <= "10";
         elsif (rxpacket_firstdw_be ="1000") then
			  bit10(1 downto 0) <= "11";
         elsif (rxpacket_firstdw_be ="0011") then
			  bit10(1 downto 0) <= "00";
         elsif (rxpacket_firstdw_be ="1100") then
			  bit10(1 downto 0) <= "10";
         elsif (rxpacket_firstdw_be ="1111") then 
			  bit10(1 downto 0) <= "00";
			else --this should never happen
			  bit10(1 downto 0) <= "00";
			end if;
       end if;
    end process;
	 
	 






	-- -----------------------------------------------------------------------------------
	-- INFO TO THE LOCAL HOST ABOUT ARRIVED WRITES AND READ COMPLETIONS ------------------
	-- Basically telling that new data is in the buffer
	
	process (trn_reset_n, user_clk_i) 
    begin
    if (trn_reset_n='0') then 
			op2p_rdcompl_localaddress_regwr_en <=  '0';
			op2p_arrivedwrite_address_regwr_en <=  '0';
			op2p_rdcompl_localaddress_regdin <= (OTHERS => '0');
			op2p_arrivedwrite_address_regdin <= (OTHERS => '0');
    else
      if (user_clk_i'event and user_clk_i = '1') then

			--if the previous state was packet decoding, and now its write-arrived:
			if (packet_state_copy = "00000001" and packet_state = "00000010") then
				if (rxpacket_type="0010") then --read completion arrived
				  op2p_rdcompl_localaddress_regwr_en <=  '1';
				  op2p_arrivedwrite_address_regwr_en <=  '0';
					op2p_rdcompl_localaddress_regdin <= rxpacket_destinationaddress;
				elsif (rxpacket_type="0000") then --write data arrived
				  op2p_rdcompl_localaddress_regwr_en <=  '0';
				  op2p_arrivedwrite_address_regwr_en <=  '1';
					op2p_arrivedwrite_address_regdin <= rxpacket_destinationaddress;
				else
				  op2p_rdcompl_localaddress_regwr_en <=  '0';
				  op2p_arrivedwrite_address_regwr_en <=  '0';
				end if;
			else
				op2p_rdcompl_localaddress_regwr_en <=  '0';
				op2p_arrivedwrite_address_regwr_en <=  '0';
			end if;   
			
       end if;        
    end if;
    end process;







	 
	-- ----------------------------------------------------------------------------------- 
	--FORWARDING BUFFER MANAGER ----------------------------------------------------------
	--
	--buffer can have max 512 entries, each 2kBytes buffer, 1MBytes total.
	
    process (trn_reset_n, user_clk_i) 
    begin
    if (trn_reset_n='0') then 
       fbm_state <= "00000000"; 
		 op2p_forw_freeupaddr_regrd_en <= '0';
		 op2p_forw_freeupaddr_regrd_en_copy <=  '0';
		 forw_packetaddr_allocated <= '0';
		 forwbus_64bit <= (OTHERS => '0');
		 which_64bit_isit <= (OTHERS => '0');
		 forwbus_8bit <= (OTHERS => '0');
		 which_8bit_isit <= (OTHERS => '0');
		 which_bit_isit <= (OTHERS => '0');
			forwbuff_position <= (OTHERS => '0');
			forwbuff_position_byteoffset <= (OTHERS => '0');
			forwbuff_position_bitoffset <= (OTHERS => '0');
			fbm_nextraddress <= (OTHERS => '0');
			forwbuf_descriptor_ddword0 <= (OTHERS => '0');
			forwbuf_descriptor_ddword1 <= (OTHERS => '0');
			forwbuf_descriptor_ddword2 <= (OTHERS => '0');
			forwbuf_descriptor_ddword3 <= (OTHERS => '0');
			forwbuf_descriptor_ddword4 <= (OTHERS => '0');
			forwbuf_descriptor_ddword5 <= (OTHERS => '0');
			forwbuf_descriptor_ddword6 <= (OTHERS => '0');
			forwbuf_descriptor_ddword7 <= (OTHERS => '0');
			free_this_location <= (OTHERS => '0');
    else
      if (user_clk_i'event and user_clk_i = '1') then
                case ( fbm_state ) is

                --********** IDLE STATE  **********
					 --Wait for vector requests from the scheduler.
					 --Also wait for new entries in the freeup FIFO. Start reading the value from it here (rd_en=1).
                when "00000000" =>   --state 0        
                  if (fbm_nextraddress_req ='1') then --request from scheduler
						  fbm_state <= "00000001"; 
						elsif (op2p_forw_freeupaddr_regempty='0') then --freeup command from local host
						  fbm_state <= "00000110";
						  op2p_forw_freeupaddr_regrd_en <= '1';
						  op2p_forw_freeupaddr_regrd_en_copy <=  '1';
						end if;
						forw_packetaddr_allocated <= '0';

                --********** find step-1 STATE ********** 
                when "00000001" =>   --state 1
						--check 64bit of the descriptor table at once. first clock cycle.
						--if buffer is full, then overwrite ddw7
						if (forwbuf_descriptor_ddword0 /= X"FFFFFFFFFFFFFFFF") then
						  forwbus_64bit <= forwbuf_descriptor_ddword0;
						  which_64bit_isit <= "000";
						elsif (forwbuf_descriptor_ddword1 /= X"FFFFFFFFFFFFFFFF") then
						  forwbus_64bit <= forwbuf_descriptor_ddword1;
						  which_64bit_isit <= "001";
						elsif (forwbuf_descriptor_ddword2 /= X"FFFFFFFFFFFFFFFF") then
						  forwbus_64bit <= forwbuf_descriptor_ddword2;
						  which_64bit_isit <= "010";
						elsif (forwbuf_descriptor_ddword3 /= X"FFFFFFFFFFFFFFFF") then
						  forwbus_64bit <= forwbuf_descriptor_ddword3;
						  which_64bit_isit <= "011";
						elsif (forwbuf_descriptor_ddword4 /= X"FFFFFFFFFFFFFFFF") then
						  forwbus_64bit <= forwbuf_descriptor_ddword4;
						  which_64bit_isit <= "100";
						elsif (forwbuf_descriptor_ddword5 /= X"FFFFFFFFFFFFFFFF") then
						  forwbus_64bit <= forwbuf_descriptor_ddword5;
						  which_64bit_isit <= "101";
						elsif (forwbuf_descriptor_ddword6 /= X"FFFFFFFFFFFFFFFF") then
						  forwbus_64bit <= forwbuf_descriptor_ddword6;
						  which_64bit_isit <= "110";
						else --elsif (forwbuf_descriptor_ddword7 /= X"FFFFFFFFFFFFFFFF") then
						  forwbus_64bit <= forwbuf_descriptor_ddword7;
						  which_64bit_isit <= "111";
						end if;
						fbm_state <= "00000010"; --next
						--fast (ststic timing path) version:
--						if (forwbuf_descriptor_ddword0 = X"FFFFFFFFFFFFFFFF" 
--							 and forwbuf_descriptor_ddword1 = X"FFFFFFFFFFFFFFFF"
--							 and forwbuf_descriptor_ddword2 = X"FFFFFFFFFFFFFFFF"
--							 and forwbuf_descriptor_ddword3 = X"FFFFFFFFFFFFFFFF") then
--							if (forwbuf_descriptor_ddword4 = X"FFFFFFFFFFFFFFFF"
--								 and forwbuf_descriptor_ddword5 = X"FFFFFFFFFFFFFFFF") then
--								if (forwbuf_descriptor_ddword6 = X"FFFFFFFFFFFFFFFF") then
--								  forwbus_64bit <= forwbuf_descriptor_ddword7;
--								  which_64bit_isit <= "111";
--								else
--								  forwbus_64bit <= forwbuf_descriptor_ddword6;
--								  which_64bit_isit <= "110";
--								end if;
--							else
--								if (forwbuf_descriptor_ddword4 = X"FFFFFFFFFFFFFFFF") then
--								  forwbus_64bit <= forwbuf_descriptor_ddword5;
--								  which_64bit_isit <= "101";
--								else
--								  forwbus_64bit <= forwbuf_descriptor_ddword4;
--								  which_64bit_isit <= "100";
--								end if;
--							end if;
--						else
--							if (and forwbuf_descriptor_ddword0 = X"FFFFFFFFFFFFFFFF"
--								 and forwbuf_descriptor_ddword1 = X"FFFFFFFFFFFFFFFF") then
--								if (forwbuf_descriptor_ddword2 = X"FFFFFFFFFFFFFFFF") then
--								  forwbus_64bit <= forwbuf_descriptor_ddword3;
--								  which_64bit_isit <= "011";
--								else
--								  forwbus_64bit <= forwbuf_descriptor_ddword2;
--								  which_64bit_isit <= "010";
--								end if;
--							else
--								if (forwbuf_descriptor_ddword0 = X"FFFFFFFFFFFFFFFF") then
--								  forwbus_64bit <= forwbuf_descriptor_ddword1;
--								  which_64bit_isit <= "001";
--								else
--								  forwbus_64bit <= forwbuf_descriptor_ddword0;
--								  which_64bit_isit <= "000";
--								end if;
--							end if;
--						end if;
						

                --********** find step-2 STATE **********     				 
                when "00000010" =>   --state 2
						--second clock cycle, analyse the 64bit, break it to a final byte:
						--if buffer full, overwrite last byte
						if (forwbuf_descriptor_byte0 /= X"FF") then
						  forwbus_8bit <= forwbuf_descriptor_byte0;
						  which_8bit_isit <= "000";
						elsif (forwbuf_descriptor_byte1 /= X"FF") then
						  forwbus_8bit <= forwbuf_descriptor_byte1;
						  which_8bit_isit <= "001";
						elsif (forwbuf_descriptor_byte2 /= X"FF") then
						  forwbus_8bit <= forwbuf_descriptor_byte2;
						  which_8bit_isit <= "010";
						elsif (forwbuf_descriptor_byte3 /= X"FF") then
						  forwbus_8bit <= forwbuf_descriptor_byte3;
						  which_8bit_isit <= "011";
						elsif (forwbuf_descriptor_byte4 /= X"FF") then
						  forwbus_8bit <= forwbuf_descriptor_byte4;
						  which_8bit_isit <= "100";
						elsif (forwbuf_descriptor_byte5 /= X"FF") then
						  forwbus_8bit <= forwbuf_descriptor_byte5;
						  which_8bit_isit <= "101";
						elsif (forwbuf_descriptor_byte6 /= X"FF") then
						  forwbus_8bit <= forwbuf_descriptor_byte6;
						  which_8bit_isit <= "110";
						else -- elsif (forwbuf_descriptor_byte7 /= X"FF") then
						  forwbus_8bit <= forwbuf_descriptor_byte7;
						  which_8bit_isit <= "111";
						end if;
						fbm_state <= "00000011"; --next
	
                --********** find step-3 STATE **********     				 
                when "00000011" =>   --state 3
						--3rd clock cycle: find a zero bit in the chosen byte: 
						if (forwbuf_descriptor_bit0 = '0') then
						  which_bit_isit <= "000";
						elsif (forwbuf_descriptor_bit1 = '0') then
						  which_bit_isit <= "001";
						elsif (forwbuf_descriptor_bit2 = '0') then
						  which_bit_isit <= "010";
						elsif (forwbuf_descriptor_bit3 = '0') then
						  which_bit_isit <= "011";
						elsif (forwbuf_descriptor_bit4 = '0') then
						  which_bit_isit <= "100";
						elsif (forwbuf_descriptor_bit5 = '0') then
						  which_bit_isit <= "101";
						elsif (forwbuf_descriptor_bit6 = '0') then
						  which_bit_isit <= "110";
						else --elsif(forwbuf_descriptor_bit7 = '0') then
						  which_bit_isit <= "111";
						end if;
						fbm_state <= "00000100"; --next
	
                --********** find step-4 STATE **********     				 
                when "00000100" =>   --state 4
						--4th clock cycle: generate the address with one clock cycle delay, for sufficient timing margin
						forwbuff_position(8 downto 6) <= which_64bit_isit;
						forwbuff_position(5 downto 3) <= which_8bit_isit;
						forwbuff_position(2 downto 0) <= which_bit_isit;
						fbm_state <= "00000101"; --next
						--address offset in DRAM:
						forwbuff_position_byteoffset(19 downto 17) <= which_64bit_isit;
						forwbuff_position_byteoffset(16 downto 14) <= which_8bit_isit;
						forwbuff_position_byteoffset(13 downto 11) <= which_bit_isit;
						forwbuff_position_byteoffset(10 downto 0) <= "00000000000"; --since we use 2kB blocks
						--location code in 64bit location registers:
						forwbuff_position_bitoffset(5 downto 3) <= which_8bit_isit;
						forwbuff_position_bitoffset(2 downto 0) <= which_bit_isit;
	
                --********** tell the result STATE ********** 
					 --Tell the vector to the scheduler, and set the bit here as used (1)   				 
                when "00000101" =>   --state 5
                    fbm_nextraddress <= forwbuff_position_byteoffset + op2p_forwarding_bufferbase_reg;
						  forw_packetaddr_allocated <= '1';
						  fbm_state <= "00001101"; --back to idle (but first wait one clock)
						  --set the bit as occupied:
						  if    (which_64bit_isit = "000") then
						    forwbuf_descriptor_ddword0 (CONV_INTEGER(forwbuff_position_bitoffset)) <= '1';
						  elsif (which_64bit_isit = "001") then
						    forwbuf_descriptor_ddword1 (CONV_INTEGER(forwbuff_position_bitoffset)) <= '1';
						  elsif (which_64bit_isit = "010") then
						    forwbuf_descriptor_ddword2 (CONV_INTEGER(forwbuff_position_bitoffset)) <= '1';
						  elsif (which_64bit_isit = "011") then
						    forwbuf_descriptor_ddword3 (CONV_INTEGER(forwbuff_position_bitoffset)) <= '1';
						  elsif (which_64bit_isit = "100") then
						    forwbuf_descriptor_ddword4 (CONV_INTEGER(forwbuff_position_bitoffset)) <= '1';
						  elsif (which_64bit_isit = "101") then
						    forwbuf_descriptor_ddword5 (CONV_INTEGER(forwbuff_position_bitoffset)) <= '1';
						  elsif (which_64bit_isit = "110") then
						    forwbuf_descriptor_ddword6 (CONV_INTEGER(forwbuff_position_bitoffset)) <= '1';
						  elsif (which_64bit_isit = "111") then
						    forwbuf_descriptor_ddword7 (CONV_INTEGER(forwbuff_position_bitoffset)) <= '1';
						  end if;

                --********** Wait STATE ********** 
					 --Tell the vector to the scheduler, and set the bit here as used (1)   				 
                when "00001101" =>   --state 13
							fbm_state <= "00000000"; --back to idle

                --********** Freeup STATE ********** 
					 --If the freeup FIFO had a new entry, free up the bit (set to zero)
					 --This state must be 2 clock cycles: 1- calculate bitposition from address value, 2-write bit and go to IDLE				 
                when "00000110" =>   --state 6
                    op2p_forw_freeupaddr_regrd_en <= '0';
						  op2p_forw_freeupaddr_regrd_en_copy <= '0';
						  fbm_state <= "00000111";
					 when "00000111" =>   --state 7
							free_this_location <= op2p_forw_freeupaddr_regdout - op2p_forwarding_bufferbase_reg;
							fbm_state <= "00001000";
					 when "00001000" =>   --state 8
							  fbm_state <= "00000000"; --back to idle
							  --set the bit as free:
							  if    (which_64bit_isit_tofreeup = "000") then
								 forwbuf_descriptor_ddword0 (CONV_INTEGER(which_bit_isit_tofreeup)) <= '0';
							  elsif (which_64bit_isit_tofreeup = "001") then
								 forwbuf_descriptor_ddword1 (CONV_INTEGER(which_bit_isit_tofreeup)) <= '0';
							  elsif (which_64bit_isit_tofreeup = "010") then
								 forwbuf_descriptor_ddword2 (CONV_INTEGER(which_bit_isit_tofreeup)) <= '0';
							  elsif (which_64bit_isit_tofreeup = "011") then
								 forwbuf_descriptor_ddword3 (CONV_INTEGER(which_bit_isit_tofreeup)) <= '0';
							  elsif (which_64bit_isit_tofreeup = "100") then
								 forwbuf_descriptor_ddword4 (CONV_INTEGER(which_bit_isit_tofreeup)) <= '0';
							  elsif (which_64bit_isit_tofreeup = "101") then
								 forwbuf_descriptor_ddword5 (CONV_INTEGER(which_bit_isit_tofreeup)) <= '0';
							  elsif (which_64bit_isit_tofreeup = "110") then
								 forwbuf_descriptor_ddword6 (CONV_INTEGER(which_bit_isit_tofreeup)) <= '0';
							  elsif (which_64bit_isit_tofreeup = "111") then
								 forwbuf_descriptor_ddword7 (CONV_INTEGER(which_bit_isit_tofreeup)) <= '0';
							  end if;
						  
                when others => --error
                      fbm_state <= "00000000"; --back to idle
                end case;     
       end if;        
    end if;
    end process;
	 
	--asynchronous: (just renaming some bits, without logic)
	forwbuf_descriptor_byte0 <= forwbus_64bit(7 downto 0);
	forwbuf_descriptor_byte1 <= forwbus_64bit(15 downto 8);
	forwbuf_descriptor_byte2 <= forwbus_64bit(23 downto 16);
	forwbuf_descriptor_byte3 <= forwbus_64bit(31 downto 24);
	forwbuf_descriptor_byte4 <= forwbus_64bit(39 downto 32);
	forwbuf_descriptor_byte5 <= forwbus_64bit(47 downto 40);
	forwbuf_descriptor_byte6 <= forwbus_64bit(55 downto 48);
	forwbuf_descriptor_byte7 <= forwbus_64bit(63 downto 56);
	forwbuf_descriptor_bit0 <= forwbus_8bit(0);
	forwbuf_descriptor_bit1 <= forwbus_8bit(1);
	forwbuf_descriptor_bit2 <= forwbus_8bit(2);
	forwbuf_descriptor_bit3 <= forwbus_8bit(3);
	forwbuf_descriptor_bit4 <= forwbus_8bit(4);
	forwbuf_descriptor_bit5 <= forwbus_8bit(5);
	forwbuf_descriptor_bit6 <= forwbus_8bit(6);
	forwbuf_descriptor_bit7 <= forwbus_8bit(7);
	which_64bit_isit_tofreeup <= free_this_location (19 downto 17);
	which_bit_isit_tofreeup <= free_this_location (16 downto 11);

	op2p_forw_freeupsize_regrd_en <= '0'; --not in use












-- -------- END OF FILE -----------------------------------------------------------
end Behavioral;







---- REQUIRED MODIFICATIONS ON THE GENERATED AURORA FILES: ------------------------------------------------------
--
----  This design includes the aurora interface core which was generated by the Xilinx 
----  CoreGenerator. All the VHD files were copied here, including the ones from the 
----  "Reference Design" folder. This file is the top level source of the module, 
----  and is not generated by CoreGen. Search for all VHD files in all subfolders, then copy all.
----  2 files had to be modified (the ones from the example design folder)
--
----  The last one has its filename and module name also modified, not only the internal logic.
----  If we use different Refclk/Linerate/widths/device-type, then we have to regenerate the
----  the Aurora core, and re-modify the files
--
----SOME MORE NOTES:
---- The file was originally generated by the Xilinx Core Generator, but
---- since that tool does not create easily useable blackbox IPs, I had to 
---- modify the top level of it. (Istvan NAgy, buenos(at)freemail.hu)
----  this is to hold all the files from the reference design sources.
----  Modification: remove the frame gen/check and chipscope and route the LocalLink ports up.
----user clock for the parallel bus:
----this is generated by external signal, and distributed up and down to every node.
----user_clk_i_local is used in this file, user_clk_i goes up one level
--
----The aurora_8b10b_v5_1_FRAME_CHECK, the aurora_8b10b_v5_1_FRAME_GEN, and the ICON core
----were removed, and their connections were eliminated.
--
----FILE COPY: 
----1.) Use search in the folder "aurora_8b10b_v5_1" for *.VHD files.
----2.) select all of them
----3.) De-select the following (ctrl+click):
----			aurora_8b10b_v5_1_example_design.vhd
----			demo_tb.vhd
----			aurora_8b10b_v5_1_frame_check.vhd
----			aurora_8b10b_v5_1_frame_gen.vhd
----4.) Copy the selected files into the project's source folder "User_Sources"
----    to overwrite all files there.
----5.) modify 2 files based on the instructions below.
--
--
----  FILE-1: 
----  aurora_8b10b_v5_1_reset_logic.vhd =========================================================================
--		REPLACE MY OLD FILE WITH A NEW ONE, AND CHANGE THE FOLLOWING:
--
--				##COMMENT THIS OUT -----------------------------------------
--							 -- Assign an IBUFG to INIT_CLK
--							 init_clk_ibufg_i : IBUFG 
--							 port map
--							 (
--								  I   =>  INIT_CLK,
--								  O   =>  init_clk_i
--							 );
--
--				##THEN COPY THIS IN -----------------------------------------
--							 init_clk_i <= INIT_CLK;
--
--
--
--
----  FILE-2: 
----  aurora_8b10b_v5_1_example_des_modified.vhd =================================================================
--		DO NOT OVERWRITE MY OLD FILE WITH A NEWLY GENERATED ONE
--		MODIFY MY OLD FILE WITH SOME DATA FROM THE NEW FILE:
--
--
--		##REPLACE THIS:  -----------------------------------------
--			  attribute core_generation_info           : string;
--			  attribute core_generation_info of MAPPED : architecture is "aurora_8b10b_v5_1,aurora_8b10b_ ...
--			-- Parameter Declarations --
--				 constant DLY : time := 1 ns;
--			-- External Register Declarations --
--		##TO THE SAME PART FROM THE NEW FILE (\example_design\aurora_8b10b_v5_1_example_design.vhd)
--
--
--		##IF NECESSARY, REPLACE THE ARCHITECTURE NAME   -----------------------------------------
--		##FROM: MAPPED
--		##TO: behavioral
--
--
--		##IF NECESSARY, REPLACE THE MODULE NAMES   -----------------------------------------
--		##FROM: aurora_8b10b_v5_1
--		##TO: THENEW NAME COMING FROM THE CORE GENERATOR. IT MIGHT USE A NEW VERSION OF THE CORE
--
--
--		##CHANGE THE GTP AND REFCLOCK PORTS IF NEEDED -----------------------------------------
--		##IN THE TOP PORT LIST AND ALSO INTERNALLY TO 
--		##THE USED PORT WIDTHS OR NAMES. BASED ON THE BOARD DESIGN
--		##FOR EXAMPLE FROM THIS:
--					  GTPD1_P   : in  std_logic;
--					  GTPD1_N   : in  std_logic;
--						RXP               : in std_logic_vector(0 to 1);
--						RXN               : in std_logic_vector(0 to 1);
--						TXP               : out std_logic_vector(0 to 1);
--						TXN               : out std_logic_vector(0 to 1)
--		##TO THIS:
--					  GTPD0_P   : in  std_logic;
--					  GTPD0_N   : in  std_logic;
--						RXP               : in std_logic_vector(0 to 4);
--						RXN               : in std_logic_vector(0 to 4);
--						TXP               : out std_logic_vector(0 to 4);
--						TXN               : out std_logic_vector(0 to 4)
--
--
--
--
--










