// Copyright (C) 2022, Andes Technology Corp. Confidential Proprietary

module kv_dsp_dec (
    instr,
    src2_sel_imm,
    src3_sel_imm,
    src4_sel_imm,
    src2_imm,
    src3_imm,
    src4_imm,
    operand_ctrl,
    function_ctrl,
    result_ctrl,
    overflow_ctrl
);
localparam OP_DSP = 7'b1111111;
localparam DSP_OCTRL_WIDTH = 44;
localparam DSP_FCTRL_WIDTH = 151;
localparam DSP_RCTRL_WIDTH = 70;
localparam DSP_HCTRL_WIDTH = 3;
input [31:0] instr;
output [DSP_OCTRL_WIDTH - 1:0] operand_ctrl;
output [DSP_FCTRL_WIDTH - 1:0] function_ctrl;
output [DSP_RCTRL_WIDTH - 1:0] result_ctrl;
output overflow_ctrl;
output src2_sel_imm;
output src3_sel_imm;
output src4_sel_imm;
output [31:0] src2_imm;
output [31:0] src3_imm;
output [31:0] src4_imm;


wire s0;
wire s1;
wire s2;
wire s3;
wire s4;
wire s5;
wire s6;
wire s7;
wire s8;
wire s9;
wire s10;
wire s11;
wire s12;
wire s13;
wire s14;
wire s15;
wire s16;
wire s17;
wire s18;
wire s19;
wire s20;
wire s21;
wire s22;
wire s23;
wire s24;
wire s25;
wire s26;
wire s27;
wire s28;
wire s29;
wire s30;
wire s31;
wire s32;
wire s33;
wire s34;
wire s35;
wire s36;
wire s37;
wire s38;
wire s39;
wire s40;
wire s41;
wire s42;
wire s43;
wire s44;
wire s45;
wire s46;
wire s47;
wire s48;
wire s49;
wire s50;
wire s51;
wire s52;
wire s53;
wire s54;
wire s55;
wire s56;
wire s57;
wire s58;
wire s59;
wire s60;
wire s61;
wire s62;
wire s63;
wire s64;
wire s65;
wire s66;
wire s67;
wire s68;
wire s69;
wire s70;
wire s71;
wire s72;
wire s73;
wire s74;
wire s75;
wire s76;
wire s77;
wire s78;
wire s79;
wire s80;
wire s81;
wire s82;
wire s83;
wire s84;
wire s85;
wire s86;
wire s87;
wire s88;
wire s89;
wire s90;
wire s91;
wire s92;
wire s93;
wire s94;
wire s95;
wire s96;
wire s97;
wire s98;
wire s99;
wire s100;
wire s101;
wire s102;
wire s103;
wire s104;
wire s105;
wire s106;
wire s107;
wire s108;
wire s109;
wire s110;
wire s111;
wire s112;
wire s113;
wire s114;
wire s115;
wire s116;
wire s117;
wire s118;
wire s119;
wire s120;
wire s121;
wire s122;
wire s123;
wire s124;
wire s125;
wire s126;
wire s127;
wire s128;
wire s129;
wire s130;
wire s131;
wire s132;
wire s133;
wire s134;
wire s135;
wire s136;
wire s137;
wire s138;
wire s139;
wire s140;
wire s141;
wire s142;
wire s143;
wire s144;
wire s145;
wire s146;
wire s147;
wire s148;
wire s149;
wire s150;
wire s151;
wire s152;
wire s153;
wire s154;
wire s155;
wire s156;
wire s157;
wire s158;
wire s159;
wire s160;
wire s161;
wire s162;
wire s163;
wire s164;
wire s165;
wire s166;
wire s167;
wire s168;
wire s169;
wire s170;
wire s171;
wire s172;
wire s173;
wire s174;
wire s175;
wire s176;
wire s177;
wire s178;
wire s179;
wire s180;
wire s181;
wire s182;
wire s183;
wire s184;
wire s185;
wire s186;
wire s187;
wire s188;
wire s189;
wire s190;
wire s191;
wire s192;
wire s193;
wire s194;
wire s195;
wire s196;
wire s197;
wire s198;
wire s199;
wire s200;
wire s201;
wire s202;
wire s203;
wire s204;
wire s205;
wire s206;
wire s207;
wire s208;
wire s209;
wire s210;
wire s211;
wire s212;
wire s213;
wire s214;
wire s215;
wire s216;
wire s217;
wire s218;
wire s219;
wire s220;
wire s221;
wire s222;
wire s223;
wire s224;
wire s225;
wire s226;
wire s227;
wire s228;
wire s229;
wire s230;
wire s231;
wire s232;
wire s233;
wire s234;
wire s235;
wire s236;
wire s237;
wire s238;
wire s239;
wire s240;
wire s241;
wire s242;
wire s243;
wire s244;
wire s245;
wire s246;
wire s247;
wire s248;
wire s249;
wire s250;
wire s251;
wire s252;
wire s253;
wire s254;
wire s255;
wire s256;
wire s257;
wire s258;
wire s259;
wire s260;
wire s261;
wire s262;
wire s263;
wire s264;
wire s265;
wire s266;
wire s267;
wire s268;
wire s269;
wire s270;
wire s271;
wire s272;
wire s273;
wire s274;
wire s275;
wire s276;
wire s277;
wire s278;
wire s279;
wire s280;
wire s281;
wire s282;
wire s283;
wire s284;
wire s285;
wire s286;
wire s287;
wire s288;
wire s289;
wire s290;
wire s291;
wire s292;
wire s293;
wire s294;
wire s295;
wire s296;
wire s297;
wire s298;
wire s299;
wire s300;
wire s301;
wire s302;
wire s303;
wire s304;
wire s305;
wire s306;
wire s307;
wire s308;
wire s309;
wire s310;
wire s311;
wire s312;
wire s313;
wire s314;
wire s315;
wire s316;
wire s317;
wire s318;
wire s319;
wire s320;
wire s321;
wire s322;
wire s323;
wire s324;
wire s325;
wire s326;
wire s327;
wire s328;
wire [31:0] s329;
wire s330;
wire s331;
wire [4:0] s332;
wire [31:0] s333;
wire [31:0] s334;
wire [31:0] s335;
wire [31:0] s336;
assign s0 = (instr[31:25] == 7'b0100100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s1 = (instr[31:25] == 7'b0100000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s2 = (instr[31:25] == 7'b1100000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s3 = (instr[31:25] == 7'b1110000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s4 = (instr[31:25] == 7'b1110011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s5 = (instr[31:26] == 6'b111010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s6 = (instr[31:30] == 2'b11) & (instr[14:12] == 3'b010) & (instr[6:0] == OP_DSP);
assign s7 = (instr[31:20] == 12'b101011100000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s8 = (instr[31:20] == 12'b101011101000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s9 = (instr[31:20] == 12'b101011111000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s10 = (instr[31:20] == 12'b101011100011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s11 = (instr[31:20] == 12'b101011101011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s12 = (instr[31:20] == 12'b101011111011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s13 = (instr[31:20] == 12'b101011100001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s14 = (instr[31:20] == 12'b101011101001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s15 = (instr[31:20] == 12'b101011111001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s16 = (instr[31:25] == 7'b0100111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s17 = (instr[31:25] == 7'b0100110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s18 = (instr[31:25] == 7'b0100010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s19 = (instr[31:25] == 7'b0100011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s20 = (instr[31:23] == 9'b101011000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s21 = (instr[31:20] == 12'b101011010000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s22 = (instr[31:20] == 12'b101011010001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s23 = (instr[31:20] == 12'b101011010100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s24 = (instr[31:25] == 7'b0001100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s25 = (instr[31:25] == 7'b0001000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s26 = (instr[31:25] == 7'b1001000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s27 = (instr[31:25] == 7'b0000010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s28 = (instr[31:25] == 7'b0000000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s29 = (instr[31:25] == 7'b0001010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s30 = (instr[31:25] == 7'b0001011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s31 = (instr[31:25] == 7'b0000101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s32 = (instr[31:25] == 7'b0001101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s33 = (instr[31:25] == 7'b0010101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s34 = (instr[31:25] == 7'b1101001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s35 = (instr[31:25] == 7'b1110001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s36 = (instr[31:25] == 7'b1111001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s37 = (instr[31:25] == 7'b1000111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s38 = (instr[31:25] == 7'b1001111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s39 = (instr[31:25] == 7'b1000011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s40 = (instr[31:25] == 7'b1001011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s41 = (instr[31:25] == 7'b0000110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s42 = (instr[31:25] == 7'b0001110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s43 = (instr[31:25] == 7'b0010110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s44 = (instr[31:25] == 7'b0101101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s45 = (instr[31:25] == 7'b0110101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s46 = (instr[31:25] == 7'b0111101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s47 = (instr[31:25] == 7'b0100100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s48 = (instr[31:25] == 7'b0100101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s49 = (instr[31:25] == 7'b0101110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s50 = (instr[31:25] == 7'b0110110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s51 = (instr[31:25] == 7'b0111110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s52 = (instr[31:25] == 7'b1001010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s53 = (instr[31:25] == 7'b0011100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s54 = (instr[31:25] == 7'b0011101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s55 = (instr[31:25] == 7'b0110000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s56 = (instr[31:25] == 7'b0111000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s57 = (instr[31:25] == 7'b0100011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s58 = (instr[31:25] == 7'b0101011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s59 = (instr[31:25] == 7'b1100111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s60 = (instr[31:25] == 7'b1101111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s61 = (instr[31:25] == 7'b0110011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s62 = (instr[31:25] == 7'b0111011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s63 = (instr[31:25] == 7'b1110111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s64 = (instr[31:25] == 7'b1111111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s65 = (instr[31:25] == 7'b0100001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s66 = (instr[31:25] == 7'b0101001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s67 = (instr[31:25] == 7'b1000111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s68 = (instr[31:25] == 7'b1001111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s69 = (instr[31:25] == 7'b1010111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s70 = (instr[31:25] == 7'b1011111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s71 = (instr[31:25] == 7'b0100110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s72 = (instr[31:25] == 7'b0100111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s73 = (instr[31:25] == 7'b1001011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s74 = (instr[31:25] == 7'b0010011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s75 = (instr[31:25] == 7'b0011011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s76 = (instr[31:25] == 7'b0110110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s77 = (instr[31:23] == 9'b011111001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s78 = (instr[31:25] == 7'b0110010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s79 = (instr[31:24] == 8'b01110101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s80 = (instr[31:25] == 7'b0101111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s81 = (instr[31:25] == 7'b0110111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s82 = (instr[31:25] == 7'b0101011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s83 = (instr[31:25] == 7'b0110011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s84 = (instr[31:25] == 7'b0110111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s85 = (instr[31:25] == 7'b0111111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s86 = (instr[31:25] == 7'b0001010) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s87 = (instr[31:25] == 7'b0001011) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s88 = (instr[31:25] == 7'b0001101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s89 = (instr[31:25] == 7'b0001001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s90 = (instr[31:25] == 7'b1001001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s91 = (instr[31:25] == 7'b0000011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s92 = (instr[31:25] == 7'b0000001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s93 = (instr[31:25] == 7'b0110001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s94 = (instr[31:25] == 7'b0111001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s95 = (instr[31:25] == 7'b1100010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s96 = (instr[31:25] == 7'b1111001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s97 = (instr[31:25] == 7'b1111000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s98 = (instr[31:25] == 7'b1100011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s99 = (instr[31:25] == 7'b1111000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s100 = (instr[31:25] == 7'b1110000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s101 = (instr[31:25] == 7'b1111110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s102 = (instr[31:25] == 7'b1111111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s103 = (instr[31:25] == 7'b0000111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s104 = (instr[31:25] == 7'b0001111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s105 = (instr[31:25] == 7'b0010111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s106 = (instr[31:25] == 7'b0011111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s107 = (instr[31:25] == 7'b0000100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s108 = (instr[31:25] == 7'b0000000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s109 = (instr[31:25] == 7'b1000000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s110 = (instr[31:25] == 7'b0010000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s111 = (instr[31:25] == 7'b0000010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s112 = (instr[31:25] == 7'b0000011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s113 = (instr[31:25] == 7'b0000010) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s114 = (instr[31:25] == 7'b0000011) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s115 = (instr[31:25] == 7'b0000101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s116 = (instr[31:25] == 7'b0000001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s117 = (instr[31:25] == 7'b1000001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s118 = (instr[31:25] == 7'b0010001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s119 = (instr[31:23] == 9'b100011000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s120 = (instr[31:24] == 8'b10000100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s121 = (instr[31:25] == 7'b1110010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s122 = (instr[31:25] == 7'b0001111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s123 = (instr[31:25] == 7'b0001110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s124 = (instr[31:25] == 7'b0000111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s125 = (instr[31:25] == 7'b0000110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s126 = (instr[31:25] == 7'b0101110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s127 = (instr[31:23] == 9'b011111000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s128 = (instr[31:25] == 7'b0101010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s129 = (instr[31:24] == 8'b01110100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s130 = (instr[31:25] == 7'b0101111) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s131 = (instr[31:25] == 7'b1000100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s132 = (instr[31:25] == 7'b1001100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s133 = (instr[31:25] == 7'b1010100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s134 = (instr[31:25] == 7'b1000110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s135 = (instr[31:25] == 7'b1001110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s136 = (instr[31:25] == 7'b1000101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s137 = (instr[31:25] == 7'b1001101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s138 = (instr[31:25] == 7'b1010101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s139 = (instr[31:25] == 7'b1000010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s140 = (instr[31:25] == 7'b1100100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s141 = (instr[31:25] == 7'b1100101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s142 = (instr[31:25] == 7'b1000101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s143 = (instr[31:25] == 7'b1000001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s144 = (instr[31:25] == 7'b0000100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s145 = (instr[31:25] == 7'b0001100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s146 = (instr[31:25] == 7'b0010100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s147 = (instr[31:25] == 7'b0101100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s148 = (instr[31:25] == 7'b0110100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s149 = (instr[31:25] == 7'b0111100) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s150 = (instr[31:25] == 7'b1000100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s151 = (instr[31:25] == 7'b1000000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s152 = (instr[31:25] == 7'b0100000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s153 = (instr[31:25] == 7'b0101000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s154 = (instr[31:25] == 7'b0100010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s155 = (instr[31:25] == 7'b0101010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s156 = (instr[31:25] == 7'b0110010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s157 = (instr[31:25] == 7'b0111010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s158 = (instr[31:25] == 7'b1010110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s159 = (instr[31:25] == 7'b1011110) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s160 = (instr[31:25] == 7'b1000011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s161 = (instr[31:25] == 7'b1010100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s162 = (instr[31:25] == 7'b1010101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s163 = (instr[31:25] == 7'b1010000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s164 = (instr[31:25] == 7'b1010001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s165 = (instr[31:25] == 7'b0010010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s166 = (instr[31:26] == 6'b110101) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s167 = (instr[31:25] == 7'b0101100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s168 = (instr[31:25] == 7'b0110100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s169 = (instr[31:23] == 9'b011110000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s170 = (instr[31:23] == 9'b011110001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s171 = (instr[31:25] == 7'b0101000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s172 = (instr[31:25] == 7'b0110000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s173 = (instr[31:24] == 8'b01110000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s174 = (instr[31:24] == 8'b01110001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s175 = (instr[31:25] == 7'b0101101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s176 = (instr[31:25] == 7'b0110101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s177 = (instr[31:23] == 9'b011110100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s178 = (instr[31:23] == 9'b011110101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s179 = (instr[31:25] == 7'b0101001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s180 = (instr[31:25] == 7'b0110001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s181 = (instr[31:24] == 8'b01110010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s182 = (instr[31:24] == 8'b01110011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s183 = (instr[31:25] == 7'b0100010) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s184 = (instr[31:25] == 7'b0100011) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s185 = (instr[31:25] == 7'b0100101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s186 = (instr[31:25] == 7'b0100001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s187 = (instr[31:25] == 7'b1100001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s188 = (instr[31:20] == 12'b101011001000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s189 = (instr[31:20] == 12'b101011001001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s190 = (instr[31:20] == 12'b101011001010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s191 = (instr[31:20] == 12'b101011001011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s192 = (instr[31:20] == 12'b101011010011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s193 = (instr[31:20] == 12'b101011011000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s194 = (instr[31:20] == 12'b101011011001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s195 = (instr[31:23] == 9'b100011010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s196 = (instr[31:24] == 8'b10000101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s197 = (instr[31:25] == 7'b1111010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s198 = (instr[31:25] == 7'b0011111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s199 = (instr[31:25] == 7'b0011110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s200 = (instr[31:25] == 7'b0010111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s201 = (instr[31:25] == 7'b0010110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s202 = (instr[31:25] == 7'b0011100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s203 = (instr[31:25] == 7'b0011000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s204 = (instr[31:25] == 7'b1011000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s205 = (instr[31:25] == 7'b0001010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s206 = (instr[31:25] == 7'b0001000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s207 = (instr[31:25] == 7'b0011010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s208 = (instr[31:25] == 7'b0011011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s209 = (instr[31:25] == 7'b1011010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s210 = (instr[31:25] == 7'b1011011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s211 = (instr[31:25] == 7'b0011010) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s212 = (instr[31:25] == 7'b0011011) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s213 = (instr[31:25] == 7'b0011101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s214 = (instr[31:25] == 7'b0011001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s215 = (instr[31:25] == 7'b1011001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s216 = (instr[31:25] == 7'b0001011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s217 = (instr[31:25] == 7'b0001001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s218 = (instr[31:25] == 7'b1010010) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s219 = (instr[31:25] == 7'b1100110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s220 = (instr[31:25] == 7'b1001101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s221 = (instr[31:25] == 7'b1001001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s222 = (instr[31:25] == 7'b1001100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s223 = (instr[31:25] == 7'b1001000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s224 = (instr[31:25] == 7'b1010011) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s225 = (instr[31:25] == 7'b1011100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s226 = (instr[31:25] == 7'b1011101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s227 = (instr[31:25] == 7'b1011000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s228 = (instr[31:25] == 7'b1011001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s229 = (instr[31:25] == 7'b0010100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s230 = (instr[31:25] == 7'b0010000) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s231 = (instr[31:25] == 7'b1010000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s232 = (instr[31:25] == 7'b0011000) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s233 = (instr[31:25] == 7'b0010010) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s234 = (instr[31:25] == 7'b0010011) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s235 = (instr[31:25] == 7'b0010010) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s236 = (instr[31:25] == 7'b0010011) & (instr[14:12] == 3'b011) & (instr[6:0] == OP_DSP);
assign s237 = (instr[31:25] == 7'b0010101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s238 = (instr[31:25] == 7'b0010001) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s239 = (instr[31:25] == 7'b1010001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s240 = (instr[31:25] == 7'b0011001) & (instr[14:12] == 3'b001) & (instr[6:0] == OP_DSP);
assign s241 = (instr[31:25] == 7'b1101111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s242 = (instr[31:25] == 7'b1100111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s243 = (instr[31:20] == 12'b101011001100) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s244 = (instr[31:20] == 12'b101011001101) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s245 = (instr[31:20] == 12'b101011001110) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s246 = (instr[31:20] == 12'b101011001111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s247 = (instr[31:20] == 12'b101011010111) & (instr[14:12] == 3'b000) & (instr[6:0] == OP_DSP);
assign s248 = 1'b0;
assign s249 = 1'b0;
assign s250 = 1'b0;
assign s251 = 1'b0;
assign s252 = 1'b0;
assign s253 = 1'b0;
assign s254 = 1'b0;
assign s255 = 1'b0;
assign s256 = 1'b0;
assign s257 = 1'b0;
assign s258 = 1'b0;
assign s259 = 1'b0;
assign s260 = 1'b0;
assign s261 = 1'b0;
assign s262 = 1'b0;
assign s263 = 1'b0;
assign s264 = 1'b0;
assign s265 = 1'b0;
assign s266 = 1'b0;
assign s267 = 1'b0;
assign s268 = 1'b0;
assign s269 = 1'b0;
assign s270 = 1'b0;
assign s271 = 1'b0;
assign s272 = 1'b0;
assign s273 = 1'b0;
assign s274 = 1'b0;
assign s275 = 1'b0;
assign s276 = 1'b0;
assign s277 = 1'b0;
assign s278 = 1'b0;
assign s279 = 1'b0;
assign s280 = 1'b0;
assign s281 = 1'b0;
assign s282 = 1'b0;
assign s283 = 1'b0;
assign s284 = 1'b0;
assign s285 = 1'b0;
assign s286 = 1'b0;
assign s287 = 1'b0;
assign s288 = 1'b0;
assign s289 = 1'b0;
assign s290 = 1'b0;
assign s291 = 1'b0;
assign s292 = 1'b0;
assign s293 = 1'b0;
assign s294 = 1'b0;
assign s295 = 1'b0;
assign s296 = 1'b0;
assign s297 = 1'b0;
assign s298 = 1'b0;
assign s299 = 1'b0;
assign s300 = 1'b0;
assign s301 = 1'b0;
assign s302 = 1'b0;
assign s303 = 1'b0;
assign s304 = 1'b0;
assign s305 = 1'b0;
assign s306 = 1'b0;
assign s307 = 1'b0;
assign s308 = 1'b0;
assign s309 = 1'b0;
assign s310 = 1'b0;
assign s311 = 1'b0;
assign s312 = 1'b0;
assign s313 = 1'b0;
assign s314 = 1'b0;
assign s315 = 1'b0;
assign s316 = 1'b0;
assign s317 = 1'b0;
assign s318 = 1'b0;
assign s319 = 1'b0;
assign s320 = 1'b0;
assign s321 = 1'b0;
assign s322 = 1'b0;
assign s323 = 1'b0;
assign s324 = 1'b0;
assign s325 = 1'b0;
assign s326 = 1'b0;
assign s327 = 1'b0;
assign s328 = 1'b0;
assign src2_sel_imm = s303 | s277 | s290 | s307 | s306 | s302 | s301 | s20 | s241 | s5 | s75 | s166 | s77 | s127 | s178 | s177 | s170 | s169 | s79 | s129 | s182 | s181 | s174 | s173;
assign src3_sel_imm = s197 | s121 | s195 | s119 | s196 | s120;
assign src4_sel_imm = s197 | s121 | s195 | s119 | s196 | s120;
assign src2_imm = s329;
assign src3_imm = ({32{s331}} & s335) | ({32{s330}} & s333);
assign src4_imm = ({32{s331}} & s336) | ({32{s330}} & s334);
assign operand_ctrl[0] = s1 | s108 | s230 | s25 | s203 | s186 | s116 | s238 | s89 | s214 | s183 | s113 | s235 | s86 | s211 | s184 | s114 | s236 | s87 | s212 | s171 | s173 | s172 | s174 | s179 | s181 | s180 | s182 | s128 | s129 | s78 | s79 | s82 | s83 | s17 | s125 | s201 | s123 | s199 | s151 | s223 | s143 | s221 | s22 | s39 | s194 | s14 | s11 | s8;
assign operand_ctrl[1] = s18 | s111 | s233 | s29 | s207 | s19 | s112 | s234 | s30 | s208 | s40;
assign operand_ctrl[2] = s120 | s196;
assign operand_ctrl[3] = s0 | s107 | s229 | s24 | s202 | s185 | s115 | s237 | s88 | s213 | s167 | s169 | s168 | s170 | s175 | s177 | s176 | s178 | s126 | s127 | s76 | s77 | s80 | s81 | s16 | s124 | s200 | s122 | s198 | s150 | s222 | s142 | s220 | s21 | s37 | s193 | s13 | s10 | s7 | s188 | s189 | s190 | s191 | s192 | s243 | s244 | s245 | s246 | s247;
assign operand_ctrl[4] = s119 | s195;
assign operand_ctrl[5] = s38;
assign operand_ctrl[6] = s110 | s232 | s118 | s240 | s97 | s96 | s23 | s15 | s12 | s9 | s152 | s153 | s55 | s56 | s65 | s66 | s93 | s94 | s95 | s98 | s99 | s100 | s269 | s295 | s267 | s271 | s274;
assign operand_ctrl[7] = s165 | s166 | s74 | s75 | s4 | s5 | s6 | s20;
assign operand_ctrl[8] = s103 | s144 | s44;
assign operand_ctrl[9] = s104 | s145 | s45;
assign operand_ctrl[10] = s106;
assign operand_ctrl[11] = s105 | s146 | s46;
assign operand_ctrl[12] = s121 | s197;
assign operand_ctrl[13] = s242 | s241;
assign operand_ctrl[14] = s154 | s155 | s57 | s58 | s67 | s68 | s59 | s60;
assign operand_ctrl[15] = s156 | s157 | s61 | s62 | s69 | s70 | s63 | s64;
assign operand_ctrl[16] = s53 | s147 | s47 | s49 | s71 | s163 | s227;
assign operand_ctrl[17] = s54 | s149 | s48 | s51 | s72 | s164 | s228;
assign operand_ctrl[18] = s148 | s50;
assign operand_ctrl[19] = s130;
assign operand_ctrl[20] = s140 | s219 | s141 | s101 | s102 | s161 | s225;
assign operand_ctrl[21] = s162 | s226;
assign operand_ctrl[22] = s2 | s109 | s231 | s26 | s204 | s187 | s117 | s239 | s90 | s215 | s139 | s218 | s52 | s209 | s160 | s224 | s73 | s210;
assign operand_ctrl[23] = s131;
assign operand_ctrl[24] = s132;
assign operand_ctrl[25] = s133;
assign operand_ctrl[26] = s134 | s136 | s158;
assign operand_ctrl[27] = s135 | s138 | s159;
assign operand_ctrl[28] = s137;
assign operand_ctrl[29] = s27 | s91 | s28 | s92;
assign operand_ctrl[30] = s205 | s216 | s206 | s217;
assign operand_ctrl[31] = s41 | s31 | s34 | s261 | s255 | s258;
assign operand_ctrl[32] = s42 | s32 | s35 | s262 | s256 | s259;
assign operand_ctrl[33] = s43 | s33 | s36 | s263 | s257 | s260;
assign operand_ctrl[34] = s84 | s85 | s303;
assign operand_ctrl[35] = s3;
assign operand_ctrl[36] = s248 | s283 | s319 | s252 | s311 | s310 | s288 | s324 | s282 | s316 | s308 | s286 | s322 | s280 | s314 | s309 | s287 | s323 | s281 | s315 | s299 | s301 | s300 | s302 | s304 | s306 | s305 | s307 | s289 | s290 | s276 | s277 | s278 | s279 | s298 | s318 | s291 | s317 | s251;
assign operand_ctrl[37] = s249 | s284 | s320 | s253 | s312 | s250 | s285 | s321 | s254 | s313;
assign operand_ctrl[38] = s292 | s264 | s325;
assign operand_ctrl[39] = s293 | s265 | s326;
assign operand_ctrl[40] = s294 | s266 | s327;
assign operand_ctrl[41] = s270 | s297 | s268 | s273 | s275;
assign operand_ctrl[42] = s296 | s272;
assign operand_ctrl[43] = s328;
assign function_ctrl[0] = s1 | s108 | s25;
assign function_ctrl[1] = s230 | s203;
assign function_ctrl[2] = s186 | s116 | s89;
assign function_ctrl[3] = s238 | s214;
assign function_ctrl[4] = s183 | s113 | s86 | s18 | s111 | s29;
assign function_ctrl[5] = s235 | s211 | s233 | s207;
assign function_ctrl[6] = s184 | s114 | s87 | s19 | s112 | s30;
assign function_ctrl[7] = s236 | s212 | s234 | s208;
assign function_ctrl[8] = s171 | s173 | s172 | s174;
assign function_ctrl[9] = s179 | s181 | s180 | s182;
assign function_ctrl[10] = s128 | s129 | s78 | s79;
assign function_ctrl[11] = s82 | s83;
assign function_ctrl[12] = s17;
assign function_ctrl[13] = s125;
assign function_ctrl[14] = s201;
assign function_ctrl[15] = s123;
assign function_ctrl[16] = s199;
assign function_ctrl[17] = s151;
assign function_ctrl[18] = s223;
assign function_ctrl[19] = s143;
assign function_ctrl[20] = s221;
assign function_ctrl[21] = s22;
assign function_ctrl[22] = s120 | s196;
assign function_ctrl[23] = s39 | s40;
assign function_ctrl[24] = s194;
assign function_ctrl[25] = s14;
assign function_ctrl[26] = s11;
assign function_ctrl[27] = s8;
assign function_ctrl[28] = s0 | s107 | s24;
assign function_ctrl[29] = s229 | s202;
assign function_ctrl[30] = s185 | s115 | s88;
assign function_ctrl[31] = s237 | s213;
assign function_ctrl[32] = s167 | s169 | s168 | s170;
assign function_ctrl[33] = s175 | s177 | s176 | s178;
assign function_ctrl[34] = s126 | s127 | s76 | s77;
assign function_ctrl[35] = s80 | s81;
assign function_ctrl[36] = s16;
assign function_ctrl[37] = s124;
assign function_ctrl[38] = s200;
assign function_ctrl[39] = s122;
assign function_ctrl[40] = s198;
assign function_ctrl[41] = s150;
assign function_ctrl[42] = s222;
assign function_ctrl[43] = s142;
assign function_ctrl[44] = s220;
assign function_ctrl[45] = s21;
assign function_ctrl[46] = s119 | s195;
assign function_ctrl[47] = s37 | s38;
assign function_ctrl[48] = s193;
assign function_ctrl[49] = s13;
assign function_ctrl[50] = s10;
assign function_ctrl[51] = s7;
assign function_ctrl[52] = s188 | s243;
assign function_ctrl[53] = s189 | s244;
assign function_ctrl[54] = s190 | s245;
assign function_ctrl[55] = s191 | s246;
assign function_ctrl[56] = s192 | s247;
assign function_ctrl[57] = s110;
assign function_ctrl[58] = s232;
assign function_ctrl[59] = s118;
assign function_ctrl[60] = s240;
assign function_ctrl[61] = s165 | s166;
assign function_ctrl[62] = s74 | s75;
assign function_ctrl[63] = s103 | s104 | s106 | s105;
assign function_ctrl[64] = s121 | s197;
assign function_ctrl[65] = s4 | s5;
assign function_ctrl[66] = s242 | s241;
assign function_ctrl[67] = s6;
assign function_ctrl[68] = s20;
assign function_ctrl[69] = s97;
assign function_ctrl[70] = s96;
assign function_ctrl[71] = s23;
assign function_ctrl[72] = s15;
assign function_ctrl[73] = s12;
assign function_ctrl[74] = s9;
assign function_ctrl[75] = s152 | s153 | s292 | s293 | s294;
assign function_ctrl[76] = s55 | s56 | s269 | s270;
assign function_ctrl[77] = s65 | s66 | s295 | s297 | s296;
assign function_ctrl[78] = s93 | s94 | s264 | s265 | s266;
assign function_ctrl[79] = s95 | s267 | s268;
assign function_ctrl[80] = s98 | s271 | s273 | s272;
assign function_ctrl[81] = s154 | s155 | s156 | s157;
assign function_ctrl[82] = s57 | s58 | s61 | s62;
assign function_ctrl[83] = s67 | s68 | s69 | s70;
assign function_ctrl[84] = s59 | s60 | s63 | s64;
assign function_ctrl[85] = s144 | s145 | s146;
assign function_ctrl[86] = s53 | s54;
assign function_ctrl[87] = s147 | s149 | s148;
assign function_ctrl[88] = s44 | s45 | s46;
assign function_ctrl[89] = s47 | s48;
assign function_ctrl[90] = s49 | s51 | s50;
assign function_ctrl[91] = s71 | s72;
assign function_ctrl[92] = s130;
assign function_ctrl[93] = s140;
assign function_ctrl[94] = s219;
assign function_ctrl[95] = s141;
assign function_ctrl[96] = s101;
assign function_ctrl[97] = s102;
assign function_ctrl[98] = s163 | s164;
assign function_ctrl[99] = s227 | s228;
assign function_ctrl[100] = s161 | s162;
assign function_ctrl[101] = s225 | s226;
assign function_ctrl[102] = s99;
assign function_ctrl[103] = s100;
assign function_ctrl[104] = s2 | s109 | s26;
assign function_ctrl[105] = s231 | s204;
assign function_ctrl[106] = s187 | s117 | s90;
assign function_ctrl[107] = s239 | s215;
assign function_ctrl[108] = s139 | s52;
assign function_ctrl[109] = s218 | s209;
assign function_ctrl[110] = s160 | s73;
assign function_ctrl[111] = s224 | s210;
assign function_ctrl[112] = s131 | s132 | s133;
assign function_ctrl[113] = s134 | s135;
assign function_ctrl[114] = s136 | s138 | s137;
assign function_ctrl[115] = s158 | s159;
assign function_ctrl[116] = s27 | s28;
assign function_ctrl[117] = s205 | s206;
assign function_ctrl[118] = s91 | s92;
assign function_ctrl[119] = s216 | s217;
assign function_ctrl[120] = s41 | s42 | s43 | s261 | s262 | s263;
assign function_ctrl[121] = s31 | s32 | s33 | s255 | s256 | s257;
assign function_ctrl[122] = s84 | s85;
assign function_ctrl[123] = s34 | s35 | s36 | s258 | s259 | s260;
assign function_ctrl[124] = s3;
assign function_ctrl[125] = s248 | s283 | s252;
assign function_ctrl[126] = s319 | s311;
assign function_ctrl[127] = s310 | s288 | s282;
assign function_ctrl[128] = s324 | s316;
assign function_ctrl[129] = s308 | s286 | s280 | s249 | s284 | s253;
assign function_ctrl[130] = s322 | s314 | s320 | s312;
assign function_ctrl[131] = s309 | s287 | s281 | s250 | s285 | s254;
assign function_ctrl[132] = s323 | s315 | s321 | s313;
assign function_ctrl[133] = s299 | s301 | s300 | s302;
assign function_ctrl[134] = s304 | s306 | s305 | s307;
assign function_ctrl[135] = s289 | s290 | s276 | s277;
assign function_ctrl[136] = s278 | s279;
assign function_ctrl[137] = s298;
assign function_ctrl[138] = s318;
assign function_ctrl[139] = s291;
assign function_ctrl[140] = s317;
assign function_ctrl[141] = s251;
assign function_ctrl[142] = s303;
assign function_ctrl[143] = s292 | s293 | s294;
assign function_ctrl[144] = s269 | s270;
assign function_ctrl[145] = s295 | s297 | s296;
assign function_ctrl[146] = s264 | s265 | s266;
assign function_ctrl[147] = s267 | s268;
assign function_ctrl[148] = s271 | s273 | s272;
assign function_ctrl[149] = s274 | s275;
assign function_ctrl[150] = s325 | s326 | s328 | s327;
assign result_ctrl[0] = s1 | s186 | s183 | s184 | s18 | s19;
assign result_ctrl[1] = s108 | s116 | s113 | s114 | s111 | s112;
assign result_ctrl[2] = s230 | s238 | s235 | s236 | s233 | s234;
assign result_ctrl[3] = s25 | s89 | s86 | s87 | s29 | s30 | s78 | s79 | s82 | s22 | s39 | s40;
assign result_ctrl[4] = s203 | s214 | s211 | s212 | s207 | s208;
assign result_ctrl[5] = s171 | s173 | s179 | s181 | s128 | s129;
assign result_ctrl[6] = s172 | s174 | s180 | s182;
assign result_ctrl[7] = s83;
assign result_ctrl[8] = s17 | s125 | s201 | s123 | s199;
assign result_ctrl[9] = s151 | s223 | s143 | s221;
assign result_ctrl[10] = s120 | s196;
assign result_ctrl[11] = s194;
assign result_ctrl[12] = s14 | s11 | s8;
assign result_ctrl[13] = s0 | s185;
assign result_ctrl[14] = s107 | s115;
assign result_ctrl[15] = s229 | s237;
assign result_ctrl[16] = s24 | s88 | s76 | s77 | s80 | s21 | s37 | s38;
assign result_ctrl[17] = s202 | s213;
assign result_ctrl[18] = s167 | s169 | s175 | s177 | s126 | s127;
assign result_ctrl[19] = s168 | s170 | s176 | s178;
assign result_ctrl[20] = s81;
assign result_ctrl[21] = s16 | s124 | s200 | s122 | s198;
assign result_ctrl[22] = s150 | s222 | s142 | s220;
assign result_ctrl[23] = s119 | s195;
assign result_ctrl[24] = s193;
assign result_ctrl[25] = s13 | s10 | s7;
assign result_ctrl[26] = s188 | s189 | s190 | s191 | s192;
assign result_ctrl[27] = s243 | s244 | s245 | s246 | s247;
assign result_ctrl[28] = s110 | s118;
assign result_ctrl[29] = s232 | s240;
assign result_ctrl[30] = s165 | s166;
assign result_ctrl[31] = s74 | s75 | s23;
assign result_ctrl[32] = s103 | s104 | s106 | s105;
assign result_ctrl[33] = s121 | s197;
assign result_ctrl[34] = s4 | s5 | s101 | s102;
assign result_ctrl[35] = s242 | s241 | s95 | s98;
assign result_ctrl[36] = s6;
assign result_ctrl[37] = s20;
assign result_ctrl[38] = s97 | s96;
assign result_ctrl[39] = s15 | s12 | s9;
assign result_ctrl[40] = s152 | s154 | s156 | s299 | s301 | s304 | s306 | s289 | s290;
assign result_ctrl[41] = s153 | s155 | s157 | s300 | s302 | s305 | s307;
assign result_ctrl[42] = s55 | s65 | s93 | s57 | s61 | s67 | s69 | s59 | s63 | s252 | s282 | s280 | s281 | s253 | s254 | s276 | s277 | s278 | s251;
assign result_ctrl[43] = s56 | s66 | s94 | s58 | s62 | s68 | s70 | s60 | s64;
assign result_ctrl[44] = s144 | s145 | s146 | s147 | s149 | s148 | s140 | s219 | s141;
assign result_ctrl[45] = s53 | s54 | s44 | s45 | s46 | s47 | s48 | s49 | s51 | s50 | s71 | s72;
assign result_ctrl[46] = s130 | s163 | s164 | s227 | s228 | s161 | s162 | s225 | s226 | s99 | s100 | s292 | s293 | s294 | s295 | s297 | s296;
assign result_ctrl[47] = s2 | s187;
assign result_ctrl[48] = s109 | s117;
assign result_ctrl[49] = s231 | s239;
assign result_ctrl[50] = s26 | s90 | s52 | s73;
assign result_ctrl[51] = s204 | s215 | s209 | s210;
assign result_ctrl[52] = s139 | s218 | s160 | s224 | s131 | s132 | s133 | s134 | s135 | s136 | s138 | s137 | s158 | s159;
assign result_ctrl[53] = s27 | s91 | s41 | s42 | s43;
assign result_ctrl[54] = s205 | s216;
assign result_ctrl[55] = s28 | s92 | s31 | s32 | s33 | s34 | s35 | s36 | s84;
assign result_ctrl[56] = s206 | s217;
assign result_ctrl[57] = s85;
assign result_ctrl[58] = s3;
assign result_ctrl[59] = s248 | s310 | s308 | s309 | s249 | s250;
assign result_ctrl[60] = s283 | s288 | s286 | s287 | s284 | s285;
assign result_ctrl[61] = s319 | s324 | s322 | s323 | s320 | s321;
assign result_ctrl[62] = s311 | s316 | s314 | s315 | s312 | s313;
assign result_ctrl[63] = s279;
assign result_ctrl[64] = s298 | s318 | s291 | s317;
assign result_ctrl[65] = s303;
assign result_ctrl[66] = s269 | s270 | s264 | s265 | s266 | s267 | s268 | s271 | s273 | s272 | s274 | s275;
assign result_ctrl[67] = s261 | s262 | s263;
assign result_ctrl[68] = s255 | s256 | s257 | s258 | s259 | s260;
assign result_ctrl[69] = s325 | s326 | s328 | s327;
assign overflow_ctrl = s25 | s203 | s89 | s214 | s86 | s211 | s87 | s212 | s29 | s207 | s30 | s208 | s78 | s79 | s82 | s83 | s22 | s120 | s196 | s39 | s40 | s24 | s202 | s88 | s213 | s76 | s77 | s80 | s81 | s21 | s119 | s195 | s37 | s38 | s74 | s75 | s121 | s197 | s23 | s55 | s56 | s65 | s66 | s93 | s94 | s95 | s98 | s57 | s58 | s61 | s62 | s67 | s68 | s69 | s70 | s59 | s60 | s63 | s64 | s53 | s54 | s44 | s45 | s46 | s47 | s48 | s49 | s51 | s50 | s71 | s72 | s26 | s204 | s90 | s215 | s52 | s209 | s73 | s210 | s27 | s205 | s91 | s216 | s41 | s42 | s43 | s28 | s206 | s92 | s217 | s31 | s32 | s33 | s84 | s85 | s34 | s35 | s36 | s252 | s311 | s282 | s316 | s280 | s314 | s281 | s315 | s253 | s312 | s254 | s313 | s276 | s277 | s278 | s279 | s251 | s269 | s270 | s264 | s265 | s266 | s267 | s268 | s271 | s273 | s272 | s274 | s275 | s261 | s262 | s263 | s255 | s256 | s257 | s258 | s259 | s260;
assign s329 = {{26{1'b0}},instr[25:20]};
assign s330 = s121 | s119 | s120;
assign s331 = s197 | s195 | s196;
assign s332 = ({5{(s121 | s197)}} & instr[24:20]) | ({5{(s120 | s196)}} & {1'd0,instr[23:20]}) | ({5{(s119 | s195)}} & {2'd0,instr[22:20]});
assign s333 = {32{1'b1}} << s332;
assign s334 = ~s333;
assign s335 = {32{1'b0}};
assign s336 = s334;
endmodule

