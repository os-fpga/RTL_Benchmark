-----------------------------------------------------------------------
----                                                               ----
---- Montgomery modular multiplier and exponentiator               ----
----                                                               ----
---- This file is part of the Montgomery modular multiplier        ----
---- and exponentiator project                                     ----
---- http://opencores.org/project,mod_mult_exp                     ----
----                                                               ----
---- Description:                                                  ----
----   This module is example implementation of the Montgomery     ----
----   modular exponentiator combined with the RS-232 communication----
----   with PC. All related to the communication logic was         ----
----   inclueded here. Input data are retrieved by serial input    ----
----   and converted into parallel data by the shift registers     ----
----   After exponentiation in similar way parallel data are       ----
----   converted into serial data. For the communication, the      ----
----   RS232RefComp module made by Digilent was used and slightly  ----
----   modified (increased data transfer speed to 115 200 bps).    ----
----                                                               ----
---- To Do:                                                        ----
----                                                               ----
---- Author(s):                                                    ----
---- - Krzysztof Gajewski, gajos@opencores.org                     ----
----                       k.gajewski@gmail.com                    ----
----                                                               ----
-----------------------------------------------------------------------
----                                                               ----
---- Copyright (C) 2019 Authors and OPENCORES.ORG                  ----
----                                                               ----
---- This source file may be used and distributed without          ----
---- restriction provided that this copyright statement is not     ----
---- removed from the file and that any derivative work contains   ----
---- the original copyright notice and the associated disclaimer.  ----
----                                                               ----
---- This source file is free software; you can redistribute it    ----
---- and-or modify it under the terms of the GNU Lesser General    ----
---- Public License as published by the Free Software Foundation;  ----
---- either version 2.1 of the License, or (at your option) any    ----
---- later version.                                                ----
----                                                               ----
---- This source is distributed in the hope that it will be        ----
---- useful, but WITHOUT ANY WARRANTY; without even the implied    ----
---- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR       ----
---- PURPOSE. See the GNU Lesser General Public License for more   ----
---- details.                                                      ----
----                                                               ----
---- You should have received a copy of the GNU Lesser General     ----
---- Public License along with this source; if not, download it    ----
---- from http://www.opencores.org/lgpl.shtml                      ----
----                                                               ----
-----------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.properties.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

-- Definition of the component
entity ModExpComm is
    generic (word_size : integer := WORD_LENGTH);
    port (
	     DATA_RXD : in  STD_LOGIC;
		  CLK      : in  STD_LOGIC;
		  RESET    : in  STD_LOGIC;
		  DATA_TXD : out STD_LOGIC
	 );
end ModExpComm;

architecture Behavioral of ModExpComm is

-- This is DCM component generated by the ISE. It was used due
-- to maximum clock speed available in the S3EBOARD served by
-- the Digilent (50 MHz) it is used in order to decrease speed
-- of exponentiator core. RS232 is working with 50 MHz and the
-- rest part of the core is working with 10 MHz. This is due
-- to timing estimation of ISE. 
component dcms is
    port ( 
	     CLKIN_IN  : in  STD_LOGIC; 
        CLKDV_OUT : out STD_LOGIC; 
        CLK0_OUT  : out STD_LOGIC
	 );
end component dcms;

-- Montgomery modular exponentiator
component ModExp is
	 generic (
        word_size   : integer := WORD_LENGTH;
        word_binary : integer := WORD_INTEGER
	 );
    Port ( 
        input         : in  STD_LOGIC_VECTOR(word_size - 1 downto 0);
        ctrl          : in  STD_LOGIC_VECTOR(2 downto 0);
        clk           : in  STD_LOGIC;
        reset         : in  STD_LOGIC;
        data_in_ready : in  STD_LOGIC;
        ready         : out STD_LOGIC;
        output        : out STD_LOGIC_VECTOR(word_size - 1 downto 0)
    );
end component ModExp;

-- RS232 component made by the Digilent
-- all checking was ignored but for communication
-- odd parity is used
component Rs232RefComp is
    port ( 
	     TXD   : out   STD_LOGIC  	:= '1';
    	  RXD   : in    STD_LOGIC;					
    	  CLK   : in    STD_LOGIC;							  --Master Clock
		  DBIN  : in    STD_LOGIC_VECTOR(7 downto 0); --Data Bus in
		  DBOUT : out   STD_LOGIC_VECTOR(7 downto 0); --Data Bus out
		  RDA	  : inout STD_LOGIC;						     --Read Data Available
		  TBE	  : inout STD_LOGIC 	:= '1';			     --Transfer Bus Empty
		  RD	  : in    STD_LOGIC;					        --Read Strobe
		  WR	  : in    STD_LOGIC;					        --Write Strobe
		  PE	  : out   STD_LOGIC;					        --Parity Error Flag
		  FE	  : out   STD_LOGIC;				           --Frame Error Flag
		  OE	  : out   STD_LOGIC;					        --Overwrite Error Flag
		  RST   : in    STD_LOGIC	   := '0'	        --Master Reset
    );
end component Rs232RefComp;

-- Register for storing control word for ModExpComm component
component Reg is
    generic(word_size : integer := 8);
	 port(
	     input  : in  STD_LOGIC_VECTOR(word_size - 1 downto 0);
		  output : out STD_LOGIC_VECTOR(word_size - 1 downto 0);
		  enable : in  STD_LOGIC;
		  clk    : in  STD_LOGIC;
		  reset  : in  STD_LOGIC
    );
end component Reg;

---- Shift registers for input and output data for the modular exponentiator 
component ShiftReg is
    generic (
	     length_1      : integer :=  BYTE;
	     length_2      : integer :=  WORD_LENGTH;
		  internal_data : integer :=  WORD_LENGTH
	 );
    port ( 
	     input  : in  STD_LOGIC_VECTOR(length_1 - 1 downto 0);
        output : out STD_LOGIC_VECTOR(length_2 - 1 downto 0);
        en     : in  STD_LOGIC;
        shift  : in  STD_LOGIC;
        clk    : in  STD_LOGIC;
        reset  : in  STD_LOGIC
	 );
end component ShiftReg;

---- some 'help' mux  at the output of the component
component AsyncMux is
    generic(
	     word_size : integer := WORD_LENGTH
	 );
    port(
	     input0 : in  STD_LOGIC_VECTOR(word_size downto 0);
	     input1 : in  STD_LOGIC_VECTOR(word_size downto 0);
		  ctrl   : in  STD_LOGIC;
		  output : out STD_LOGIC_VECTOR(word_size downto 0)
    );
end component AsyncMux;

---- State machine
component ModExpDataCtrlSM is
    port(
        clk                : in  STD_LOGIC;
		  reset              : in  STD_LOGIC;
        RDAsig             : in  STD_LOGIC;
        TBEsig             : in  STD_LOGIC;
        RDsig              : out STD_LOGIC;
        WRsig              : out STD_LOGIC;
		  data_in_ready      : out STD_LOGIC;
        readySig           : in  STD_LOGIC;
        modExpCtrlRegEn    : out STD_LOGIC;
        dataToModExpEn     : out STD_LOGIC;
        dataToModExpShift     : out STD_LOGIC;
        dataFromModExpEn      : out STD_LOGIC;
        dataFromModExpShift   : out STD_LOGIC;
        muxCtrl            : out STD_LOGIC;
		  opcodes            : in  STD_LOGIC_VECTOR(2 downto 0);
        controlStateOut    : out STD_LOGIC_VECTOR(2 downto 0)
);
end component ModExpDataCtrlSM;

-- All signals needed in the implementation
signal clk_div : STD_LOGIC;
signal clk_0   : STD_LOGIC;

signal dataTXD : STD_LOGIC_VECTOR(7 downto 0);
signal dataRXD : STD_LOGIC_VECTOR(7 downto 0);
signal RDAsig  : STD_LOGIC;
signal TBEsig  : STD_LOGIC;
signal RDsig   : STD_LOGIC;
signal WRsig   : STD_LOGIC;
signal PEsig   : STD_LOGIC;
signal FEsig   : STD_LOGIC;
signal OEsig   : STD_LOGIC;

signal modExpInput     : STD_LOGIC_VECTOR(word_size - 1 downto 0);
signal modExpCtrl      : STD_LOGIC_VECTOR(2 downto 0);
signal modExpCtrlRegEn : STD_LOGIC;
signal data_in_ready   : STD_LOGIC;
signal readySig        : STD_LOGIC;
signal modExpOutput    : STD_LOGIC_VECTOR(word_size - 1 downto 0);

signal dataToModExpEn    : STD_LOGIC;
signal dataToModExpShift : STD_LOGIC;

signal dataFromModExpEn    : STD_LOGIC;
signal dataFromModExpShift : STD_LOGIC;

signal inputToMux       : STD_LOGIC_VECTOR(BYTE - 1 downto 0);
signal controlStateOut  : STD_LOGIC_VECTOR(2 downto 0);
signal muxCtrl          : STD_LOGIC;

signal ctrl_zero            : STD_LOGIC_VECTOR(4 downto 0) := "00000";
signal control_state_to_out : STD_LOGIC_VECTOR(7 downto 0);
		
begin
-- Architecture definition
	 ctrl_zero <= (others => '0');
	 control_state_to_out <= controlStateOut & ctrl_zero;
	 
	 -- DCM
	 dcm_module : dcms 
	     port map( 
	         CLKIN_IN  => CLK,
            CLKDV_OUT => clk_div, --clk_null,
            CLK0_OUT  => clk_0
	     );
	 
	 -- RS232 component
    serialPort : Rs232RefComp 
	     port map ( 
		      TXD   => DATA_TXD,
    	      RXD   => DATA_RXD,
    	      CLK   => clk_0,
		      DBIN  => dataTXD,
		      DBOUT => dataRXD,
		      RDA   => RDAsig, --Read Data Available
		      TBE   => TBEsig, --Transfer Bus Empty
		      RD	   => RDsig,  --Read Strobe
		      WR    => WRsig,  --Write Strobe
		      PE	   => PEsig,  --Parity Error Flag
		      FE	   => FEsig,  --Frame Error Flag
		      OE    => OEsig,  --Overwrite Error Flag
		      RST   => RESET   --Master Reset
        );
	 
	 -- Shift register at input of the modular exponentiator
	 -- (convert data from 8 bit to 32 bit, 64 bit, 512 bit, etc.)
	 modExpCompIn : ShiftReg 
	     generic map(
	         length_1      => BYTE, 
				length_2      => WORD_LENGTH, 
				internal_data => WORD_LENGTH
		  )
        port map ( 
	         input  => dataRXD,
            output => modExpInput,
            en     => dataToModExpEn,
            shift  => dataToModExpShift,
            clk    => CLK_div,
            reset  => RESET
	     );
	 
	 -- Control register
	 modCtrl : Reg
        generic map(
				word_size => 3
		  )	 
	     port map (
	         input  => dataRXD(2 downto 0),
		      output => modExpCtrl,
		      enable => modExpCtrlRegEn,
		      clk    => CLK_div,
		      reset  => RESET
        );

	 -- Modular exponentiator component
	 ModExpComp : ModExp 
	     port map ( 
		      input         => modExpInput,
		      ctrl          => modExpCtrl,
		      clk           => CLK_div,
		      reset         => RESET,
		      data_in_ready => data_in_ready,
		      ready         => readySig,
		      output        => modExpOutput
	     );	 
	 
	 -- Shift register at output of the modular exponentiator
	 -- (convert data from 32 bit, 64 bit, 512 bit, etc. to 8 bit)
	 dataFromModExpComponent : ShiftReg 
	     generic map(
	         length_1      => WORD_LENGTH, 
				length_2      => BYTE, 
				internal_data => WORD_LENGTH
		  )
        port map ( 
            input  => modExpOutput,
				output => inputToMux,
            en     => dataFromModExpEn,
            shift  => dataFromModExpShift,
            clk    => CLK_div,
            reset  => RESET
	     );
    
	 -- Multiplexer at the output of the component
    outMux : AsyncMux
        generic map(
		      word_size => BYTE - 1
		  )
        port map(
	         input0 => inputToMux,
	         input1 => control_state_to_out,
	         ctrl   => muxCtrl,
	         output => dataTXD
        );

    -- State machine
    stateMachine : ModExpDataCtrlSM 
	     port map(
	         clk                 => CLK_div,
		      reset               => RESET,
            RDAsig              => RDAsig,
            TBEsig              => TBEsig,
            RDsig               => RDsig,
            WRsig               => WRsig,
		      data_in_ready       => data_in_ready,
            readySig            => readySig,
            modExpCtrlRegEn     => modExpCtrlRegEn,
            dataToModExpEn      => dataToModExpEn,
            dataToModExpShift   => dataToModExpShift,
            dataFromModExpEn    => dataFromModExpEn,
            dataFromModExpShift => dataFromModExpShift,
            muxCtrl             => muxCtrl,
		      opcodes             => dataRXD(2 downto 0),
            controlStateOut     => controlStateOut
        );

end Behavioral;