library ieee;
use ieee.std_logic_1164.all;

entity top is
port( a: in std_logic_vector(127 downto 0);
asqrt: out std_logic_vector(63 downto 0));
end top;

ARCHITECTURE Behavioral of top is

signal one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617: std_logic;

begin

w0 <= not a(126) and not a(127);
w1 <= a(126) and a(127);
w2 <= a(126) and not w0;
w3 <= not a(124) and not a(125);
w4 <= not w2 and not w3;
w5 <= not w1 and not w4;
w6 <= a(124) and not w5;
w7 <= not a(122) and not a(123);
w8 <= not a(124) and w7;
w9 <= not w6 and not w8;
w10 <= not a(124) and not w5;
w11 <= a(125) and not w10;
w12 <= w3 and not w5;
w13 <= not w11 and not w12;
w14 <= not w9 and w13;
w15 <= w0 and not w14;
w16 <= w9 and not w13;
w17 <= a(126) and w3;
w18 <= not a(126) and not w3;
w19 <= a(127) and not w18;
w20 <= not w17 and w19;
w21 <= not w16 and not w20;
w22 <= not w15 and w21;
w23 <= a(122) and not w22;
w24 <= not a(120) and not a(121);
w25 <= not a(122) and w24;
w26 <= not w23 and not w25;
w27 <= not w5 and not w26;
w28 <= not w1 and not w25;
w29 <= not w4 and w28;
w30 <= not w23 and w29;
w31 <= w7 and not w22;
w32 <= not a(122) and not w22;
w33 <= a(123) and not w32;
w34 <= not w31 and not w33;
w35 <= not w30 and w34;
w36 <= not w27 and not w35;
w37 <= not w5 and not w20;
w38 <= not w16 and w37;
w39 <= not w15 and w38;
w40 <= not w31 and not w39;
w41 <= a(124) and not w40;
w42 <= not a(124) and not w39;
w43 <= not w31 and w42;
w44 <= not w41 and not w43;
w45 <= w14 and not w22;
w46 <= not w16 and not w45;
w47 <= not w44 and w46;
w48 <= not w36 and w47;
w49 <= w0 and not w48;
w50 <= w36 and w44;
w51 <= w13 and not w22;
w52 <= w9 and not w51;
w53 <= not w0 and not w14;
w54 <= not w52 and w53;
w55 <= not w13 and not w20;
w56 <= not w16 and w55;
w57 <= not w15 and w56;
w58 <= not w54 and not w57;
w59 <= not w50 and w58;
w60 <= not w49 and w59;
w61 <= a(120) and not w60;
w62 <= not a(118) and not a(119);
w63 <= not a(120) and w62;
w64 <= not w61 and not w63;
w65 <= not w22 and not w64;
w66 <= not a(120) and not w60;
w67 <= a(121) and not w66;
w68 <= w24 and not w60;
w69 <= not w67 and not w68;
w70 <= not w20 and not w63;
w71 <= not w16 and w70;
w72 <= not w15 and w71;
w73 <= not w61 and w72;
w74 <= w69 and not w73;
w75 <= not w65 and not w74;
w76 <= not w5 and not w75;
w77 <= w5 and not w65;
w78 <= not w74 and w77;
w79 <= not w22 and not w57;
w80 <= not w54 and w79;
w81 <= not w50 and w80;
w82 <= not w49 and w81;
w83 <= not w68 and not w82;
w84 <= a(122) and not w83;
w85 <= not a(122) and not w82;
w86 <= not w68 and w85;
w87 <= not w84 and not w86;
w88 <= not w78 and not w87;
w89 <= not w76 and not w88;
w90 <= not w27 and not w30;
w91 <= not w34 and w90;
w92 <= not w60 and w91;
w93 <= not w60 and w90;
w94 <= w34 and not w93;
w95 <= not w92 and not w94;
w96 <= not w36 and not w44;
w97 <= not w60 and w96;
w98 <= not w50 and not w97;
w99 <= not w95 and w98;
w100 <= not w89 and w99;
w101 <= w0 and not w100;
w102 <= not w76 and w95;
w103 <= not w88 and w102;
w104 <= w36 and not w60;
w105 <= not w44 and not w104;
w106 <= not w0 and not w50;
w107 <= not w105 and w106;
w108 <= not w43 and not w57;
w109 <= not w41 and w108;
w110 <= not w54 and w109;
w111 <= not w50 and w110;
w112 <= not w49 and w111;
w113 <= not w107 and not w112;
w114 <= not w103 and w113;
w115 <= not w101 and w114;
w116 <= a(118) and not w115;
w117 <= not a(116) and not a(117);
w118 <= not a(118) and w117;
w119 <= not w116 and not w118;
w120 <= not w60 and not w119;
w121 <= not w57 and not w118;
w122 <= not w54 and w121;
w123 <= not w50 and w122;
w124 <= not w49 and w123;
w125 <= not w116 and w124;
w126 <= not a(118) and not w115;
w127 <= a(119) and not w126;
w128 <= w62 and not w115;
w129 <= not w127 and not w128;
w130 <= not w125 and w129;
w131 <= not w120 and not w130;
w132 <= not w22 and not w131;
w133 <= w22 and not w120;
w134 <= not w130 and w133;
w135 <= not w60 and not w112;
w136 <= not w107 and w135;
w137 <= not w103 and w136;
w138 <= not w101 and w137;
w139 <= not w128 and not w138;
w140 <= a(120) and not w139;
w141 <= not a(120) and not w138;
w142 <= not w128 and w141;
w143 <= not w140 and not w142;
w144 <= not w134 and not w143;
w145 <= not w132 and not w144;
w146 <= not w5 and not w145;
w147 <= w5 and not w132;
w148 <= not w144 and w147;
w149 <= not w69 and not w73;
w150 <= not w65 and w149;
w151 <= not w115 and w150;
w152 <= not w65 and not w73;
w153 <= not w115 and w152;
w154 <= w69 and not w153;
w155 <= not w151 and not w154;
w156 <= not w148 and not w155;
w157 <= not w146 and not w156;
w158 <= not w78 and w87;
w159 <= not w76 and w158;
w160 <= not w115 and w159;
w161 <= not w76 and not w78;
w162 <= not w115 and w161;
w163 <= not w87 and not w162;
w164 <= not w160 and not w163;
w165 <= not w89 and not w95;
w166 <= not w115 and w165;
w167 <= not w103 and not w166;
w168 <= not w164 and w167;
w169 <= not w157 and w168;
w170 <= w0 and not w169;
w171 <= not w146 and w164;
w172 <= not w156 and w171;
w173 <= w89 and not w115;
w174 <= not w95 and not w173;
w175 <= not w0 and not w103;
w176 <= not w174 and w175;
w177 <= not w92 and not w112;
w178 <= not w94 and w177;
w179 <= not w107 and w178;
w180 <= not w103 and w179;
w181 <= not w101 and w180;
w182 <= not w176 and not w181;
w183 <= not w172 and w182;
w184 <= not w170 and w183;
w185 <= a(116) and not w184;
w186 <= not a(114) and not a(115);
w187 <= not a(116) and w186;
w188 <= not w185 and not w187;
w189 <= not w115 and not w188;
w190 <= not w112 and not w187;
w191 <= not w107 and w190;
w192 <= not w103 and w191;
w193 <= not w101 and w192;
w194 <= not w185 and w193;
w195 <= not a(116) and not w184;
w196 <= a(117) and not w195;
w197 <= w117 and not w184;
w198 <= not w196 and not w197;
w199 <= not w194 and w198;
w200 <= not w189 and not w199;
w201 <= not w60 and not w200;
w202 <= w60 and not w189;
w203 <= not w199 and w202;
w204 <= not w115 and not w181;
w205 <= not w176 and w204;
w206 <= not w172 and w205;
w207 <= not w170 and w206;
w208 <= not w197 and not w207;
w209 <= a(118) and not w208;
w210 <= not a(118) and not w207;
w211 <= not w197 and w210;
w212 <= not w209 and not w211;
w213 <= not w203 and not w212;
w214 <= not w201 and not w213;
w215 <= not w22 and not w214;
w216 <= not w120 and not w125;
w217 <= not w129 and w216;
w218 <= not w184 and w217;
w219 <= not w184 and w216;
w220 <= w129 and not w219;
w221 <= not w218 and not w220;
w222 <= w22 and not w201;
w223 <= not w213 and w222;
w224 <= not w221 and not w223;
w225 <= not w215 and not w224;
w226 <= not w5 and not w225;
w227 <= not w134 and w143;
w228 <= not w132 and w227;
w229 <= not w184 and w228;
w230 <= not w132 and not w134;
w231 <= not w184 and w230;
w232 <= not w143 and not w231;
w233 <= not w229 and not w232;
w234 <= w5 and not w215;
w235 <= not w224 and w234;
w236 <= not w233 and not w235;
w237 <= not w226 and not w236;
w238 <= not w146 and w155;
w239 <= not w148 and w238;
w240 <= not w184 and w239;
w241 <= not w146 and not w148;
w242 <= not w184 and w241;
w243 <= not w155 and not w242;
w244 <= not w240 and not w243;
w245 <= not w157 and not w164;
w246 <= not w184 and w245;
w247 <= not w172 and not w246;
w248 <= not w244 and w247;
w249 <= not w237 and w248;
w250 <= w0 and not w249;
w251 <= not w226 and w244;
w252 <= not w236 and w251;
w253 <= not w164 and not w184;
w254 <= w157 and not w253;
w255 <= not w0 and not w245;
w256 <= not w254 and w255;
w257 <= not w160 and not w181;
w258 <= not w163 and w257;
w259 <= not w176 and w258;
w260 <= not w172 and w259;
w261 <= not w170 and w260;
w262 <= not w256 and not w261;
w263 <= not w252 and w262;
w264 <= not w250 and w263;
w265 <= a(114) and not w264;
w266 <= not a(112) and not a(113);
w267 <= not a(114) and w266;
w268 <= not w265 and not w267;
w269 <= not w184 and not w268;
w270 <= not w181 and not w267;
w271 <= not w176 and w270;
w272 <= not w172 and w271;
w273 <= not w170 and w272;
w274 <= not w265 and w273;
w275 <= not a(114) and not w264;
w276 <= a(115) and not w275;
w277 <= w186 and not w264;
w278 <= not w276 and not w277;
w279 <= not w274 and w278;
w280 <= not w269 and not w279;
w281 <= not w115 and not w280;
w282 <= w115 and not w269;
w283 <= not w279 and w282;
w284 <= not w184 and not w261;
w285 <= not w256 and w284;
w286 <= not w252 and w285;
w287 <= not w250 and w286;
w288 <= not w277 and not w287;
w289 <= a(116) and not w288;
w290 <= not a(116) and not w287;
w291 <= not w277 and w290;
w292 <= not w289 and not w291;
w293 <= not w283 and not w292;
w294 <= not w281 and not w293;
w295 <= not w60 and not w294;
w296 <= not w189 and not w194;
w297 <= not w198 and w296;
w298 <= not w264 and w297;
w299 <= not w264 and w296;
w300 <= w198 and not w299;
w301 <= not w298 and not w300;
w302 <= w60 and not w281;
w303 <= not w293 and w302;
w304 <= not w301 and not w303;
w305 <= not w295 and not w304;
w306 <= not w22 and not w305;
w307 <= not w203 and w212;
w308 <= not w201 and w307;
w309 <= not w264 and w308;
w310 <= not w201 and not w203;
w311 <= not w264 and w310;
w312 <= not w212 and not w311;
w313 <= not w309 and not w312;
w314 <= w22 and not w295;
w315 <= not w304 and w314;
w316 <= not w313 and not w315;
w317 <= not w306 and not w316;
w318 <= not w5 and not w317;
w319 <= not w215 and w221;
w320 <= not w223 and w319;
w321 <= not w264 and w320;
w322 <= not w215 and not w223;
w323 <= not w264 and w322;
w324 <= not w221 and not w323;
w325 <= not w321 and not w324;
w326 <= w5 and not w306;
w327 <= not w316 and w326;
w328 <= not w325 and not w327;
w329 <= not w318 and not w328;
w330 <= w233 and not w235;
w331 <= not w226 and w330;
w332 <= not w264 and w331;
w333 <= not w226 and not w235;
w334 <= not w264 and w333;
w335 <= not w233 and not w334;
w336 <= not w332 and not w335;
w337 <= not w237 and not w244;
w338 <= not w264 and w337;
w339 <= not w252 and not w338;
w340 <= not w336 and w339;
w341 <= not w329 and w340;
w342 <= w0 and not w341;
w343 <= not w318 and w336;
w344 <= not w328 and w343;
w345 <= not w244 and not w264;
w346 <= w237 and not w345;
w347 <= not w0 and not w337;
w348 <= not w346 and w347;
w349 <= not w240 and not w261;
w350 <= not w243 and w349;
w351 <= not w256 and w350;
w352 <= not w252 and w351;
w353 <= not w250 and w352;
w354 <= not w348 and not w353;
w355 <= not w344 and w354;
w356 <= not w342 and w355;
w357 <= a(112) and not w356;
w358 <= not a(110) and not a(111);
w359 <= not a(112) and w358;
w360 <= not w357 and not w359;
w361 <= not w264 and not w360;
w362 <= not a(112) and not w356;
w363 <= a(113) and not w362;
w364 <= w266 and not w356;
w365 <= not w363 and not w364;
w366 <= not w261 and not w359;
w367 <= not w256 and w366;
w368 <= not w252 and w367;
w369 <= not w250 and w368;
w370 <= not w357 and w369;
w371 <= w365 and not w370;
w372 <= not w361 and not w371;
w373 <= not w184 and not w372;
w374 <= w184 and not w361;
w375 <= not w371 and w374;
w376 <= not w264 and not w353;
w377 <= not w348 and w376;
w378 <= not w344 and w377;
w379 <= not w342 and w378;
w380 <= not w364 and not w379;
w381 <= a(114) and not w380;
w382 <= not a(114) and not w379;
w383 <= not w364 and w382;
w384 <= not w381 and not w383;
w385 <= not w375 and not w384;
w386 <= not w373 and not w385;
w387 <= not w115 and not w386;
w388 <= not w269 and not w274;
w389 <= not w278 and w388;
w390 <= not w356 and w389;
w391 <= not w356 and w388;
w392 <= w278 and not w391;
w393 <= not w390 and not w392;
w394 <= w115 and not w373;
w395 <= not w385 and w394;
w396 <= not w393 and not w395;
w397 <= not w387 and not w396;
w398 <= not w60 and not w397;
w399 <= not w283 and w292;
w400 <= not w281 and w399;
w401 <= not w356 and w400;
w402 <= not w281 and not w283;
w403 <= not w356 and w402;
w404 <= not w292 and not w403;
w405 <= not w401 and not w404;
w406 <= w60 and not w387;
w407 <= not w396 and w406;
w408 <= not w405 and not w407;
w409 <= not w398 and not w408;
w410 <= not w22 and not w409;
w411 <= not w295 and w301;
w412 <= not w303 and w411;
w413 <= not w356 and w412;
w414 <= not w295 and not w303;
w415 <= not w356 and w414;
w416 <= not w301 and not w415;
w417 <= not w413 and not w416;
w418 <= w22 and not w398;
w419 <= not w408 and w418;
w420 <= not w417 and not w419;
w421 <= not w410 and not w420;
w422 <= not w5 and not w421;
w423 <= w313 and not w315;
w424 <= not w306 and w423;
w425 <= not w356 and w424;
w426 <= not w306 and not w315;
w427 <= not w356 and w426;
w428 <= not w313 and not w427;
w429 <= not w425 and not w428;
w430 <= w5 and not w410;
w431 <= not w420 and w430;
w432 <= not w429 and not w431;
w433 <= not w422 and not w432;
w434 <= not w318 and w325;
w435 <= not w327 and w434;
w436 <= not w356 and w435;
w437 <= not w318 and not w327;
w438 <= not w356 and w437;
w439 <= not w325 and not w438;
w440 <= not w436 and not w439;
w441 <= not w329 and not w336;
w442 <= not w356 and w441;
w443 <= not w344 and not w442;
w444 <= not w440 and w443;
w445 <= not w433 and w444;
w446 <= w0 and not w445;
w447 <= not w422 and w440;
w448 <= not w432 and w447;
w449 <= not w336 and not w356;
w450 <= w329 and not w449;
w451 <= not w0 and not w441;
w452 <= not w450 and w451;
w453 <= not w332 and not w353;
w454 <= not w335 and w453;
w455 <= not w348 and w454;
w456 <= not w344 and w455;
w457 <= not w342 and w456;
w458 <= not w452 and not w457;
w459 <= not w448 and w458;
w460 <= not w446 and w459;
w461 <= a(110) and not w460;
w462 <= not a(108) and not a(109);
w463 <= not a(110) and w462;
w464 <= not w461 and not w463;
w465 <= not w356 and not w464;
w466 <= not w353 and not w463;
w467 <= not w348 and w466;
w468 <= not w344 and w467;
w469 <= not w342 and w468;
w470 <= not w461 and w469;
w471 <= not a(110) and not w460;
w472 <= a(111) and not w471;
w473 <= w358 and not w460;
w474 <= not w472 and not w473;
w475 <= not w470 and w474;
w476 <= not w465 and not w475;
w477 <= not w264 and not w476;
w478 <= w264 and not w465;
w479 <= not w475 and w478;
w480 <= not w356 and not w457;
w481 <= not w452 and w480;
w482 <= not w448 and w481;
w483 <= not w446 and w482;
w484 <= not w473 and not w483;
w485 <= a(112) and not w484;
w486 <= not a(112) and not w483;
w487 <= not w473 and w486;
w488 <= not w485 and not w487;
w489 <= not w479 and not w488;
w490 <= not w477 and not w489;
w491 <= not w184 and not w490;
w492 <= w184 and not w477;
w493 <= not w489 and w492;
w494 <= not w365 and not w370;
w495 <= not w361 and w494;
w496 <= not w460 and w495;
w497 <= not w361 and not w370;
w498 <= not w460 and w497;
w499 <= w365 and not w498;
w500 <= not w496 and not w499;
w501 <= not w493 and not w500;
w502 <= not w491 and not w501;
w503 <= not w115 and not w502;
w504 <= not w375 and w384;
w505 <= not w373 and w504;
w506 <= not w460 and w505;
w507 <= not w373 and not w375;
w508 <= not w460 and w507;
w509 <= not w384 and not w508;
w510 <= not w506 and not w509;
w511 <= w115 and not w491;
w512 <= not w501 and w511;
w513 <= not w510 and not w512;
w514 <= not w503 and not w513;
w515 <= not w60 and not w514;
w516 <= not w387 and w393;
w517 <= not w395 and w516;
w518 <= not w460 and w517;
w519 <= not w387 and not w395;
w520 <= not w460 and w519;
w521 <= not w393 and not w520;
w522 <= not w518 and not w521;
w523 <= w60 and not w503;
w524 <= not w513 and w523;
w525 <= not w522 and not w524;
w526 <= not w515 and not w525;
w527 <= not w22 and not w526;
w528 <= w405 and not w407;
w529 <= not w398 and w528;
w530 <= not w460 and w529;
w531 <= not w398 and not w407;
w532 <= not w460 and w531;
w533 <= not w405 and not w532;
w534 <= not w530 and not w533;
w535 <= w22 and not w515;
w536 <= not w525 and w535;
w537 <= not w534 and not w536;
w538 <= not w527 and not w537;
w539 <= not w5 and not w538;
w540 <= not w410 and w417;
w541 <= not w419 and w540;
w542 <= not w460 and w541;
w543 <= not w410 and not w419;
w544 <= not w460 and w543;
w545 <= not w417 and not w544;
w546 <= not w542 and not w545;
w547 <= w5 and not w527;
w548 <= not w537 and w547;
w549 <= not w546 and not w548;
w550 <= not w539 and not w549;
w551 <= w429 and not w431;
w552 <= not w422 and w551;
w553 <= not w460 and w552;
w554 <= not w422 and not w431;
w555 <= not w460 and w554;
w556 <= not w429 and not w555;
w557 <= not w553 and not w556;
w558 <= not w433 and not w440;
w559 <= not w460 and w558;
w560 <= not w448 and not w559;
w561 <= not w557 and w560;
w562 <= not w550 and w561;
w563 <= w0 and not w562;
w564 <= not w539 and w557;
w565 <= not w549 and w564;
w566 <= not w440 and not w460;
w567 <= w433 and not w566;
w568 <= not w0 and not w558;
w569 <= not w567 and w568;
w570 <= not w436 and not w457;
w571 <= not w439 and w570;
w572 <= not w452 and w571;
w573 <= not w448 and w572;
w574 <= not w446 and w573;
w575 <= not w569 and not w574;
w576 <= not w565 and w575;
w577 <= not w563 and w576;
w578 <= a(108) and not w577;
w579 <= not a(106) and not a(107);
w580 <= not a(108) and w579;
w581 <= not w578 and not w580;
w582 <= not w460 and not w581;
w583 <= not w457 and not w580;
w584 <= not w452 and w583;
w585 <= not w448 and w584;
w586 <= not w446 and w585;
w587 <= not w578 and w586;
w588 <= not a(108) and not w577;
w589 <= a(109) and not w588;
w590 <= w462 and not w577;
w591 <= not w589 and not w590;
w592 <= not w587 and w591;
w593 <= not w582 and not w592;
w594 <= not w356 and not w593;
w595 <= w356 and not w582;
w596 <= not w592 and w595;
w597 <= not w460 and not w574;
w598 <= not w569 and w597;
w599 <= not w565 and w598;
w600 <= not w563 and w599;
w601 <= not w590 and not w600;
w602 <= a(110) and not w601;
w603 <= not a(110) and not w600;
w604 <= not w590 and w603;
w605 <= not w602 and not w604;
w606 <= not w596 and not w605;
w607 <= not w594 and not w606;
w608 <= not w264 and not w607;
w609 <= not w465 and not w470;
w610 <= not w474 and w609;
w611 <= not w577 and w610;
w612 <= not w577 and w609;
w613 <= w474 and not w612;
w614 <= not w611 and not w613;
w615 <= w264 and not w594;
w616 <= not w606 and w615;
w617 <= not w614 and not w616;
w618 <= not w608 and not w617;
w619 <= not w184 and not w618;
w620 <= not w479 and w488;
w621 <= not w477 and w620;
w622 <= not w577 and w621;
w623 <= not w477 and not w479;
w624 <= not w577 and w623;
w625 <= not w488 and not w624;
w626 <= not w622 and not w625;
w627 <= w184 and not w608;
w628 <= not w617 and w627;
w629 <= not w626 and not w628;
w630 <= not w619 and not w629;
w631 <= not w115 and not w630;
w632 <= w115 and not w619;
w633 <= not w629 and w632;
w634 <= not w491 and w500;
w635 <= not w493 and w634;
w636 <= not w577 and w635;
w637 <= not w491 and not w493;
w638 <= not w577 and w637;
w639 <= not w500 and not w638;
w640 <= not w636 and not w639;
w641 <= not w633 and not w640;
w642 <= not w631 and not w641;
w643 <= not w60 and not w642;
w644 <= w510 and not w512;
w645 <= not w503 and w644;
w646 <= not w577 and w645;
w647 <= not w503 and not w512;
w648 <= not w577 and w647;
w649 <= not w510 and not w648;
w650 <= not w646 and not w649;
w651 <= w60 and not w631;
w652 <= not w641 and w651;
w653 <= not w650 and not w652;
w654 <= not w643 and not w653;
w655 <= not w22 and not w654;
w656 <= not w515 and w522;
w657 <= not w524 and w656;
w658 <= not w577 and w657;
w659 <= not w515 and not w524;
w660 <= not w577 and w659;
w661 <= not w522 and not w660;
w662 <= not w658 and not w661;
w663 <= w22 and not w643;
w664 <= not w653 and w663;
w665 <= not w662 and not w664;
w666 <= not w655 and not w665;
w667 <= not w5 and not w666;
w668 <= w534 and not w536;
w669 <= not w527 and w668;
w670 <= not w577 and w669;
w671 <= not w527 and not w536;
w672 <= not w577 and w671;
w673 <= not w534 and not w672;
w674 <= not w670 and not w673;
w675 <= w5 and not w655;
w676 <= not w665 and w675;
w677 <= not w674 and not w676;
w678 <= not w667 and not w677;
w679 <= not w539 and w546;
w680 <= not w548 and w679;
w681 <= not w577 and w680;
w682 <= not w539 and not w548;
w683 <= not w577 and w682;
w684 <= not w546 and not w683;
w685 <= not w681 and not w684;
w686 <= not w550 and not w557;
w687 <= not w577 and w686;
w688 <= not w565 and not w687;
w689 <= not w685 and w688;
w690 <= not w678 and w689;
w691 <= w0 and not w690;
w692 <= not w667 and w685;
w693 <= not w677 and w692;
w694 <= not w557 and not w577;
w695 <= w550 and not w694;
w696 <= not w0 and not w686;
w697 <= not w695 and w696;
w698 <= not w553 and not w574;
w699 <= not w556 and w698;
w700 <= not w569 and w699;
w701 <= not w565 and w700;
w702 <= not w563 and w701;
w703 <= not w697 and not w702;
w704 <= not w693 and w703;
w705 <= not w691 and w704;
w706 <= a(106) and not w705;
w707 <= not a(104) and not a(105);
w708 <= not a(106) and w707;
w709 <= not w706 and not w708;
w710 <= not w577 and not w709;
w711 <= not w574 and not w708;
w712 <= not w569 and w711;
w713 <= not w565 and w712;
w714 <= not w563 and w713;
w715 <= not w706 and w714;
w716 <= not a(106) and not w705;
w717 <= a(107) and not w716;
w718 <= w579 and not w705;
w719 <= not w717 and not w718;
w720 <= not w715 and w719;
w721 <= not w710 and not w720;
w722 <= not w460 and not w721;
w723 <= w460 and not w710;
w724 <= not w720 and w723;
w725 <= not w577 and not w702;
w726 <= not w697 and w725;
w727 <= not w693 and w726;
w728 <= not w691 and w727;
w729 <= not w718 and not w728;
w730 <= a(108) and not w729;
w731 <= not a(108) and not w728;
w732 <= not w718 and w731;
w733 <= not w730 and not w732;
w734 <= not w724 and not w733;
w735 <= not w722 and not w734;
w736 <= not w356 and not w735;
w737 <= not w582 and not w587;
w738 <= not w591 and w737;
w739 <= not w705 and w738;
w740 <= not w705 and w737;
w741 <= w591 and not w740;
w742 <= not w739 and not w741;
w743 <= w356 and not w722;
w744 <= not w734 and w743;
w745 <= not w742 and not w744;
w746 <= not w736 and not w745;
w747 <= not w264 and not w746;
w748 <= not w596 and w605;
w749 <= not w594 and w748;
w750 <= not w705 and w749;
w751 <= not w594 and not w596;
w752 <= not w705 and w751;
w753 <= not w605 and not w752;
w754 <= not w750 and not w753;
w755 <= w264 and not w736;
w756 <= not w745 and w755;
w757 <= not w754 and not w756;
w758 <= not w747 and not w757;
w759 <= not w184 and not w758;
w760 <= not w608 and w614;
w761 <= not w616 and w760;
w762 <= not w705 and w761;
w763 <= not w608 and not w616;
w764 <= not w705 and w763;
w765 <= not w614 and not w764;
w766 <= not w762 and not w765;
w767 <= w184 and not w747;
w768 <= not w757 and w767;
w769 <= not w766 and not w768;
w770 <= not w759 and not w769;
w771 <= not w115 and not w770;
w772 <= w626 and not w628;
w773 <= not w619 and w772;
w774 <= not w705 and w773;
w775 <= not w619 and not w628;
w776 <= not w705 and w775;
w777 <= not w626 and not w776;
w778 <= not w774 and not w777;
w779 <= w115 and not w759;
w780 <= not w769 and w779;
w781 <= not w778 and not w780;
w782 <= not w771 and not w781;
w783 <= not w60 and not w782;
w784 <= w60 and not w771;
w785 <= not w781 and w784;
w786 <= not w631 and w640;
w787 <= not w633 and w786;
w788 <= not w705 and w787;
w789 <= not w631 and not w633;
w790 <= not w705 and w789;
w791 <= not w640 and not w790;
w792 <= not w788 and not w791;
w793 <= not w785 and not w792;
w794 <= not w783 and not w793;
w795 <= not w22 and not w794;
w796 <= w650 and not w652;
w797 <= not w643 and w796;
w798 <= not w705 and w797;
w799 <= not w643 and not w652;
w800 <= not w705 and w799;
w801 <= not w650 and not w800;
w802 <= not w798 and not w801;
w803 <= w22 and not w783;
w804 <= not w793 and w803;
w805 <= not w802 and not w804;
w806 <= not w795 and not w805;
w807 <= not w5 and not w806;
w808 <= not w655 and w662;
w809 <= not w664 and w808;
w810 <= not w705 and w809;
w811 <= not w655 and not w664;
w812 <= not w705 and w811;
w813 <= not w662 and not w812;
w814 <= not w810 and not w813;
w815 <= w5 and not w795;
w816 <= not w805 and w815;
w817 <= not w814 and not w816;
w818 <= not w807 and not w817;
w819 <= w674 and not w676;
w820 <= not w667 and w819;
w821 <= not w705 and w820;
w822 <= not w667 and not w676;
w823 <= not w705 and w822;
w824 <= not w674 and not w823;
w825 <= not w821 and not w824;
w826 <= not w678 and not w685;
w827 <= not w705 and w826;
w828 <= not w693 and not w827;
w829 <= not w825 and w828;
w830 <= not w818 and w829;
w831 <= w0 and not w830;
w832 <= not w807 and w825;
w833 <= not w817 and w832;
w834 <= not w685 and not w705;
w835 <= w678 and not w834;
w836 <= not w0 and not w826;
w837 <= not w835 and w836;
w838 <= not w681 and not w702;
w839 <= not w684 and w838;
w840 <= not w697 and w839;
w841 <= not w693 and w840;
w842 <= not w691 and w841;
w843 <= not w837 and not w842;
w844 <= not w833 and w843;
w845 <= not w831 and w844;
w846 <= a(104) and not w845;
w847 <= not a(102) and not a(103);
w848 <= not a(104) and w847;
w849 <= not w846 and not w848;
w850 <= not w705 and not w849;
w851 <= not w702 and not w848;
w852 <= not w697 and w851;
w853 <= not w693 and w852;
w854 <= not w691 and w853;
w855 <= not w846 and w854;
w856 <= not a(104) and not w845;
w857 <= a(105) and not w856;
w858 <= w707 and not w845;
w859 <= not w857 and not w858;
w860 <= not w855 and w859;
w861 <= not w850 and not w860;
w862 <= not w577 and not w861;
w863 <= w577 and not w850;
w864 <= not w860 and w863;
w865 <= not w705 and not w842;
w866 <= not w837 and w865;
w867 <= not w833 and w866;
w868 <= not w831 and w867;
w869 <= not w858 and not w868;
w870 <= a(106) and not w869;
w871 <= not a(106) and not w868;
w872 <= not w858 and w871;
w873 <= not w870 and not w872;
w874 <= not w864 and not w873;
w875 <= not w862 and not w874;
w876 <= not w460 and not w875;
w877 <= not w710 and not w715;
w878 <= not w719 and w877;
w879 <= not w845 and w878;
w880 <= not w845 and w877;
w881 <= w719 and not w880;
w882 <= not w879 and not w881;
w883 <= w460 and not w862;
w884 <= not w874 and w883;
w885 <= not w882 and not w884;
w886 <= not w876 and not w885;
w887 <= not w356 and not w886;
w888 <= not w724 and w733;
w889 <= not w722 and w888;
w890 <= not w845 and w889;
w891 <= not w722 and not w724;
w892 <= not w845 and w891;
w893 <= not w733 and not w892;
w894 <= not w890 and not w893;
w895 <= w356 and not w876;
w896 <= not w885 and w895;
w897 <= not w894 and not w896;
w898 <= not w887 and not w897;
w899 <= not w264 and not w898;
w900 <= not w736 and w742;
w901 <= not w744 and w900;
w902 <= not w845 and w901;
w903 <= not w736 and not w744;
w904 <= not w845 and w903;
w905 <= not w742 and not w904;
w906 <= not w902 and not w905;
w907 <= w264 and not w887;
w908 <= not w897 and w907;
w909 <= not w906 and not w908;
w910 <= not w899 and not w909;
w911 <= not w184 and not w910;
w912 <= w754 and not w756;
w913 <= not w747 and w912;
w914 <= not w845 and w913;
w915 <= not w747 and not w756;
w916 <= not w845 and w915;
w917 <= not w754 and not w916;
w918 <= not w914 and not w917;
w919 <= w184 and not w899;
w920 <= not w909 and w919;
w921 <= not w918 and not w920;
w922 <= not w911 and not w921;
w923 <= not w115 and not w922;
w924 <= not w759 and w766;
w925 <= not w768 and w924;
w926 <= not w845 and w925;
w927 <= not w759 and not w768;
w928 <= not w845 and w927;
w929 <= not w766 and not w928;
w930 <= not w926 and not w929;
w931 <= w115 and not w911;
w932 <= not w921 and w931;
w933 <= not w930 and not w932;
w934 <= not w923 and not w933;
w935 <= not w60 and not w934;
w936 <= w778 and not w780;
w937 <= not w771 and w936;
w938 <= not w845 and w937;
w939 <= not w771 and not w780;
w940 <= not w845 and w939;
w941 <= not w778 and not w940;
w942 <= not w938 and not w941;
w943 <= w60 and not w923;
w944 <= not w933 and w943;
w945 <= not w942 and not w944;
w946 <= not w935 and not w945;
w947 <= not w22 and not w946;
w948 <= w22 and not w935;
w949 <= not w945 and w948;
w950 <= not w783 and w792;
w951 <= not w785 and w950;
w952 <= not w845 and w951;
w953 <= not w783 and not w785;
w954 <= not w845 and w953;
w955 <= not w792 and not w954;
w956 <= not w952 and not w955;
w957 <= not w949 and not w956;
w958 <= not w947 and not w957;
w959 <= not w5 and not w958;
w960 <= w802 and not w804;
w961 <= not w795 and w960;
w962 <= not w845 and w961;
w963 <= not w795 and not w804;
w964 <= not w845 and w963;
w965 <= not w802 and not w964;
w966 <= not w962 and not w965;
w967 <= w5 and not w947;
w968 <= not w957 and w967;
w969 <= not w966 and not w968;
w970 <= not w959 and not w969;
w971 <= not w807 and w814;
w972 <= not w816 and w971;
w973 <= not w845 and w972;
w974 <= not w807 and not w816;
w975 <= not w845 and w974;
w976 <= not w814 and not w975;
w977 <= not w973 and not w976;
w978 <= not w818 and not w825;
w979 <= not w845 and w978;
w980 <= not w833 and not w979;
w981 <= not w977 and w980;
w982 <= not w970 and w981;
w983 <= w0 and not w982;
w984 <= not w959 and w977;
w985 <= not w969 and w984;
w986 <= not w825 and not w845;
w987 <= w818 and not w986;
w988 <= not w0 and not w978;
w989 <= not w987 and w988;
w990 <= not w821 and not w842;
w991 <= not w824 and w990;
w992 <= not w837 and w991;
w993 <= not w833 and w992;
w994 <= not w831 and w993;
w995 <= not w989 and not w994;
w996 <= not w985 and w995;
w997 <= not w983 and w996;
w998 <= a(102) and not w997;
w999 <= not a(100) and not a(101);
w1000 <= not a(102) and w999;
w1001 <= not w998 and not w1000;
w1002 <= not w845 and not w1001;
w1003 <= not w842 and not w1000;
w1004 <= not w837 and w1003;
w1005 <= not w833 and w1004;
w1006 <= not w831 and w1005;
w1007 <= not w998 and w1006;
w1008 <= not a(102) and not w997;
w1009 <= a(103) and not w1008;
w1010 <= w847 and not w997;
w1011 <= not w1009 and not w1010;
w1012 <= not w1007 and w1011;
w1013 <= not w1002 and not w1012;
w1014 <= not w705 and not w1013;
w1015 <= w705 and not w1002;
w1016 <= not w1012 and w1015;
w1017 <= not w845 and not w994;
w1018 <= not w989 and w1017;
w1019 <= not w985 and w1018;
w1020 <= not w983 and w1019;
w1021 <= not w1010 and not w1020;
w1022 <= a(104) and not w1021;
w1023 <= not a(104) and not w1020;
w1024 <= not w1010 and w1023;
w1025 <= not w1022 and not w1024;
w1026 <= not w1016 and not w1025;
w1027 <= not w1014 and not w1026;
w1028 <= not w577 and not w1027;
w1029 <= not w850 and not w855;
w1030 <= not w859 and w1029;
w1031 <= not w997 and w1030;
w1032 <= not w997 and w1029;
w1033 <= w859 and not w1032;
w1034 <= not w1031 and not w1033;
w1035 <= w577 and not w1014;
w1036 <= not w1026 and w1035;
w1037 <= not w1034 and not w1036;
w1038 <= not w1028 and not w1037;
w1039 <= not w460 and not w1038;
w1040 <= not w864 and w873;
w1041 <= not w862 and w1040;
w1042 <= not w997 and w1041;
w1043 <= not w862 and not w864;
w1044 <= not w997 and w1043;
w1045 <= not w873 and not w1044;
w1046 <= not w1042 and not w1045;
w1047 <= w460 and not w1028;
w1048 <= not w1037 and w1047;
w1049 <= not w1046 and not w1048;
w1050 <= not w1039 and not w1049;
w1051 <= not w356 and not w1050;
w1052 <= not w876 and w882;
w1053 <= not w884 and w1052;
w1054 <= not w997 and w1053;
w1055 <= not w876 and not w884;
w1056 <= not w997 and w1055;
w1057 <= not w882 and not w1056;
w1058 <= not w1054 and not w1057;
w1059 <= w356 and not w1039;
w1060 <= not w1049 and w1059;
w1061 <= not w1058 and not w1060;
w1062 <= not w1051 and not w1061;
w1063 <= not w264 and not w1062;
w1064 <= w894 and not w896;
w1065 <= not w887 and w1064;
w1066 <= not w997 and w1065;
w1067 <= not w887 and not w896;
w1068 <= not w997 and w1067;
w1069 <= not w894 and not w1068;
w1070 <= not w1066 and not w1069;
w1071 <= w264 and not w1051;
w1072 <= not w1061 and w1071;
w1073 <= not w1070 and not w1072;
w1074 <= not w1063 and not w1073;
w1075 <= not w184 and not w1074;
w1076 <= not w899 and w906;
w1077 <= not w908 and w1076;
w1078 <= not w997 and w1077;
w1079 <= not w899 and not w908;
w1080 <= not w997 and w1079;
w1081 <= not w906 and not w1080;
w1082 <= not w1078 and not w1081;
w1083 <= w184 and not w1063;
w1084 <= not w1073 and w1083;
w1085 <= not w1082 and not w1084;
w1086 <= not w1075 and not w1085;
w1087 <= not w115 and not w1086;
w1088 <= w918 and not w920;
w1089 <= not w911 and w1088;
w1090 <= not w997 and w1089;
w1091 <= not w911 and not w920;
w1092 <= not w997 and w1091;
w1093 <= not w918 and not w1092;
w1094 <= not w1090 and not w1093;
w1095 <= w115 and not w1075;
w1096 <= not w1085 and w1095;
w1097 <= not w1094 and not w1096;
w1098 <= not w1087 and not w1097;
w1099 <= not w60 and not w1098;
w1100 <= not w923 and w930;
w1101 <= not w932 and w1100;
w1102 <= not w997 and w1101;
w1103 <= not w923 and not w932;
w1104 <= not w997 and w1103;
w1105 <= not w930 and not w1104;
w1106 <= not w1102 and not w1105;
w1107 <= w60 and not w1087;
w1108 <= not w1097 and w1107;
w1109 <= not w1106 and not w1108;
w1110 <= not w1099 and not w1109;
w1111 <= not w22 and not w1110;
w1112 <= w942 and not w944;
w1113 <= not w935 and w1112;
w1114 <= not w997 and w1113;
w1115 <= not w935 and not w944;
w1116 <= not w997 and w1115;
w1117 <= not w942 and not w1116;
w1118 <= not w1114 and not w1117;
w1119 <= w22 and not w1099;
w1120 <= not w1109 and w1119;
w1121 <= not w1118 and not w1120;
w1122 <= not w1111 and not w1121;
w1123 <= not w5 and not w1122;
w1124 <= w5 and not w1111;
w1125 <= not w1121 and w1124;
w1126 <= not w947 and w956;
w1127 <= not w949 and w1126;
w1128 <= not w997 and w1127;
w1129 <= not w947 and not w949;
w1130 <= not w997 and w1129;
w1131 <= not w956 and not w1130;
w1132 <= not w1128 and not w1131;
w1133 <= not w1125 and not w1132;
w1134 <= not w1123 and not w1133;
w1135 <= w966 and not w968;
w1136 <= not w959 and w1135;
w1137 <= not w997 and w1136;
w1138 <= not w959 and not w968;
w1139 <= not w997 and w1138;
w1140 <= not w966 and not w1139;
w1141 <= not w1137 and not w1140;
w1142 <= not w970 and not w977;
w1143 <= not w997 and w1142;
w1144 <= not w985 and not w1143;
w1145 <= not w1141 and w1144;
w1146 <= not w1134 and w1145;
w1147 <= w0 and not w1146;
w1148 <= not w1123 and w1141;
w1149 <= not w1133 and w1148;
w1150 <= not w977 and not w997;
w1151 <= w970 and not w1150;
w1152 <= not w0 and not w1142;
w1153 <= not w1151 and w1152;
w1154 <= not w973 and not w994;
w1155 <= not w976 and w1154;
w1156 <= not w989 and w1155;
w1157 <= not w985 and w1156;
w1158 <= not w983 and w1157;
w1159 <= not w1153 and not w1158;
w1160 <= not w1149 and w1159;
w1161 <= not w1147 and w1160;
w1162 <= a(100) and not w1161;
w1163 <= not a(98) and not a(99);
w1164 <= not a(100) and w1163;
w1165 <= not w1162 and not w1164;
w1166 <= not w997 and not w1165;
w1167 <= not w994 and not w1164;
w1168 <= not w989 and w1167;
w1169 <= not w985 and w1168;
w1170 <= not w983 and w1169;
w1171 <= not w1162 and w1170;
w1172 <= not a(100) and not w1161;
w1173 <= a(101) and not w1172;
w1174 <= w999 and not w1161;
w1175 <= not w1173 and not w1174;
w1176 <= not w1171 and w1175;
w1177 <= not w1166 and not w1176;
w1178 <= not w845 and not w1177;
w1179 <= w845 and not w1166;
w1180 <= not w1176 and w1179;
w1181 <= not w997 and not w1158;
w1182 <= not w1153 and w1181;
w1183 <= not w1149 and w1182;
w1184 <= not w1147 and w1183;
w1185 <= not w1174 and not w1184;
w1186 <= a(102) and not w1185;
w1187 <= not a(102) and not w1184;
w1188 <= not w1174 and w1187;
w1189 <= not w1186 and not w1188;
w1190 <= not w1180 and not w1189;
w1191 <= not w1178 and not w1190;
w1192 <= not w705 and not w1191;
w1193 <= not w1002 and not w1007;
w1194 <= not w1011 and w1193;
w1195 <= not w1161 and w1194;
w1196 <= not w1161 and w1193;
w1197 <= w1011 and not w1196;
w1198 <= not w1195 and not w1197;
w1199 <= w705 and not w1178;
w1200 <= not w1190 and w1199;
w1201 <= not w1198 and not w1200;
w1202 <= not w1192 and not w1201;
w1203 <= not w577 and not w1202;
w1204 <= not w1016 and w1025;
w1205 <= not w1014 and w1204;
w1206 <= not w1161 and w1205;
w1207 <= not w1014 and not w1016;
w1208 <= not w1161 and w1207;
w1209 <= not w1025 and not w1208;
w1210 <= not w1206 and not w1209;
w1211 <= w577 and not w1192;
w1212 <= not w1201 and w1211;
w1213 <= not w1210 and not w1212;
w1214 <= not w1203 and not w1213;
w1215 <= not w460 and not w1214;
w1216 <= not w1028 and w1034;
w1217 <= not w1036 and w1216;
w1218 <= not w1161 and w1217;
w1219 <= not w1028 and not w1036;
w1220 <= not w1161 and w1219;
w1221 <= not w1034 and not w1220;
w1222 <= not w1218 and not w1221;
w1223 <= w460 and not w1203;
w1224 <= not w1213 and w1223;
w1225 <= not w1222 and not w1224;
w1226 <= not w1215 and not w1225;
w1227 <= not w356 and not w1226;
w1228 <= w1046 and not w1048;
w1229 <= not w1039 and w1228;
w1230 <= not w1161 and w1229;
w1231 <= not w1039 and not w1048;
w1232 <= not w1161 and w1231;
w1233 <= not w1046 and not w1232;
w1234 <= not w1230 and not w1233;
w1235 <= w356 and not w1215;
w1236 <= not w1225 and w1235;
w1237 <= not w1234 and not w1236;
w1238 <= not w1227 and not w1237;
w1239 <= not w264 and not w1238;
w1240 <= not w1051 and w1058;
w1241 <= not w1060 and w1240;
w1242 <= not w1161 and w1241;
w1243 <= not w1051 and not w1060;
w1244 <= not w1161 and w1243;
w1245 <= not w1058 and not w1244;
w1246 <= not w1242 and not w1245;
w1247 <= w264 and not w1227;
w1248 <= not w1237 and w1247;
w1249 <= not w1246 and not w1248;
w1250 <= not w1239 and not w1249;
w1251 <= not w184 and not w1250;
w1252 <= w1070 and not w1072;
w1253 <= not w1063 and w1252;
w1254 <= not w1161 and w1253;
w1255 <= not w1063 and not w1072;
w1256 <= not w1161 and w1255;
w1257 <= not w1070 and not w1256;
w1258 <= not w1254 and not w1257;
w1259 <= w184 and not w1239;
w1260 <= not w1249 and w1259;
w1261 <= not w1258 and not w1260;
w1262 <= not w1251 and not w1261;
w1263 <= not w115 and not w1262;
w1264 <= not w1075 and w1082;
w1265 <= not w1084 and w1264;
w1266 <= not w1161 and w1265;
w1267 <= not w1075 and not w1084;
w1268 <= not w1161 and w1267;
w1269 <= not w1082 and not w1268;
w1270 <= not w1266 and not w1269;
w1271 <= w115 and not w1251;
w1272 <= not w1261 and w1271;
w1273 <= not w1270 and not w1272;
w1274 <= not w1263 and not w1273;
w1275 <= not w60 and not w1274;
w1276 <= w1094 and not w1096;
w1277 <= not w1087 and w1276;
w1278 <= not w1161 and w1277;
w1279 <= not w1087 and not w1096;
w1280 <= not w1161 and w1279;
w1281 <= not w1094 and not w1280;
w1282 <= not w1278 and not w1281;
w1283 <= w60 and not w1263;
w1284 <= not w1273 and w1283;
w1285 <= not w1282 and not w1284;
w1286 <= not w1275 and not w1285;
w1287 <= not w22 and not w1286;
w1288 <= not w1099 and w1106;
w1289 <= not w1108 and w1288;
w1290 <= not w1161 and w1289;
w1291 <= not w1099 and not w1108;
w1292 <= not w1161 and w1291;
w1293 <= not w1106 and not w1292;
w1294 <= not w1290 and not w1293;
w1295 <= w22 and not w1275;
w1296 <= not w1285 and w1295;
w1297 <= not w1294 and not w1296;
w1298 <= not w1287 and not w1297;
w1299 <= not w5 and not w1298;
w1300 <= w1118 and not w1120;
w1301 <= not w1111 and w1300;
w1302 <= not w1161 and w1301;
w1303 <= not w1111 and not w1120;
w1304 <= not w1161 and w1303;
w1305 <= not w1118 and not w1304;
w1306 <= not w1302 and not w1305;
w1307 <= w5 and not w1287;
w1308 <= not w1297 and w1307;
w1309 <= not w1306 and not w1308;
w1310 <= not w1299 and not w1309;
w1311 <= not w1123 and w1132;
w1312 <= not w1125 and w1311;
w1313 <= not w1161 and w1312;
w1314 <= not w1123 and not w1125;
w1315 <= not w1161 and w1314;
w1316 <= not w1132 and not w1315;
w1317 <= not w1313 and not w1316;
w1318 <= not w1134 and not w1141;
w1319 <= not w1161 and w1318;
w1320 <= not w1149 and not w1319;
w1321 <= not w1317 and w1320;
w1322 <= not w1310 and w1321;
w1323 <= w0 and not w1322;
w1324 <= not w1299 and w1317;
w1325 <= not w1309 and w1324;
w1326 <= not w1141 and not w1161;
w1327 <= w1134 and not w1326;
w1328 <= not w0 and not w1318;
w1329 <= not w1327 and w1328;
w1330 <= not w1137 and not w1158;
w1331 <= not w1140 and w1330;
w1332 <= not w1153 and w1331;
w1333 <= not w1149 and w1332;
w1334 <= not w1147 and w1333;
w1335 <= not w1329 and not w1334;
w1336 <= not w1325 and w1335;
w1337 <= not w1323 and w1336;
w1338 <= a(98) and not w1337;
w1339 <= not a(96) and not a(97);
w1340 <= not a(98) and w1339;
w1341 <= not w1338 and not w1340;
w1342 <= not w1161 and not w1341;
w1343 <= not w1158 and not w1340;
w1344 <= not w1153 and w1343;
w1345 <= not w1149 and w1344;
w1346 <= not w1147 and w1345;
w1347 <= not w1338 and w1346;
w1348 <= not a(98) and not w1337;
w1349 <= a(99) and not w1348;
w1350 <= w1163 and not w1337;
w1351 <= not w1349 and not w1350;
w1352 <= not w1347 and w1351;
w1353 <= not w1342 and not w1352;
w1354 <= not w997 and not w1353;
w1355 <= w997 and not w1342;
w1356 <= not w1352 and w1355;
w1357 <= not w1161 and not w1334;
w1358 <= not w1329 and w1357;
w1359 <= not w1325 and w1358;
w1360 <= not w1323 and w1359;
w1361 <= not w1350 and not w1360;
w1362 <= a(100) and not w1361;
w1363 <= not a(100) and not w1360;
w1364 <= not w1350 and w1363;
w1365 <= not w1362 and not w1364;
w1366 <= not w1356 and not w1365;
w1367 <= not w1354 and not w1366;
w1368 <= not w845 and not w1367;
w1369 <= not w1166 and not w1171;
w1370 <= not w1175 and w1369;
w1371 <= not w1337 and w1370;
w1372 <= not w1337 and w1369;
w1373 <= w1175 and not w1372;
w1374 <= not w1371 and not w1373;
w1375 <= w845 and not w1354;
w1376 <= not w1366 and w1375;
w1377 <= not w1374 and not w1376;
w1378 <= not w1368 and not w1377;
w1379 <= not w705 and not w1378;
w1380 <= not w1180 and w1189;
w1381 <= not w1178 and w1380;
w1382 <= not w1337 and w1381;
w1383 <= not w1178 and not w1180;
w1384 <= not w1337 and w1383;
w1385 <= not w1189 and not w1384;
w1386 <= not w1382 and not w1385;
w1387 <= w705 and not w1368;
w1388 <= not w1377 and w1387;
w1389 <= not w1386 and not w1388;
w1390 <= not w1379 and not w1389;
w1391 <= not w577 and not w1390;
w1392 <= not w1192 and w1198;
w1393 <= not w1200 and w1392;
w1394 <= not w1337 and w1393;
w1395 <= not w1192 and not w1200;
w1396 <= not w1337 and w1395;
w1397 <= not w1198 and not w1396;
w1398 <= not w1394 and not w1397;
w1399 <= w577 and not w1379;
w1400 <= not w1389 and w1399;
w1401 <= not w1398 and not w1400;
w1402 <= not w1391 and not w1401;
w1403 <= not w460 and not w1402;
w1404 <= w1210 and not w1212;
w1405 <= not w1203 and w1404;
w1406 <= not w1337 and w1405;
w1407 <= not w1203 and not w1212;
w1408 <= not w1337 and w1407;
w1409 <= not w1210 and not w1408;
w1410 <= not w1406 and not w1409;
w1411 <= w460 and not w1391;
w1412 <= not w1401 and w1411;
w1413 <= not w1410 and not w1412;
w1414 <= not w1403 and not w1413;
w1415 <= not w356 and not w1414;
w1416 <= not w1215 and w1222;
w1417 <= not w1224 and w1416;
w1418 <= not w1337 and w1417;
w1419 <= not w1215 and not w1224;
w1420 <= not w1337 and w1419;
w1421 <= not w1222 and not w1420;
w1422 <= not w1418 and not w1421;
w1423 <= w356 and not w1403;
w1424 <= not w1413 and w1423;
w1425 <= not w1422 and not w1424;
w1426 <= not w1415 and not w1425;
w1427 <= not w264 and not w1426;
w1428 <= w1234 and not w1236;
w1429 <= not w1227 and w1428;
w1430 <= not w1337 and w1429;
w1431 <= not w1227 and not w1236;
w1432 <= not w1337 and w1431;
w1433 <= not w1234 and not w1432;
w1434 <= not w1430 and not w1433;
w1435 <= w264 and not w1415;
w1436 <= not w1425 and w1435;
w1437 <= not w1434 and not w1436;
w1438 <= not w1427 and not w1437;
w1439 <= not w184 and not w1438;
w1440 <= not w1239 and w1246;
w1441 <= not w1248 and w1440;
w1442 <= not w1337 and w1441;
w1443 <= not w1239 and not w1248;
w1444 <= not w1337 and w1443;
w1445 <= not w1246 and not w1444;
w1446 <= not w1442 and not w1445;
w1447 <= w184 and not w1427;
w1448 <= not w1437 and w1447;
w1449 <= not w1446 and not w1448;
w1450 <= not w1439 and not w1449;
w1451 <= not w115 and not w1450;
w1452 <= w1258 and not w1260;
w1453 <= not w1251 and w1452;
w1454 <= not w1337 and w1453;
w1455 <= not w1251 and not w1260;
w1456 <= not w1337 and w1455;
w1457 <= not w1258 and not w1456;
w1458 <= not w1454 and not w1457;
w1459 <= w115 and not w1439;
w1460 <= not w1449 and w1459;
w1461 <= not w1458 and not w1460;
w1462 <= not w1451 and not w1461;
w1463 <= not w60 and not w1462;
w1464 <= not w1263 and w1270;
w1465 <= not w1272 and w1464;
w1466 <= not w1337 and w1465;
w1467 <= not w1263 and not w1272;
w1468 <= not w1337 and w1467;
w1469 <= not w1270 and not w1468;
w1470 <= not w1466 and not w1469;
w1471 <= w60 and not w1451;
w1472 <= not w1461 and w1471;
w1473 <= not w1470 and not w1472;
w1474 <= not w1463 and not w1473;
w1475 <= not w22 and not w1474;
w1476 <= w1282 and not w1284;
w1477 <= not w1275 and w1476;
w1478 <= not w1337 and w1477;
w1479 <= not w1275 and not w1284;
w1480 <= not w1337 and w1479;
w1481 <= not w1282 and not w1480;
w1482 <= not w1478 and not w1481;
w1483 <= w22 and not w1463;
w1484 <= not w1473 and w1483;
w1485 <= not w1482 and not w1484;
w1486 <= not w1475 and not w1485;
w1487 <= not w5 and not w1486;
w1488 <= not w1287 and w1294;
w1489 <= not w1296 and w1488;
w1490 <= not w1337 and w1489;
w1491 <= not w1287 and not w1296;
w1492 <= not w1337 and w1491;
w1493 <= not w1294 and not w1492;
w1494 <= not w1490 and not w1493;
w1495 <= w5 and not w1475;
w1496 <= not w1485 and w1495;
w1497 <= not w1494 and not w1496;
w1498 <= not w1487 and not w1497;
w1499 <= w1306 and not w1308;
w1500 <= not w1299 and w1499;
w1501 <= not w1337 and w1500;
w1502 <= not w1299 and not w1308;
w1503 <= not w1337 and w1502;
w1504 <= not w1306 and not w1503;
w1505 <= not w1501 and not w1504;
w1506 <= not w1310 and not w1317;
w1507 <= not w1337 and w1506;
w1508 <= not w1325 and not w1507;
w1509 <= not w1505 and w1508;
w1510 <= not w1498 and w1509;
w1511 <= w0 and not w1510;
w1512 <= not w1487 and w1505;
w1513 <= not w1497 and w1512;
w1514 <= not w1317 and not w1337;
w1515 <= w1310 and not w1514;
w1516 <= not w0 and not w1506;
w1517 <= not w1515 and w1516;
w1518 <= not w1313 and not w1334;
w1519 <= not w1316 and w1518;
w1520 <= not w1329 and w1519;
w1521 <= not w1325 and w1520;
w1522 <= not w1323 and w1521;
w1523 <= not w1517 and not w1522;
w1524 <= not w1513 and w1523;
w1525 <= not w1511 and w1524;
w1526 <= a(96) and not w1525;
w1527 <= not a(94) and not a(95);
w1528 <= not a(96) and w1527;
w1529 <= not w1526 and not w1528;
w1530 <= not w1337 and not w1529;
w1531 <= not a(96) and not w1525;
w1532 <= a(97) and not w1531;
w1533 <= w1339 and not w1525;
w1534 <= not w1532 and not w1533;
w1535 <= not w1334 and not w1528;
w1536 <= not w1329 and w1535;
w1537 <= not w1325 and w1536;
w1538 <= not w1323 and w1537;
w1539 <= not w1526 and w1538;
w1540 <= w1534 and not w1539;
w1541 <= not w1530 and not w1540;
w1542 <= not w1161 and not w1541;
w1543 <= w1161 and not w1530;
w1544 <= not w1540 and w1543;
w1545 <= not w1337 and not w1522;
w1546 <= not w1517 and w1545;
w1547 <= not w1513 and w1546;
w1548 <= not w1511 and w1547;
w1549 <= not w1533 and not w1548;
w1550 <= a(98) and not w1549;
w1551 <= not a(98) and not w1548;
w1552 <= not w1533 and w1551;
w1553 <= not w1550 and not w1552;
w1554 <= not w1544 and not w1553;
w1555 <= not w1542 and not w1554;
w1556 <= not w997 and not w1555;
w1557 <= not w1342 and not w1347;
w1558 <= not w1351 and w1557;
w1559 <= not w1525 and w1558;
w1560 <= not w1525 and w1557;
w1561 <= w1351 and not w1560;
w1562 <= not w1559 and not w1561;
w1563 <= w997 and not w1542;
w1564 <= not w1554 and w1563;
w1565 <= not w1562 and not w1564;
w1566 <= not w1556 and not w1565;
w1567 <= not w845 and not w1566;
w1568 <= not w1356 and w1365;
w1569 <= not w1354 and w1568;
w1570 <= not w1525 and w1569;
w1571 <= not w1354 and not w1356;
w1572 <= not w1525 and w1571;
w1573 <= not w1365 and not w1572;
w1574 <= not w1570 and not w1573;
w1575 <= w845 and not w1556;
w1576 <= not w1565 and w1575;
w1577 <= not w1574 and not w1576;
w1578 <= not w1567 and not w1577;
w1579 <= not w705 and not w1578;
w1580 <= not w1368 and w1374;
w1581 <= not w1376 and w1580;
w1582 <= not w1525 and w1581;
w1583 <= not w1368 and not w1376;
w1584 <= not w1525 and w1583;
w1585 <= not w1374 and not w1584;
w1586 <= not w1582 and not w1585;
w1587 <= w705 and not w1567;
w1588 <= not w1577 and w1587;
w1589 <= not w1586 and not w1588;
w1590 <= not w1579 and not w1589;
w1591 <= not w577 and not w1590;
w1592 <= w1386 and not w1388;
w1593 <= not w1379 and w1592;
w1594 <= not w1525 and w1593;
w1595 <= not w1379 and not w1388;
w1596 <= not w1525 and w1595;
w1597 <= not w1386 and not w1596;
w1598 <= not w1594 and not w1597;
w1599 <= w577 and not w1579;
w1600 <= not w1589 and w1599;
w1601 <= not w1598 and not w1600;
w1602 <= not w1591 and not w1601;
w1603 <= not w460 and not w1602;
w1604 <= not w1391 and w1398;
w1605 <= not w1400 and w1604;
w1606 <= not w1525 and w1605;
w1607 <= not w1391 and not w1400;
w1608 <= not w1525 and w1607;
w1609 <= not w1398 and not w1608;
w1610 <= not w1606 and not w1609;
w1611 <= w460 and not w1591;
w1612 <= not w1601 and w1611;
w1613 <= not w1610 and not w1612;
w1614 <= not w1603 and not w1613;
w1615 <= not w356 and not w1614;
w1616 <= w1410 and not w1412;
w1617 <= not w1403 and w1616;
w1618 <= not w1525 and w1617;
w1619 <= not w1403 and not w1412;
w1620 <= not w1525 and w1619;
w1621 <= not w1410 and not w1620;
w1622 <= not w1618 and not w1621;
w1623 <= w356 and not w1603;
w1624 <= not w1613 and w1623;
w1625 <= not w1622 and not w1624;
w1626 <= not w1615 and not w1625;
w1627 <= not w264 and not w1626;
w1628 <= not w1415 and w1422;
w1629 <= not w1424 and w1628;
w1630 <= not w1525 and w1629;
w1631 <= not w1415 and not w1424;
w1632 <= not w1525 and w1631;
w1633 <= not w1422 and not w1632;
w1634 <= not w1630 and not w1633;
w1635 <= w264 and not w1615;
w1636 <= not w1625 and w1635;
w1637 <= not w1634 and not w1636;
w1638 <= not w1627 and not w1637;
w1639 <= not w184 and not w1638;
w1640 <= w1434 and not w1436;
w1641 <= not w1427 and w1640;
w1642 <= not w1525 and w1641;
w1643 <= not w1427 and not w1436;
w1644 <= not w1525 and w1643;
w1645 <= not w1434 and not w1644;
w1646 <= not w1642 and not w1645;
w1647 <= w184 and not w1627;
w1648 <= not w1637 and w1647;
w1649 <= not w1646 and not w1648;
w1650 <= not w1639 and not w1649;
w1651 <= not w115 and not w1650;
w1652 <= not w1439 and w1446;
w1653 <= not w1448 and w1652;
w1654 <= not w1525 and w1653;
w1655 <= not w1439 and not w1448;
w1656 <= not w1525 and w1655;
w1657 <= not w1446 and not w1656;
w1658 <= not w1654 and not w1657;
w1659 <= w115 and not w1639;
w1660 <= not w1649 and w1659;
w1661 <= not w1658 and not w1660;
w1662 <= not w1651 and not w1661;
w1663 <= not w60 and not w1662;
w1664 <= w1458 and not w1460;
w1665 <= not w1451 and w1664;
w1666 <= not w1525 and w1665;
w1667 <= not w1451 and not w1460;
w1668 <= not w1525 and w1667;
w1669 <= not w1458 and not w1668;
w1670 <= not w1666 and not w1669;
w1671 <= w60 and not w1651;
w1672 <= not w1661 and w1671;
w1673 <= not w1670 and not w1672;
w1674 <= not w1663 and not w1673;
w1675 <= not w22 and not w1674;
w1676 <= not w1463 and w1470;
w1677 <= not w1472 and w1676;
w1678 <= not w1525 and w1677;
w1679 <= not w1463 and not w1472;
w1680 <= not w1525 and w1679;
w1681 <= not w1470 and not w1680;
w1682 <= not w1678 and not w1681;
w1683 <= w22 and not w1663;
w1684 <= not w1673 and w1683;
w1685 <= not w1682 and not w1684;
w1686 <= not w1675 and not w1685;
w1687 <= not w5 and not w1686;
w1688 <= w1482 and not w1484;
w1689 <= not w1475 and w1688;
w1690 <= not w1525 and w1689;
w1691 <= not w1475 and not w1484;
w1692 <= not w1525 and w1691;
w1693 <= not w1482 and not w1692;
w1694 <= not w1690 and not w1693;
w1695 <= w5 and not w1675;
w1696 <= not w1685 and w1695;
w1697 <= not w1694 and not w1696;
w1698 <= not w1687 and not w1697;
w1699 <= not w1487 and w1494;
w1700 <= not w1496 and w1699;
w1701 <= not w1525 and w1700;
w1702 <= not w1487 and not w1496;
w1703 <= not w1525 and w1702;
w1704 <= not w1494 and not w1703;
w1705 <= not w1701 and not w1704;
w1706 <= not w1498 and not w1505;
w1707 <= not w1525 and w1706;
w1708 <= not w1513 and not w1707;
w1709 <= not w1705 and w1708;
w1710 <= not w1698 and w1709;
w1711 <= w0 and not w1710;
w1712 <= not w1687 and w1705;
w1713 <= not w1697 and w1712;
w1714 <= not w1505 and not w1525;
w1715 <= w1498 and not w1714;
w1716 <= not w0 and not w1706;
w1717 <= not w1715 and w1716;
w1718 <= not w1501 and not w1522;
w1719 <= not w1504 and w1718;
w1720 <= not w1517 and w1719;
w1721 <= not w1513 and w1720;
w1722 <= not w1511 and w1721;
w1723 <= not w1717 and not w1722;
w1724 <= not w1713 and w1723;
w1725 <= not w1711 and w1724;
w1726 <= a(94) and not w1725;
w1727 <= not a(92) and not a(93);
w1728 <= not a(94) and w1727;
w1729 <= not w1726 and not w1728;
w1730 <= not w1525 and not w1729;
w1731 <= not w1522 and not w1728;
w1732 <= not w1517 and w1731;
w1733 <= not w1513 and w1732;
w1734 <= not w1511 and w1733;
w1735 <= not w1726 and w1734;
w1736 <= not a(94) and not w1725;
w1737 <= a(95) and not w1736;
w1738 <= w1527 and not w1725;
w1739 <= not w1737 and not w1738;
w1740 <= not w1735 and w1739;
w1741 <= not w1730 and not w1740;
w1742 <= not w1337 and not w1741;
w1743 <= w1337 and not w1730;
w1744 <= not w1740 and w1743;
w1745 <= not w1525 and not w1722;
w1746 <= not w1717 and w1745;
w1747 <= not w1713 and w1746;
w1748 <= not w1711 and w1747;
w1749 <= not w1738 and not w1748;
w1750 <= a(96) and not w1749;
w1751 <= not a(96) and not w1748;
w1752 <= not w1738 and w1751;
w1753 <= not w1750 and not w1752;
w1754 <= not w1744 and not w1753;
w1755 <= not w1742 and not w1754;
w1756 <= not w1161 and not w1755;
w1757 <= w1161 and not w1742;
w1758 <= not w1754 and w1757;
w1759 <= not w1534 and not w1539;
w1760 <= not w1530 and w1759;
w1761 <= not w1725 and w1760;
w1762 <= not w1530 and not w1539;
w1763 <= not w1725 and w1762;
w1764 <= w1534 and not w1763;
w1765 <= not w1761 and not w1764;
w1766 <= not w1758 and not w1765;
w1767 <= not w1756 and not w1766;
w1768 <= not w997 and not w1767;
w1769 <= not w1544 and w1553;
w1770 <= not w1542 and w1769;
w1771 <= not w1725 and w1770;
w1772 <= not w1542 and not w1544;
w1773 <= not w1725 and w1772;
w1774 <= not w1553 and not w1773;
w1775 <= not w1771 and not w1774;
w1776 <= w997 and not w1756;
w1777 <= not w1766 and w1776;
w1778 <= not w1775 and not w1777;
w1779 <= not w1768 and not w1778;
w1780 <= not w845 and not w1779;
w1781 <= not w1556 and w1562;
w1782 <= not w1564 and w1781;
w1783 <= not w1725 and w1782;
w1784 <= not w1556 and not w1564;
w1785 <= not w1725 and w1784;
w1786 <= not w1562 and not w1785;
w1787 <= not w1783 and not w1786;
w1788 <= w845 and not w1768;
w1789 <= not w1778 and w1788;
w1790 <= not w1787 and not w1789;
w1791 <= not w1780 and not w1790;
w1792 <= not w705 and not w1791;
w1793 <= w1574 and not w1576;
w1794 <= not w1567 and w1793;
w1795 <= not w1725 and w1794;
w1796 <= not w1567 and not w1576;
w1797 <= not w1725 and w1796;
w1798 <= not w1574 and not w1797;
w1799 <= not w1795 and not w1798;
w1800 <= w705 and not w1780;
w1801 <= not w1790 and w1800;
w1802 <= not w1799 and not w1801;
w1803 <= not w1792 and not w1802;
w1804 <= not w577 and not w1803;
w1805 <= not w1579 and w1586;
w1806 <= not w1588 and w1805;
w1807 <= not w1725 and w1806;
w1808 <= not w1579 and not w1588;
w1809 <= not w1725 and w1808;
w1810 <= not w1586 and not w1809;
w1811 <= not w1807 and not w1810;
w1812 <= w577 and not w1792;
w1813 <= not w1802 and w1812;
w1814 <= not w1811 and not w1813;
w1815 <= not w1804 and not w1814;
w1816 <= not w460 and not w1815;
w1817 <= w1598 and not w1600;
w1818 <= not w1591 and w1817;
w1819 <= not w1725 and w1818;
w1820 <= not w1591 and not w1600;
w1821 <= not w1725 and w1820;
w1822 <= not w1598 and not w1821;
w1823 <= not w1819 and not w1822;
w1824 <= w460 and not w1804;
w1825 <= not w1814 and w1824;
w1826 <= not w1823 and not w1825;
w1827 <= not w1816 and not w1826;
w1828 <= not w356 and not w1827;
w1829 <= not w1603 and w1610;
w1830 <= not w1612 and w1829;
w1831 <= not w1725 and w1830;
w1832 <= not w1603 and not w1612;
w1833 <= not w1725 and w1832;
w1834 <= not w1610 and not w1833;
w1835 <= not w1831 and not w1834;
w1836 <= w356 and not w1816;
w1837 <= not w1826 and w1836;
w1838 <= not w1835 and not w1837;
w1839 <= not w1828 and not w1838;
w1840 <= not w264 and not w1839;
w1841 <= w1622 and not w1624;
w1842 <= not w1615 and w1841;
w1843 <= not w1725 and w1842;
w1844 <= not w1615 and not w1624;
w1845 <= not w1725 and w1844;
w1846 <= not w1622 and not w1845;
w1847 <= not w1843 and not w1846;
w1848 <= w264 and not w1828;
w1849 <= not w1838 and w1848;
w1850 <= not w1847 and not w1849;
w1851 <= not w1840 and not w1850;
w1852 <= not w184 and not w1851;
w1853 <= not w1627 and w1634;
w1854 <= not w1636 and w1853;
w1855 <= not w1725 and w1854;
w1856 <= not w1627 and not w1636;
w1857 <= not w1725 and w1856;
w1858 <= not w1634 and not w1857;
w1859 <= not w1855 and not w1858;
w1860 <= w184 and not w1840;
w1861 <= not w1850 and w1860;
w1862 <= not w1859 and not w1861;
w1863 <= not w1852 and not w1862;
w1864 <= not w115 and not w1863;
w1865 <= w1646 and not w1648;
w1866 <= not w1639 and w1865;
w1867 <= not w1725 and w1866;
w1868 <= not w1639 and not w1648;
w1869 <= not w1725 and w1868;
w1870 <= not w1646 and not w1869;
w1871 <= not w1867 and not w1870;
w1872 <= w115 and not w1852;
w1873 <= not w1862 and w1872;
w1874 <= not w1871 and not w1873;
w1875 <= not w1864 and not w1874;
w1876 <= not w60 and not w1875;
w1877 <= not w1651 and w1658;
w1878 <= not w1660 and w1877;
w1879 <= not w1725 and w1878;
w1880 <= not w1651 and not w1660;
w1881 <= not w1725 and w1880;
w1882 <= not w1658 and not w1881;
w1883 <= not w1879 and not w1882;
w1884 <= w60 and not w1864;
w1885 <= not w1874 and w1884;
w1886 <= not w1883 and not w1885;
w1887 <= not w1876 and not w1886;
w1888 <= not w22 and not w1887;
w1889 <= w1670 and not w1672;
w1890 <= not w1663 and w1889;
w1891 <= not w1725 and w1890;
w1892 <= not w1663 and not w1672;
w1893 <= not w1725 and w1892;
w1894 <= not w1670 and not w1893;
w1895 <= not w1891 and not w1894;
w1896 <= w22 and not w1876;
w1897 <= not w1886 and w1896;
w1898 <= not w1895 and not w1897;
w1899 <= not w1888 and not w1898;
w1900 <= not w5 and not w1899;
w1901 <= not w1675 and w1682;
w1902 <= not w1684 and w1901;
w1903 <= not w1725 and w1902;
w1904 <= not w1675 and not w1684;
w1905 <= not w1725 and w1904;
w1906 <= not w1682 and not w1905;
w1907 <= not w1903 and not w1906;
w1908 <= w5 and not w1888;
w1909 <= not w1898 and w1908;
w1910 <= not w1907 and not w1909;
w1911 <= not w1900 and not w1910;
w1912 <= w1694 and not w1696;
w1913 <= not w1687 and w1912;
w1914 <= not w1725 and w1913;
w1915 <= not w1687 and not w1696;
w1916 <= not w1725 and w1915;
w1917 <= not w1694 and not w1916;
w1918 <= not w1914 and not w1917;
w1919 <= not w1698 and not w1705;
w1920 <= not w1725 and w1919;
w1921 <= not w1713 and not w1920;
w1922 <= not w1918 and w1921;
w1923 <= not w1911 and w1922;
w1924 <= w0 and not w1923;
w1925 <= not w1900 and w1918;
w1926 <= not w1910 and w1925;
w1927 <= not w1705 and not w1725;
w1928 <= w1698 and not w1927;
w1929 <= not w0 and not w1919;
w1930 <= not w1928 and w1929;
w1931 <= not w1701 and not w1722;
w1932 <= not w1704 and w1931;
w1933 <= not w1717 and w1932;
w1934 <= not w1713 and w1933;
w1935 <= not w1711 and w1934;
w1936 <= not w1930 and not w1935;
w1937 <= not w1926 and w1936;
w1938 <= not w1924 and w1937;
w1939 <= a(92) and not w1938;
w1940 <= not a(90) and not a(91);
w1941 <= not a(92) and w1940;
w1942 <= not w1939 and not w1941;
w1943 <= not w1725 and not w1942;
w1944 <= not w1722 and not w1941;
w1945 <= not w1717 and w1944;
w1946 <= not w1713 and w1945;
w1947 <= not w1711 and w1946;
w1948 <= not w1939 and w1947;
w1949 <= not a(92) and not w1938;
w1950 <= a(93) and not w1949;
w1951 <= w1727 and not w1938;
w1952 <= not w1950 and not w1951;
w1953 <= not w1948 and w1952;
w1954 <= not w1943 and not w1953;
w1955 <= not w1525 and not w1954;
w1956 <= w1525 and not w1943;
w1957 <= not w1953 and w1956;
w1958 <= not w1725 and not w1935;
w1959 <= not w1930 and w1958;
w1960 <= not w1926 and w1959;
w1961 <= not w1924 and w1960;
w1962 <= not w1951 and not w1961;
w1963 <= a(94) and not w1962;
w1964 <= not a(94) and not w1961;
w1965 <= not w1951 and w1964;
w1966 <= not w1963 and not w1965;
w1967 <= not w1957 and not w1966;
w1968 <= not w1955 and not w1967;
w1969 <= not w1337 and not w1968;
w1970 <= not w1730 and not w1735;
w1971 <= not w1739 and w1970;
w1972 <= not w1938 and w1971;
w1973 <= not w1938 and w1970;
w1974 <= w1739 and not w1973;
w1975 <= not w1972 and not w1974;
w1976 <= w1337 and not w1955;
w1977 <= not w1967 and w1976;
w1978 <= not w1975 and not w1977;
w1979 <= not w1969 and not w1978;
w1980 <= not w1161 and not w1979;
w1981 <= not w1744 and w1753;
w1982 <= not w1742 and w1981;
w1983 <= not w1938 and w1982;
w1984 <= not w1742 and not w1744;
w1985 <= not w1938 and w1984;
w1986 <= not w1753 and not w1985;
w1987 <= not w1983 and not w1986;
w1988 <= w1161 and not w1969;
w1989 <= not w1978 and w1988;
w1990 <= not w1987 and not w1989;
w1991 <= not w1980 and not w1990;
w1992 <= not w997 and not w1991;
w1993 <= w997 and not w1980;
w1994 <= not w1990 and w1993;
w1995 <= not w1756 and w1765;
w1996 <= not w1758 and w1995;
w1997 <= not w1938 and w1996;
w1998 <= not w1756 and not w1758;
w1999 <= not w1938 and w1998;
w2000 <= not w1765 and not w1999;
w2001 <= not w1997 and not w2000;
w2002 <= not w1994 and not w2001;
w2003 <= not w1992 and not w2002;
w2004 <= not w845 and not w2003;
w2005 <= w1775 and not w1777;
w2006 <= not w1768 and w2005;
w2007 <= not w1938 and w2006;
w2008 <= not w1768 and not w1777;
w2009 <= not w1938 and w2008;
w2010 <= not w1775 and not w2009;
w2011 <= not w2007 and not w2010;
w2012 <= w845 and not w1992;
w2013 <= not w2002 and w2012;
w2014 <= not w2011 and not w2013;
w2015 <= not w2004 and not w2014;
w2016 <= not w705 and not w2015;
w2017 <= not w1780 and w1787;
w2018 <= not w1789 and w2017;
w2019 <= not w1938 and w2018;
w2020 <= not w1780 and not w1789;
w2021 <= not w1938 and w2020;
w2022 <= not w1787 and not w2021;
w2023 <= not w2019 and not w2022;
w2024 <= w705 and not w2004;
w2025 <= not w2014 and w2024;
w2026 <= not w2023 and not w2025;
w2027 <= not w2016 and not w2026;
w2028 <= not w577 and not w2027;
w2029 <= w1799 and not w1801;
w2030 <= not w1792 and w2029;
w2031 <= not w1938 and w2030;
w2032 <= not w1792 and not w1801;
w2033 <= not w1938 and w2032;
w2034 <= not w1799 and not w2033;
w2035 <= not w2031 and not w2034;
w2036 <= w577 and not w2016;
w2037 <= not w2026 and w2036;
w2038 <= not w2035 and not w2037;
w2039 <= not w2028 and not w2038;
w2040 <= not w460 and not w2039;
w2041 <= not w1804 and w1811;
w2042 <= not w1813 and w2041;
w2043 <= not w1938 and w2042;
w2044 <= not w1804 and not w1813;
w2045 <= not w1938 and w2044;
w2046 <= not w1811 and not w2045;
w2047 <= not w2043 and not w2046;
w2048 <= w460 and not w2028;
w2049 <= not w2038 and w2048;
w2050 <= not w2047 and not w2049;
w2051 <= not w2040 and not w2050;
w2052 <= not w356 and not w2051;
w2053 <= w1823 and not w1825;
w2054 <= not w1816 and w2053;
w2055 <= not w1938 and w2054;
w2056 <= not w1816 and not w1825;
w2057 <= not w1938 and w2056;
w2058 <= not w1823 and not w2057;
w2059 <= not w2055 and not w2058;
w2060 <= w356 and not w2040;
w2061 <= not w2050 and w2060;
w2062 <= not w2059 and not w2061;
w2063 <= not w2052 and not w2062;
w2064 <= not w264 and not w2063;
w2065 <= not w1828 and w1835;
w2066 <= not w1837 and w2065;
w2067 <= not w1938 and w2066;
w2068 <= not w1828 and not w1837;
w2069 <= not w1938 and w2068;
w2070 <= not w1835 and not w2069;
w2071 <= not w2067 and not w2070;
w2072 <= w264 and not w2052;
w2073 <= not w2062 and w2072;
w2074 <= not w2071 and not w2073;
w2075 <= not w2064 and not w2074;
w2076 <= not w184 and not w2075;
w2077 <= w1847 and not w1849;
w2078 <= not w1840 and w2077;
w2079 <= not w1938 and w2078;
w2080 <= not w1840 and not w1849;
w2081 <= not w1938 and w2080;
w2082 <= not w1847 and not w2081;
w2083 <= not w2079 and not w2082;
w2084 <= w184 and not w2064;
w2085 <= not w2074 and w2084;
w2086 <= not w2083 and not w2085;
w2087 <= not w2076 and not w2086;
w2088 <= not w115 and not w2087;
w2089 <= not w1852 and w1859;
w2090 <= not w1861 and w2089;
w2091 <= not w1938 and w2090;
w2092 <= not w1852 and not w1861;
w2093 <= not w1938 and w2092;
w2094 <= not w1859 and not w2093;
w2095 <= not w2091 and not w2094;
w2096 <= w115 and not w2076;
w2097 <= not w2086 and w2096;
w2098 <= not w2095 and not w2097;
w2099 <= not w2088 and not w2098;
w2100 <= not w60 and not w2099;
w2101 <= w1871 and not w1873;
w2102 <= not w1864 and w2101;
w2103 <= not w1938 and w2102;
w2104 <= not w1864 and not w1873;
w2105 <= not w1938 and w2104;
w2106 <= not w1871 and not w2105;
w2107 <= not w2103 and not w2106;
w2108 <= w60 and not w2088;
w2109 <= not w2098 and w2108;
w2110 <= not w2107 and not w2109;
w2111 <= not w2100 and not w2110;
w2112 <= not w22 and not w2111;
w2113 <= not w1876 and w1883;
w2114 <= not w1885 and w2113;
w2115 <= not w1938 and w2114;
w2116 <= not w1876 and not w1885;
w2117 <= not w1938 and w2116;
w2118 <= not w1883 and not w2117;
w2119 <= not w2115 and not w2118;
w2120 <= w22 and not w2100;
w2121 <= not w2110 and w2120;
w2122 <= not w2119 and not w2121;
w2123 <= not w2112 and not w2122;
w2124 <= not w5 and not w2123;
w2125 <= w1895 and not w1897;
w2126 <= not w1888 and w2125;
w2127 <= not w1938 and w2126;
w2128 <= not w1888 and not w1897;
w2129 <= not w1938 and w2128;
w2130 <= not w1895 and not w2129;
w2131 <= not w2127 and not w2130;
w2132 <= w5 and not w2112;
w2133 <= not w2122 and w2132;
w2134 <= not w2131 and not w2133;
w2135 <= not w2124 and not w2134;
w2136 <= not w1900 and w1907;
w2137 <= not w1909 and w2136;
w2138 <= not w1938 and w2137;
w2139 <= not w1900 and not w1909;
w2140 <= not w1938 and w2139;
w2141 <= not w1907 and not w2140;
w2142 <= not w2138 and not w2141;
w2143 <= not w1911 and not w1918;
w2144 <= not w1938 and w2143;
w2145 <= not w1926 and not w2144;
w2146 <= not w2142 and w2145;
w2147 <= not w2135 and w2146;
w2148 <= w0 and not w2147;
w2149 <= not w2124 and w2142;
w2150 <= not w2134 and w2149;
w2151 <= not w1918 and not w1938;
w2152 <= w1911 and not w2151;
w2153 <= not w0 and not w2143;
w2154 <= not w2152 and w2153;
w2155 <= not w1914 and not w1935;
w2156 <= not w1917 and w2155;
w2157 <= not w1930 and w2156;
w2158 <= not w1926 and w2157;
w2159 <= not w1924 and w2158;
w2160 <= not w2154 and not w2159;
w2161 <= not w2150 and w2160;
w2162 <= not w2148 and w2161;
w2163 <= a(90) and not w2162;
w2164 <= not a(88) and not a(89);
w2165 <= not a(90) and w2164;
w2166 <= not w2163 and not w2165;
w2167 <= not w1938 and not w2166;
w2168 <= not w1935 and not w2165;
w2169 <= not w1930 and w2168;
w2170 <= not w1926 and w2169;
w2171 <= not w1924 and w2170;
w2172 <= not w2163 and w2171;
w2173 <= not a(90) and not w2162;
w2174 <= a(91) and not w2173;
w2175 <= w1940 and not w2162;
w2176 <= not w2174 and not w2175;
w2177 <= not w2172 and w2176;
w2178 <= not w2167 and not w2177;
w2179 <= not w1725 and not w2178;
w2180 <= w1725 and not w2167;
w2181 <= not w2177 and w2180;
w2182 <= not w1938 and not w2159;
w2183 <= not w2154 and w2182;
w2184 <= not w2150 and w2183;
w2185 <= not w2148 and w2184;
w2186 <= not w2175 and not w2185;
w2187 <= a(92) and not w2186;
w2188 <= not a(92) and not w2185;
w2189 <= not w2175 and w2188;
w2190 <= not w2187 and not w2189;
w2191 <= not w2181 and not w2190;
w2192 <= not w2179 and not w2191;
w2193 <= not w1525 and not w2192;
w2194 <= not w1943 and not w1948;
w2195 <= not w1952 and w2194;
w2196 <= not w2162 and w2195;
w2197 <= not w2162 and w2194;
w2198 <= w1952 and not w2197;
w2199 <= not w2196 and not w2198;
w2200 <= w1525 and not w2179;
w2201 <= not w2191 and w2200;
w2202 <= not w2199 and not w2201;
w2203 <= not w2193 and not w2202;
w2204 <= not w1337 and not w2203;
w2205 <= not w1957 and w1966;
w2206 <= not w1955 and w2205;
w2207 <= not w2162 and w2206;
w2208 <= not w1955 and not w1957;
w2209 <= not w2162 and w2208;
w2210 <= not w1966 and not w2209;
w2211 <= not w2207 and not w2210;
w2212 <= w1337 and not w2193;
w2213 <= not w2202 and w2212;
w2214 <= not w2211 and not w2213;
w2215 <= not w2204 and not w2214;
w2216 <= not w1161 and not w2215;
w2217 <= not w1969 and w1975;
w2218 <= not w1977 and w2217;
w2219 <= not w2162 and w2218;
w2220 <= not w1969 and not w1977;
w2221 <= not w2162 and w2220;
w2222 <= not w1975 and not w2221;
w2223 <= not w2219 and not w2222;
w2224 <= w1161 and not w2204;
w2225 <= not w2214 and w2224;
w2226 <= not w2223 and not w2225;
w2227 <= not w2216 and not w2226;
w2228 <= not w997 and not w2227;
w2229 <= w1987 and not w1989;
w2230 <= not w1980 and w2229;
w2231 <= not w2162 and w2230;
w2232 <= not w1980 and not w1989;
w2233 <= not w2162 and w2232;
w2234 <= not w1987 and not w2233;
w2235 <= not w2231 and not w2234;
w2236 <= w997 and not w2216;
w2237 <= not w2226 and w2236;
w2238 <= not w2235 and not w2237;
w2239 <= not w2228 and not w2238;
w2240 <= not w845 and not w2239;
w2241 <= w845 and not w2228;
w2242 <= not w2238 and w2241;
w2243 <= not w1992 and w2001;
w2244 <= not w1994 and w2243;
w2245 <= not w2162 and w2244;
w2246 <= not w1992 and not w1994;
w2247 <= not w2162 and w2246;
w2248 <= not w2001 and not w2247;
w2249 <= not w2245 and not w2248;
w2250 <= not w2242 and not w2249;
w2251 <= not w2240 and not w2250;
w2252 <= not w705 and not w2251;
w2253 <= w2011 and not w2013;
w2254 <= not w2004 and w2253;
w2255 <= not w2162 and w2254;
w2256 <= not w2004 and not w2013;
w2257 <= not w2162 and w2256;
w2258 <= not w2011 and not w2257;
w2259 <= not w2255 and not w2258;
w2260 <= w705 and not w2240;
w2261 <= not w2250 and w2260;
w2262 <= not w2259 and not w2261;
w2263 <= not w2252 and not w2262;
w2264 <= not w577 and not w2263;
w2265 <= not w2016 and w2023;
w2266 <= not w2025 and w2265;
w2267 <= not w2162 and w2266;
w2268 <= not w2016 and not w2025;
w2269 <= not w2162 and w2268;
w2270 <= not w2023 and not w2269;
w2271 <= not w2267 and not w2270;
w2272 <= w577 and not w2252;
w2273 <= not w2262 and w2272;
w2274 <= not w2271 and not w2273;
w2275 <= not w2264 and not w2274;
w2276 <= not w460 and not w2275;
w2277 <= w2035 and not w2037;
w2278 <= not w2028 and w2277;
w2279 <= not w2162 and w2278;
w2280 <= not w2028 and not w2037;
w2281 <= not w2162 and w2280;
w2282 <= not w2035 and not w2281;
w2283 <= not w2279 and not w2282;
w2284 <= w460 and not w2264;
w2285 <= not w2274 and w2284;
w2286 <= not w2283 and not w2285;
w2287 <= not w2276 and not w2286;
w2288 <= not w356 and not w2287;
w2289 <= not w2040 and w2047;
w2290 <= not w2049 and w2289;
w2291 <= not w2162 and w2290;
w2292 <= not w2040 and not w2049;
w2293 <= not w2162 and w2292;
w2294 <= not w2047 and not w2293;
w2295 <= not w2291 and not w2294;
w2296 <= w356 and not w2276;
w2297 <= not w2286 and w2296;
w2298 <= not w2295 and not w2297;
w2299 <= not w2288 and not w2298;
w2300 <= not w264 and not w2299;
w2301 <= w2059 and not w2061;
w2302 <= not w2052 and w2301;
w2303 <= not w2162 and w2302;
w2304 <= not w2052 and not w2061;
w2305 <= not w2162 and w2304;
w2306 <= not w2059 and not w2305;
w2307 <= not w2303 and not w2306;
w2308 <= w264 and not w2288;
w2309 <= not w2298 and w2308;
w2310 <= not w2307 and not w2309;
w2311 <= not w2300 and not w2310;
w2312 <= not w184 and not w2311;
w2313 <= not w2064 and w2071;
w2314 <= not w2073 and w2313;
w2315 <= not w2162 and w2314;
w2316 <= not w2064 and not w2073;
w2317 <= not w2162 and w2316;
w2318 <= not w2071 and not w2317;
w2319 <= not w2315 and not w2318;
w2320 <= w184 and not w2300;
w2321 <= not w2310 and w2320;
w2322 <= not w2319 and not w2321;
w2323 <= not w2312 and not w2322;
w2324 <= not w115 and not w2323;
w2325 <= w2083 and not w2085;
w2326 <= not w2076 and w2325;
w2327 <= not w2162 and w2326;
w2328 <= not w2076 and not w2085;
w2329 <= not w2162 and w2328;
w2330 <= not w2083 and not w2329;
w2331 <= not w2327 and not w2330;
w2332 <= w115 and not w2312;
w2333 <= not w2322 and w2332;
w2334 <= not w2331 and not w2333;
w2335 <= not w2324 and not w2334;
w2336 <= not w60 and not w2335;
w2337 <= not w2088 and w2095;
w2338 <= not w2097 and w2337;
w2339 <= not w2162 and w2338;
w2340 <= not w2088 and not w2097;
w2341 <= not w2162 and w2340;
w2342 <= not w2095 and not w2341;
w2343 <= not w2339 and not w2342;
w2344 <= w60 and not w2324;
w2345 <= not w2334 and w2344;
w2346 <= not w2343 and not w2345;
w2347 <= not w2336 and not w2346;
w2348 <= not w22 and not w2347;
w2349 <= w2107 and not w2109;
w2350 <= not w2100 and w2349;
w2351 <= not w2162 and w2350;
w2352 <= not w2100 and not w2109;
w2353 <= not w2162 and w2352;
w2354 <= not w2107 and not w2353;
w2355 <= not w2351 and not w2354;
w2356 <= w22 and not w2336;
w2357 <= not w2346 and w2356;
w2358 <= not w2355 and not w2357;
w2359 <= not w2348 and not w2358;
w2360 <= not w5 and not w2359;
w2361 <= not w2112 and w2119;
w2362 <= not w2121 and w2361;
w2363 <= not w2162 and w2362;
w2364 <= not w2112 and not w2121;
w2365 <= not w2162 and w2364;
w2366 <= not w2119 and not w2365;
w2367 <= not w2363 and not w2366;
w2368 <= w5 and not w2348;
w2369 <= not w2358 and w2368;
w2370 <= not w2367 and not w2369;
w2371 <= not w2360 and not w2370;
w2372 <= w2131 and not w2133;
w2373 <= not w2124 and w2372;
w2374 <= not w2162 and w2373;
w2375 <= not w2124 and not w2133;
w2376 <= not w2162 and w2375;
w2377 <= not w2131 and not w2376;
w2378 <= not w2374 and not w2377;
w2379 <= not w2135 and not w2142;
w2380 <= not w2162 and w2379;
w2381 <= not w2150 and not w2380;
w2382 <= not w2378 and w2381;
w2383 <= not w2371 and w2382;
w2384 <= w0 and not w2383;
w2385 <= not w2360 and w2378;
w2386 <= not w2370 and w2385;
w2387 <= not w2142 and not w2162;
w2388 <= w2135 and not w2387;
w2389 <= not w0 and not w2379;
w2390 <= not w2388 and w2389;
w2391 <= not w2138 and not w2159;
w2392 <= not w2141 and w2391;
w2393 <= not w2154 and w2392;
w2394 <= not w2150 and w2393;
w2395 <= not w2148 and w2394;
w2396 <= not w2390 and not w2395;
w2397 <= not w2386 and w2396;
w2398 <= not w2384 and w2397;
w2399 <= a(88) and not w2398;
w2400 <= not a(86) and not a(87);
w2401 <= not a(88) and w2400;
w2402 <= not w2399 and not w2401;
w2403 <= not w2162 and not w2402;
w2404 <= not w2159 and not w2401;
w2405 <= not w2154 and w2404;
w2406 <= not w2150 and w2405;
w2407 <= not w2148 and w2406;
w2408 <= not w2399 and w2407;
w2409 <= not a(88) and not w2398;
w2410 <= a(89) and not w2409;
w2411 <= w2164 and not w2398;
w2412 <= not w2410 and not w2411;
w2413 <= not w2408 and w2412;
w2414 <= not w2403 and not w2413;
w2415 <= not w1938 and not w2414;
w2416 <= w1938 and not w2403;
w2417 <= not w2413 and w2416;
w2418 <= not w2162 and not w2395;
w2419 <= not w2390 and w2418;
w2420 <= not w2386 and w2419;
w2421 <= not w2384 and w2420;
w2422 <= not w2411 and not w2421;
w2423 <= a(90) and not w2422;
w2424 <= not a(90) and not w2421;
w2425 <= not w2411 and w2424;
w2426 <= not w2423 and not w2425;
w2427 <= not w2417 and not w2426;
w2428 <= not w2415 and not w2427;
w2429 <= not w1725 and not w2428;
w2430 <= not w2167 and not w2172;
w2431 <= not w2176 and w2430;
w2432 <= not w2398 and w2431;
w2433 <= not w2398 and w2430;
w2434 <= w2176 and not w2433;
w2435 <= not w2432 and not w2434;
w2436 <= w1725 and not w2415;
w2437 <= not w2427 and w2436;
w2438 <= not w2435 and not w2437;
w2439 <= not w2429 and not w2438;
w2440 <= not w1525 and not w2439;
w2441 <= not w2181 and w2190;
w2442 <= not w2179 and w2441;
w2443 <= not w2398 and w2442;
w2444 <= not w2179 and not w2181;
w2445 <= not w2398 and w2444;
w2446 <= not w2190 and not w2445;
w2447 <= not w2443 and not w2446;
w2448 <= w1525 and not w2429;
w2449 <= not w2438 and w2448;
w2450 <= not w2447 and not w2449;
w2451 <= not w2440 and not w2450;
w2452 <= not w1337 and not w2451;
w2453 <= not w2193 and w2199;
w2454 <= not w2201 and w2453;
w2455 <= not w2398 and w2454;
w2456 <= not w2193 and not w2201;
w2457 <= not w2398 and w2456;
w2458 <= not w2199 and not w2457;
w2459 <= not w2455 and not w2458;
w2460 <= w1337 and not w2440;
w2461 <= not w2450 and w2460;
w2462 <= not w2459 and not w2461;
w2463 <= not w2452 and not w2462;
w2464 <= not w1161 and not w2463;
w2465 <= w2211 and not w2213;
w2466 <= not w2204 and w2465;
w2467 <= not w2398 and w2466;
w2468 <= not w2204 and not w2213;
w2469 <= not w2398 and w2468;
w2470 <= not w2211 and not w2469;
w2471 <= not w2467 and not w2470;
w2472 <= w1161 and not w2452;
w2473 <= not w2462 and w2472;
w2474 <= not w2471 and not w2473;
w2475 <= not w2464 and not w2474;
w2476 <= not w997 and not w2475;
w2477 <= not w2216 and w2223;
w2478 <= not w2225 and w2477;
w2479 <= not w2398 and w2478;
w2480 <= not w2216 and not w2225;
w2481 <= not w2398 and w2480;
w2482 <= not w2223 and not w2481;
w2483 <= not w2479 and not w2482;
w2484 <= w997 and not w2464;
w2485 <= not w2474 and w2484;
w2486 <= not w2483 and not w2485;
w2487 <= not w2476 and not w2486;
w2488 <= not w845 and not w2487;
w2489 <= w2235 and not w2237;
w2490 <= not w2228 and w2489;
w2491 <= not w2398 and w2490;
w2492 <= not w2228 and not w2237;
w2493 <= not w2398 and w2492;
w2494 <= not w2235 and not w2493;
w2495 <= not w2491 and not w2494;
w2496 <= w845 and not w2476;
w2497 <= not w2486 and w2496;
w2498 <= not w2495 and not w2497;
w2499 <= not w2488 and not w2498;
w2500 <= not w705 and not w2499;
w2501 <= w705 and not w2488;
w2502 <= not w2498 and w2501;
w2503 <= not w2240 and w2249;
w2504 <= not w2242 and w2503;
w2505 <= not w2398 and w2504;
w2506 <= not w2240 and not w2242;
w2507 <= not w2398 and w2506;
w2508 <= not w2249 and not w2507;
w2509 <= not w2505 and not w2508;
w2510 <= not w2502 and not w2509;
w2511 <= not w2500 and not w2510;
w2512 <= not w577 and not w2511;
w2513 <= w2259 and not w2261;
w2514 <= not w2252 and w2513;
w2515 <= not w2398 and w2514;
w2516 <= not w2252 and not w2261;
w2517 <= not w2398 and w2516;
w2518 <= not w2259 and not w2517;
w2519 <= not w2515 and not w2518;
w2520 <= w577 and not w2500;
w2521 <= not w2510 and w2520;
w2522 <= not w2519 and not w2521;
w2523 <= not w2512 and not w2522;
w2524 <= not w460 and not w2523;
w2525 <= not w2264 and w2271;
w2526 <= not w2273 and w2525;
w2527 <= not w2398 and w2526;
w2528 <= not w2264 and not w2273;
w2529 <= not w2398 and w2528;
w2530 <= not w2271 and not w2529;
w2531 <= not w2527 and not w2530;
w2532 <= w460 and not w2512;
w2533 <= not w2522 and w2532;
w2534 <= not w2531 and not w2533;
w2535 <= not w2524 and not w2534;
w2536 <= not w356 and not w2535;
w2537 <= w2283 and not w2285;
w2538 <= not w2276 and w2537;
w2539 <= not w2398 and w2538;
w2540 <= not w2276 and not w2285;
w2541 <= not w2398 and w2540;
w2542 <= not w2283 and not w2541;
w2543 <= not w2539 and not w2542;
w2544 <= w356 and not w2524;
w2545 <= not w2534 and w2544;
w2546 <= not w2543 and not w2545;
w2547 <= not w2536 and not w2546;
w2548 <= not w264 and not w2547;
w2549 <= not w2288 and w2295;
w2550 <= not w2297 and w2549;
w2551 <= not w2398 and w2550;
w2552 <= not w2288 and not w2297;
w2553 <= not w2398 and w2552;
w2554 <= not w2295 and not w2553;
w2555 <= not w2551 and not w2554;
w2556 <= w264 and not w2536;
w2557 <= not w2546 and w2556;
w2558 <= not w2555 and not w2557;
w2559 <= not w2548 and not w2558;
w2560 <= not w184 and not w2559;
w2561 <= w2307 and not w2309;
w2562 <= not w2300 and w2561;
w2563 <= not w2398 and w2562;
w2564 <= not w2300 and not w2309;
w2565 <= not w2398 and w2564;
w2566 <= not w2307 and not w2565;
w2567 <= not w2563 and not w2566;
w2568 <= w184 and not w2548;
w2569 <= not w2558 and w2568;
w2570 <= not w2567 and not w2569;
w2571 <= not w2560 and not w2570;
w2572 <= not w115 and not w2571;
w2573 <= not w2312 and w2319;
w2574 <= not w2321 and w2573;
w2575 <= not w2398 and w2574;
w2576 <= not w2312 and not w2321;
w2577 <= not w2398 and w2576;
w2578 <= not w2319 and not w2577;
w2579 <= not w2575 and not w2578;
w2580 <= w115 and not w2560;
w2581 <= not w2570 and w2580;
w2582 <= not w2579 and not w2581;
w2583 <= not w2572 and not w2582;
w2584 <= not w60 and not w2583;
w2585 <= w2331 and not w2333;
w2586 <= not w2324 and w2585;
w2587 <= not w2398 and w2586;
w2588 <= not w2324 and not w2333;
w2589 <= not w2398 and w2588;
w2590 <= not w2331 and not w2589;
w2591 <= not w2587 and not w2590;
w2592 <= w60 and not w2572;
w2593 <= not w2582 and w2592;
w2594 <= not w2591 and not w2593;
w2595 <= not w2584 and not w2594;
w2596 <= not w22 and not w2595;
w2597 <= not w2336 and w2343;
w2598 <= not w2345 and w2597;
w2599 <= not w2398 and w2598;
w2600 <= not w2336 and not w2345;
w2601 <= not w2398 and w2600;
w2602 <= not w2343 and not w2601;
w2603 <= not w2599 and not w2602;
w2604 <= w22 and not w2584;
w2605 <= not w2594 and w2604;
w2606 <= not w2603 and not w2605;
w2607 <= not w2596 and not w2606;
w2608 <= not w5 and not w2607;
w2609 <= w2355 and not w2357;
w2610 <= not w2348 and w2609;
w2611 <= not w2398 and w2610;
w2612 <= not w2348 and not w2357;
w2613 <= not w2398 and w2612;
w2614 <= not w2355 and not w2613;
w2615 <= not w2611 and not w2614;
w2616 <= w5 and not w2596;
w2617 <= not w2606 and w2616;
w2618 <= not w2615 and not w2617;
w2619 <= not w2608 and not w2618;
w2620 <= not w2360 and w2367;
w2621 <= not w2369 and w2620;
w2622 <= not w2398 and w2621;
w2623 <= not w2360 and not w2369;
w2624 <= not w2398 and w2623;
w2625 <= not w2367 and not w2624;
w2626 <= not w2622 and not w2625;
w2627 <= not w2371 and not w2378;
w2628 <= not w2398 and w2627;
w2629 <= not w2386 and not w2628;
w2630 <= not w2626 and w2629;
w2631 <= not w2619 and w2630;
w2632 <= w0 and not w2631;
w2633 <= not w2608 and w2626;
w2634 <= not w2618 and w2633;
w2635 <= not w2378 and not w2398;
w2636 <= w2371 and not w2635;
w2637 <= not w0 and not w2627;
w2638 <= not w2636 and w2637;
w2639 <= not w2374 and not w2395;
w2640 <= not w2377 and w2639;
w2641 <= not w2390 and w2640;
w2642 <= not w2386 and w2641;
w2643 <= not w2384 and w2642;
w2644 <= not w2638 and not w2643;
w2645 <= not w2634 and w2644;
w2646 <= not w2632 and w2645;
w2647 <= a(86) and not w2646;
w2648 <= not a(84) and not a(85);
w2649 <= not a(86) and w2648;
w2650 <= not w2647 and not w2649;
w2651 <= not w2398 and not w2650;
w2652 <= not w2395 and not w2649;
w2653 <= not w2390 and w2652;
w2654 <= not w2386 and w2653;
w2655 <= not w2384 and w2654;
w2656 <= not w2647 and w2655;
w2657 <= not a(86) and not w2646;
w2658 <= a(87) and not w2657;
w2659 <= w2400 and not w2646;
w2660 <= not w2658 and not w2659;
w2661 <= not w2656 and w2660;
w2662 <= not w2651 and not w2661;
w2663 <= not w2162 and not w2662;
w2664 <= w2162 and not w2651;
w2665 <= not w2661 and w2664;
w2666 <= not w2398 and not w2643;
w2667 <= not w2638 and w2666;
w2668 <= not w2634 and w2667;
w2669 <= not w2632 and w2668;
w2670 <= not w2659 and not w2669;
w2671 <= a(88) and not w2670;
w2672 <= not a(88) and not w2669;
w2673 <= not w2659 and w2672;
w2674 <= not w2671 and not w2673;
w2675 <= not w2665 and not w2674;
w2676 <= not w2663 and not w2675;
w2677 <= not w1938 and not w2676;
w2678 <= not w2403 and not w2408;
w2679 <= not w2412 and w2678;
w2680 <= not w2646 and w2679;
w2681 <= not w2646 and w2678;
w2682 <= w2412 and not w2681;
w2683 <= not w2680 and not w2682;
w2684 <= w1938 and not w2663;
w2685 <= not w2675 and w2684;
w2686 <= not w2683 and not w2685;
w2687 <= not w2677 and not w2686;
w2688 <= not w1725 and not w2687;
w2689 <= not w2417 and w2426;
w2690 <= not w2415 and w2689;
w2691 <= not w2646 and w2690;
w2692 <= not w2415 and not w2417;
w2693 <= not w2646 and w2692;
w2694 <= not w2426 and not w2693;
w2695 <= not w2691 and not w2694;
w2696 <= w1725 and not w2677;
w2697 <= not w2686 and w2696;
w2698 <= not w2695 and not w2697;
w2699 <= not w2688 and not w2698;
w2700 <= not w1525 and not w2699;
w2701 <= not w2429 and w2435;
w2702 <= not w2437 and w2701;
w2703 <= not w2646 and w2702;
w2704 <= not w2429 and not w2437;
w2705 <= not w2646 and w2704;
w2706 <= not w2435 and not w2705;
w2707 <= not w2703 and not w2706;
w2708 <= w1525 and not w2688;
w2709 <= not w2698 and w2708;
w2710 <= not w2707 and not w2709;
w2711 <= not w2700 and not w2710;
w2712 <= not w1337 and not w2711;
w2713 <= w2447 and not w2449;
w2714 <= not w2440 and w2713;
w2715 <= not w2646 and w2714;
w2716 <= not w2440 and not w2449;
w2717 <= not w2646 and w2716;
w2718 <= not w2447 and not w2717;
w2719 <= not w2715 and not w2718;
w2720 <= w1337 and not w2700;
w2721 <= not w2710 and w2720;
w2722 <= not w2719 and not w2721;
w2723 <= not w2712 and not w2722;
w2724 <= not w1161 and not w2723;
w2725 <= not w2452 and w2459;
w2726 <= not w2461 and w2725;
w2727 <= not w2646 and w2726;
w2728 <= not w2452 and not w2461;
w2729 <= not w2646 and w2728;
w2730 <= not w2459 and not w2729;
w2731 <= not w2727 and not w2730;
w2732 <= w1161 and not w2712;
w2733 <= not w2722 and w2732;
w2734 <= not w2731 and not w2733;
w2735 <= not w2724 and not w2734;
w2736 <= not w997 and not w2735;
w2737 <= w2471 and not w2473;
w2738 <= not w2464 and w2737;
w2739 <= not w2646 and w2738;
w2740 <= not w2464 and not w2473;
w2741 <= not w2646 and w2740;
w2742 <= not w2471 and not w2741;
w2743 <= not w2739 and not w2742;
w2744 <= w997 and not w2724;
w2745 <= not w2734 and w2744;
w2746 <= not w2743 and not w2745;
w2747 <= not w2736 and not w2746;
w2748 <= not w845 and not w2747;
w2749 <= not w2476 and w2483;
w2750 <= not w2485 and w2749;
w2751 <= not w2646 and w2750;
w2752 <= not w2476 and not w2485;
w2753 <= not w2646 and w2752;
w2754 <= not w2483 and not w2753;
w2755 <= not w2751 and not w2754;
w2756 <= w845 and not w2736;
w2757 <= not w2746 and w2756;
w2758 <= not w2755 and not w2757;
w2759 <= not w2748 and not w2758;
w2760 <= not w705 and not w2759;
w2761 <= w2495 and not w2497;
w2762 <= not w2488 and w2761;
w2763 <= not w2646 and w2762;
w2764 <= not w2488 and not w2497;
w2765 <= not w2646 and w2764;
w2766 <= not w2495 and not w2765;
w2767 <= not w2763 and not w2766;
w2768 <= w705 and not w2748;
w2769 <= not w2758 and w2768;
w2770 <= not w2767 and not w2769;
w2771 <= not w2760 and not w2770;
w2772 <= not w577 and not w2771;
w2773 <= w577 and not w2760;
w2774 <= not w2770 and w2773;
w2775 <= not w2500 and w2509;
w2776 <= not w2502 and w2775;
w2777 <= not w2646 and w2776;
w2778 <= not w2500 and not w2502;
w2779 <= not w2646 and w2778;
w2780 <= not w2509 and not w2779;
w2781 <= not w2777 and not w2780;
w2782 <= not w2774 and not w2781;
w2783 <= not w2772 and not w2782;
w2784 <= not w460 and not w2783;
w2785 <= w2519 and not w2521;
w2786 <= not w2512 and w2785;
w2787 <= not w2646 and w2786;
w2788 <= not w2512 and not w2521;
w2789 <= not w2646 and w2788;
w2790 <= not w2519 and not w2789;
w2791 <= not w2787 and not w2790;
w2792 <= w460 and not w2772;
w2793 <= not w2782 and w2792;
w2794 <= not w2791 and not w2793;
w2795 <= not w2784 and not w2794;
w2796 <= not w356 and not w2795;
w2797 <= not w2524 and w2531;
w2798 <= not w2533 and w2797;
w2799 <= not w2646 and w2798;
w2800 <= not w2524 and not w2533;
w2801 <= not w2646 and w2800;
w2802 <= not w2531 and not w2801;
w2803 <= not w2799 and not w2802;
w2804 <= w356 and not w2784;
w2805 <= not w2794 and w2804;
w2806 <= not w2803 and not w2805;
w2807 <= not w2796 and not w2806;
w2808 <= not w264 and not w2807;
w2809 <= w2543 and not w2545;
w2810 <= not w2536 and w2809;
w2811 <= not w2646 and w2810;
w2812 <= not w2536 and not w2545;
w2813 <= not w2646 and w2812;
w2814 <= not w2543 and not w2813;
w2815 <= not w2811 and not w2814;
w2816 <= w264 and not w2796;
w2817 <= not w2806 and w2816;
w2818 <= not w2815 and not w2817;
w2819 <= not w2808 and not w2818;
w2820 <= not w184 and not w2819;
w2821 <= not w2548 and w2555;
w2822 <= not w2557 and w2821;
w2823 <= not w2646 and w2822;
w2824 <= not w2548 and not w2557;
w2825 <= not w2646 and w2824;
w2826 <= not w2555 and not w2825;
w2827 <= not w2823 and not w2826;
w2828 <= w184 and not w2808;
w2829 <= not w2818 and w2828;
w2830 <= not w2827 and not w2829;
w2831 <= not w2820 and not w2830;
w2832 <= not w115 and not w2831;
w2833 <= w2567 and not w2569;
w2834 <= not w2560 and w2833;
w2835 <= not w2646 and w2834;
w2836 <= not w2560 and not w2569;
w2837 <= not w2646 and w2836;
w2838 <= not w2567 and not w2837;
w2839 <= not w2835 and not w2838;
w2840 <= w115 and not w2820;
w2841 <= not w2830 and w2840;
w2842 <= not w2839 and not w2841;
w2843 <= not w2832 and not w2842;
w2844 <= not w60 and not w2843;
w2845 <= not w2572 and w2579;
w2846 <= not w2581 and w2845;
w2847 <= not w2646 and w2846;
w2848 <= not w2572 and not w2581;
w2849 <= not w2646 and w2848;
w2850 <= not w2579 and not w2849;
w2851 <= not w2847 and not w2850;
w2852 <= w60 and not w2832;
w2853 <= not w2842 and w2852;
w2854 <= not w2851 and not w2853;
w2855 <= not w2844 and not w2854;
w2856 <= not w22 and not w2855;
w2857 <= w2591 and not w2593;
w2858 <= not w2584 and w2857;
w2859 <= not w2646 and w2858;
w2860 <= not w2584 and not w2593;
w2861 <= not w2646 and w2860;
w2862 <= not w2591 and not w2861;
w2863 <= not w2859 and not w2862;
w2864 <= w22 and not w2844;
w2865 <= not w2854 and w2864;
w2866 <= not w2863 and not w2865;
w2867 <= not w2856 and not w2866;
w2868 <= not w5 and not w2867;
w2869 <= not w2596 and w2603;
w2870 <= not w2605 and w2869;
w2871 <= not w2646 and w2870;
w2872 <= not w2596 and not w2605;
w2873 <= not w2646 and w2872;
w2874 <= not w2603 and not w2873;
w2875 <= not w2871 and not w2874;
w2876 <= w5 and not w2856;
w2877 <= not w2866 and w2876;
w2878 <= not w2875 and not w2877;
w2879 <= not w2868 and not w2878;
w2880 <= w2615 and not w2617;
w2881 <= not w2608 and w2880;
w2882 <= not w2646 and w2881;
w2883 <= not w2608 and not w2617;
w2884 <= not w2646 and w2883;
w2885 <= not w2615 and not w2884;
w2886 <= not w2882 and not w2885;
w2887 <= not w2619 and not w2626;
w2888 <= not w2646 and w2887;
w2889 <= not w2634 and not w2888;
w2890 <= not w2886 and w2889;
w2891 <= not w2879 and w2890;
w2892 <= w0 and not w2891;
w2893 <= not w2868 and w2886;
w2894 <= not w2878 and w2893;
w2895 <= not w2626 and not w2646;
w2896 <= w2619 and not w2895;
w2897 <= not w0 and not w2887;
w2898 <= not w2896 and w2897;
w2899 <= not w2622 and not w2643;
w2900 <= not w2625 and w2899;
w2901 <= not w2638 and w2900;
w2902 <= not w2634 and w2901;
w2903 <= not w2632 and w2902;
w2904 <= not w2898 and not w2903;
w2905 <= not w2894 and w2904;
w2906 <= not w2892 and w2905;
w2907 <= a(84) and not w2906;
w2908 <= not a(82) and not a(83);
w2909 <= not a(84) and w2908;
w2910 <= not w2907 and not w2909;
w2911 <= not w2646 and not w2910;
w2912 <= not w2643 and not w2909;
w2913 <= not w2638 and w2912;
w2914 <= not w2634 and w2913;
w2915 <= not w2632 and w2914;
w2916 <= not w2907 and w2915;
w2917 <= not a(84) and not w2906;
w2918 <= a(85) and not w2917;
w2919 <= w2648 and not w2906;
w2920 <= not w2918 and not w2919;
w2921 <= not w2916 and w2920;
w2922 <= not w2911 and not w2921;
w2923 <= not w2398 and not w2922;
w2924 <= w2398 and not w2911;
w2925 <= not w2921 and w2924;
w2926 <= not w2646 and not w2903;
w2927 <= not w2898 and w2926;
w2928 <= not w2894 and w2927;
w2929 <= not w2892 and w2928;
w2930 <= not w2919 and not w2929;
w2931 <= a(86) and not w2930;
w2932 <= not a(86) and not w2929;
w2933 <= not w2919 and w2932;
w2934 <= not w2931 and not w2933;
w2935 <= not w2925 and not w2934;
w2936 <= not w2923 and not w2935;
w2937 <= not w2162 and not w2936;
w2938 <= not w2651 and not w2656;
w2939 <= not w2660 and w2938;
w2940 <= not w2906 and w2939;
w2941 <= not w2906 and w2938;
w2942 <= w2660 and not w2941;
w2943 <= not w2940 and not w2942;
w2944 <= w2162 and not w2923;
w2945 <= not w2935 and w2944;
w2946 <= not w2943 and not w2945;
w2947 <= not w2937 and not w2946;
w2948 <= not w1938 and not w2947;
w2949 <= not w2665 and w2674;
w2950 <= not w2663 and w2949;
w2951 <= not w2906 and w2950;
w2952 <= not w2663 and not w2665;
w2953 <= not w2906 and w2952;
w2954 <= not w2674 and not w2953;
w2955 <= not w2951 and not w2954;
w2956 <= w1938 and not w2937;
w2957 <= not w2946 and w2956;
w2958 <= not w2955 and not w2957;
w2959 <= not w2948 and not w2958;
w2960 <= not w1725 and not w2959;
w2961 <= not w2677 and w2683;
w2962 <= not w2685 and w2961;
w2963 <= not w2906 and w2962;
w2964 <= not w2677 and not w2685;
w2965 <= not w2906 and w2964;
w2966 <= not w2683 and not w2965;
w2967 <= not w2963 and not w2966;
w2968 <= w1725 and not w2948;
w2969 <= not w2958 and w2968;
w2970 <= not w2967 and not w2969;
w2971 <= not w2960 and not w2970;
w2972 <= not w1525 and not w2971;
w2973 <= w2695 and not w2697;
w2974 <= not w2688 and w2973;
w2975 <= not w2906 and w2974;
w2976 <= not w2688 and not w2697;
w2977 <= not w2906 and w2976;
w2978 <= not w2695 and not w2977;
w2979 <= not w2975 and not w2978;
w2980 <= w1525 and not w2960;
w2981 <= not w2970 and w2980;
w2982 <= not w2979 and not w2981;
w2983 <= not w2972 and not w2982;
w2984 <= not w1337 and not w2983;
w2985 <= not w2700 and w2707;
w2986 <= not w2709 and w2985;
w2987 <= not w2906 and w2986;
w2988 <= not w2700 and not w2709;
w2989 <= not w2906 and w2988;
w2990 <= not w2707 and not w2989;
w2991 <= not w2987 and not w2990;
w2992 <= w1337 and not w2972;
w2993 <= not w2982 and w2992;
w2994 <= not w2991 and not w2993;
w2995 <= not w2984 and not w2994;
w2996 <= not w1161 and not w2995;
w2997 <= w2719 and not w2721;
w2998 <= not w2712 and w2997;
w2999 <= not w2906 and w2998;
w3000 <= not w2712 and not w2721;
w3001 <= not w2906 and w3000;
w3002 <= not w2719 and not w3001;
w3003 <= not w2999 and not w3002;
w3004 <= w1161 and not w2984;
w3005 <= not w2994 and w3004;
w3006 <= not w3003 and not w3005;
w3007 <= not w2996 and not w3006;
w3008 <= not w997 and not w3007;
w3009 <= not w2724 and w2731;
w3010 <= not w2733 and w3009;
w3011 <= not w2906 and w3010;
w3012 <= not w2724 and not w2733;
w3013 <= not w2906 and w3012;
w3014 <= not w2731 and not w3013;
w3015 <= not w3011 and not w3014;
w3016 <= w997 and not w2996;
w3017 <= not w3006 and w3016;
w3018 <= not w3015 and not w3017;
w3019 <= not w3008 and not w3018;
w3020 <= not w845 and not w3019;
w3021 <= w2743 and not w2745;
w3022 <= not w2736 and w3021;
w3023 <= not w2906 and w3022;
w3024 <= not w2736 and not w2745;
w3025 <= not w2906 and w3024;
w3026 <= not w2743 and not w3025;
w3027 <= not w3023 and not w3026;
w3028 <= w845 and not w3008;
w3029 <= not w3018 and w3028;
w3030 <= not w3027 and not w3029;
w3031 <= not w3020 and not w3030;
w3032 <= not w705 and not w3031;
w3033 <= not w2748 and w2755;
w3034 <= not w2757 and w3033;
w3035 <= not w2906 and w3034;
w3036 <= not w2748 and not w2757;
w3037 <= not w2906 and w3036;
w3038 <= not w2755 and not w3037;
w3039 <= not w3035 and not w3038;
w3040 <= w705 and not w3020;
w3041 <= not w3030 and w3040;
w3042 <= not w3039 and not w3041;
w3043 <= not w3032 and not w3042;
w3044 <= not w577 and not w3043;
w3045 <= w2767 and not w2769;
w3046 <= not w2760 and w3045;
w3047 <= not w2906 and w3046;
w3048 <= not w2760 and not w2769;
w3049 <= not w2906 and w3048;
w3050 <= not w2767 and not w3049;
w3051 <= not w3047 and not w3050;
w3052 <= w577 and not w3032;
w3053 <= not w3042 and w3052;
w3054 <= not w3051 and not w3053;
w3055 <= not w3044 and not w3054;
w3056 <= not w460 and not w3055;
w3057 <= w460 and not w3044;
w3058 <= not w3054 and w3057;
w3059 <= not w2772 and w2781;
w3060 <= not w2774 and w3059;
w3061 <= not w2906 and w3060;
w3062 <= not w2772 and not w2774;
w3063 <= not w2906 and w3062;
w3064 <= not w2781 and not w3063;
w3065 <= not w3061 and not w3064;
w3066 <= not w3058 and not w3065;
w3067 <= not w3056 and not w3066;
w3068 <= not w356 and not w3067;
w3069 <= w2791 and not w2793;
w3070 <= not w2784 and w3069;
w3071 <= not w2906 and w3070;
w3072 <= not w2784 and not w2793;
w3073 <= not w2906 and w3072;
w3074 <= not w2791 and not w3073;
w3075 <= not w3071 and not w3074;
w3076 <= w356 and not w3056;
w3077 <= not w3066 and w3076;
w3078 <= not w3075 and not w3077;
w3079 <= not w3068 and not w3078;
w3080 <= not w264 and not w3079;
w3081 <= not w2796 and w2803;
w3082 <= not w2805 and w3081;
w3083 <= not w2906 and w3082;
w3084 <= not w2796 and not w2805;
w3085 <= not w2906 and w3084;
w3086 <= not w2803 and not w3085;
w3087 <= not w3083 and not w3086;
w3088 <= w264 and not w3068;
w3089 <= not w3078 and w3088;
w3090 <= not w3087 and not w3089;
w3091 <= not w3080 and not w3090;
w3092 <= not w184 and not w3091;
w3093 <= w2815 and not w2817;
w3094 <= not w2808 and w3093;
w3095 <= not w2906 and w3094;
w3096 <= not w2808 and not w2817;
w3097 <= not w2906 and w3096;
w3098 <= not w2815 and not w3097;
w3099 <= not w3095 and not w3098;
w3100 <= w184 and not w3080;
w3101 <= not w3090 and w3100;
w3102 <= not w3099 and not w3101;
w3103 <= not w3092 and not w3102;
w3104 <= not w115 and not w3103;
w3105 <= not w2820 and w2827;
w3106 <= not w2829 and w3105;
w3107 <= not w2906 and w3106;
w3108 <= not w2820 and not w2829;
w3109 <= not w2906 and w3108;
w3110 <= not w2827 and not w3109;
w3111 <= not w3107 and not w3110;
w3112 <= w115 and not w3092;
w3113 <= not w3102 and w3112;
w3114 <= not w3111 and not w3113;
w3115 <= not w3104 and not w3114;
w3116 <= not w60 and not w3115;
w3117 <= w2839 and not w2841;
w3118 <= not w2832 and w3117;
w3119 <= not w2906 and w3118;
w3120 <= not w2832 and not w2841;
w3121 <= not w2906 and w3120;
w3122 <= not w2839 and not w3121;
w3123 <= not w3119 and not w3122;
w3124 <= w60 and not w3104;
w3125 <= not w3114 and w3124;
w3126 <= not w3123 and not w3125;
w3127 <= not w3116 and not w3126;
w3128 <= not w22 and not w3127;
w3129 <= not w2844 and w2851;
w3130 <= not w2853 and w3129;
w3131 <= not w2906 and w3130;
w3132 <= not w2844 and not w2853;
w3133 <= not w2906 and w3132;
w3134 <= not w2851 and not w3133;
w3135 <= not w3131 and not w3134;
w3136 <= w22 and not w3116;
w3137 <= not w3126 and w3136;
w3138 <= not w3135 and not w3137;
w3139 <= not w3128 and not w3138;
w3140 <= not w5 and not w3139;
w3141 <= w2863 and not w2865;
w3142 <= not w2856 and w3141;
w3143 <= not w2906 and w3142;
w3144 <= not w2856 and not w2865;
w3145 <= not w2906 and w3144;
w3146 <= not w2863 and not w3145;
w3147 <= not w3143 and not w3146;
w3148 <= w5 and not w3128;
w3149 <= not w3138 and w3148;
w3150 <= not w3147 and not w3149;
w3151 <= not w3140 and not w3150;
w3152 <= not w2868 and w2875;
w3153 <= not w2877 and w3152;
w3154 <= not w2906 and w3153;
w3155 <= not w2868 and not w2877;
w3156 <= not w2906 and w3155;
w3157 <= not w2875 and not w3156;
w3158 <= not w3154 and not w3157;
w3159 <= not w2879 and not w2886;
w3160 <= not w2906 and w3159;
w3161 <= not w2894 and not w3160;
w3162 <= not w3158 and w3161;
w3163 <= not w3151 and w3162;
w3164 <= w0 and not w3163;
w3165 <= not w3140 and w3158;
w3166 <= not w3150 and w3165;
w3167 <= not w2886 and not w2906;
w3168 <= w2879 and not w3167;
w3169 <= not w0 and not w3159;
w3170 <= not w3168 and w3169;
w3171 <= not w2882 and not w2903;
w3172 <= not w2885 and w3171;
w3173 <= not w2898 and w3172;
w3174 <= not w2894 and w3173;
w3175 <= not w2892 and w3174;
w3176 <= not w3170 and not w3175;
w3177 <= not w3166 and w3176;
w3178 <= not w3164 and w3177;
w3179 <= a(82) and not w3178;
w3180 <= not a(80) and not a(81);
w3181 <= not a(82) and w3180;
w3182 <= not w3179 and not w3181;
w3183 <= not w2906 and not w3182;
w3184 <= not w2903 and not w3181;
w3185 <= not w2898 and w3184;
w3186 <= not w2894 and w3185;
w3187 <= not w2892 and w3186;
w3188 <= not w3179 and w3187;
w3189 <= not a(82) and not w3178;
w3190 <= a(83) and not w3189;
w3191 <= w2908 and not w3178;
w3192 <= not w3190 and not w3191;
w3193 <= not w3188 and w3192;
w3194 <= not w3183 and not w3193;
w3195 <= not w2646 and not w3194;
w3196 <= w2646 and not w3183;
w3197 <= not w3193 and w3196;
w3198 <= not w2906 and not w3175;
w3199 <= not w3170 and w3198;
w3200 <= not w3166 and w3199;
w3201 <= not w3164 and w3200;
w3202 <= not w3191 and not w3201;
w3203 <= a(84) and not w3202;
w3204 <= not a(84) and not w3201;
w3205 <= not w3191 and w3204;
w3206 <= not w3203 and not w3205;
w3207 <= not w3197 and not w3206;
w3208 <= not w3195 and not w3207;
w3209 <= not w2398 and not w3208;
w3210 <= not w2911 and not w2916;
w3211 <= not w2920 and w3210;
w3212 <= not w3178 and w3211;
w3213 <= not w3178 and w3210;
w3214 <= w2920 and not w3213;
w3215 <= not w3212 and not w3214;
w3216 <= w2398 and not w3195;
w3217 <= not w3207 and w3216;
w3218 <= not w3215 and not w3217;
w3219 <= not w3209 and not w3218;
w3220 <= not w2162 and not w3219;
w3221 <= not w2925 and w2934;
w3222 <= not w2923 and w3221;
w3223 <= not w3178 and w3222;
w3224 <= not w2923 and not w2925;
w3225 <= not w3178 and w3224;
w3226 <= not w2934 and not w3225;
w3227 <= not w3223 and not w3226;
w3228 <= w2162 and not w3209;
w3229 <= not w3218 and w3228;
w3230 <= not w3227 and not w3229;
w3231 <= not w3220 and not w3230;
w3232 <= not w1938 and not w3231;
w3233 <= not w2937 and w2943;
w3234 <= not w2945 and w3233;
w3235 <= not w3178 and w3234;
w3236 <= not w2937 and not w2945;
w3237 <= not w3178 and w3236;
w3238 <= not w2943 and not w3237;
w3239 <= not w3235 and not w3238;
w3240 <= w1938 and not w3220;
w3241 <= not w3230 and w3240;
w3242 <= not w3239 and not w3241;
w3243 <= not w3232 and not w3242;
w3244 <= not w1725 and not w3243;
w3245 <= w2955 and not w2957;
w3246 <= not w2948 and w3245;
w3247 <= not w3178 and w3246;
w3248 <= not w2948 and not w2957;
w3249 <= not w3178 and w3248;
w3250 <= not w2955 and not w3249;
w3251 <= not w3247 and not w3250;
w3252 <= w1725 and not w3232;
w3253 <= not w3242 and w3252;
w3254 <= not w3251 and not w3253;
w3255 <= not w3244 and not w3254;
w3256 <= not w1525 and not w3255;
w3257 <= not w2960 and w2967;
w3258 <= not w2969 and w3257;
w3259 <= not w3178 and w3258;
w3260 <= not w2960 and not w2969;
w3261 <= not w3178 and w3260;
w3262 <= not w2967 and not w3261;
w3263 <= not w3259 and not w3262;
w3264 <= w1525 and not w3244;
w3265 <= not w3254 and w3264;
w3266 <= not w3263 and not w3265;
w3267 <= not w3256 and not w3266;
w3268 <= not w1337 and not w3267;
w3269 <= w2979 and not w2981;
w3270 <= not w2972 and w3269;
w3271 <= not w3178 and w3270;
w3272 <= not w2972 and not w2981;
w3273 <= not w3178 and w3272;
w3274 <= not w2979 and not w3273;
w3275 <= not w3271 and not w3274;
w3276 <= w1337 and not w3256;
w3277 <= not w3266 and w3276;
w3278 <= not w3275 and not w3277;
w3279 <= not w3268 and not w3278;
w3280 <= not w1161 and not w3279;
w3281 <= not w2984 and w2991;
w3282 <= not w2993 and w3281;
w3283 <= not w3178 and w3282;
w3284 <= not w2984 and not w2993;
w3285 <= not w3178 and w3284;
w3286 <= not w2991 and not w3285;
w3287 <= not w3283 and not w3286;
w3288 <= w1161 and not w3268;
w3289 <= not w3278 and w3288;
w3290 <= not w3287 and not w3289;
w3291 <= not w3280 and not w3290;
w3292 <= not w997 and not w3291;
w3293 <= w3003 and not w3005;
w3294 <= not w2996 and w3293;
w3295 <= not w3178 and w3294;
w3296 <= not w2996 and not w3005;
w3297 <= not w3178 and w3296;
w3298 <= not w3003 and not w3297;
w3299 <= not w3295 and not w3298;
w3300 <= w997 and not w3280;
w3301 <= not w3290 and w3300;
w3302 <= not w3299 and not w3301;
w3303 <= not w3292 and not w3302;
w3304 <= not w845 and not w3303;
w3305 <= not w3008 and w3015;
w3306 <= not w3017 and w3305;
w3307 <= not w3178 and w3306;
w3308 <= not w3008 and not w3017;
w3309 <= not w3178 and w3308;
w3310 <= not w3015 and not w3309;
w3311 <= not w3307 and not w3310;
w3312 <= w845 and not w3292;
w3313 <= not w3302 and w3312;
w3314 <= not w3311 and not w3313;
w3315 <= not w3304 and not w3314;
w3316 <= not w705 and not w3315;
w3317 <= w3027 and not w3029;
w3318 <= not w3020 and w3317;
w3319 <= not w3178 and w3318;
w3320 <= not w3020 and not w3029;
w3321 <= not w3178 and w3320;
w3322 <= not w3027 and not w3321;
w3323 <= not w3319 and not w3322;
w3324 <= w705 and not w3304;
w3325 <= not w3314 and w3324;
w3326 <= not w3323 and not w3325;
w3327 <= not w3316 and not w3326;
w3328 <= not w577 and not w3327;
w3329 <= not w3032 and w3039;
w3330 <= not w3041 and w3329;
w3331 <= not w3178 and w3330;
w3332 <= not w3032 and not w3041;
w3333 <= not w3178 and w3332;
w3334 <= not w3039 and not w3333;
w3335 <= not w3331 and not w3334;
w3336 <= w577 and not w3316;
w3337 <= not w3326 and w3336;
w3338 <= not w3335 and not w3337;
w3339 <= not w3328 and not w3338;
w3340 <= not w460 and not w3339;
w3341 <= w3051 and not w3053;
w3342 <= not w3044 and w3341;
w3343 <= not w3178 and w3342;
w3344 <= not w3044 and not w3053;
w3345 <= not w3178 and w3344;
w3346 <= not w3051 and not w3345;
w3347 <= not w3343 and not w3346;
w3348 <= w460 and not w3328;
w3349 <= not w3338 and w3348;
w3350 <= not w3347 and not w3349;
w3351 <= not w3340 and not w3350;
w3352 <= not w356 and not w3351;
w3353 <= w356 and not w3340;
w3354 <= not w3350 and w3353;
w3355 <= not w3056 and w3065;
w3356 <= not w3058 and w3355;
w3357 <= not w3178 and w3356;
w3358 <= not w3056 and not w3058;
w3359 <= not w3178 and w3358;
w3360 <= not w3065 and not w3359;
w3361 <= not w3357 and not w3360;
w3362 <= not w3354 and not w3361;
w3363 <= not w3352 and not w3362;
w3364 <= not w264 and not w3363;
w3365 <= w3075 and not w3077;
w3366 <= not w3068 and w3365;
w3367 <= not w3178 and w3366;
w3368 <= not w3068 and not w3077;
w3369 <= not w3178 and w3368;
w3370 <= not w3075 and not w3369;
w3371 <= not w3367 and not w3370;
w3372 <= w264 and not w3352;
w3373 <= not w3362 and w3372;
w3374 <= not w3371 and not w3373;
w3375 <= not w3364 and not w3374;
w3376 <= not w184 and not w3375;
w3377 <= not w3080 and w3087;
w3378 <= not w3089 and w3377;
w3379 <= not w3178 and w3378;
w3380 <= not w3080 and not w3089;
w3381 <= not w3178 and w3380;
w3382 <= not w3087 and not w3381;
w3383 <= not w3379 and not w3382;
w3384 <= w184 and not w3364;
w3385 <= not w3374 and w3384;
w3386 <= not w3383 and not w3385;
w3387 <= not w3376 and not w3386;
w3388 <= not w115 and not w3387;
w3389 <= w3099 and not w3101;
w3390 <= not w3092 and w3389;
w3391 <= not w3178 and w3390;
w3392 <= not w3092 and not w3101;
w3393 <= not w3178 and w3392;
w3394 <= not w3099 and not w3393;
w3395 <= not w3391 and not w3394;
w3396 <= w115 and not w3376;
w3397 <= not w3386 and w3396;
w3398 <= not w3395 and not w3397;
w3399 <= not w3388 and not w3398;
w3400 <= not w60 and not w3399;
w3401 <= not w3104 and w3111;
w3402 <= not w3113 and w3401;
w3403 <= not w3178 and w3402;
w3404 <= not w3104 and not w3113;
w3405 <= not w3178 and w3404;
w3406 <= not w3111 and not w3405;
w3407 <= not w3403 and not w3406;
w3408 <= w60 and not w3388;
w3409 <= not w3398 and w3408;
w3410 <= not w3407 and not w3409;
w3411 <= not w3400 and not w3410;
w3412 <= not w22 and not w3411;
w3413 <= w3123 and not w3125;
w3414 <= not w3116 and w3413;
w3415 <= not w3178 and w3414;
w3416 <= not w3116 and not w3125;
w3417 <= not w3178 and w3416;
w3418 <= not w3123 and not w3417;
w3419 <= not w3415 and not w3418;
w3420 <= w22 and not w3400;
w3421 <= not w3410 and w3420;
w3422 <= not w3419 and not w3421;
w3423 <= not w3412 and not w3422;
w3424 <= not w5 and not w3423;
w3425 <= not w3128 and w3135;
w3426 <= not w3137 and w3425;
w3427 <= not w3178 and w3426;
w3428 <= not w3128 and not w3137;
w3429 <= not w3178 and w3428;
w3430 <= not w3135 and not w3429;
w3431 <= not w3427 and not w3430;
w3432 <= w5 and not w3412;
w3433 <= not w3422 and w3432;
w3434 <= not w3431 and not w3433;
w3435 <= not w3424 and not w3434;
w3436 <= w3147 and not w3149;
w3437 <= not w3140 and w3436;
w3438 <= not w3178 and w3437;
w3439 <= not w3140 and not w3149;
w3440 <= not w3178 and w3439;
w3441 <= not w3147 and not w3440;
w3442 <= not w3438 and not w3441;
w3443 <= not w3151 and not w3158;
w3444 <= not w3178 and w3443;
w3445 <= not w3166 and not w3444;
w3446 <= not w3442 and w3445;
w3447 <= not w3435 and w3446;
w3448 <= w0 and not w3447;
w3449 <= not w3424 and w3442;
w3450 <= not w3434 and w3449;
w3451 <= not w3158 and not w3178;
w3452 <= w3151 and not w3451;
w3453 <= not w0 and not w3443;
w3454 <= not w3452 and w3453;
w3455 <= not w3154 and not w3175;
w3456 <= not w3157 and w3455;
w3457 <= not w3170 and w3456;
w3458 <= not w3166 and w3457;
w3459 <= not w3164 and w3458;
w3460 <= not w3454 and not w3459;
w3461 <= not w3450 and w3460;
w3462 <= not w3448 and w3461;
w3463 <= a(80) and not w3462;
w3464 <= not a(78) and not a(79);
w3465 <= not a(80) and w3464;
w3466 <= not w3463 and not w3465;
w3467 <= not w3178 and not w3466;
w3468 <= not w3175 and not w3465;
w3469 <= not w3170 and w3468;
w3470 <= not w3166 and w3469;
w3471 <= not w3164 and w3470;
w3472 <= not w3463 and w3471;
w3473 <= not a(80) and not w3462;
w3474 <= a(81) and not w3473;
w3475 <= w3180 and not w3462;
w3476 <= not w3474 and not w3475;
w3477 <= not w3472 and w3476;
w3478 <= not w3467 and not w3477;
w3479 <= not w2906 and not w3478;
w3480 <= w2906 and not w3467;
w3481 <= not w3477 and w3480;
w3482 <= not w3178 and not w3459;
w3483 <= not w3454 and w3482;
w3484 <= not w3450 and w3483;
w3485 <= not w3448 and w3484;
w3486 <= not w3475 and not w3485;
w3487 <= a(82) and not w3486;
w3488 <= not a(82) and not w3485;
w3489 <= not w3475 and w3488;
w3490 <= not w3487 and not w3489;
w3491 <= not w3481 and not w3490;
w3492 <= not w3479 and not w3491;
w3493 <= not w2646 and not w3492;
w3494 <= not w3183 and not w3188;
w3495 <= not w3192 and w3494;
w3496 <= not w3462 and w3495;
w3497 <= not w3462 and w3494;
w3498 <= w3192 and not w3497;
w3499 <= not w3496 and not w3498;
w3500 <= w2646 and not w3479;
w3501 <= not w3491 and w3500;
w3502 <= not w3499 and not w3501;
w3503 <= not w3493 and not w3502;
w3504 <= not w2398 and not w3503;
w3505 <= not w3197 and w3206;
w3506 <= not w3195 and w3505;
w3507 <= not w3462 and w3506;
w3508 <= not w3195 and not w3197;
w3509 <= not w3462 and w3508;
w3510 <= not w3206 and not w3509;
w3511 <= not w3507 and not w3510;
w3512 <= w2398 and not w3493;
w3513 <= not w3502 and w3512;
w3514 <= not w3511 and not w3513;
w3515 <= not w3504 and not w3514;
w3516 <= not w2162 and not w3515;
w3517 <= not w3209 and w3215;
w3518 <= not w3217 and w3517;
w3519 <= not w3462 and w3518;
w3520 <= not w3209 and not w3217;
w3521 <= not w3462 and w3520;
w3522 <= not w3215 and not w3521;
w3523 <= not w3519 and not w3522;
w3524 <= w2162 and not w3504;
w3525 <= not w3514 and w3524;
w3526 <= not w3523 and not w3525;
w3527 <= not w3516 and not w3526;
w3528 <= not w1938 and not w3527;
w3529 <= w3227 and not w3229;
w3530 <= not w3220 and w3529;
w3531 <= not w3462 and w3530;
w3532 <= not w3220 and not w3229;
w3533 <= not w3462 and w3532;
w3534 <= not w3227 and not w3533;
w3535 <= not w3531 and not w3534;
w3536 <= w1938 and not w3516;
w3537 <= not w3526 and w3536;
w3538 <= not w3535 and not w3537;
w3539 <= not w3528 and not w3538;
w3540 <= not w1725 and not w3539;
w3541 <= not w3232 and w3239;
w3542 <= not w3241 and w3541;
w3543 <= not w3462 and w3542;
w3544 <= not w3232 and not w3241;
w3545 <= not w3462 and w3544;
w3546 <= not w3239 and not w3545;
w3547 <= not w3543 and not w3546;
w3548 <= w1725 and not w3528;
w3549 <= not w3538 and w3548;
w3550 <= not w3547 and not w3549;
w3551 <= not w3540 and not w3550;
w3552 <= not w1525 and not w3551;
w3553 <= w3251 and not w3253;
w3554 <= not w3244 and w3553;
w3555 <= not w3462 and w3554;
w3556 <= not w3244 and not w3253;
w3557 <= not w3462 and w3556;
w3558 <= not w3251 and not w3557;
w3559 <= not w3555 and not w3558;
w3560 <= w1525 and not w3540;
w3561 <= not w3550 and w3560;
w3562 <= not w3559 and not w3561;
w3563 <= not w3552 and not w3562;
w3564 <= not w1337 and not w3563;
w3565 <= not w3256 and w3263;
w3566 <= not w3265 and w3565;
w3567 <= not w3462 and w3566;
w3568 <= not w3256 and not w3265;
w3569 <= not w3462 and w3568;
w3570 <= not w3263 and not w3569;
w3571 <= not w3567 and not w3570;
w3572 <= w1337 and not w3552;
w3573 <= not w3562 and w3572;
w3574 <= not w3571 and not w3573;
w3575 <= not w3564 and not w3574;
w3576 <= not w1161 and not w3575;
w3577 <= w3275 and not w3277;
w3578 <= not w3268 and w3577;
w3579 <= not w3462 and w3578;
w3580 <= not w3268 and not w3277;
w3581 <= not w3462 and w3580;
w3582 <= not w3275 and not w3581;
w3583 <= not w3579 and not w3582;
w3584 <= w1161 and not w3564;
w3585 <= not w3574 and w3584;
w3586 <= not w3583 and not w3585;
w3587 <= not w3576 and not w3586;
w3588 <= not w997 and not w3587;
w3589 <= not w3280 and w3287;
w3590 <= not w3289 and w3589;
w3591 <= not w3462 and w3590;
w3592 <= not w3280 and not w3289;
w3593 <= not w3462 and w3592;
w3594 <= not w3287 and not w3593;
w3595 <= not w3591 and not w3594;
w3596 <= w997 and not w3576;
w3597 <= not w3586 and w3596;
w3598 <= not w3595 and not w3597;
w3599 <= not w3588 and not w3598;
w3600 <= not w845 and not w3599;
w3601 <= w3299 and not w3301;
w3602 <= not w3292 and w3601;
w3603 <= not w3462 and w3602;
w3604 <= not w3292 and not w3301;
w3605 <= not w3462 and w3604;
w3606 <= not w3299 and not w3605;
w3607 <= not w3603 and not w3606;
w3608 <= w845 and not w3588;
w3609 <= not w3598 and w3608;
w3610 <= not w3607 and not w3609;
w3611 <= not w3600 and not w3610;
w3612 <= not w705 and not w3611;
w3613 <= not w3304 and w3311;
w3614 <= not w3313 and w3613;
w3615 <= not w3462 and w3614;
w3616 <= not w3304 and not w3313;
w3617 <= not w3462 and w3616;
w3618 <= not w3311 and not w3617;
w3619 <= not w3615 and not w3618;
w3620 <= w705 and not w3600;
w3621 <= not w3610 and w3620;
w3622 <= not w3619 and not w3621;
w3623 <= not w3612 and not w3622;
w3624 <= not w577 and not w3623;
w3625 <= w3323 and not w3325;
w3626 <= not w3316 and w3625;
w3627 <= not w3462 and w3626;
w3628 <= not w3316 and not w3325;
w3629 <= not w3462 and w3628;
w3630 <= not w3323 and not w3629;
w3631 <= not w3627 and not w3630;
w3632 <= w577 and not w3612;
w3633 <= not w3622 and w3632;
w3634 <= not w3631 and not w3633;
w3635 <= not w3624 and not w3634;
w3636 <= not w460 and not w3635;
w3637 <= not w3328 and w3335;
w3638 <= not w3337 and w3637;
w3639 <= not w3462 and w3638;
w3640 <= not w3328 and not w3337;
w3641 <= not w3462 and w3640;
w3642 <= not w3335 and not w3641;
w3643 <= not w3639 and not w3642;
w3644 <= w460 and not w3624;
w3645 <= not w3634 and w3644;
w3646 <= not w3643 and not w3645;
w3647 <= not w3636 and not w3646;
w3648 <= not w356 and not w3647;
w3649 <= w3347 and not w3349;
w3650 <= not w3340 and w3649;
w3651 <= not w3462 and w3650;
w3652 <= not w3340 and not w3349;
w3653 <= not w3462 and w3652;
w3654 <= not w3347 and not w3653;
w3655 <= not w3651 and not w3654;
w3656 <= w356 and not w3636;
w3657 <= not w3646 and w3656;
w3658 <= not w3655 and not w3657;
w3659 <= not w3648 and not w3658;
w3660 <= not w264 and not w3659;
w3661 <= w264 and not w3648;
w3662 <= not w3658 and w3661;
w3663 <= not w3352 and w3361;
w3664 <= not w3354 and w3663;
w3665 <= not w3462 and w3664;
w3666 <= not w3352 and not w3354;
w3667 <= not w3462 and w3666;
w3668 <= not w3361 and not w3667;
w3669 <= not w3665 and not w3668;
w3670 <= not w3662 and not w3669;
w3671 <= not w3660 and not w3670;
w3672 <= not w184 and not w3671;
w3673 <= w3371 and not w3373;
w3674 <= not w3364 and w3673;
w3675 <= not w3462 and w3674;
w3676 <= not w3364 and not w3373;
w3677 <= not w3462 and w3676;
w3678 <= not w3371 and not w3677;
w3679 <= not w3675 and not w3678;
w3680 <= w184 and not w3660;
w3681 <= not w3670 and w3680;
w3682 <= not w3679 and not w3681;
w3683 <= not w3672 and not w3682;
w3684 <= not w115 and not w3683;
w3685 <= not w3376 and w3383;
w3686 <= not w3385 and w3685;
w3687 <= not w3462 and w3686;
w3688 <= not w3376 and not w3385;
w3689 <= not w3462 and w3688;
w3690 <= not w3383 and not w3689;
w3691 <= not w3687 and not w3690;
w3692 <= w115 and not w3672;
w3693 <= not w3682 and w3692;
w3694 <= not w3691 and not w3693;
w3695 <= not w3684 and not w3694;
w3696 <= not w60 and not w3695;
w3697 <= w3395 and not w3397;
w3698 <= not w3388 and w3697;
w3699 <= not w3462 and w3698;
w3700 <= not w3388 and not w3397;
w3701 <= not w3462 and w3700;
w3702 <= not w3395 and not w3701;
w3703 <= not w3699 and not w3702;
w3704 <= w60 and not w3684;
w3705 <= not w3694 and w3704;
w3706 <= not w3703 and not w3705;
w3707 <= not w3696 and not w3706;
w3708 <= not w22 and not w3707;
w3709 <= not w3400 and w3407;
w3710 <= not w3409 and w3709;
w3711 <= not w3462 and w3710;
w3712 <= not w3400 and not w3409;
w3713 <= not w3462 and w3712;
w3714 <= not w3407 and not w3713;
w3715 <= not w3711 and not w3714;
w3716 <= w22 and not w3696;
w3717 <= not w3706 and w3716;
w3718 <= not w3715 and not w3717;
w3719 <= not w3708 and not w3718;
w3720 <= not w5 and not w3719;
w3721 <= w3419 and not w3421;
w3722 <= not w3412 and w3721;
w3723 <= not w3462 and w3722;
w3724 <= not w3412 and not w3421;
w3725 <= not w3462 and w3724;
w3726 <= not w3419 and not w3725;
w3727 <= not w3723 and not w3726;
w3728 <= w5 and not w3708;
w3729 <= not w3718 and w3728;
w3730 <= not w3727 and not w3729;
w3731 <= not w3720 and not w3730;
w3732 <= not w3424 and w3431;
w3733 <= not w3433 and w3732;
w3734 <= not w3462 and w3733;
w3735 <= not w3424 and not w3433;
w3736 <= not w3462 and w3735;
w3737 <= not w3431 and not w3736;
w3738 <= not w3734 and not w3737;
w3739 <= not w3435 and not w3442;
w3740 <= not w3462 and w3739;
w3741 <= not w3450 and not w3740;
w3742 <= not w3738 and w3741;
w3743 <= not w3731 and w3742;
w3744 <= w0 and not w3743;
w3745 <= not w3720 and w3738;
w3746 <= not w3730 and w3745;
w3747 <= not w3442 and not w3462;
w3748 <= w3435 and not w3747;
w3749 <= not w0 and not w3739;
w3750 <= not w3748 and w3749;
w3751 <= not w3438 and not w3459;
w3752 <= not w3441 and w3751;
w3753 <= not w3454 and w3752;
w3754 <= not w3450 and w3753;
w3755 <= not w3448 and w3754;
w3756 <= not w3750 and not w3755;
w3757 <= not w3746 and w3756;
w3758 <= not w3744 and w3757;
w3759 <= a(78) and not w3758;
w3760 <= not a(76) and not a(77);
w3761 <= not a(78) and w3760;
w3762 <= not w3759 and not w3761;
w3763 <= not w3462 and not w3762;
w3764 <= not w3459 and not w3761;
w3765 <= not w3454 and w3764;
w3766 <= not w3450 and w3765;
w3767 <= not w3448 and w3766;
w3768 <= not w3759 and w3767;
w3769 <= not a(78) and not w3758;
w3770 <= a(79) and not w3769;
w3771 <= w3464 and not w3758;
w3772 <= not w3770 and not w3771;
w3773 <= not w3768 and w3772;
w3774 <= not w3763 and not w3773;
w3775 <= not w3178 and not w3774;
w3776 <= w3178 and not w3763;
w3777 <= not w3773 and w3776;
w3778 <= not w3462 and not w3755;
w3779 <= not w3750 and w3778;
w3780 <= not w3746 and w3779;
w3781 <= not w3744 and w3780;
w3782 <= not w3771 and not w3781;
w3783 <= a(80) and not w3782;
w3784 <= not a(80) and not w3781;
w3785 <= not w3771 and w3784;
w3786 <= not w3783 and not w3785;
w3787 <= not w3777 and not w3786;
w3788 <= not w3775 and not w3787;
w3789 <= not w2906 and not w3788;
w3790 <= not w3467 and not w3472;
w3791 <= not w3476 and w3790;
w3792 <= not w3758 and w3791;
w3793 <= not w3758 and w3790;
w3794 <= w3476 and not w3793;
w3795 <= not w3792 and not w3794;
w3796 <= w2906 and not w3775;
w3797 <= not w3787 and w3796;
w3798 <= not w3795 and not w3797;
w3799 <= not w3789 and not w3798;
w3800 <= not w2646 and not w3799;
w3801 <= not w3481 and w3490;
w3802 <= not w3479 and w3801;
w3803 <= not w3758 and w3802;
w3804 <= not w3479 and not w3481;
w3805 <= not w3758 and w3804;
w3806 <= not w3490 and not w3805;
w3807 <= not w3803 and not w3806;
w3808 <= w2646 and not w3789;
w3809 <= not w3798 and w3808;
w3810 <= not w3807 and not w3809;
w3811 <= not w3800 and not w3810;
w3812 <= not w2398 and not w3811;
w3813 <= not w3493 and w3499;
w3814 <= not w3501 and w3813;
w3815 <= not w3758 and w3814;
w3816 <= not w3493 and not w3501;
w3817 <= not w3758 and w3816;
w3818 <= not w3499 and not w3817;
w3819 <= not w3815 and not w3818;
w3820 <= w2398 and not w3800;
w3821 <= not w3810 and w3820;
w3822 <= not w3819 and not w3821;
w3823 <= not w3812 and not w3822;
w3824 <= not w2162 and not w3823;
w3825 <= w3511 and not w3513;
w3826 <= not w3504 and w3825;
w3827 <= not w3758 and w3826;
w3828 <= not w3504 and not w3513;
w3829 <= not w3758 and w3828;
w3830 <= not w3511 and not w3829;
w3831 <= not w3827 and not w3830;
w3832 <= w2162 and not w3812;
w3833 <= not w3822 and w3832;
w3834 <= not w3831 and not w3833;
w3835 <= not w3824 and not w3834;
w3836 <= not w1938 and not w3835;
w3837 <= not w3516 and w3523;
w3838 <= not w3525 and w3837;
w3839 <= not w3758 and w3838;
w3840 <= not w3516 and not w3525;
w3841 <= not w3758 and w3840;
w3842 <= not w3523 and not w3841;
w3843 <= not w3839 and not w3842;
w3844 <= w1938 and not w3824;
w3845 <= not w3834 and w3844;
w3846 <= not w3843 and not w3845;
w3847 <= not w3836 and not w3846;
w3848 <= not w1725 and not w3847;
w3849 <= w3535 and not w3537;
w3850 <= not w3528 and w3849;
w3851 <= not w3758 and w3850;
w3852 <= not w3528 and not w3537;
w3853 <= not w3758 and w3852;
w3854 <= not w3535 and not w3853;
w3855 <= not w3851 and not w3854;
w3856 <= w1725 and not w3836;
w3857 <= not w3846 and w3856;
w3858 <= not w3855 and not w3857;
w3859 <= not w3848 and not w3858;
w3860 <= not w1525 and not w3859;
w3861 <= not w3540 and w3547;
w3862 <= not w3549 and w3861;
w3863 <= not w3758 and w3862;
w3864 <= not w3540 and not w3549;
w3865 <= not w3758 and w3864;
w3866 <= not w3547 and not w3865;
w3867 <= not w3863 and not w3866;
w3868 <= w1525 and not w3848;
w3869 <= not w3858 and w3868;
w3870 <= not w3867 and not w3869;
w3871 <= not w3860 and not w3870;
w3872 <= not w1337 and not w3871;
w3873 <= w3559 and not w3561;
w3874 <= not w3552 and w3873;
w3875 <= not w3758 and w3874;
w3876 <= not w3552 and not w3561;
w3877 <= not w3758 and w3876;
w3878 <= not w3559 and not w3877;
w3879 <= not w3875 and not w3878;
w3880 <= w1337 and not w3860;
w3881 <= not w3870 and w3880;
w3882 <= not w3879 and not w3881;
w3883 <= not w3872 and not w3882;
w3884 <= not w1161 and not w3883;
w3885 <= not w3564 and w3571;
w3886 <= not w3573 and w3885;
w3887 <= not w3758 and w3886;
w3888 <= not w3564 and not w3573;
w3889 <= not w3758 and w3888;
w3890 <= not w3571 and not w3889;
w3891 <= not w3887 and not w3890;
w3892 <= w1161 and not w3872;
w3893 <= not w3882 and w3892;
w3894 <= not w3891 and not w3893;
w3895 <= not w3884 and not w3894;
w3896 <= not w997 and not w3895;
w3897 <= w3583 and not w3585;
w3898 <= not w3576 and w3897;
w3899 <= not w3758 and w3898;
w3900 <= not w3576 and not w3585;
w3901 <= not w3758 and w3900;
w3902 <= not w3583 and not w3901;
w3903 <= not w3899 and not w3902;
w3904 <= w997 and not w3884;
w3905 <= not w3894 and w3904;
w3906 <= not w3903 and not w3905;
w3907 <= not w3896 and not w3906;
w3908 <= not w845 and not w3907;
w3909 <= not w3588 and w3595;
w3910 <= not w3597 and w3909;
w3911 <= not w3758 and w3910;
w3912 <= not w3588 and not w3597;
w3913 <= not w3758 and w3912;
w3914 <= not w3595 and not w3913;
w3915 <= not w3911 and not w3914;
w3916 <= w845 and not w3896;
w3917 <= not w3906 and w3916;
w3918 <= not w3915 and not w3917;
w3919 <= not w3908 and not w3918;
w3920 <= not w705 and not w3919;
w3921 <= w3607 and not w3609;
w3922 <= not w3600 and w3921;
w3923 <= not w3758 and w3922;
w3924 <= not w3600 and not w3609;
w3925 <= not w3758 and w3924;
w3926 <= not w3607 and not w3925;
w3927 <= not w3923 and not w3926;
w3928 <= w705 and not w3908;
w3929 <= not w3918 and w3928;
w3930 <= not w3927 and not w3929;
w3931 <= not w3920 and not w3930;
w3932 <= not w577 and not w3931;
w3933 <= not w3612 and w3619;
w3934 <= not w3621 and w3933;
w3935 <= not w3758 and w3934;
w3936 <= not w3612 and not w3621;
w3937 <= not w3758 and w3936;
w3938 <= not w3619 and not w3937;
w3939 <= not w3935 and not w3938;
w3940 <= w577 and not w3920;
w3941 <= not w3930 and w3940;
w3942 <= not w3939 and not w3941;
w3943 <= not w3932 and not w3942;
w3944 <= not w460 and not w3943;
w3945 <= w3631 and not w3633;
w3946 <= not w3624 and w3945;
w3947 <= not w3758 and w3946;
w3948 <= not w3624 and not w3633;
w3949 <= not w3758 and w3948;
w3950 <= not w3631 and not w3949;
w3951 <= not w3947 and not w3950;
w3952 <= w460 and not w3932;
w3953 <= not w3942 and w3952;
w3954 <= not w3951 and not w3953;
w3955 <= not w3944 and not w3954;
w3956 <= not w356 and not w3955;
w3957 <= not w3636 and w3643;
w3958 <= not w3645 and w3957;
w3959 <= not w3758 and w3958;
w3960 <= not w3636 and not w3645;
w3961 <= not w3758 and w3960;
w3962 <= not w3643 and not w3961;
w3963 <= not w3959 and not w3962;
w3964 <= w356 and not w3944;
w3965 <= not w3954 and w3964;
w3966 <= not w3963 and not w3965;
w3967 <= not w3956 and not w3966;
w3968 <= not w264 and not w3967;
w3969 <= w3655 and not w3657;
w3970 <= not w3648 and w3969;
w3971 <= not w3758 and w3970;
w3972 <= not w3648 and not w3657;
w3973 <= not w3758 and w3972;
w3974 <= not w3655 and not w3973;
w3975 <= not w3971 and not w3974;
w3976 <= w264 and not w3956;
w3977 <= not w3966 and w3976;
w3978 <= not w3975 and not w3977;
w3979 <= not w3968 and not w3978;
w3980 <= not w184 and not w3979;
w3981 <= w184 and not w3968;
w3982 <= not w3978 and w3981;
w3983 <= not w3660 and w3669;
w3984 <= not w3662 and w3983;
w3985 <= not w3758 and w3984;
w3986 <= not w3660 and not w3662;
w3987 <= not w3758 and w3986;
w3988 <= not w3669 and not w3987;
w3989 <= not w3985 and not w3988;
w3990 <= not w3982 and not w3989;
w3991 <= not w3980 and not w3990;
w3992 <= not w115 and not w3991;
w3993 <= w3679 and not w3681;
w3994 <= not w3672 and w3993;
w3995 <= not w3758 and w3994;
w3996 <= not w3672 and not w3681;
w3997 <= not w3758 and w3996;
w3998 <= not w3679 and not w3997;
w3999 <= not w3995 and not w3998;
w4000 <= w115 and not w3980;
w4001 <= not w3990 and w4000;
w4002 <= not w3999 and not w4001;
w4003 <= not w3992 and not w4002;
w4004 <= not w60 and not w4003;
w4005 <= not w3684 and w3691;
w4006 <= not w3693 and w4005;
w4007 <= not w3758 and w4006;
w4008 <= not w3684 and not w3693;
w4009 <= not w3758 and w4008;
w4010 <= not w3691 and not w4009;
w4011 <= not w4007 and not w4010;
w4012 <= w60 and not w3992;
w4013 <= not w4002 and w4012;
w4014 <= not w4011 and not w4013;
w4015 <= not w4004 and not w4014;
w4016 <= not w22 and not w4015;
w4017 <= w3703 and not w3705;
w4018 <= not w3696 and w4017;
w4019 <= not w3758 and w4018;
w4020 <= not w3696 and not w3705;
w4021 <= not w3758 and w4020;
w4022 <= not w3703 and not w4021;
w4023 <= not w4019 and not w4022;
w4024 <= w22 and not w4004;
w4025 <= not w4014 and w4024;
w4026 <= not w4023 and not w4025;
w4027 <= not w4016 and not w4026;
w4028 <= not w5 and not w4027;
w4029 <= not w3708 and w3715;
w4030 <= not w3717 and w4029;
w4031 <= not w3758 and w4030;
w4032 <= not w3708 and not w3717;
w4033 <= not w3758 and w4032;
w4034 <= not w3715 and not w4033;
w4035 <= not w4031 and not w4034;
w4036 <= w5 and not w4016;
w4037 <= not w4026 and w4036;
w4038 <= not w4035 and not w4037;
w4039 <= not w4028 and not w4038;
w4040 <= w3727 and not w3729;
w4041 <= not w3720 and w4040;
w4042 <= not w3758 and w4041;
w4043 <= not w3720 and not w3729;
w4044 <= not w3758 and w4043;
w4045 <= not w3727 and not w4044;
w4046 <= not w4042 and not w4045;
w4047 <= not w3731 and not w3738;
w4048 <= not w3758 and w4047;
w4049 <= not w3746 and not w4048;
w4050 <= not w4046 and w4049;
w4051 <= not w4039 and w4050;
w4052 <= w0 and not w4051;
w4053 <= not w4028 and w4046;
w4054 <= not w4038 and w4053;
w4055 <= not w3738 and not w3758;
w4056 <= w3731 and not w4055;
w4057 <= not w0 and not w4047;
w4058 <= not w4056 and w4057;
w4059 <= not w3734 and not w3755;
w4060 <= not w3737 and w4059;
w4061 <= not w3750 and w4060;
w4062 <= not w3746 and w4061;
w4063 <= not w3744 and w4062;
w4064 <= not w4058 and not w4063;
w4065 <= not w4054 and w4064;
w4066 <= not w4052 and w4065;
w4067 <= a(76) and not w4066;
w4068 <= not a(74) and not a(75);
w4069 <= not a(76) and w4068;
w4070 <= not w4067 and not w4069;
w4071 <= not w3758 and not w4070;
w4072 <= not w3755 and not w4069;
w4073 <= not w3750 and w4072;
w4074 <= not w3746 and w4073;
w4075 <= not w3744 and w4074;
w4076 <= not w4067 and w4075;
w4077 <= not a(76) and not w4066;
w4078 <= a(77) and not w4077;
w4079 <= w3760 and not w4066;
w4080 <= not w4078 and not w4079;
w4081 <= not w4076 and w4080;
w4082 <= not w4071 and not w4081;
w4083 <= not w3462 and not w4082;
w4084 <= w3462 and not w4071;
w4085 <= not w4081 and w4084;
w4086 <= not w3758 and not w4063;
w4087 <= not w4058 and w4086;
w4088 <= not w4054 and w4087;
w4089 <= not w4052 and w4088;
w4090 <= not w4079 and not w4089;
w4091 <= a(78) and not w4090;
w4092 <= not a(78) and not w4089;
w4093 <= not w4079 and w4092;
w4094 <= not w4091 and not w4093;
w4095 <= not w4085 and not w4094;
w4096 <= not w4083 and not w4095;
w4097 <= not w3178 and not w4096;
w4098 <= not w3763 and not w3768;
w4099 <= not w3772 and w4098;
w4100 <= not w4066 and w4099;
w4101 <= not w4066 and w4098;
w4102 <= w3772 and not w4101;
w4103 <= not w4100 and not w4102;
w4104 <= w3178 and not w4083;
w4105 <= not w4095 and w4104;
w4106 <= not w4103 and not w4105;
w4107 <= not w4097 and not w4106;
w4108 <= not w2906 and not w4107;
w4109 <= not w3777 and w3786;
w4110 <= not w3775 and w4109;
w4111 <= not w4066 and w4110;
w4112 <= not w3775 and not w3777;
w4113 <= not w4066 and w4112;
w4114 <= not w3786 and not w4113;
w4115 <= not w4111 and not w4114;
w4116 <= w2906 and not w4097;
w4117 <= not w4106 and w4116;
w4118 <= not w4115 and not w4117;
w4119 <= not w4108 and not w4118;
w4120 <= not w2646 and not w4119;
w4121 <= not w3789 and w3795;
w4122 <= not w3797 and w4121;
w4123 <= not w4066 and w4122;
w4124 <= not w3789 and not w3797;
w4125 <= not w4066 and w4124;
w4126 <= not w3795 and not w4125;
w4127 <= not w4123 and not w4126;
w4128 <= w2646 and not w4108;
w4129 <= not w4118 and w4128;
w4130 <= not w4127 and not w4129;
w4131 <= not w4120 and not w4130;
w4132 <= not w2398 and not w4131;
w4133 <= w3807 and not w3809;
w4134 <= not w3800 and w4133;
w4135 <= not w4066 and w4134;
w4136 <= not w3800 and not w3809;
w4137 <= not w4066 and w4136;
w4138 <= not w3807 and not w4137;
w4139 <= not w4135 and not w4138;
w4140 <= w2398 and not w4120;
w4141 <= not w4130 and w4140;
w4142 <= not w4139 and not w4141;
w4143 <= not w4132 and not w4142;
w4144 <= not w2162 and not w4143;
w4145 <= not w3812 and w3819;
w4146 <= not w3821 and w4145;
w4147 <= not w4066 and w4146;
w4148 <= not w3812 and not w3821;
w4149 <= not w4066 and w4148;
w4150 <= not w3819 and not w4149;
w4151 <= not w4147 and not w4150;
w4152 <= w2162 and not w4132;
w4153 <= not w4142 and w4152;
w4154 <= not w4151 and not w4153;
w4155 <= not w4144 and not w4154;
w4156 <= not w1938 and not w4155;
w4157 <= w3831 and not w3833;
w4158 <= not w3824 and w4157;
w4159 <= not w4066 and w4158;
w4160 <= not w3824 and not w3833;
w4161 <= not w4066 and w4160;
w4162 <= not w3831 and not w4161;
w4163 <= not w4159 and not w4162;
w4164 <= w1938 and not w4144;
w4165 <= not w4154 and w4164;
w4166 <= not w4163 and not w4165;
w4167 <= not w4156 and not w4166;
w4168 <= not w1725 and not w4167;
w4169 <= not w3836 and w3843;
w4170 <= not w3845 and w4169;
w4171 <= not w4066 and w4170;
w4172 <= not w3836 and not w3845;
w4173 <= not w4066 and w4172;
w4174 <= not w3843 and not w4173;
w4175 <= not w4171 and not w4174;
w4176 <= w1725 and not w4156;
w4177 <= not w4166 and w4176;
w4178 <= not w4175 and not w4177;
w4179 <= not w4168 and not w4178;
w4180 <= not w1525 and not w4179;
w4181 <= w3855 and not w3857;
w4182 <= not w3848 and w4181;
w4183 <= not w4066 and w4182;
w4184 <= not w3848 and not w3857;
w4185 <= not w4066 and w4184;
w4186 <= not w3855 and not w4185;
w4187 <= not w4183 and not w4186;
w4188 <= w1525 and not w4168;
w4189 <= not w4178 and w4188;
w4190 <= not w4187 and not w4189;
w4191 <= not w4180 and not w4190;
w4192 <= not w1337 and not w4191;
w4193 <= not w3860 and w3867;
w4194 <= not w3869 and w4193;
w4195 <= not w4066 and w4194;
w4196 <= not w3860 and not w3869;
w4197 <= not w4066 and w4196;
w4198 <= not w3867 and not w4197;
w4199 <= not w4195 and not w4198;
w4200 <= w1337 and not w4180;
w4201 <= not w4190 and w4200;
w4202 <= not w4199 and not w4201;
w4203 <= not w4192 and not w4202;
w4204 <= not w1161 and not w4203;
w4205 <= w3879 and not w3881;
w4206 <= not w3872 and w4205;
w4207 <= not w4066 and w4206;
w4208 <= not w3872 and not w3881;
w4209 <= not w4066 and w4208;
w4210 <= not w3879 and not w4209;
w4211 <= not w4207 and not w4210;
w4212 <= w1161 and not w4192;
w4213 <= not w4202 and w4212;
w4214 <= not w4211 and not w4213;
w4215 <= not w4204 and not w4214;
w4216 <= not w997 and not w4215;
w4217 <= not w3884 and w3891;
w4218 <= not w3893 and w4217;
w4219 <= not w4066 and w4218;
w4220 <= not w3884 and not w3893;
w4221 <= not w4066 and w4220;
w4222 <= not w3891 and not w4221;
w4223 <= not w4219 and not w4222;
w4224 <= w997 and not w4204;
w4225 <= not w4214 and w4224;
w4226 <= not w4223 and not w4225;
w4227 <= not w4216 and not w4226;
w4228 <= not w845 and not w4227;
w4229 <= w3903 and not w3905;
w4230 <= not w3896 and w4229;
w4231 <= not w4066 and w4230;
w4232 <= not w3896 and not w3905;
w4233 <= not w4066 and w4232;
w4234 <= not w3903 and not w4233;
w4235 <= not w4231 and not w4234;
w4236 <= w845 and not w4216;
w4237 <= not w4226 and w4236;
w4238 <= not w4235 and not w4237;
w4239 <= not w4228 and not w4238;
w4240 <= not w705 and not w4239;
w4241 <= not w3908 and w3915;
w4242 <= not w3917 and w4241;
w4243 <= not w4066 and w4242;
w4244 <= not w3908 and not w3917;
w4245 <= not w4066 and w4244;
w4246 <= not w3915 and not w4245;
w4247 <= not w4243 and not w4246;
w4248 <= w705 and not w4228;
w4249 <= not w4238 and w4248;
w4250 <= not w4247 and not w4249;
w4251 <= not w4240 and not w4250;
w4252 <= not w577 and not w4251;
w4253 <= w3927 and not w3929;
w4254 <= not w3920 and w4253;
w4255 <= not w4066 and w4254;
w4256 <= not w3920 and not w3929;
w4257 <= not w4066 and w4256;
w4258 <= not w3927 and not w4257;
w4259 <= not w4255 and not w4258;
w4260 <= w577 and not w4240;
w4261 <= not w4250 and w4260;
w4262 <= not w4259 and not w4261;
w4263 <= not w4252 and not w4262;
w4264 <= not w460 and not w4263;
w4265 <= not w3932 and w3939;
w4266 <= not w3941 and w4265;
w4267 <= not w4066 and w4266;
w4268 <= not w3932 and not w3941;
w4269 <= not w4066 and w4268;
w4270 <= not w3939 and not w4269;
w4271 <= not w4267 and not w4270;
w4272 <= w460 and not w4252;
w4273 <= not w4262 and w4272;
w4274 <= not w4271 and not w4273;
w4275 <= not w4264 and not w4274;
w4276 <= not w356 and not w4275;
w4277 <= w3951 and not w3953;
w4278 <= not w3944 and w4277;
w4279 <= not w4066 and w4278;
w4280 <= not w3944 and not w3953;
w4281 <= not w4066 and w4280;
w4282 <= not w3951 and not w4281;
w4283 <= not w4279 and not w4282;
w4284 <= w356 and not w4264;
w4285 <= not w4274 and w4284;
w4286 <= not w4283 and not w4285;
w4287 <= not w4276 and not w4286;
w4288 <= not w264 and not w4287;
w4289 <= not w3956 and w3963;
w4290 <= not w3965 and w4289;
w4291 <= not w4066 and w4290;
w4292 <= not w3956 and not w3965;
w4293 <= not w4066 and w4292;
w4294 <= not w3963 and not w4293;
w4295 <= not w4291 and not w4294;
w4296 <= w264 and not w4276;
w4297 <= not w4286 and w4296;
w4298 <= not w4295 and not w4297;
w4299 <= not w4288 and not w4298;
w4300 <= not w184 and not w4299;
w4301 <= w3975 and not w3977;
w4302 <= not w3968 and w4301;
w4303 <= not w4066 and w4302;
w4304 <= not w3968 and not w3977;
w4305 <= not w4066 and w4304;
w4306 <= not w3975 and not w4305;
w4307 <= not w4303 and not w4306;
w4308 <= w184 and not w4288;
w4309 <= not w4298 and w4308;
w4310 <= not w4307 and not w4309;
w4311 <= not w4300 and not w4310;
w4312 <= not w115 and not w4311;
w4313 <= w115 and not w4300;
w4314 <= not w4310 and w4313;
w4315 <= not w3980 and w3989;
w4316 <= not w3982 and w4315;
w4317 <= not w4066 and w4316;
w4318 <= not w3980 and not w3982;
w4319 <= not w4066 and w4318;
w4320 <= not w3989 and not w4319;
w4321 <= not w4317 and not w4320;
w4322 <= not w4314 and not w4321;
w4323 <= not w4312 and not w4322;
w4324 <= not w60 and not w4323;
w4325 <= w3999 and not w4001;
w4326 <= not w3992 and w4325;
w4327 <= not w4066 and w4326;
w4328 <= not w3992 and not w4001;
w4329 <= not w4066 and w4328;
w4330 <= not w3999 and not w4329;
w4331 <= not w4327 and not w4330;
w4332 <= w60 and not w4312;
w4333 <= not w4322 and w4332;
w4334 <= not w4331 and not w4333;
w4335 <= not w4324 and not w4334;
w4336 <= not w22 and not w4335;
w4337 <= not w4004 and w4011;
w4338 <= not w4013 and w4337;
w4339 <= not w4066 and w4338;
w4340 <= not w4004 and not w4013;
w4341 <= not w4066 and w4340;
w4342 <= not w4011 and not w4341;
w4343 <= not w4339 and not w4342;
w4344 <= w22 and not w4324;
w4345 <= not w4334 and w4344;
w4346 <= not w4343 and not w4345;
w4347 <= not w4336 and not w4346;
w4348 <= not w5 and not w4347;
w4349 <= w4023 and not w4025;
w4350 <= not w4016 and w4349;
w4351 <= not w4066 and w4350;
w4352 <= not w4016 and not w4025;
w4353 <= not w4066 and w4352;
w4354 <= not w4023 and not w4353;
w4355 <= not w4351 and not w4354;
w4356 <= w5 and not w4336;
w4357 <= not w4346 and w4356;
w4358 <= not w4355 and not w4357;
w4359 <= not w4348 and not w4358;
w4360 <= not w4028 and w4035;
w4361 <= not w4037 and w4360;
w4362 <= not w4066 and w4361;
w4363 <= not w4028 and not w4037;
w4364 <= not w4066 and w4363;
w4365 <= not w4035 and not w4364;
w4366 <= not w4362 and not w4365;
w4367 <= not w4039 and not w4046;
w4368 <= not w4066 and w4367;
w4369 <= not w4054 and not w4368;
w4370 <= not w4366 and w4369;
w4371 <= not w4359 and w4370;
w4372 <= w0 and not w4371;
w4373 <= not w4348 and w4366;
w4374 <= not w4358 and w4373;
w4375 <= not w4046 and not w4066;
w4376 <= w4039 and not w4375;
w4377 <= not w0 and not w4367;
w4378 <= not w4376 and w4377;
w4379 <= not w4042 and not w4063;
w4380 <= not w4045 and w4379;
w4381 <= not w4058 and w4380;
w4382 <= not w4054 and w4381;
w4383 <= not w4052 and w4382;
w4384 <= not w4378 and not w4383;
w4385 <= not w4374 and w4384;
w4386 <= not w4372 and w4385;
w4387 <= a(74) and not w4386;
w4388 <= not a(72) and not a(73);
w4389 <= not a(74) and w4388;
w4390 <= not w4387 and not w4389;
w4391 <= not w4066 and not w4390;
w4392 <= not w4063 and not w4389;
w4393 <= not w4058 and w4392;
w4394 <= not w4054 and w4393;
w4395 <= not w4052 and w4394;
w4396 <= not w4387 and w4395;
w4397 <= not a(74) and not w4386;
w4398 <= a(75) and not w4397;
w4399 <= w4068 and not w4386;
w4400 <= not w4398 and not w4399;
w4401 <= not w4396 and w4400;
w4402 <= not w4391 and not w4401;
w4403 <= not w3758 and not w4402;
w4404 <= w3758 and not w4391;
w4405 <= not w4401 and w4404;
w4406 <= not w4066 and not w4383;
w4407 <= not w4378 and w4406;
w4408 <= not w4374 and w4407;
w4409 <= not w4372 and w4408;
w4410 <= not w4399 and not w4409;
w4411 <= a(76) and not w4410;
w4412 <= not a(76) and not w4409;
w4413 <= not w4399 and w4412;
w4414 <= not w4411 and not w4413;
w4415 <= not w4405 and not w4414;
w4416 <= not w4403 and not w4415;
w4417 <= not w3462 and not w4416;
w4418 <= not w4071 and not w4076;
w4419 <= not w4080 and w4418;
w4420 <= not w4386 and w4419;
w4421 <= not w4386 and w4418;
w4422 <= w4080 and not w4421;
w4423 <= not w4420 and not w4422;
w4424 <= w3462 and not w4403;
w4425 <= not w4415 and w4424;
w4426 <= not w4423 and not w4425;
w4427 <= not w4417 and not w4426;
w4428 <= not w3178 and not w4427;
w4429 <= not w4085 and w4094;
w4430 <= not w4083 and w4429;
w4431 <= not w4386 and w4430;
w4432 <= not w4083 and not w4085;
w4433 <= not w4386 and w4432;
w4434 <= not w4094 and not w4433;
w4435 <= not w4431 and not w4434;
w4436 <= w3178 and not w4417;
w4437 <= not w4426 and w4436;
w4438 <= not w4435 and not w4437;
w4439 <= not w4428 and not w4438;
w4440 <= not w2906 and not w4439;
w4441 <= not w4097 and w4103;
w4442 <= not w4105 and w4441;
w4443 <= not w4386 and w4442;
w4444 <= not w4097 and not w4105;
w4445 <= not w4386 and w4444;
w4446 <= not w4103 and not w4445;
w4447 <= not w4443 and not w4446;
w4448 <= w2906 and not w4428;
w4449 <= not w4438 and w4448;
w4450 <= not w4447 and not w4449;
w4451 <= not w4440 and not w4450;
w4452 <= not w2646 and not w4451;
w4453 <= w4115 and not w4117;
w4454 <= not w4108 and w4453;
w4455 <= not w4386 and w4454;
w4456 <= not w4108 and not w4117;
w4457 <= not w4386 and w4456;
w4458 <= not w4115 and not w4457;
w4459 <= not w4455 and not w4458;
w4460 <= w2646 and not w4440;
w4461 <= not w4450 and w4460;
w4462 <= not w4459 and not w4461;
w4463 <= not w4452 and not w4462;
w4464 <= not w2398 and not w4463;
w4465 <= not w4120 and w4127;
w4466 <= not w4129 and w4465;
w4467 <= not w4386 and w4466;
w4468 <= not w4120 and not w4129;
w4469 <= not w4386 and w4468;
w4470 <= not w4127 and not w4469;
w4471 <= not w4467 and not w4470;
w4472 <= w2398 and not w4452;
w4473 <= not w4462 and w4472;
w4474 <= not w4471 and not w4473;
w4475 <= not w4464 and not w4474;
w4476 <= not w2162 and not w4475;
w4477 <= w4139 and not w4141;
w4478 <= not w4132 and w4477;
w4479 <= not w4386 and w4478;
w4480 <= not w4132 and not w4141;
w4481 <= not w4386 and w4480;
w4482 <= not w4139 and not w4481;
w4483 <= not w4479 and not w4482;
w4484 <= w2162 and not w4464;
w4485 <= not w4474 and w4484;
w4486 <= not w4483 and not w4485;
w4487 <= not w4476 and not w4486;
w4488 <= not w1938 and not w4487;
w4489 <= not w4144 and w4151;
w4490 <= not w4153 and w4489;
w4491 <= not w4386 and w4490;
w4492 <= not w4144 and not w4153;
w4493 <= not w4386 and w4492;
w4494 <= not w4151 and not w4493;
w4495 <= not w4491 and not w4494;
w4496 <= w1938 and not w4476;
w4497 <= not w4486 and w4496;
w4498 <= not w4495 and not w4497;
w4499 <= not w4488 and not w4498;
w4500 <= not w1725 and not w4499;
w4501 <= w4163 and not w4165;
w4502 <= not w4156 and w4501;
w4503 <= not w4386 and w4502;
w4504 <= not w4156 and not w4165;
w4505 <= not w4386 and w4504;
w4506 <= not w4163 and not w4505;
w4507 <= not w4503 and not w4506;
w4508 <= w1725 and not w4488;
w4509 <= not w4498 and w4508;
w4510 <= not w4507 and not w4509;
w4511 <= not w4500 and not w4510;
w4512 <= not w1525 and not w4511;
w4513 <= not w4168 and w4175;
w4514 <= not w4177 and w4513;
w4515 <= not w4386 and w4514;
w4516 <= not w4168 and not w4177;
w4517 <= not w4386 and w4516;
w4518 <= not w4175 and not w4517;
w4519 <= not w4515 and not w4518;
w4520 <= w1525 and not w4500;
w4521 <= not w4510 and w4520;
w4522 <= not w4519 and not w4521;
w4523 <= not w4512 and not w4522;
w4524 <= not w1337 and not w4523;
w4525 <= w4187 and not w4189;
w4526 <= not w4180 and w4525;
w4527 <= not w4386 and w4526;
w4528 <= not w4180 and not w4189;
w4529 <= not w4386 and w4528;
w4530 <= not w4187 and not w4529;
w4531 <= not w4527 and not w4530;
w4532 <= w1337 and not w4512;
w4533 <= not w4522 and w4532;
w4534 <= not w4531 and not w4533;
w4535 <= not w4524 and not w4534;
w4536 <= not w1161 and not w4535;
w4537 <= not w4192 and w4199;
w4538 <= not w4201 and w4537;
w4539 <= not w4386 and w4538;
w4540 <= not w4192 and not w4201;
w4541 <= not w4386 and w4540;
w4542 <= not w4199 and not w4541;
w4543 <= not w4539 and not w4542;
w4544 <= w1161 and not w4524;
w4545 <= not w4534 and w4544;
w4546 <= not w4543 and not w4545;
w4547 <= not w4536 and not w4546;
w4548 <= not w997 and not w4547;
w4549 <= w4211 and not w4213;
w4550 <= not w4204 and w4549;
w4551 <= not w4386 and w4550;
w4552 <= not w4204 and not w4213;
w4553 <= not w4386 and w4552;
w4554 <= not w4211 and not w4553;
w4555 <= not w4551 and not w4554;
w4556 <= w997 and not w4536;
w4557 <= not w4546 and w4556;
w4558 <= not w4555 and not w4557;
w4559 <= not w4548 and not w4558;
w4560 <= not w845 and not w4559;
w4561 <= not w4216 and w4223;
w4562 <= not w4225 and w4561;
w4563 <= not w4386 and w4562;
w4564 <= not w4216 and not w4225;
w4565 <= not w4386 and w4564;
w4566 <= not w4223 and not w4565;
w4567 <= not w4563 and not w4566;
w4568 <= w845 and not w4548;
w4569 <= not w4558 and w4568;
w4570 <= not w4567 and not w4569;
w4571 <= not w4560 and not w4570;
w4572 <= not w705 and not w4571;
w4573 <= w4235 and not w4237;
w4574 <= not w4228 and w4573;
w4575 <= not w4386 and w4574;
w4576 <= not w4228 and not w4237;
w4577 <= not w4386 and w4576;
w4578 <= not w4235 and not w4577;
w4579 <= not w4575 and not w4578;
w4580 <= w705 and not w4560;
w4581 <= not w4570 and w4580;
w4582 <= not w4579 and not w4581;
w4583 <= not w4572 and not w4582;
w4584 <= not w577 and not w4583;
w4585 <= not w4240 and w4247;
w4586 <= not w4249 and w4585;
w4587 <= not w4386 and w4586;
w4588 <= not w4240 and not w4249;
w4589 <= not w4386 and w4588;
w4590 <= not w4247 and not w4589;
w4591 <= not w4587 and not w4590;
w4592 <= w577 and not w4572;
w4593 <= not w4582 and w4592;
w4594 <= not w4591 and not w4593;
w4595 <= not w4584 and not w4594;
w4596 <= not w460 and not w4595;
w4597 <= w4259 and not w4261;
w4598 <= not w4252 and w4597;
w4599 <= not w4386 and w4598;
w4600 <= not w4252 and not w4261;
w4601 <= not w4386 and w4600;
w4602 <= not w4259 and not w4601;
w4603 <= not w4599 and not w4602;
w4604 <= w460 and not w4584;
w4605 <= not w4594 and w4604;
w4606 <= not w4603 and not w4605;
w4607 <= not w4596 and not w4606;
w4608 <= not w356 and not w4607;
w4609 <= not w4264 and w4271;
w4610 <= not w4273 and w4609;
w4611 <= not w4386 and w4610;
w4612 <= not w4264 and not w4273;
w4613 <= not w4386 and w4612;
w4614 <= not w4271 and not w4613;
w4615 <= not w4611 and not w4614;
w4616 <= w356 and not w4596;
w4617 <= not w4606 and w4616;
w4618 <= not w4615 and not w4617;
w4619 <= not w4608 and not w4618;
w4620 <= not w264 and not w4619;
w4621 <= w4283 and not w4285;
w4622 <= not w4276 and w4621;
w4623 <= not w4386 and w4622;
w4624 <= not w4276 and not w4285;
w4625 <= not w4386 and w4624;
w4626 <= not w4283 and not w4625;
w4627 <= not w4623 and not w4626;
w4628 <= w264 and not w4608;
w4629 <= not w4618 and w4628;
w4630 <= not w4627 and not w4629;
w4631 <= not w4620 and not w4630;
w4632 <= not w184 and not w4631;
w4633 <= not w4288 and w4295;
w4634 <= not w4297 and w4633;
w4635 <= not w4386 and w4634;
w4636 <= not w4288 and not w4297;
w4637 <= not w4386 and w4636;
w4638 <= not w4295 and not w4637;
w4639 <= not w4635 and not w4638;
w4640 <= w184 and not w4620;
w4641 <= not w4630 and w4640;
w4642 <= not w4639 and not w4641;
w4643 <= not w4632 and not w4642;
w4644 <= not w115 and not w4643;
w4645 <= w4307 and not w4309;
w4646 <= not w4300 and w4645;
w4647 <= not w4386 and w4646;
w4648 <= not w4300 and not w4309;
w4649 <= not w4386 and w4648;
w4650 <= not w4307 and not w4649;
w4651 <= not w4647 and not w4650;
w4652 <= w115 and not w4632;
w4653 <= not w4642 and w4652;
w4654 <= not w4651 and not w4653;
w4655 <= not w4644 and not w4654;
w4656 <= not w60 and not w4655;
w4657 <= w60 and not w4644;
w4658 <= not w4654 and w4657;
w4659 <= not w4312 and w4321;
w4660 <= not w4314 and w4659;
w4661 <= not w4386 and w4660;
w4662 <= not w4312 and not w4314;
w4663 <= not w4386 and w4662;
w4664 <= not w4321 and not w4663;
w4665 <= not w4661 and not w4664;
w4666 <= not w4658 and not w4665;
w4667 <= not w4656 and not w4666;
w4668 <= not w22 and not w4667;
w4669 <= w4331 and not w4333;
w4670 <= not w4324 and w4669;
w4671 <= not w4386 and w4670;
w4672 <= not w4324 and not w4333;
w4673 <= not w4386 and w4672;
w4674 <= not w4331 and not w4673;
w4675 <= not w4671 and not w4674;
w4676 <= w22 and not w4656;
w4677 <= not w4666 and w4676;
w4678 <= not w4675 and not w4677;
w4679 <= not w4668 and not w4678;
w4680 <= not w5 and not w4679;
w4681 <= not w4336 and w4343;
w4682 <= not w4345 and w4681;
w4683 <= not w4386 and w4682;
w4684 <= not w4336 and not w4345;
w4685 <= not w4386 and w4684;
w4686 <= not w4343 and not w4685;
w4687 <= not w4683 and not w4686;
w4688 <= w5 and not w4668;
w4689 <= not w4678 and w4688;
w4690 <= not w4687 and not w4689;
w4691 <= not w4680 and not w4690;
w4692 <= w4355 and not w4357;
w4693 <= not w4348 and w4692;
w4694 <= not w4386 and w4693;
w4695 <= not w4348 and not w4357;
w4696 <= not w4386 and w4695;
w4697 <= not w4355 and not w4696;
w4698 <= not w4694 and not w4697;
w4699 <= not w4359 and not w4366;
w4700 <= not w4386 and w4699;
w4701 <= not w4374 and not w4700;
w4702 <= not w4698 and w4701;
w4703 <= not w4691 and w4702;
w4704 <= w0 and not w4703;
w4705 <= not w4680 and w4698;
w4706 <= not w4690 and w4705;
w4707 <= not w4366 and not w4386;
w4708 <= w4359 and not w4707;
w4709 <= not w0 and not w4699;
w4710 <= not w4708 and w4709;
w4711 <= not w4362 and not w4383;
w4712 <= not w4365 and w4711;
w4713 <= not w4378 and w4712;
w4714 <= not w4374 and w4713;
w4715 <= not w4372 and w4714;
w4716 <= not w4710 and not w4715;
w4717 <= not w4706 and w4716;
w4718 <= not w4704 and w4717;
w4719 <= a(72) and not w4718;
w4720 <= not a(70) and not a(71);
w4721 <= not a(72) and w4720;
w4722 <= not w4719 and not w4721;
w4723 <= not w4386 and not w4722;
w4724 <= not w4383 and not w4721;
w4725 <= not w4378 and w4724;
w4726 <= not w4374 and w4725;
w4727 <= not w4372 and w4726;
w4728 <= not w4719 and w4727;
w4729 <= not a(72) and not w4718;
w4730 <= a(73) and not w4729;
w4731 <= w4388 and not w4718;
w4732 <= not w4730 and not w4731;
w4733 <= not w4728 and w4732;
w4734 <= not w4723 and not w4733;
w4735 <= not w4066 and not w4734;
w4736 <= w4066 and not w4723;
w4737 <= not w4733 and w4736;
w4738 <= not w4386 and not w4715;
w4739 <= not w4710 and w4738;
w4740 <= not w4706 and w4739;
w4741 <= not w4704 and w4740;
w4742 <= not w4731 and not w4741;
w4743 <= a(74) and not w4742;
w4744 <= not a(74) and not w4741;
w4745 <= not w4731 and w4744;
w4746 <= not w4743 and not w4745;
w4747 <= not w4737 and not w4746;
w4748 <= not w4735 and not w4747;
w4749 <= not w3758 and not w4748;
w4750 <= not w4391 and not w4396;
w4751 <= not w4400 and w4750;
w4752 <= not w4718 and w4751;
w4753 <= not w4718 and w4750;
w4754 <= w4400 and not w4753;
w4755 <= not w4752 and not w4754;
w4756 <= w3758 and not w4735;
w4757 <= not w4747 and w4756;
w4758 <= not w4755 and not w4757;
w4759 <= not w4749 and not w4758;
w4760 <= not w3462 and not w4759;
w4761 <= not w4405 and w4414;
w4762 <= not w4403 and w4761;
w4763 <= not w4718 and w4762;
w4764 <= not w4403 and not w4405;
w4765 <= not w4718 and w4764;
w4766 <= not w4414 and not w4765;
w4767 <= not w4763 and not w4766;
w4768 <= w3462 and not w4749;
w4769 <= not w4758 and w4768;
w4770 <= not w4767 and not w4769;
w4771 <= not w4760 and not w4770;
w4772 <= not w3178 and not w4771;
w4773 <= not w4417 and w4423;
w4774 <= not w4425 and w4773;
w4775 <= not w4718 and w4774;
w4776 <= not w4417 and not w4425;
w4777 <= not w4718 and w4776;
w4778 <= not w4423 and not w4777;
w4779 <= not w4775 and not w4778;
w4780 <= w3178 and not w4760;
w4781 <= not w4770 and w4780;
w4782 <= not w4779 and not w4781;
w4783 <= not w4772 and not w4782;
w4784 <= not w2906 and not w4783;
w4785 <= w4435 and not w4437;
w4786 <= not w4428 and w4785;
w4787 <= not w4718 and w4786;
w4788 <= not w4428 and not w4437;
w4789 <= not w4718 and w4788;
w4790 <= not w4435 and not w4789;
w4791 <= not w4787 and not w4790;
w4792 <= w2906 and not w4772;
w4793 <= not w4782 and w4792;
w4794 <= not w4791 and not w4793;
w4795 <= not w4784 and not w4794;
w4796 <= not w2646 and not w4795;
w4797 <= not w4440 and w4447;
w4798 <= not w4449 and w4797;
w4799 <= not w4718 and w4798;
w4800 <= not w4440 and not w4449;
w4801 <= not w4718 and w4800;
w4802 <= not w4447 and not w4801;
w4803 <= not w4799 and not w4802;
w4804 <= w2646 and not w4784;
w4805 <= not w4794 and w4804;
w4806 <= not w4803 and not w4805;
w4807 <= not w4796 and not w4806;
w4808 <= not w2398 and not w4807;
w4809 <= w4459 and not w4461;
w4810 <= not w4452 and w4809;
w4811 <= not w4718 and w4810;
w4812 <= not w4452 and not w4461;
w4813 <= not w4718 and w4812;
w4814 <= not w4459 and not w4813;
w4815 <= not w4811 and not w4814;
w4816 <= w2398 and not w4796;
w4817 <= not w4806 and w4816;
w4818 <= not w4815 and not w4817;
w4819 <= not w4808 and not w4818;
w4820 <= not w2162 and not w4819;
w4821 <= not w4464 and w4471;
w4822 <= not w4473 and w4821;
w4823 <= not w4718 and w4822;
w4824 <= not w4464 and not w4473;
w4825 <= not w4718 and w4824;
w4826 <= not w4471 and not w4825;
w4827 <= not w4823 and not w4826;
w4828 <= w2162 and not w4808;
w4829 <= not w4818 and w4828;
w4830 <= not w4827 and not w4829;
w4831 <= not w4820 and not w4830;
w4832 <= not w1938 and not w4831;
w4833 <= w4483 and not w4485;
w4834 <= not w4476 and w4833;
w4835 <= not w4718 and w4834;
w4836 <= not w4476 and not w4485;
w4837 <= not w4718 and w4836;
w4838 <= not w4483 and not w4837;
w4839 <= not w4835 and not w4838;
w4840 <= w1938 and not w4820;
w4841 <= not w4830 and w4840;
w4842 <= not w4839 and not w4841;
w4843 <= not w4832 and not w4842;
w4844 <= not w1725 and not w4843;
w4845 <= not w4488 and w4495;
w4846 <= not w4497 and w4845;
w4847 <= not w4718 and w4846;
w4848 <= not w4488 and not w4497;
w4849 <= not w4718 and w4848;
w4850 <= not w4495 and not w4849;
w4851 <= not w4847 and not w4850;
w4852 <= w1725 and not w4832;
w4853 <= not w4842 and w4852;
w4854 <= not w4851 and not w4853;
w4855 <= not w4844 and not w4854;
w4856 <= not w1525 and not w4855;
w4857 <= w4507 and not w4509;
w4858 <= not w4500 and w4857;
w4859 <= not w4718 and w4858;
w4860 <= not w4500 and not w4509;
w4861 <= not w4718 and w4860;
w4862 <= not w4507 and not w4861;
w4863 <= not w4859 and not w4862;
w4864 <= w1525 and not w4844;
w4865 <= not w4854 and w4864;
w4866 <= not w4863 and not w4865;
w4867 <= not w4856 and not w4866;
w4868 <= not w1337 and not w4867;
w4869 <= not w4512 and w4519;
w4870 <= not w4521 and w4869;
w4871 <= not w4718 and w4870;
w4872 <= not w4512 and not w4521;
w4873 <= not w4718 and w4872;
w4874 <= not w4519 and not w4873;
w4875 <= not w4871 and not w4874;
w4876 <= w1337 and not w4856;
w4877 <= not w4866 and w4876;
w4878 <= not w4875 and not w4877;
w4879 <= not w4868 and not w4878;
w4880 <= not w1161 and not w4879;
w4881 <= w4531 and not w4533;
w4882 <= not w4524 and w4881;
w4883 <= not w4718 and w4882;
w4884 <= not w4524 and not w4533;
w4885 <= not w4718 and w4884;
w4886 <= not w4531 and not w4885;
w4887 <= not w4883 and not w4886;
w4888 <= w1161 and not w4868;
w4889 <= not w4878 and w4888;
w4890 <= not w4887 and not w4889;
w4891 <= not w4880 and not w4890;
w4892 <= not w997 and not w4891;
w4893 <= not w4536 and w4543;
w4894 <= not w4545 and w4893;
w4895 <= not w4718 and w4894;
w4896 <= not w4536 and not w4545;
w4897 <= not w4718 and w4896;
w4898 <= not w4543 and not w4897;
w4899 <= not w4895 and not w4898;
w4900 <= w997 and not w4880;
w4901 <= not w4890 and w4900;
w4902 <= not w4899 and not w4901;
w4903 <= not w4892 and not w4902;
w4904 <= not w845 and not w4903;
w4905 <= w4555 and not w4557;
w4906 <= not w4548 and w4905;
w4907 <= not w4718 and w4906;
w4908 <= not w4548 and not w4557;
w4909 <= not w4718 and w4908;
w4910 <= not w4555 and not w4909;
w4911 <= not w4907 and not w4910;
w4912 <= w845 and not w4892;
w4913 <= not w4902 and w4912;
w4914 <= not w4911 and not w4913;
w4915 <= not w4904 and not w4914;
w4916 <= not w705 and not w4915;
w4917 <= not w4560 and w4567;
w4918 <= not w4569 and w4917;
w4919 <= not w4718 and w4918;
w4920 <= not w4560 and not w4569;
w4921 <= not w4718 and w4920;
w4922 <= not w4567 and not w4921;
w4923 <= not w4919 and not w4922;
w4924 <= w705 and not w4904;
w4925 <= not w4914 and w4924;
w4926 <= not w4923 and not w4925;
w4927 <= not w4916 and not w4926;
w4928 <= not w577 and not w4927;
w4929 <= w4579 and not w4581;
w4930 <= not w4572 and w4929;
w4931 <= not w4718 and w4930;
w4932 <= not w4572 and not w4581;
w4933 <= not w4718 and w4932;
w4934 <= not w4579 and not w4933;
w4935 <= not w4931 and not w4934;
w4936 <= w577 and not w4916;
w4937 <= not w4926 and w4936;
w4938 <= not w4935 and not w4937;
w4939 <= not w4928 and not w4938;
w4940 <= not w460 and not w4939;
w4941 <= not w4584 and w4591;
w4942 <= not w4593 and w4941;
w4943 <= not w4718 and w4942;
w4944 <= not w4584 and not w4593;
w4945 <= not w4718 and w4944;
w4946 <= not w4591 and not w4945;
w4947 <= not w4943 and not w4946;
w4948 <= w460 and not w4928;
w4949 <= not w4938 and w4948;
w4950 <= not w4947 and not w4949;
w4951 <= not w4940 and not w4950;
w4952 <= not w356 and not w4951;
w4953 <= w4603 and not w4605;
w4954 <= not w4596 and w4953;
w4955 <= not w4718 and w4954;
w4956 <= not w4596 and not w4605;
w4957 <= not w4718 and w4956;
w4958 <= not w4603 and not w4957;
w4959 <= not w4955 and not w4958;
w4960 <= w356 and not w4940;
w4961 <= not w4950 and w4960;
w4962 <= not w4959 and not w4961;
w4963 <= not w4952 and not w4962;
w4964 <= not w264 and not w4963;
w4965 <= not w4608 and w4615;
w4966 <= not w4617 and w4965;
w4967 <= not w4718 and w4966;
w4968 <= not w4608 and not w4617;
w4969 <= not w4718 and w4968;
w4970 <= not w4615 and not w4969;
w4971 <= not w4967 and not w4970;
w4972 <= w264 and not w4952;
w4973 <= not w4962 and w4972;
w4974 <= not w4971 and not w4973;
w4975 <= not w4964 and not w4974;
w4976 <= not w184 and not w4975;
w4977 <= w4627 and not w4629;
w4978 <= not w4620 and w4977;
w4979 <= not w4718 and w4978;
w4980 <= not w4620 and not w4629;
w4981 <= not w4718 and w4980;
w4982 <= not w4627 and not w4981;
w4983 <= not w4979 and not w4982;
w4984 <= w184 and not w4964;
w4985 <= not w4974 and w4984;
w4986 <= not w4983 and not w4985;
w4987 <= not w4976 and not w4986;
w4988 <= not w115 and not w4987;
w4989 <= not w4632 and w4639;
w4990 <= not w4641 and w4989;
w4991 <= not w4718 and w4990;
w4992 <= not w4632 and not w4641;
w4993 <= not w4718 and w4992;
w4994 <= not w4639 and not w4993;
w4995 <= not w4991 and not w4994;
w4996 <= w115 and not w4976;
w4997 <= not w4986 and w4996;
w4998 <= not w4995 and not w4997;
w4999 <= not w4988 and not w4998;
w5000 <= not w60 and not w4999;
w5001 <= w4651 and not w4653;
w5002 <= not w4644 and w5001;
w5003 <= not w4718 and w5002;
w5004 <= not w4644 and not w4653;
w5005 <= not w4718 and w5004;
w5006 <= not w4651 and not w5005;
w5007 <= not w5003 and not w5006;
w5008 <= w60 and not w4988;
w5009 <= not w4998 and w5008;
w5010 <= not w5007 and not w5009;
w5011 <= not w5000 and not w5010;
w5012 <= not w22 and not w5011;
w5013 <= w22 and not w5000;
w5014 <= not w5010 and w5013;
w5015 <= not w4656 and w4665;
w5016 <= not w4658 and w5015;
w5017 <= not w4718 and w5016;
w5018 <= not w4656 and not w4658;
w5019 <= not w4718 and w5018;
w5020 <= not w4665 and not w5019;
w5021 <= not w5017 and not w5020;
w5022 <= not w5014 and not w5021;
w5023 <= not w5012 and not w5022;
w5024 <= not w5 and not w5023;
w5025 <= w4675 and not w4677;
w5026 <= not w4668 and w5025;
w5027 <= not w4718 and w5026;
w5028 <= not w4668 and not w4677;
w5029 <= not w4718 and w5028;
w5030 <= not w4675 and not w5029;
w5031 <= not w5027 and not w5030;
w5032 <= w5 and not w5012;
w5033 <= not w5022 and w5032;
w5034 <= not w5031 and not w5033;
w5035 <= not w5024 and not w5034;
w5036 <= not w4680 and w4687;
w5037 <= not w4689 and w5036;
w5038 <= not w4718 and w5037;
w5039 <= not w4680 and not w4689;
w5040 <= not w4718 and w5039;
w5041 <= not w4687 and not w5040;
w5042 <= not w5038 and not w5041;
w5043 <= not w4691 and not w4698;
w5044 <= not w4718 and w5043;
w5045 <= not w4706 and not w5044;
w5046 <= not w5042 and w5045;
w5047 <= not w5035 and w5046;
w5048 <= w0 and not w5047;
w5049 <= not w5024 and w5042;
w5050 <= not w5034 and w5049;
w5051 <= not w4698 and not w4718;
w5052 <= w4691 and not w5051;
w5053 <= not w0 and not w5043;
w5054 <= not w5052 and w5053;
w5055 <= not w4694 and not w4715;
w5056 <= not w4697 and w5055;
w5057 <= not w4710 and w5056;
w5058 <= not w4706 and w5057;
w5059 <= not w4704 and w5058;
w5060 <= not w5054 and not w5059;
w5061 <= not w5050 and w5060;
w5062 <= not w5048 and w5061;
w5063 <= a(70) and not w5062;
w5064 <= not a(68) and not a(69);
w5065 <= not a(70) and w5064;
w5066 <= not w5063 and not w5065;
w5067 <= not w4718 and not w5066;
w5068 <= not w4715 and not w5065;
w5069 <= not w4710 and w5068;
w5070 <= not w4706 and w5069;
w5071 <= not w4704 and w5070;
w5072 <= not w5063 and w5071;
w5073 <= not a(70) and not w5062;
w5074 <= a(71) and not w5073;
w5075 <= w4720 and not w5062;
w5076 <= not w5074 and not w5075;
w5077 <= not w5072 and w5076;
w5078 <= not w5067 and not w5077;
w5079 <= not w4386 and not w5078;
w5080 <= w4386 and not w5067;
w5081 <= not w5077 and w5080;
w5082 <= not w4718 and not w5059;
w5083 <= not w5054 and w5082;
w5084 <= not w5050 and w5083;
w5085 <= not w5048 and w5084;
w5086 <= not w5075 and not w5085;
w5087 <= a(72) and not w5086;
w5088 <= not a(72) and not w5085;
w5089 <= not w5075 and w5088;
w5090 <= not w5087 and not w5089;
w5091 <= not w5081 and not w5090;
w5092 <= not w5079 and not w5091;
w5093 <= not w4066 and not w5092;
w5094 <= not w4723 and not w4728;
w5095 <= not w4732 and w5094;
w5096 <= not w5062 and w5095;
w5097 <= not w5062 and w5094;
w5098 <= w4732 and not w5097;
w5099 <= not w5096 and not w5098;
w5100 <= w4066 and not w5079;
w5101 <= not w5091 and w5100;
w5102 <= not w5099 and not w5101;
w5103 <= not w5093 and not w5102;
w5104 <= not w3758 and not w5103;
w5105 <= not w4737 and w4746;
w5106 <= not w4735 and w5105;
w5107 <= not w5062 and w5106;
w5108 <= not w4735 and not w4737;
w5109 <= not w5062 and w5108;
w5110 <= not w4746 and not w5109;
w5111 <= not w5107 and not w5110;
w5112 <= w3758 and not w5093;
w5113 <= not w5102 and w5112;
w5114 <= not w5111 and not w5113;
w5115 <= not w5104 and not w5114;
w5116 <= not w3462 and not w5115;
w5117 <= not w4749 and w4755;
w5118 <= not w4757 and w5117;
w5119 <= not w5062 and w5118;
w5120 <= not w4749 and not w4757;
w5121 <= not w5062 and w5120;
w5122 <= not w4755 and not w5121;
w5123 <= not w5119 and not w5122;
w5124 <= w3462 and not w5104;
w5125 <= not w5114 and w5124;
w5126 <= not w5123 and not w5125;
w5127 <= not w5116 and not w5126;
w5128 <= not w3178 and not w5127;
w5129 <= w4767 and not w4769;
w5130 <= not w4760 and w5129;
w5131 <= not w5062 and w5130;
w5132 <= not w4760 and not w4769;
w5133 <= not w5062 and w5132;
w5134 <= not w4767 and not w5133;
w5135 <= not w5131 and not w5134;
w5136 <= w3178 and not w5116;
w5137 <= not w5126 and w5136;
w5138 <= not w5135 and not w5137;
w5139 <= not w5128 and not w5138;
w5140 <= not w2906 and not w5139;
w5141 <= not w4772 and w4779;
w5142 <= not w4781 and w5141;
w5143 <= not w5062 and w5142;
w5144 <= not w4772 and not w4781;
w5145 <= not w5062 and w5144;
w5146 <= not w4779 and not w5145;
w5147 <= not w5143 and not w5146;
w5148 <= w2906 and not w5128;
w5149 <= not w5138 and w5148;
w5150 <= not w5147 and not w5149;
w5151 <= not w5140 and not w5150;
w5152 <= not w2646 and not w5151;
w5153 <= w4791 and not w4793;
w5154 <= not w4784 and w5153;
w5155 <= not w5062 and w5154;
w5156 <= not w4784 and not w4793;
w5157 <= not w5062 and w5156;
w5158 <= not w4791 and not w5157;
w5159 <= not w5155 and not w5158;
w5160 <= w2646 and not w5140;
w5161 <= not w5150 and w5160;
w5162 <= not w5159 and not w5161;
w5163 <= not w5152 and not w5162;
w5164 <= not w2398 and not w5163;
w5165 <= not w4796 and w4803;
w5166 <= not w4805 and w5165;
w5167 <= not w5062 and w5166;
w5168 <= not w4796 and not w4805;
w5169 <= not w5062 and w5168;
w5170 <= not w4803 and not w5169;
w5171 <= not w5167 and not w5170;
w5172 <= w2398 and not w5152;
w5173 <= not w5162 and w5172;
w5174 <= not w5171 and not w5173;
w5175 <= not w5164 and not w5174;
w5176 <= not w2162 and not w5175;
w5177 <= w4815 and not w4817;
w5178 <= not w4808 and w5177;
w5179 <= not w5062 and w5178;
w5180 <= not w4808 and not w4817;
w5181 <= not w5062 and w5180;
w5182 <= not w4815 and not w5181;
w5183 <= not w5179 and not w5182;
w5184 <= w2162 and not w5164;
w5185 <= not w5174 and w5184;
w5186 <= not w5183 and not w5185;
w5187 <= not w5176 and not w5186;
w5188 <= not w1938 and not w5187;
w5189 <= not w4820 and w4827;
w5190 <= not w4829 and w5189;
w5191 <= not w5062 and w5190;
w5192 <= not w4820 and not w4829;
w5193 <= not w5062 and w5192;
w5194 <= not w4827 and not w5193;
w5195 <= not w5191 and not w5194;
w5196 <= w1938 and not w5176;
w5197 <= not w5186 and w5196;
w5198 <= not w5195 and not w5197;
w5199 <= not w5188 and not w5198;
w5200 <= not w1725 and not w5199;
w5201 <= w4839 and not w4841;
w5202 <= not w4832 and w5201;
w5203 <= not w5062 and w5202;
w5204 <= not w4832 and not w4841;
w5205 <= not w5062 and w5204;
w5206 <= not w4839 and not w5205;
w5207 <= not w5203 and not w5206;
w5208 <= w1725 and not w5188;
w5209 <= not w5198 and w5208;
w5210 <= not w5207 and not w5209;
w5211 <= not w5200 and not w5210;
w5212 <= not w1525 and not w5211;
w5213 <= not w4844 and w4851;
w5214 <= not w4853 and w5213;
w5215 <= not w5062 and w5214;
w5216 <= not w4844 and not w4853;
w5217 <= not w5062 and w5216;
w5218 <= not w4851 and not w5217;
w5219 <= not w5215 and not w5218;
w5220 <= w1525 and not w5200;
w5221 <= not w5210 and w5220;
w5222 <= not w5219 and not w5221;
w5223 <= not w5212 and not w5222;
w5224 <= not w1337 and not w5223;
w5225 <= w4863 and not w4865;
w5226 <= not w4856 and w5225;
w5227 <= not w5062 and w5226;
w5228 <= not w4856 and not w4865;
w5229 <= not w5062 and w5228;
w5230 <= not w4863 and not w5229;
w5231 <= not w5227 and not w5230;
w5232 <= w1337 and not w5212;
w5233 <= not w5222 and w5232;
w5234 <= not w5231 and not w5233;
w5235 <= not w5224 and not w5234;
w5236 <= not w1161 and not w5235;
w5237 <= not w4868 and w4875;
w5238 <= not w4877 and w5237;
w5239 <= not w5062 and w5238;
w5240 <= not w4868 and not w4877;
w5241 <= not w5062 and w5240;
w5242 <= not w4875 and not w5241;
w5243 <= not w5239 and not w5242;
w5244 <= w1161 and not w5224;
w5245 <= not w5234 and w5244;
w5246 <= not w5243 and not w5245;
w5247 <= not w5236 and not w5246;
w5248 <= not w997 and not w5247;
w5249 <= w4887 and not w4889;
w5250 <= not w4880 and w5249;
w5251 <= not w5062 and w5250;
w5252 <= not w4880 and not w4889;
w5253 <= not w5062 and w5252;
w5254 <= not w4887 and not w5253;
w5255 <= not w5251 and not w5254;
w5256 <= w997 and not w5236;
w5257 <= not w5246 and w5256;
w5258 <= not w5255 and not w5257;
w5259 <= not w5248 and not w5258;
w5260 <= not w845 and not w5259;
w5261 <= not w4892 and w4899;
w5262 <= not w4901 and w5261;
w5263 <= not w5062 and w5262;
w5264 <= not w4892 and not w4901;
w5265 <= not w5062 and w5264;
w5266 <= not w4899 and not w5265;
w5267 <= not w5263 and not w5266;
w5268 <= w845 and not w5248;
w5269 <= not w5258 and w5268;
w5270 <= not w5267 and not w5269;
w5271 <= not w5260 and not w5270;
w5272 <= not w705 and not w5271;
w5273 <= w4911 and not w4913;
w5274 <= not w4904 and w5273;
w5275 <= not w5062 and w5274;
w5276 <= not w4904 and not w4913;
w5277 <= not w5062 and w5276;
w5278 <= not w4911 and not w5277;
w5279 <= not w5275 and not w5278;
w5280 <= w705 and not w5260;
w5281 <= not w5270 and w5280;
w5282 <= not w5279 and not w5281;
w5283 <= not w5272 and not w5282;
w5284 <= not w577 and not w5283;
w5285 <= not w4916 and w4923;
w5286 <= not w4925 and w5285;
w5287 <= not w5062 and w5286;
w5288 <= not w4916 and not w4925;
w5289 <= not w5062 and w5288;
w5290 <= not w4923 and not w5289;
w5291 <= not w5287 and not w5290;
w5292 <= w577 and not w5272;
w5293 <= not w5282 and w5292;
w5294 <= not w5291 and not w5293;
w5295 <= not w5284 and not w5294;
w5296 <= not w460 and not w5295;
w5297 <= w4935 and not w4937;
w5298 <= not w4928 and w5297;
w5299 <= not w5062 and w5298;
w5300 <= not w4928 and not w4937;
w5301 <= not w5062 and w5300;
w5302 <= not w4935 and not w5301;
w5303 <= not w5299 and not w5302;
w5304 <= w460 and not w5284;
w5305 <= not w5294 and w5304;
w5306 <= not w5303 and not w5305;
w5307 <= not w5296 and not w5306;
w5308 <= not w356 and not w5307;
w5309 <= not w4940 and w4947;
w5310 <= not w4949 and w5309;
w5311 <= not w5062 and w5310;
w5312 <= not w4940 and not w4949;
w5313 <= not w5062 and w5312;
w5314 <= not w4947 and not w5313;
w5315 <= not w5311 and not w5314;
w5316 <= w356 and not w5296;
w5317 <= not w5306 and w5316;
w5318 <= not w5315 and not w5317;
w5319 <= not w5308 and not w5318;
w5320 <= not w264 and not w5319;
w5321 <= w4959 and not w4961;
w5322 <= not w4952 and w5321;
w5323 <= not w5062 and w5322;
w5324 <= not w4952 and not w4961;
w5325 <= not w5062 and w5324;
w5326 <= not w4959 and not w5325;
w5327 <= not w5323 and not w5326;
w5328 <= w264 and not w5308;
w5329 <= not w5318 and w5328;
w5330 <= not w5327 and not w5329;
w5331 <= not w5320 and not w5330;
w5332 <= not w184 and not w5331;
w5333 <= not w4964 and w4971;
w5334 <= not w4973 and w5333;
w5335 <= not w5062 and w5334;
w5336 <= not w4964 and not w4973;
w5337 <= not w5062 and w5336;
w5338 <= not w4971 and not w5337;
w5339 <= not w5335 and not w5338;
w5340 <= w184 and not w5320;
w5341 <= not w5330 and w5340;
w5342 <= not w5339 and not w5341;
w5343 <= not w5332 and not w5342;
w5344 <= not w115 and not w5343;
w5345 <= w4983 and not w4985;
w5346 <= not w4976 and w5345;
w5347 <= not w5062 and w5346;
w5348 <= not w4976 and not w4985;
w5349 <= not w5062 and w5348;
w5350 <= not w4983 and not w5349;
w5351 <= not w5347 and not w5350;
w5352 <= w115 and not w5332;
w5353 <= not w5342 and w5352;
w5354 <= not w5351 and not w5353;
w5355 <= not w5344 and not w5354;
w5356 <= not w60 and not w5355;
w5357 <= not w4988 and w4995;
w5358 <= not w4997 and w5357;
w5359 <= not w5062 and w5358;
w5360 <= not w4988 and not w4997;
w5361 <= not w5062 and w5360;
w5362 <= not w4995 and not w5361;
w5363 <= not w5359 and not w5362;
w5364 <= w60 and not w5344;
w5365 <= not w5354 and w5364;
w5366 <= not w5363 and not w5365;
w5367 <= not w5356 and not w5366;
w5368 <= not w22 and not w5367;
w5369 <= w5007 and not w5009;
w5370 <= not w5000 and w5369;
w5371 <= not w5062 and w5370;
w5372 <= not w5000 and not w5009;
w5373 <= not w5062 and w5372;
w5374 <= not w5007 and not w5373;
w5375 <= not w5371 and not w5374;
w5376 <= w22 and not w5356;
w5377 <= not w5366 and w5376;
w5378 <= not w5375 and not w5377;
w5379 <= not w5368 and not w5378;
w5380 <= not w5 and not w5379;
w5381 <= w5 and not w5368;
w5382 <= not w5378 and w5381;
w5383 <= not w5012 and w5021;
w5384 <= not w5014 and w5383;
w5385 <= not w5062 and w5384;
w5386 <= not w5012 and not w5014;
w5387 <= not w5062 and w5386;
w5388 <= not w5021 and not w5387;
w5389 <= not w5385 and not w5388;
w5390 <= not w5382 and not w5389;
w5391 <= not w5380 and not w5390;
w5392 <= w5031 and not w5033;
w5393 <= not w5024 and w5392;
w5394 <= not w5062 and w5393;
w5395 <= not w5024 and not w5033;
w5396 <= not w5062 and w5395;
w5397 <= not w5031 and not w5396;
w5398 <= not w5394 and not w5397;
w5399 <= not w5035 and not w5042;
w5400 <= not w5062 and w5399;
w5401 <= not w5050 and not w5400;
w5402 <= not w5398 and w5401;
w5403 <= not w5391 and w5402;
w5404 <= w0 and not w5403;
w5405 <= not w5380 and w5398;
w5406 <= not w5390 and w5405;
w5407 <= not w5042 and not w5062;
w5408 <= w5035 and not w5407;
w5409 <= not w0 and not w5399;
w5410 <= not w5408 and w5409;
w5411 <= not w5038 and not w5059;
w5412 <= not w5041 and w5411;
w5413 <= not w5054 and w5412;
w5414 <= not w5050 and w5413;
w5415 <= not w5048 and w5414;
w5416 <= not w5410 and not w5415;
w5417 <= not w5406 and w5416;
w5418 <= not w5404 and w5417;
w5419 <= a(68) and not w5418;
w5420 <= not a(66) and not a(67);
w5421 <= not a(68) and w5420;
w5422 <= not w5419 and not w5421;
w5423 <= not w5062 and not w5422;
w5424 <= not w5059 and not w5421;
w5425 <= not w5054 and w5424;
w5426 <= not w5050 and w5425;
w5427 <= not w5048 and w5426;
w5428 <= not w5419 and w5427;
w5429 <= not a(68) and not w5418;
w5430 <= a(69) and not w5429;
w5431 <= w5064 and not w5418;
w5432 <= not w5430 and not w5431;
w5433 <= not w5428 and w5432;
w5434 <= not w5423 and not w5433;
w5435 <= not w4718 and not w5434;
w5436 <= w4718 and not w5423;
w5437 <= not w5433 and w5436;
w5438 <= not w5062 and not w5415;
w5439 <= not w5410 and w5438;
w5440 <= not w5406 and w5439;
w5441 <= not w5404 and w5440;
w5442 <= not w5431 and not w5441;
w5443 <= a(70) and not w5442;
w5444 <= not a(70) and not w5441;
w5445 <= not w5431 and w5444;
w5446 <= not w5443 and not w5445;
w5447 <= not w5437 and not w5446;
w5448 <= not w5435 and not w5447;
w5449 <= not w4386 and not w5448;
w5450 <= not w5067 and not w5072;
w5451 <= not w5076 and w5450;
w5452 <= not w5418 and w5451;
w5453 <= not w5418 and w5450;
w5454 <= w5076 and not w5453;
w5455 <= not w5452 and not w5454;
w5456 <= w4386 and not w5435;
w5457 <= not w5447 and w5456;
w5458 <= not w5455 and not w5457;
w5459 <= not w5449 and not w5458;
w5460 <= not w4066 and not w5459;
w5461 <= not w5081 and w5090;
w5462 <= not w5079 and w5461;
w5463 <= not w5418 and w5462;
w5464 <= not w5079 and not w5081;
w5465 <= not w5418 and w5464;
w5466 <= not w5090 and not w5465;
w5467 <= not w5463 and not w5466;
w5468 <= w4066 and not w5449;
w5469 <= not w5458 and w5468;
w5470 <= not w5467 and not w5469;
w5471 <= not w5460 and not w5470;
w5472 <= not w3758 and not w5471;
w5473 <= not w5093 and w5099;
w5474 <= not w5101 and w5473;
w5475 <= not w5418 and w5474;
w5476 <= not w5093 and not w5101;
w5477 <= not w5418 and w5476;
w5478 <= not w5099 and not w5477;
w5479 <= not w5475 and not w5478;
w5480 <= w3758 and not w5460;
w5481 <= not w5470 and w5480;
w5482 <= not w5479 and not w5481;
w5483 <= not w5472 and not w5482;
w5484 <= not w3462 and not w5483;
w5485 <= w5111 and not w5113;
w5486 <= not w5104 and w5485;
w5487 <= not w5418 and w5486;
w5488 <= not w5104 and not w5113;
w5489 <= not w5418 and w5488;
w5490 <= not w5111 and not w5489;
w5491 <= not w5487 and not w5490;
w5492 <= w3462 and not w5472;
w5493 <= not w5482 and w5492;
w5494 <= not w5491 and not w5493;
w5495 <= not w5484 and not w5494;
w5496 <= not w3178 and not w5495;
w5497 <= not w5116 and w5123;
w5498 <= not w5125 and w5497;
w5499 <= not w5418 and w5498;
w5500 <= not w5116 and not w5125;
w5501 <= not w5418 and w5500;
w5502 <= not w5123 and not w5501;
w5503 <= not w5499 and not w5502;
w5504 <= w3178 and not w5484;
w5505 <= not w5494 and w5504;
w5506 <= not w5503 and not w5505;
w5507 <= not w5496 and not w5506;
w5508 <= not w2906 and not w5507;
w5509 <= w5135 and not w5137;
w5510 <= not w5128 and w5509;
w5511 <= not w5418 and w5510;
w5512 <= not w5128 and not w5137;
w5513 <= not w5418 and w5512;
w5514 <= not w5135 and not w5513;
w5515 <= not w5511 and not w5514;
w5516 <= w2906 and not w5496;
w5517 <= not w5506 and w5516;
w5518 <= not w5515 and not w5517;
w5519 <= not w5508 and not w5518;
w5520 <= not w2646 and not w5519;
w5521 <= not w5140 and w5147;
w5522 <= not w5149 and w5521;
w5523 <= not w5418 and w5522;
w5524 <= not w5140 and not w5149;
w5525 <= not w5418 and w5524;
w5526 <= not w5147 and not w5525;
w5527 <= not w5523 and not w5526;
w5528 <= w2646 and not w5508;
w5529 <= not w5518 and w5528;
w5530 <= not w5527 and not w5529;
w5531 <= not w5520 and not w5530;
w5532 <= not w2398 and not w5531;
w5533 <= w5159 and not w5161;
w5534 <= not w5152 and w5533;
w5535 <= not w5418 and w5534;
w5536 <= not w5152 and not w5161;
w5537 <= not w5418 and w5536;
w5538 <= not w5159 and not w5537;
w5539 <= not w5535 and not w5538;
w5540 <= w2398 and not w5520;
w5541 <= not w5530 and w5540;
w5542 <= not w5539 and not w5541;
w5543 <= not w5532 and not w5542;
w5544 <= not w2162 and not w5543;
w5545 <= not w5164 and w5171;
w5546 <= not w5173 and w5545;
w5547 <= not w5418 and w5546;
w5548 <= not w5164 and not w5173;
w5549 <= not w5418 and w5548;
w5550 <= not w5171 and not w5549;
w5551 <= not w5547 and not w5550;
w5552 <= w2162 and not w5532;
w5553 <= not w5542 and w5552;
w5554 <= not w5551 and not w5553;
w5555 <= not w5544 and not w5554;
w5556 <= not w1938 and not w5555;
w5557 <= w5183 and not w5185;
w5558 <= not w5176 and w5557;
w5559 <= not w5418 and w5558;
w5560 <= not w5176 and not w5185;
w5561 <= not w5418 and w5560;
w5562 <= not w5183 and not w5561;
w5563 <= not w5559 and not w5562;
w5564 <= w1938 and not w5544;
w5565 <= not w5554 and w5564;
w5566 <= not w5563 and not w5565;
w5567 <= not w5556 and not w5566;
w5568 <= not w1725 and not w5567;
w5569 <= not w5188 and w5195;
w5570 <= not w5197 and w5569;
w5571 <= not w5418 and w5570;
w5572 <= not w5188 and not w5197;
w5573 <= not w5418 and w5572;
w5574 <= not w5195 and not w5573;
w5575 <= not w5571 and not w5574;
w5576 <= w1725 and not w5556;
w5577 <= not w5566 and w5576;
w5578 <= not w5575 and not w5577;
w5579 <= not w5568 and not w5578;
w5580 <= not w1525 and not w5579;
w5581 <= w5207 and not w5209;
w5582 <= not w5200 and w5581;
w5583 <= not w5418 and w5582;
w5584 <= not w5200 and not w5209;
w5585 <= not w5418 and w5584;
w5586 <= not w5207 and not w5585;
w5587 <= not w5583 and not w5586;
w5588 <= w1525 and not w5568;
w5589 <= not w5578 and w5588;
w5590 <= not w5587 and not w5589;
w5591 <= not w5580 and not w5590;
w5592 <= not w1337 and not w5591;
w5593 <= not w5212 and w5219;
w5594 <= not w5221 and w5593;
w5595 <= not w5418 and w5594;
w5596 <= not w5212 and not w5221;
w5597 <= not w5418 and w5596;
w5598 <= not w5219 and not w5597;
w5599 <= not w5595 and not w5598;
w5600 <= w1337 and not w5580;
w5601 <= not w5590 and w5600;
w5602 <= not w5599 and not w5601;
w5603 <= not w5592 and not w5602;
w5604 <= not w1161 and not w5603;
w5605 <= w5231 and not w5233;
w5606 <= not w5224 and w5605;
w5607 <= not w5418 and w5606;
w5608 <= not w5224 and not w5233;
w5609 <= not w5418 and w5608;
w5610 <= not w5231 and not w5609;
w5611 <= not w5607 and not w5610;
w5612 <= w1161 and not w5592;
w5613 <= not w5602 and w5612;
w5614 <= not w5611 and not w5613;
w5615 <= not w5604 and not w5614;
w5616 <= not w997 and not w5615;
w5617 <= not w5236 and w5243;
w5618 <= not w5245 and w5617;
w5619 <= not w5418 and w5618;
w5620 <= not w5236 and not w5245;
w5621 <= not w5418 and w5620;
w5622 <= not w5243 and not w5621;
w5623 <= not w5619 and not w5622;
w5624 <= w997 and not w5604;
w5625 <= not w5614 and w5624;
w5626 <= not w5623 and not w5625;
w5627 <= not w5616 and not w5626;
w5628 <= not w845 and not w5627;
w5629 <= w5255 and not w5257;
w5630 <= not w5248 and w5629;
w5631 <= not w5418 and w5630;
w5632 <= not w5248 and not w5257;
w5633 <= not w5418 and w5632;
w5634 <= not w5255 and not w5633;
w5635 <= not w5631 and not w5634;
w5636 <= w845 and not w5616;
w5637 <= not w5626 and w5636;
w5638 <= not w5635 and not w5637;
w5639 <= not w5628 and not w5638;
w5640 <= not w705 and not w5639;
w5641 <= not w5260 and w5267;
w5642 <= not w5269 and w5641;
w5643 <= not w5418 and w5642;
w5644 <= not w5260 and not w5269;
w5645 <= not w5418 and w5644;
w5646 <= not w5267 and not w5645;
w5647 <= not w5643 and not w5646;
w5648 <= w705 and not w5628;
w5649 <= not w5638 and w5648;
w5650 <= not w5647 and not w5649;
w5651 <= not w5640 and not w5650;
w5652 <= not w577 and not w5651;
w5653 <= w5279 and not w5281;
w5654 <= not w5272 and w5653;
w5655 <= not w5418 and w5654;
w5656 <= not w5272 and not w5281;
w5657 <= not w5418 and w5656;
w5658 <= not w5279 and not w5657;
w5659 <= not w5655 and not w5658;
w5660 <= w577 and not w5640;
w5661 <= not w5650 and w5660;
w5662 <= not w5659 and not w5661;
w5663 <= not w5652 and not w5662;
w5664 <= not w460 and not w5663;
w5665 <= not w5284 and w5291;
w5666 <= not w5293 and w5665;
w5667 <= not w5418 and w5666;
w5668 <= not w5284 and not w5293;
w5669 <= not w5418 and w5668;
w5670 <= not w5291 and not w5669;
w5671 <= not w5667 and not w5670;
w5672 <= w460 and not w5652;
w5673 <= not w5662 and w5672;
w5674 <= not w5671 and not w5673;
w5675 <= not w5664 and not w5674;
w5676 <= not w356 and not w5675;
w5677 <= w5303 and not w5305;
w5678 <= not w5296 and w5677;
w5679 <= not w5418 and w5678;
w5680 <= not w5296 and not w5305;
w5681 <= not w5418 and w5680;
w5682 <= not w5303 and not w5681;
w5683 <= not w5679 and not w5682;
w5684 <= w356 and not w5664;
w5685 <= not w5674 and w5684;
w5686 <= not w5683 and not w5685;
w5687 <= not w5676 and not w5686;
w5688 <= not w264 and not w5687;
w5689 <= not w5308 and w5315;
w5690 <= not w5317 and w5689;
w5691 <= not w5418 and w5690;
w5692 <= not w5308 and not w5317;
w5693 <= not w5418 and w5692;
w5694 <= not w5315 and not w5693;
w5695 <= not w5691 and not w5694;
w5696 <= w264 and not w5676;
w5697 <= not w5686 and w5696;
w5698 <= not w5695 and not w5697;
w5699 <= not w5688 and not w5698;
w5700 <= not w184 and not w5699;
w5701 <= w5327 and not w5329;
w5702 <= not w5320 and w5701;
w5703 <= not w5418 and w5702;
w5704 <= not w5320 and not w5329;
w5705 <= not w5418 and w5704;
w5706 <= not w5327 and not w5705;
w5707 <= not w5703 and not w5706;
w5708 <= w184 and not w5688;
w5709 <= not w5698 and w5708;
w5710 <= not w5707 and not w5709;
w5711 <= not w5700 and not w5710;
w5712 <= not w115 and not w5711;
w5713 <= not w5332 and w5339;
w5714 <= not w5341 and w5713;
w5715 <= not w5418 and w5714;
w5716 <= not w5332 and not w5341;
w5717 <= not w5418 and w5716;
w5718 <= not w5339 and not w5717;
w5719 <= not w5715 and not w5718;
w5720 <= w115 and not w5700;
w5721 <= not w5710 and w5720;
w5722 <= not w5719 and not w5721;
w5723 <= not w5712 and not w5722;
w5724 <= not w60 and not w5723;
w5725 <= w5351 and not w5353;
w5726 <= not w5344 and w5725;
w5727 <= not w5418 and w5726;
w5728 <= not w5344 and not w5353;
w5729 <= not w5418 and w5728;
w5730 <= not w5351 and not w5729;
w5731 <= not w5727 and not w5730;
w5732 <= w60 and not w5712;
w5733 <= not w5722 and w5732;
w5734 <= not w5731 and not w5733;
w5735 <= not w5724 and not w5734;
w5736 <= not w22 and not w5735;
w5737 <= not w5356 and w5363;
w5738 <= not w5365 and w5737;
w5739 <= not w5418 and w5738;
w5740 <= not w5356 and not w5365;
w5741 <= not w5418 and w5740;
w5742 <= not w5363 and not w5741;
w5743 <= not w5739 and not w5742;
w5744 <= w22 and not w5724;
w5745 <= not w5734 and w5744;
w5746 <= not w5743 and not w5745;
w5747 <= not w5736 and not w5746;
w5748 <= not w5 and not w5747;
w5749 <= w5375 and not w5377;
w5750 <= not w5368 and w5749;
w5751 <= not w5418 and w5750;
w5752 <= not w5368 and not w5377;
w5753 <= not w5418 and w5752;
w5754 <= not w5375 and not w5753;
w5755 <= not w5751 and not w5754;
w5756 <= w5 and not w5736;
w5757 <= not w5746 and w5756;
w5758 <= not w5755 and not w5757;
w5759 <= not w5748 and not w5758;
w5760 <= not w5380 and w5389;
w5761 <= not w5382 and w5760;
w5762 <= not w5418 and w5761;
w5763 <= not w5380 and not w5382;
w5764 <= not w5418 and w5763;
w5765 <= not w5389 and not w5764;
w5766 <= not w5762 and not w5765;
w5767 <= not w5391 and not w5398;
w5768 <= not w5418 and w5767;
w5769 <= not w5406 and not w5768;
w5770 <= not w5766 and w5769;
w5771 <= not w5759 and w5770;
w5772 <= w0 and not w5771;
w5773 <= not w5748 and w5766;
w5774 <= not w5758 and w5773;
w5775 <= not w5398 and not w5418;
w5776 <= w5391 and not w5775;
w5777 <= not w0 and not w5767;
w5778 <= not w5776 and w5777;
w5779 <= not w5394 and not w5415;
w5780 <= not w5397 and w5779;
w5781 <= not w5410 and w5780;
w5782 <= not w5406 and w5781;
w5783 <= not w5404 and w5782;
w5784 <= not w5778 and not w5783;
w5785 <= not w5774 and w5784;
w5786 <= not w5772 and w5785;
w5787 <= a(66) and not w5786;
w5788 <= not a(64) and not a(65);
w5789 <= not a(66) and w5788;
w5790 <= not w5787 and not w5789;
w5791 <= not w5418 and not w5790;
w5792 <= not w5415 and not w5789;
w5793 <= not w5410 and w5792;
w5794 <= not w5406 and w5793;
w5795 <= not w5404 and w5794;
w5796 <= not w5787 and w5795;
w5797 <= not a(66) and not w5786;
w5798 <= a(67) and not w5797;
w5799 <= w5420 and not w5786;
w5800 <= not w5798 and not w5799;
w5801 <= not w5796 and w5800;
w5802 <= not w5791 and not w5801;
w5803 <= not w5062 and not w5802;
w5804 <= w5062 and not w5791;
w5805 <= not w5801 and w5804;
w5806 <= not w5418 and not w5783;
w5807 <= not w5778 and w5806;
w5808 <= not w5774 and w5807;
w5809 <= not w5772 and w5808;
w5810 <= not w5799 and not w5809;
w5811 <= a(68) and not w5810;
w5812 <= not a(68) and not w5809;
w5813 <= not w5799 and w5812;
w5814 <= not w5811 and not w5813;
w5815 <= not w5805 and not w5814;
w5816 <= not w5803 and not w5815;
w5817 <= not w4718 and not w5816;
w5818 <= not w5423 and not w5428;
w5819 <= not w5432 and w5818;
w5820 <= not w5786 and w5819;
w5821 <= not w5786 and w5818;
w5822 <= w5432 and not w5821;
w5823 <= not w5820 and not w5822;
w5824 <= w4718 and not w5803;
w5825 <= not w5815 and w5824;
w5826 <= not w5823 and not w5825;
w5827 <= not w5817 and not w5826;
w5828 <= not w4386 and not w5827;
w5829 <= not w5437 and w5446;
w5830 <= not w5435 and w5829;
w5831 <= not w5786 and w5830;
w5832 <= not w5435 and not w5437;
w5833 <= not w5786 and w5832;
w5834 <= not w5446 and not w5833;
w5835 <= not w5831 and not w5834;
w5836 <= w4386 and not w5817;
w5837 <= not w5826 and w5836;
w5838 <= not w5835 and not w5837;
w5839 <= not w5828 and not w5838;
w5840 <= not w4066 and not w5839;
w5841 <= not w5449 and w5455;
w5842 <= not w5457 and w5841;
w5843 <= not w5786 and w5842;
w5844 <= not w5449 and not w5457;
w5845 <= not w5786 and w5844;
w5846 <= not w5455 and not w5845;
w5847 <= not w5843 and not w5846;
w5848 <= w4066 and not w5828;
w5849 <= not w5838 and w5848;
w5850 <= not w5847 and not w5849;
w5851 <= not w5840 and not w5850;
w5852 <= not w3758 and not w5851;
w5853 <= w5467 and not w5469;
w5854 <= not w5460 and w5853;
w5855 <= not w5786 and w5854;
w5856 <= not w5460 and not w5469;
w5857 <= not w5786 and w5856;
w5858 <= not w5467 and not w5857;
w5859 <= not w5855 and not w5858;
w5860 <= w3758 and not w5840;
w5861 <= not w5850 and w5860;
w5862 <= not w5859 and not w5861;
w5863 <= not w5852 and not w5862;
w5864 <= not w3462 and not w5863;
w5865 <= not w5472 and w5479;
w5866 <= not w5481 and w5865;
w5867 <= not w5786 and w5866;
w5868 <= not w5472 and not w5481;
w5869 <= not w5786 and w5868;
w5870 <= not w5479 and not w5869;
w5871 <= not w5867 and not w5870;
w5872 <= w3462 and not w5852;
w5873 <= not w5862 and w5872;
w5874 <= not w5871 and not w5873;
w5875 <= not w5864 and not w5874;
w5876 <= not w3178 and not w5875;
w5877 <= w5491 and not w5493;
w5878 <= not w5484 and w5877;
w5879 <= not w5786 and w5878;
w5880 <= not w5484 and not w5493;
w5881 <= not w5786 and w5880;
w5882 <= not w5491 and not w5881;
w5883 <= not w5879 and not w5882;
w5884 <= w3178 and not w5864;
w5885 <= not w5874 and w5884;
w5886 <= not w5883 and not w5885;
w5887 <= not w5876 and not w5886;
w5888 <= not w2906 and not w5887;
w5889 <= not w5496 and w5503;
w5890 <= not w5505 and w5889;
w5891 <= not w5786 and w5890;
w5892 <= not w5496 and not w5505;
w5893 <= not w5786 and w5892;
w5894 <= not w5503 and not w5893;
w5895 <= not w5891 and not w5894;
w5896 <= w2906 and not w5876;
w5897 <= not w5886 and w5896;
w5898 <= not w5895 and not w5897;
w5899 <= not w5888 and not w5898;
w5900 <= not w2646 and not w5899;
w5901 <= w5515 and not w5517;
w5902 <= not w5508 and w5901;
w5903 <= not w5786 and w5902;
w5904 <= not w5508 and not w5517;
w5905 <= not w5786 and w5904;
w5906 <= not w5515 and not w5905;
w5907 <= not w5903 and not w5906;
w5908 <= w2646 and not w5888;
w5909 <= not w5898 and w5908;
w5910 <= not w5907 and not w5909;
w5911 <= not w5900 and not w5910;
w5912 <= not w2398 and not w5911;
w5913 <= not w5520 and w5527;
w5914 <= not w5529 and w5913;
w5915 <= not w5786 and w5914;
w5916 <= not w5520 and not w5529;
w5917 <= not w5786 and w5916;
w5918 <= not w5527 and not w5917;
w5919 <= not w5915 and not w5918;
w5920 <= w2398 and not w5900;
w5921 <= not w5910 and w5920;
w5922 <= not w5919 and not w5921;
w5923 <= not w5912 and not w5922;
w5924 <= not w2162 and not w5923;
w5925 <= w5539 and not w5541;
w5926 <= not w5532 and w5925;
w5927 <= not w5786 and w5926;
w5928 <= not w5532 and not w5541;
w5929 <= not w5786 and w5928;
w5930 <= not w5539 and not w5929;
w5931 <= not w5927 and not w5930;
w5932 <= w2162 and not w5912;
w5933 <= not w5922 and w5932;
w5934 <= not w5931 and not w5933;
w5935 <= not w5924 and not w5934;
w5936 <= not w1938 and not w5935;
w5937 <= not w5544 and w5551;
w5938 <= not w5553 and w5937;
w5939 <= not w5786 and w5938;
w5940 <= not w5544 and not w5553;
w5941 <= not w5786 and w5940;
w5942 <= not w5551 and not w5941;
w5943 <= not w5939 and not w5942;
w5944 <= w1938 and not w5924;
w5945 <= not w5934 and w5944;
w5946 <= not w5943 and not w5945;
w5947 <= not w5936 and not w5946;
w5948 <= not w1725 and not w5947;
w5949 <= w5563 and not w5565;
w5950 <= not w5556 and w5949;
w5951 <= not w5786 and w5950;
w5952 <= not w5556 and not w5565;
w5953 <= not w5786 and w5952;
w5954 <= not w5563 and not w5953;
w5955 <= not w5951 and not w5954;
w5956 <= w1725 and not w5936;
w5957 <= not w5946 and w5956;
w5958 <= not w5955 and not w5957;
w5959 <= not w5948 and not w5958;
w5960 <= not w1525 and not w5959;
w5961 <= not w5568 and w5575;
w5962 <= not w5577 and w5961;
w5963 <= not w5786 and w5962;
w5964 <= not w5568 and not w5577;
w5965 <= not w5786 and w5964;
w5966 <= not w5575 and not w5965;
w5967 <= not w5963 and not w5966;
w5968 <= w1525 and not w5948;
w5969 <= not w5958 and w5968;
w5970 <= not w5967 and not w5969;
w5971 <= not w5960 and not w5970;
w5972 <= not w1337 and not w5971;
w5973 <= w5587 and not w5589;
w5974 <= not w5580 and w5973;
w5975 <= not w5786 and w5974;
w5976 <= not w5580 and not w5589;
w5977 <= not w5786 and w5976;
w5978 <= not w5587 and not w5977;
w5979 <= not w5975 and not w5978;
w5980 <= w1337 and not w5960;
w5981 <= not w5970 and w5980;
w5982 <= not w5979 and not w5981;
w5983 <= not w5972 and not w5982;
w5984 <= not w1161 and not w5983;
w5985 <= not w5592 and w5599;
w5986 <= not w5601 and w5985;
w5987 <= not w5786 and w5986;
w5988 <= not w5592 and not w5601;
w5989 <= not w5786 and w5988;
w5990 <= not w5599 and not w5989;
w5991 <= not w5987 and not w5990;
w5992 <= w1161 and not w5972;
w5993 <= not w5982 and w5992;
w5994 <= not w5991 and not w5993;
w5995 <= not w5984 and not w5994;
w5996 <= not w997 and not w5995;
w5997 <= w5611 and not w5613;
w5998 <= not w5604 and w5997;
w5999 <= not w5786 and w5998;
w6000 <= not w5604 and not w5613;
w6001 <= not w5786 and w6000;
w6002 <= not w5611 and not w6001;
w6003 <= not w5999 and not w6002;
w6004 <= w997 and not w5984;
w6005 <= not w5994 and w6004;
w6006 <= not w6003 and not w6005;
w6007 <= not w5996 and not w6006;
w6008 <= not w845 and not w6007;
w6009 <= not w5616 and w5623;
w6010 <= not w5625 and w6009;
w6011 <= not w5786 and w6010;
w6012 <= not w5616 and not w5625;
w6013 <= not w5786 and w6012;
w6014 <= not w5623 and not w6013;
w6015 <= not w6011 and not w6014;
w6016 <= w845 and not w5996;
w6017 <= not w6006 and w6016;
w6018 <= not w6015 and not w6017;
w6019 <= not w6008 and not w6018;
w6020 <= not w705 and not w6019;
w6021 <= w5635 and not w5637;
w6022 <= not w5628 and w6021;
w6023 <= not w5786 and w6022;
w6024 <= not w5628 and not w5637;
w6025 <= not w5786 and w6024;
w6026 <= not w5635 and not w6025;
w6027 <= not w6023 and not w6026;
w6028 <= w705 and not w6008;
w6029 <= not w6018 and w6028;
w6030 <= not w6027 and not w6029;
w6031 <= not w6020 and not w6030;
w6032 <= not w577 and not w6031;
w6033 <= not w5640 and w5647;
w6034 <= not w5649 and w6033;
w6035 <= not w5786 and w6034;
w6036 <= not w5640 and not w5649;
w6037 <= not w5786 and w6036;
w6038 <= not w5647 and not w6037;
w6039 <= not w6035 and not w6038;
w6040 <= w577 and not w6020;
w6041 <= not w6030 and w6040;
w6042 <= not w6039 and not w6041;
w6043 <= not w6032 and not w6042;
w6044 <= not w460 and not w6043;
w6045 <= w5659 and not w5661;
w6046 <= not w5652 and w6045;
w6047 <= not w5786 and w6046;
w6048 <= not w5652 and not w5661;
w6049 <= not w5786 and w6048;
w6050 <= not w5659 and not w6049;
w6051 <= not w6047 and not w6050;
w6052 <= w460 and not w6032;
w6053 <= not w6042 and w6052;
w6054 <= not w6051 and not w6053;
w6055 <= not w6044 and not w6054;
w6056 <= not w356 and not w6055;
w6057 <= not w5664 and w5671;
w6058 <= not w5673 and w6057;
w6059 <= not w5786 and w6058;
w6060 <= not w5664 and not w5673;
w6061 <= not w5786 and w6060;
w6062 <= not w5671 and not w6061;
w6063 <= not w6059 and not w6062;
w6064 <= w356 and not w6044;
w6065 <= not w6054 and w6064;
w6066 <= not w6063 and not w6065;
w6067 <= not w6056 and not w6066;
w6068 <= not w264 and not w6067;
w6069 <= w5683 and not w5685;
w6070 <= not w5676 and w6069;
w6071 <= not w5786 and w6070;
w6072 <= not w5676 and not w5685;
w6073 <= not w5786 and w6072;
w6074 <= not w5683 and not w6073;
w6075 <= not w6071 and not w6074;
w6076 <= w264 and not w6056;
w6077 <= not w6066 and w6076;
w6078 <= not w6075 and not w6077;
w6079 <= not w6068 and not w6078;
w6080 <= not w184 and not w6079;
w6081 <= not w5688 and w5695;
w6082 <= not w5697 and w6081;
w6083 <= not w5786 and w6082;
w6084 <= not w5688 and not w5697;
w6085 <= not w5786 and w6084;
w6086 <= not w5695 and not w6085;
w6087 <= not w6083 and not w6086;
w6088 <= w184 and not w6068;
w6089 <= not w6078 and w6088;
w6090 <= not w6087 and not w6089;
w6091 <= not w6080 and not w6090;
w6092 <= not w115 and not w6091;
w6093 <= w5707 and not w5709;
w6094 <= not w5700 and w6093;
w6095 <= not w5786 and w6094;
w6096 <= not w5700 and not w5709;
w6097 <= not w5786 and w6096;
w6098 <= not w5707 and not w6097;
w6099 <= not w6095 and not w6098;
w6100 <= w115 and not w6080;
w6101 <= not w6090 and w6100;
w6102 <= not w6099 and not w6101;
w6103 <= not w6092 and not w6102;
w6104 <= not w60 and not w6103;
w6105 <= not w5712 and w5719;
w6106 <= not w5721 and w6105;
w6107 <= not w5786 and w6106;
w6108 <= not w5712 and not w5721;
w6109 <= not w5786 and w6108;
w6110 <= not w5719 and not w6109;
w6111 <= not w6107 and not w6110;
w6112 <= w60 and not w6092;
w6113 <= not w6102 and w6112;
w6114 <= not w6111 and not w6113;
w6115 <= not w6104 and not w6114;
w6116 <= not w22 and not w6115;
w6117 <= w5731 and not w5733;
w6118 <= not w5724 and w6117;
w6119 <= not w5786 and w6118;
w6120 <= not w5724 and not w5733;
w6121 <= not w5786 and w6120;
w6122 <= not w5731 and not w6121;
w6123 <= not w6119 and not w6122;
w6124 <= w22 and not w6104;
w6125 <= not w6114 and w6124;
w6126 <= not w6123 and not w6125;
w6127 <= not w6116 and not w6126;
w6128 <= not w5 and not w6127;
w6129 <= not w5736 and w5743;
w6130 <= not w5745 and w6129;
w6131 <= not w5786 and w6130;
w6132 <= not w5736 and not w5745;
w6133 <= not w5786 and w6132;
w6134 <= not w5743 and not w6133;
w6135 <= not w6131 and not w6134;
w6136 <= w5 and not w6116;
w6137 <= not w6126 and w6136;
w6138 <= not w6135 and not w6137;
w6139 <= not w6128 and not w6138;
w6140 <= w5755 and not w5757;
w6141 <= not w5748 and w6140;
w6142 <= not w5786 and w6141;
w6143 <= not w5748 and not w5757;
w6144 <= not w5786 and w6143;
w6145 <= not w5755 and not w6144;
w6146 <= not w6142 and not w6145;
w6147 <= not w5759 and not w5766;
w6148 <= not w5786 and w6147;
w6149 <= not w5774 and not w6148;
w6150 <= not w6146 and w6149;
w6151 <= not w6139 and w6150;
w6152 <= w0 and not w6151;
w6153 <= not w6128 and w6146;
w6154 <= not w6138 and w6153;
w6155 <= not w5766 and not w5786;
w6156 <= w5759 and not w6155;
w6157 <= not w0 and not w6147;
w6158 <= not w6156 and w6157;
w6159 <= not w5762 and not w5783;
w6160 <= not w5765 and w6159;
w6161 <= not w5778 and w6160;
w6162 <= not w5774 and w6161;
w6163 <= not w5772 and w6162;
w6164 <= not w6158 and not w6163;
w6165 <= not w6154 and w6164;
w6166 <= not w6152 and w6165;
w6167 <= a(64) and not w6166;
w6168 <= not a(62) and not a(63);
w6169 <= not a(64) and w6168;
w6170 <= not w6167 and not w6169;
w6171 <= not w5786 and not w6170;
w6172 <= not a(64) and not w6166;
w6173 <= a(65) and not w6172;
w6174 <= w5788 and not w6166;
w6175 <= not w6173 and not w6174;
w6176 <= not w5783 and not w6169;
w6177 <= not w5778 and w6176;
w6178 <= not w5774 and w6177;
w6179 <= not w5772 and w6178;
w6180 <= not w6167 and w6179;
w6181 <= w6175 and not w6180;
w6182 <= not w6171 and not w6181;
w6183 <= not w5418 and not w6182;
w6184 <= w5418 and not w6171;
w6185 <= not w6181 and w6184;
w6186 <= not w5786 and not w6163;
w6187 <= not w6158 and w6186;
w6188 <= not w6154 and w6187;
w6189 <= not w6152 and w6188;
w6190 <= not w6174 and not w6189;
w6191 <= a(66) and not w6190;
w6192 <= not a(66) and not w6189;
w6193 <= not w6174 and w6192;
w6194 <= not w6191 and not w6193;
w6195 <= not w6185 and not w6194;
w6196 <= not w6183 and not w6195;
w6197 <= not w5062 and not w6196;
w6198 <= not w5791 and not w5796;
w6199 <= not w5800 and w6198;
w6200 <= not w6166 and w6199;
w6201 <= not w6166 and w6198;
w6202 <= w5800 and not w6201;
w6203 <= not w6200 and not w6202;
w6204 <= w5062 and not w6183;
w6205 <= not w6195 and w6204;
w6206 <= not w6203 and not w6205;
w6207 <= not w6197 and not w6206;
w6208 <= not w4718 and not w6207;
w6209 <= not w5805 and w5814;
w6210 <= not w5803 and w6209;
w6211 <= not w6166 and w6210;
w6212 <= not w5803 and not w5805;
w6213 <= not w6166 and w6212;
w6214 <= not w5814 and not w6213;
w6215 <= not w6211 and not w6214;
w6216 <= w4718 and not w6197;
w6217 <= not w6206 and w6216;
w6218 <= not w6215 and not w6217;
w6219 <= not w6208 and not w6218;
w6220 <= not w4386 and not w6219;
w6221 <= not w5817 and w5823;
w6222 <= not w5825 and w6221;
w6223 <= not w6166 and w6222;
w6224 <= not w5817 and not w5825;
w6225 <= not w6166 and w6224;
w6226 <= not w5823 and not w6225;
w6227 <= not w6223 and not w6226;
w6228 <= w4386 and not w6208;
w6229 <= not w6218 and w6228;
w6230 <= not w6227 and not w6229;
w6231 <= not w6220 and not w6230;
w6232 <= not w4066 and not w6231;
w6233 <= w5835 and not w5837;
w6234 <= not w5828 and w6233;
w6235 <= not w6166 and w6234;
w6236 <= not w5828 and not w5837;
w6237 <= not w6166 and w6236;
w6238 <= not w5835 and not w6237;
w6239 <= not w6235 and not w6238;
w6240 <= w4066 and not w6220;
w6241 <= not w6230 and w6240;
w6242 <= not w6239 and not w6241;
w6243 <= not w6232 and not w6242;
w6244 <= not w3758 and not w6243;
w6245 <= not w5840 and w5847;
w6246 <= not w5849 and w6245;
w6247 <= not w6166 and w6246;
w6248 <= not w5840 and not w5849;
w6249 <= not w6166 and w6248;
w6250 <= not w5847 and not w6249;
w6251 <= not w6247 and not w6250;
w6252 <= w3758 and not w6232;
w6253 <= not w6242 and w6252;
w6254 <= not w6251 and not w6253;
w6255 <= not w6244 and not w6254;
w6256 <= not w3462 and not w6255;
w6257 <= w5859 and not w5861;
w6258 <= not w5852 and w6257;
w6259 <= not w6166 and w6258;
w6260 <= not w5852 and not w5861;
w6261 <= not w6166 and w6260;
w6262 <= not w5859 and not w6261;
w6263 <= not w6259 and not w6262;
w6264 <= w3462 and not w6244;
w6265 <= not w6254 and w6264;
w6266 <= not w6263 and not w6265;
w6267 <= not w6256 and not w6266;
w6268 <= not w3178 and not w6267;
w6269 <= not w5864 and w5871;
w6270 <= not w5873 and w6269;
w6271 <= not w6166 and w6270;
w6272 <= not w5864 and not w5873;
w6273 <= not w6166 and w6272;
w6274 <= not w5871 and not w6273;
w6275 <= not w6271 and not w6274;
w6276 <= w3178 and not w6256;
w6277 <= not w6266 and w6276;
w6278 <= not w6275 and not w6277;
w6279 <= not w6268 and not w6278;
w6280 <= not w2906 and not w6279;
w6281 <= w5883 and not w5885;
w6282 <= not w5876 and w6281;
w6283 <= not w6166 and w6282;
w6284 <= not w5876 and not w5885;
w6285 <= not w6166 and w6284;
w6286 <= not w5883 and not w6285;
w6287 <= not w6283 and not w6286;
w6288 <= w2906 and not w6268;
w6289 <= not w6278 and w6288;
w6290 <= not w6287 and not w6289;
w6291 <= not w6280 and not w6290;
w6292 <= not w2646 and not w6291;
w6293 <= not w5888 and w5895;
w6294 <= not w5897 and w6293;
w6295 <= not w6166 and w6294;
w6296 <= not w5888 and not w5897;
w6297 <= not w6166 and w6296;
w6298 <= not w5895 and not w6297;
w6299 <= not w6295 and not w6298;
w6300 <= w2646 and not w6280;
w6301 <= not w6290 and w6300;
w6302 <= not w6299 and not w6301;
w6303 <= not w6292 and not w6302;
w6304 <= not w2398 and not w6303;
w6305 <= w5907 and not w5909;
w6306 <= not w5900 and w6305;
w6307 <= not w6166 and w6306;
w6308 <= not w5900 and not w5909;
w6309 <= not w6166 and w6308;
w6310 <= not w5907 and not w6309;
w6311 <= not w6307 and not w6310;
w6312 <= w2398 and not w6292;
w6313 <= not w6302 and w6312;
w6314 <= not w6311 and not w6313;
w6315 <= not w6304 and not w6314;
w6316 <= not w2162 and not w6315;
w6317 <= not w5912 and w5919;
w6318 <= not w5921 and w6317;
w6319 <= not w6166 and w6318;
w6320 <= not w5912 and not w5921;
w6321 <= not w6166 and w6320;
w6322 <= not w5919 and not w6321;
w6323 <= not w6319 and not w6322;
w6324 <= w2162 and not w6304;
w6325 <= not w6314 and w6324;
w6326 <= not w6323 and not w6325;
w6327 <= not w6316 and not w6326;
w6328 <= not w1938 and not w6327;
w6329 <= w5931 and not w5933;
w6330 <= not w5924 and w6329;
w6331 <= not w6166 and w6330;
w6332 <= not w5924 and not w5933;
w6333 <= not w6166 and w6332;
w6334 <= not w5931 and not w6333;
w6335 <= not w6331 and not w6334;
w6336 <= w1938 and not w6316;
w6337 <= not w6326 and w6336;
w6338 <= not w6335 and not w6337;
w6339 <= not w6328 and not w6338;
w6340 <= not w1725 and not w6339;
w6341 <= not w5936 and w5943;
w6342 <= not w5945 and w6341;
w6343 <= not w6166 and w6342;
w6344 <= not w5936 and not w5945;
w6345 <= not w6166 and w6344;
w6346 <= not w5943 and not w6345;
w6347 <= not w6343 and not w6346;
w6348 <= w1725 and not w6328;
w6349 <= not w6338 and w6348;
w6350 <= not w6347 and not w6349;
w6351 <= not w6340 and not w6350;
w6352 <= not w1525 and not w6351;
w6353 <= w5955 and not w5957;
w6354 <= not w5948 and w6353;
w6355 <= not w6166 and w6354;
w6356 <= not w5948 and not w5957;
w6357 <= not w6166 and w6356;
w6358 <= not w5955 and not w6357;
w6359 <= not w6355 and not w6358;
w6360 <= w1525 and not w6340;
w6361 <= not w6350 and w6360;
w6362 <= not w6359 and not w6361;
w6363 <= not w6352 and not w6362;
w6364 <= not w1337 and not w6363;
w6365 <= not w5960 and w5967;
w6366 <= not w5969 and w6365;
w6367 <= not w6166 and w6366;
w6368 <= not w5960 and not w5969;
w6369 <= not w6166 and w6368;
w6370 <= not w5967 and not w6369;
w6371 <= not w6367 and not w6370;
w6372 <= w1337 and not w6352;
w6373 <= not w6362 and w6372;
w6374 <= not w6371 and not w6373;
w6375 <= not w6364 and not w6374;
w6376 <= not w1161 and not w6375;
w6377 <= w5979 and not w5981;
w6378 <= not w5972 and w6377;
w6379 <= not w6166 and w6378;
w6380 <= not w5972 and not w5981;
w6381 <= not w6166 and w6380;
w6382 <= not w5979 and not w6381;
w6383 <= not w6379 and not w6382;
w6384 <= w1161 and not w6364;
w6385 <= not w6374 and w6384;
w6386 <= not w6383 and not w6385;
w6387 <= not w6376 and not w6386;
w6388 <= not w997 and not w6387;
w6389 <= not w5984 and w5991;
w6390 <= not w5993 and w6389;
w6391 <= not w6166 and w6390;
w6392 <= not w5984 and not w5993;
w6393 <= not w6166 and w6392;
w6394 <= not w5991 and not w6393;
w6395 <= not w6391 and not w6394;
w6396 <= w997 and not w6376;
w6397 <= not w6386 and w6396;
w6398 <= not w6395 and not w6397;
w6399 <= not w6388 and not w6398;
w6400 <= not w845 and not w6399;
w6401 <= w6003 and not w6005;
w6402 <= not w5996 and w6401;
w6403 <= not w6166 and w6402;
w6404 <= not w5996 and not w6005;
w6405 <= not w6166 and w6404;
w6406 <= not w6003 and not w6405;
w6407 <= not w6403 and not w6406;
w6408 <= w845 and not w6388;
w6409 <= not w6398 and w6408;
w6410 <= not w6407 and not w6409;
w6411 <= not w6400 and not w6410;
w6412 <= not w705 and not w6411;
w6413 <= not w6008 and w6015;
w6414 <= not w6017 and w6413;
w6415 <= not w6166 and w6414;
w6416 <= not w6008 and not w6017;
w6417 <= not w6166 and w6416;
w6418 <= not w6015 and not w6417;
w6419 <= not w6415 and not w6418;
w6420 <= w705 and not w6400;
w6421 <= not w6410 and w6420;
w6422 <= not w6419 and not w6421;
w6423 <= not w6412 and not w6422;
w6424 <= not w577 and not w6423;
w6425 <= w6027 and not w6029;
w6426 <= not w6020 and w6425;
w6427 <= not w6166 and w6426;
w6428 <= not w6020 and not w6029;
w6429 <= not w6166 and w6428;
w6430 <= not w6027 and not w6429;
w6431 <= not w6427 and not w6430;
w6432 <= w577 and not w6412;
w6433 <= not w6422 and w6432;
w6434 <= not w6431 and not w6433;
w6435 <= not w6424 and not w6434;
w6436 <= not w460 and not w6435;
w6437 <= not w6032 and w6039;
w6438 <= not w6041 and w6437;
w6439 <= not w6166 and w6438;
w6440 <= not w6032 and not w6041;
w6441 <= not w6166 and w6440;
w6442 <= not w6039 and not w6441;
w6443 <= not w6439 and not w6442;
w6444 <= w460 and not w6424;
w6445 <= not w6434 and w6444;
w6446 <= not w6443 and not w6445;
w6447 <= not w6436 and not w6446;
w6448 <= not w356 and not w6447;
w6449 <= w6051 and not w6053;
w6450 <= not w6044 and w6449;
w6451 <= not w6166 and w6450;
w6452 <= not w6044 and not w6053;
w6453 <= not w6166 and w6452;
w6454 <= not w6051 and not w6453;
w6455 <= not w6451 and not w6454;
w6456 <= w356 and not w6436;
w6457 <= not w6446 and w6456;
w6458 <= not w6455 and not w6457;
w6459 <= not w6448 and not w6458;
w6460 <= not w264 and not w6459;
w6461 <= not w6056 and w6063;
w6462 <= not w6065 and w6461;
w6463 <= not w6166 and w6462;
w6464 <= not w6056 and not w6065;
w6465 <= not w6166 and w6464;
w6466 <= not w6063 and not w6465;
w6467 <= not w6463 and not w6466;
w6468 <= w264 and not w6448;
w6469 <= not w6458 and w6468;
w6470 <= not w6467 and not w6469;
w6471 <= not w6460 and not w6470;
w6472 <= not w184 and not w6471;
w6473 <= w6075 and not w6077;
w6474 <= not w6068 and w6473;
w6475 <= not w6166 and w6474;
w6476 <= not w6068 and not w6077;
w6477 <= not w6166 and w6476;
w6478 <= not w6075 and not w6477;
w6479 <= not w6475 and not w6478;
w6480 <= w184 and not w6460;
w6481 <= not w6470 and w6480;
w6482 <= not w6479 and not w6481;
w6483 <= not w6472 and not w6482;
w6484 <= not w115 and not w6483;
w6485 <= not w6080 and w6087;
w6486 <= not w6089 and w6485;
w6487 <= not w6166 and w6486;
w6488 <= not w6080 and not w6089;
w6489 <= not w6166 and w6488;
w6490 <= not w6087 and not w6489;
w6491 <= not w6487 and not w6490;
w6492 <= w115 and not w6472;
w6493 <= not w6482 and w6492;
w6494 <= not w6491 and not w6493;
w6495 <= not w6484 and not w6494;
w6496 <= not w60 and not w6495;
w6497 <= w6099 and not w6101;
w6498 <= not w6092 and w6497;
w6499 <= not w6166 and w6498;
w6500 <= not w6092 and not w6101;
w6501 <= not w6166 and w6500;
w6502 <= not w6099 and not w6501;
w6503 <= not w6499 and not w6502;
w6504 <= w60 and not w6484;
w6505 <= not w6494 and w6504;
w6506 <= not w6503 and not w6505;
w6507 <= not w6496 and not w6506;
w6508 <= not w22 and not w6507;
w6509 <= not w6104 and w6111;
w6510 <= not w6113 and w6509;
w6511 <= not w6166 and w6510;
w6512 <= not w6104 and not w6113;
w6513 <= not w6166 and w6512;
w6514 <= not w6111 and not w6513;
w6515 <= not w6511 and not w6514;
w6516 <= w22 and not w6496;
w6517 <= not w6506 and w6516;
w6518 <= not w6515 and not w6517;
w6519 <= not w6508 and not w6518;
w6520 <= not w5 and not w6519;
w6521 <= w6123 and not w6125;
w6522 <= not w6116 and w6521;
w6523 <= not w6166 and w6522;
w6524 <= not w6116 and not w6125;
w6525 <= not w6166 and w6524;
w6526 <= not w6123 and not w6525;
w6527 <= not w6523 and not w6526;
w6528 <= w5 and not w6508;
w6529 <= not w6518 and w6528;
w6530 <= not w6527 and not w6529;
w6531 <= not w6520 and not w6530;
w6532 <= not w6128 and w6135;
w6533 <= not w6137 and w6532;
w6534 <= not w6166 and w6533;
w6535 <= not w6128 and not w6137;
w6536 <= not w6166 and w6535;
w6537 <= not w6135 and not w6536;
w6538 <= not w6534 and not w6537;
w6539 <= not w6139 and not w6146;
w6540 <= not w6166 and w6539;
w6541 <= not w6154 and not w6540;
w6542 <= not w6538 and w6541;
w6543 <= not w6531 and w6542;
w6544 <= w0 and not w6543;
w6545 <= not w6520 and w6538;
w6546 <= not w6530 and w6545;
w6547 <= not w6146 and not w6166;
w6548 <= w6139 and not w6547;
w6549 <= not w0 and not w6539;
w6550 <= not w6548 and w6549;
w6551 <= not w6142 and not w6163;
w6552 <= not w6145 and w6551;
w6553 <= not w6158 and w6552;
w6554 <= not w6154 and w6553;
w6555 <= not w6152 and w6554;
w6556 <= not w6550 and not w6555;
w6557 <= not w6546 and w6556;
w6558 <= not w6544 and w6557;
w6559 <= a(62) and not w6558;
w6560 <= not a(60) and not a(61);
w6561 <= not a(62) and w6560;
w6562 <= not w6559 and not w6561;
w6563 <= not w6166 and not w6562;
w6564 <= not w6163 and not w6561;
w6565 <= not w6158 and w6564;
w6566 <= not w6154 and w6565;
w6567 <= not w6152 and w6566;
w6568 <= not w6559 and w6567;
w6569 <= not a(62) and not w6558;
w6570 <= a(63) and not w6569;
w6571 <= w6168 and not w6558;
w6572 <= not w6570 and not w6571;
w6573 <= not w6568 and w6572;
w6574 <= not w6563 and not w6573;
w6575 <= not w5786 and not w6574;
w6576 <= w5786 and not w6563;
w6577 <= not w6573 and w6576;
w6578 <= not w6166 and not w6555;
w6579 <= not w6550 and w6578;
w6580 <= not w6546 and w6579;
w6581 <= not w6544 and w6580;
w6582 <= not w6571 and not w6581;
w6583 <= a(64) and not w6582;
w6584 <= not a(64) and not w6581;
w6585 <= not w6571 and w6584;
w6586 <= not w6583 and not w6585;
w6587 <= not w6577 and not w6586;
w6588 <= not w6575 and not w6587;
w6589 <= not w5418 and not w6588;
w6590 <= w5418 and not w6575;
w6591 <= not w6587 and w6590;
w6592 <= not w6175 and not w6180;
w6593 <= not w6171 and w6592;
w6594 <= not w6558 and w6593;
w6595 <= not w6171 and not w6180;
w6596 <= not w6558 and w6595;
w6597 <= w6175 and not w6596;
w6598 <= not w6594 and not w6597;
w6599 <= not w6591 and not w6598;
w6600 <= not w6589 and not w6599;
w6601 <= not w5062 and not w6600;
w6602 <= not w6185 and w6194;
w6603 <= not w6183 and w6602;
w6604 <= not w6558 and w6603;
w6605 <= not w6183 and not w6185;
w6606 <= not w6558 and w6605;
w6607 <= not w6194 and not w6606;
w6608 <= not w6604 and not w6607;
w6609 <= w5062 and not w6589;
w6610 <= not w6599 and w6609;
w6611 <= not w6608 and not w6610;
w6612 <= not w6601 and not w6611;
w6613 <= not w4718 and not w6612;
w6614 <= not w6197 and w6203;
w6615 <= not w6205 and w6614;
w6616 <= not w6558 and w6615;
w6617 <= not w6197 and not w6205;
w6618 <= not w6558 and w6617;
w6619 <= not w6203 and not w6618;
w6620 <= not w6616 and not w6619;
w6621 <= w4718 and not w6601;
w6622 <= not w6611 and w6621;
w6623 <= not w6620 and not w6622;
w6624 <= not w6613 and not w6623;
w6625 <= not w4386 and not w6624;
w6626 <= w6215 and not w6217;
w6627 <= not w6208 and w6626;
w6628 <= not w6558 and w6627;
w6629 <= not w6208 and not w6217;
w6630 <= not w6558 and w6629;
w6631 <= not w6215 and not w6630;
w6632 <= not w6628 and not w6631;
w6633 <= w4386 and not w6613;
w6634 <= not w6623 and w6633;
w6635 <= not w6632 and not w6634;
w6636 <= not w6625 and not w6635;
w6637 <= not w4066 and not w6636;
w6638 <= not w6220 and w6227;
w6639 <= not w6229 and w6638;
w6640 <= not w6558 and w6639;
w6641 <= not w6220 and not w6229;
w6642 <= not w6558 and w6641;
w6643 <= not w6227 and not w6642;
w6644 <= not w6640 and not w6643;
w6645 <= w4066 and not w6625;
w6646 <= not w6635 and w6645;
w6647 <= not w6644 and not w6646;
w6648 <= not w6637 and not w6647;
w6649 <= not w3758 and not w6648;
w6650 <= w6239 and not w6241;
w6651 <= not w6232 and w6650;
w6652 <= not w6558 and w6651;
w6653 <= not w6232 and not w6241;
w6654 <= not w6558 and w6653;
w6655 <= not w6239 and not w6654;
w6656 <= not w6652 and not w6655;
w6657 <= w3758 and not w6637;
w6658 <= not w6647 and w6657;
w6659 <= not w6656 and not w6658;
w6660 <= not w6649 and not w6659;
w6661 <= not w3462 and not w6660;
w6662 <= not w6244 and w6251;
w6663 <= not w6253 and w6662;
w6664 <= not w6558 and w6663;
w6665 <= not w6244 and not w6253;
w6666 <= not w6558 and w6665;
w6667 <= not w6251 and not w6666;
w6668 <= not w6664 and not w6667;
w6669 <= w3462 and not w6649;
w6670 <= not w6659 and w6669;
w6671 <= not w6668 and not w6670;
w6672 <= not w6661 and not w6671;
w6673 <= not w3178 and not w6672;
w6674 <= w6263 and not w6265;
w6675 <= not w6256 and w6674;
w6676 <= not w6558 and w6675;
w6677 <= not w6256 and not w6265;
w6678 <= not w6558 and w6677;
w6679 <= not w6263 and not w6678;
w6680 <= not w6676 and not w6679;
w6681 <= w3178 and not w6661;
w6682 <= not w6671 and w6681;
w6683 <= not w6680 and not w6682;
w6684 <= not w6673 and not w6683;
w6685 <= not w2906 and not w6684;
w6686 <= not w6268 and w6275;
w6687 <= not w6277 and w6686;
w6688 <= not w6558 and w6687;
w6689 <= not w6268 and not w6277;
w6690 <= not w6558 and w6689;
w6691 <= not w6275 and not w6690;
w6692 <= not w6688 and not w6691;
w6693 <= w2906 and not w6673;
w6694 <= not w6683 and w6693;
w6695 <= not w6692 and not w6694;
w6696 <= not w6685 and not w6695;
w6697 <= not w2646 and not w6696;
w6698 <= w6287 and not w6289;
w6699 <= not w6280 and w6698;
w6700 <= not w6558 and w6699;
w6701 <= not w6280 and not w6289;
w6702 <= not w6558 and w6701;
w6703 <= not w6287 and not w6702;
w6704 <= not w6700 and not w6703;
w6705 <= w2646 and not w6685;
w6706 <= not w6695 and w6705;
w6707 <= not w6704 and not w6706;
w6708 <= not w6697 and not w6707;
w6709 <= not w2398 and not w6708;
w6710 <= not w6292 and w6299;
w6711 <= not w6301 and w6710;
w6712 <= not w6558 and w6711;
w6713 <= not w6292 and not w6301;
w6714 <= not w6558 and w6713;
w6715 <= not w6299 and not w6714;
w6716 <= not w6712 and not w6715;
w6717 <= w2398 and not w6697;
w6718 <= not w6707 and w6717;
w6719 <= not w6716 and not w6718;
w6720 <= not w6709 and not w6719;
w6721 <= not w2162 and not w6720;
w6722 <= w6311 and not w6313;
w6723 <= not w6304 and w6722;
w6724 <= not w6558 and w6723;
w6725 <= not w6304 and not w6313;
w6726 <= not w6558 and w6725;
w6727 <= not w6311 and not w6726;
w6728 <= not w6724 and not w6727;
w6729 <= w2162 and not w6709;
w6730 <= not w6719 and w6729;
w6731 <= not w6728 and not w6730;
w6732 <= not w6721 and not w6731;
w6733 <= not w1938 and not w6732;
w6734 <= not w6316 and w6323;
w6735 <= not w6325 and w6734;
w6736 <= not w6558 and w6735;
w6737 <= not w6316 and not w6325;
w6738 <= not w6558 and w6737;
w6739 <= not w6323 and not w6738;
w6740 <= not w6736 and not w6739;
w6741 <= w1938 and not w6721;
w6742 <= not w6731 and w6741;
w6743 <= not w6740 and not w6742;
w6744 <= not w6733 and not w6743;
w6745 <= not w1725 and not w6744;
w6746 <= w6335 and not w6337;
w6747 <= not w6328 and w6746;
w6748 <= not w6558 and w6747;
w6749 <= not w6328 and not w6337;
w6750 <= not w6558 and w6749;
w6751 <= not w6335 and not w6750;
w6752 <= not w6748 and not w6751;
w6753 <= w1725 and not w6733;
w6754 <= not w6743 and w6753;
w6755 <= not w6752 and not w6754;
w6756 <= not w6745 and not w6755;
w6757 <= not w1525 and not w6756;
w6758 <= not w6340 and w6347;
w6759 <= not w6349 and w6758;
w6760 <= not w6558 and w6759;
w6761 <= not w6340 and not w6349;
w6762 <= not w6558 and w6761;
w6763 <= not w6347 and not w6762;
w6764 <= not w6760 and not w6763;
w6765 <= w1525 and not w6745;
w6766 <= not w6755 and w6765;
w6767 <= not w6764 and not w6766;
w6768 <= not w6757 and not w6767;
w6769 <= not w1337 and not w6768;
w6770 <= w6359 and not w6361;
w6771 <= not w6352 and w6770;
w6772 <= not w6558 and w6771;
w6773 <= not w6352 and not w6361;
w6774 <= not w6558 and w6773;
w6775 <= not w6359 and not w6774;
w6776 <= not w6772 and not w6775;
w6777 <= w1337 and not w6757;
w6778 <= not w6767 and w6777;
w6779 <= not w6776 and not w6778;
w6780 <= not w6769 and not w6779;
w6781 <= not w1161 and not w6780;
w6782 <= not w6364 and w6371;
w6783 <= not w6373 and w6782;
w6784 <= not w6558 and w6783;
w6785 <= not w6364 and not w6373;
w6786 <= not w6558 and w6785;
w6787 <= not w6371 and not w6786;
w6788 <= not w6784 and not w6787;
w6789 <= w1161 and not w6769;
w6790 <= not w6779 and w6789;
w6791 <= not w6788 and not w6790;
w6792 <= not w6781 and not w6791;
w6793 <= not w997 and not w6792;
w6794 <= w6383 and not w6385;
w6795 <= not w6376 and w6794;
w6796 <= not w6558 and w6795;
w6797 <= not w6376 and not w6385;
w6798 <= not w6558 and w6797;
w6799 <= not w6383 and not w6798;
w6800 <= not w6796 and not w6799;
w6801 <= w997 and not w6781;
w6802 <= not w6791 and w6801;
w6803 <= not w6800 and not w6802;
w6804 <= not w6793 and not w6803;
w6805 <= not w845 and not w6804;
w6806 <= not w6388 and w6395;
w6807 <= not w6397 and w6806;
w6808 <= not w6558 and w6807;
w6809 <= not w6388 and not w6397;
w6810 <= not w6558 and w6809;
w6811 <= not w6395 and not w6810;
w6812 <= not w6808 and not w6811;
w6813 <= w845 and not w6793;
w6814 <= not w6803 and w6813;
w6815 <= not w6812 and not w6814;
w6816 <= not w6805 and not w6815;
w6817 <= not w705 and not w6816;
w6818 <= w6407 and not w6409;
w6819 <= not w6400 and w6818;
w6820 <= not w6558 and w6819;
w6821 <= not w6400 and not w6409;
w6822 <= not w6558 and w6821;
w6823 <= not w6407 and not w6822;
w6824 <= not w6820 and not w6823;
w6825 <= w705 and not w6805;
w6826 <= not w6815 and w6825;
w6827 <= not w6824 and not w6826;
w6828 <= not w6817 and not w6827;
w6829 <= not w577 and not w6828;
w6830 <= not w6412 and w6419;
w6831 <= not w6421 and w6830;
w6832 <= not w6558 and w6831;
w6833 <= not w6412 and not w6421;
w6834 <= not w6558 and w6833;
w6835 <= not w6419 and not w6834;
w6836 <= not w6832 and not w6835;
w6837 <= w577 and not w6817;
w6838 <= not w6827 and w6837;
w6839 <= not w6836 and not w6838;
w6840 <= not w6829 and not w6839;
w6841 <= not w460 and not w6840;
w6842 <= w6431 and not w6433;
w6843 <= not w6424 and w6842;
w6844 <= not w6558 and w6843;
w6845 <= not w6424 and not w6433;
w6846 <= not w6558 and w6845;
w6847 <= not w6431 and not w6846;
w6848 <= not w6844 and not w6847;
w6849 <= w460 and not w6829;
w6850 <= not w6839 and w6849;
w6851 <= not w6848 and not w6850;
w6852 <= not w6841 and not w6851;
w6853 <= not w356 and not w6852;
w6854 <= not w6436 and w6443;
w6855 <= not w6445 and w6854;
w6856 <= not w6558 and w6855;
w6857 <= not w6436 and not w6445;
w6858 <= not w6558 and w6857;
w6859 <= not w6443 and not w6858;
w6860 <= not w6856 and not w6859;
w6861 <= w356 and not w6841;
w6862 <= not w6851 and w6861;
w6863 <= not w6860 and not w6862;
w6864 <= not w6853 and not w6863;
w6865 <= not w264 and not w6864;
w6866 <= w6455 and not w6457;
w6867 <= not w6448 and w6866;
w6868 <= not w6558 and w6867;
w6869 <= not w6448 and not w6457;
w6870 <= not w6558 and w6869;
w6871 <= not w6455 and not w6870;
w6872 <= not w6868 and not w6871;
w6873 <= w264 and not w6853;
w6874 <= not w6863 and w6873;
w6875 <= not w6872 and not w6874;
w6876 <= not w6865 and not w6875;
w6877 <= not w184 and not w6876;
w6878 <= not w6460 and w6467;
w6879 <= not w6469 and w6878;
w6880 <= not w6558 and w6879;
w6881 <= not w6460 and not w6469;
w6882 <= not w6558 and w6881;
w6883 <= not w6467 and not w6882;
w6884 <= not w6880 and not w6883;
w6885 <= w184 and not w6865;
w6886 <= not w6875 and w6885;
w6887 <= not w6884 and not w6886;
w6888 <= not w6877 and not w6887;
w6889 <= not w115 and not w6888;
w6890 <= w6479 and not w6481;
w6891 <= not w6472 and w6890;
w6892 <= not w6558 and w6891;
w6893 <= not w6472 and not w6481;
w6894 <= not w6558 and w6893;
w6895 <= not w6479 and not w6894;
w6896 <= not w6892 and not w6895;
w6897 <= w115 and not w6877;
w6898 <= not w6887 and w6897;
w6899 <= not w6896 and not w6898;
w6900 <= not w6889 and not w6899;
w6901 <= not w60 and not w6900;
w6902 <= not w6484 and w6491;
w6903 <= not w6493 and w6902;
w6904 <= not w6558 and w6903;
w6905 <= not w6484 and not w6493;
w6906 <= not w6558 and w6905;
w6907 <= not w6491 and not w6906;
w6908 <= not w6904 and not w6907;
w6909 <= w60 and not w6889;
w6910 <= not w6899 and w6909;
w6911 <= not w6908 and not w6910;
w6912 <= not w6901 and not w6911;
w6913 <= not w22 and not w6912;
w6914 <= w6503 and not w6505;
w6915 <= not w6496 and w6914;
w6916 <= not w6558 and w6915;
w6917 <= not w6496 and not w6505;
w6918 <= not w6558 and w6917;
w6919 <= not w6503 and not w6918;
w6920 <= not w6916 and not w6919;
w6921 <= w22 and not w6901;
w6922 <= not w6911 and w6921;
w6923 <= not w6920 and not w6922;
w6924 <= not w6913 and not w6923;
w6925 <= not w5 and not w6924;
w6926 <= not w6508 and w6515;
w6927 <= not w6517 and w6926;
w6928 <= not w6558 and w6927;
w6929 <= not w6508 and not w6517;
w6930 <= not w6558 and w6929;
w6931 <= not w6515 and not w6930;
w6932 <= not w6928 and not w6931;
w6933 <= w5 and not w6913;
w6934 <= not w6923 and w6933;
w6935 <= not w6932 and not w6934;
w6936 <= not w6925 and not w6935;
w6937 <= w6527 and not w6529;
w6938 <= not w6520 and w6937;
w6939 <= not w6558 and w6938;
w6940 <= not w6520 and not w6529;
w6941 <= not w6558 and w6940;
w6942 <= not w6527 and not w6941;
w6943 <= not w6939 and not w6942;
w6944 <= not w6531 and not w6538;
w6945 <= not w6558 and w6944;
w6946 <= not w6546 and not w6945;
w6947 <= not w6943 and w6946;
w6948 <= not w6936 and w6947;
w6949 <= w0 and not w6948;
w6950 <= not w6925 and w6943;
w6951 <= not w6935 and w6950;
w6952 <= not w6538 and not w6558;
w6953 <= w6531 and not w6952;
w6954 <= not w0 and not w6944;
w6955 <= not w6953 and w6954;
w6956 <= not w6534 and not w6555;
w6957 <= not w6537 and w6956;
w6958 <= not w6550 and w6957;
w6959 <= not w6546 and w6958;
w6960 <= not w6544 and w6959;
w6961 <= not w6955 and not w6960;
w6962 <= not w6951 and w6961;
w6963 <= not w6949 and w6962;
w6964 <= a(60) and not w6963;
w6965 <= not a(58) and not a(59);
w6966 <= not a(60) and w6965;
w6967 <= not w6964 and not w6966;
w6968 <= not w6558 and not w6967;
w6969 <= not w6555 and not w6966;
w6970 <= not w6550 and w6969;
w6971 <= not w6546 and w6970;
w6972 <= not w6544 and w6971;
w6973 <= not w6964 and w6972;
w6974 <= not a(60) and not w6963;
w6975 <= a(61) and not w6974;
w6976 <= w6560 and not w6963;
w6977 <= not w6975 and not w6976;
w6978 <= not w6973 and w6977;
w6979 <= not w6968 and not w6978;
w6980 <= not w6166 and not w6979;
w6981 <= w6166 and not w6968;
w6982 <= not w6978 and w6981;
w6983 <= not w6558 and not w6960;
w6984 <= not w6955 and w6983;
w6985 <= not w6951 and w6984;
w6986 <= not w6949 and w6985;
w6987 <= not w6976 and not w6986;
w6988 <= a(62) and not w6987;
w6989 <= not a(62) and not w6986;
w6990 <= not w6976 and w6989;
w6991 <= not w6988 and not w6990;
w6992 <= not w6982 and not w6991;
w6993 <= not w6980 and not w6992;
w6994 <= not w5786 and not w6993;
w6995 <= not w6563 and not w6568;
w6996 <= not w6572 and w6995;
w6997 <= not w6963 and w6996;
w6998 <= not w6963 and w6995;
w6999 <= w6572 and not w6998;
w7000 <= not w6997 and not w6999;
w7001 <= w5786 and not w6980;
w7002 <= not w6992 and w7001;
w7003 <= not w7000 and not w7002;
w7004 <= not w6994 and not w7003;
w7005 <= not w5418 and not w7004;
w7006 <= not w6577 and w6586;
w7007 <= not w6575 and w7006;
w7008 <= not w6963 and w7007;
w7009 <= not w6575 and not w6577;
w7010 <= not w6963 and w7009;
w7011 <= not w6586 and not w7010;
w7012 <= not w7008 and not w7011;
w7013 <= w5418 and not w6994;
w7014 <= not w7003 and w7013;
w7015 <= not w7012 and not w7014;
w7016 <= not w7005 and not w7015;
w7017 <= not w5062 and not w7016;
w7018 <= w5062 and not w7005;
w7019 <= not w7015 and w7018;
w7020 <= not w6589 and w6598;
w7021 <= not w6591 and w7020;
w7022 <= not w6963 and w7021;
w7023 <= not w6589 and not w6591;
w7024 <= not w6963 and w7023;
w7025 <= not w6598 and not w7024;
w7026 <= not w7022 and not w7025;
w7027 <= not w7019 and not w7026;
w7028 <= not w7017 and not w7027;
w7029 <= not w4718 and not w7028;
w7030 <= w6608 and not w6610;
w7031 <= not w6601 and w7030;
w7032 <= not w6963 and w7031;
w7033 <= not w6601 and not w6610;
w7034 <= not w6963 and w7033;
w7035 <= not w6608 and not w7034;
w7036 <= not w7032 and not w7035;
w7037 <= w4718 and not w7017;
w7038 <= not w7027 and w7037;
w7039 <= not w7036 and not w7038;
w7040 <= not w7029 and not w7039;
w7041 <= not w4386 and not w7040;
w7042 <= not w6613 and w6620;
w7043 <= not w6622 and w7042;
w7044 <= not w6963 and w7043;
w7045 <= not w6613 and not w6622;
w7046 <= not w6963 and w7045;
w7047 <= not w6620 and not w7046;
w7048 <= not w7044 and not w7047;
w7049 <= w4386 and not w7029;
w7050 <= not w7039 and w7049;
w7051 <= not w7048 and not w7050;
w7052 <= not w7041 and not w7051;
w7053 <= not w4066 and not w7052;
w7054 <= w6632 and not w6634;
w7055 <= not w6625 and w7054;
w7056 <= not w6963 and w7055;
w7057 <= not w6625 and not w6634;
w7058 <= not w6963 and w7057;
w7059 <= not w6632 and not w7058;
w7060 <= not w7056 and not w7059;
w7061 <= w4066 and not w7041;
w7062 <= not w7051 and w7061;
w7063 <= not w7060 and not w7062;
w7064 <= not w7053 and not w7063;
w7065 <= not w3758 and not w7064;
w7066 <= not w6637 and w6644;
w7067 <= not w6646 and w7066;
w7068 <= not w6963 and w7067;
w7069 <= not w6637 and not w6646;
w7070 <= not w6963 and w7069;
w7071 <= not w6644 and not w7070;
w7072 <= not w7068 and not w7071;
w7073 <= w3758 and not w7053;
w7074 <= not w7063 and w7073;
w7075 <= not w7072 and not w7074;
w7076 <= not w7065 and not w7075;
w7077 <= not w3462 and not w7076;
w7078 <= w6656 and not w6658;
w7079 <= not w6649 and w7078;
w7080 <= not w6963 and w7079;
w7081 <= not w6649 and not w6658;
w7082 <= not w6963 and w7081;
w7083 <= not w6656 and not w7082;
w7084 <= not w7080 and not w7083;
w7085 <= w3462 and not w7065;
w7086 <= not w7075 and w7085;
w7087 <= not w7084 and not w7086;
w7088 <= not w7077 and not w7087;
w7089 <= not w3178 and not w7088;
w7090 <= not w6661 and w6668;
w7091 <= not w6670 and w7090;
w7092 <= not w6963 and w7091;
w7093 <= not w6661 and not w6670;
w7094 <= not w6963 and w7093;
w7095 <= not w6668 and not w7094;
w7096 <= not w7092 and not w7095;
w7097 <= w3178 and not w7077;
w7098 <= not w7087 and w7097;
w7099 <= not w7096 and not w7098;
w7100 <= not w7089 and not w7099;
w7101 <= not w2906 and not w7100;
w7102 <= w6680 and not w6682;
w7103 <= not w6673 and w7102;
w7104 <= not w6963 and w7103;
w7105 <= not w6673 and not w6682;
w7106 <= not w6963 and w7105;
w7107 <= not w6680 and not w7106;
w7108 <= not w7104 and not w7107;
w7109 <= w2906 and not w7089;
w7110 <= not w7099 and w7109;
w7111 <= not w7108 and not w7110;
w7112 <= not w7101 and not w7111;
w7113 <= not w2646 and not w7112;
w7114 <= not w6685 and w6692;
w7115 <= not w6694 and w7114;
w7116 <= not w6963 and w7115;
w7117 <= not w6685 and not w6694;
w7118 <= not w6963 and w7117;
w7119 <= not w6692 and not w7118;
w7120 <= not w7116 and not w7119;
w7121 <= w2646 and not w7101;
w7122 <= not w7111 and w7121;
w7123 <= not w7120 and not w7122;
w7124 <= not w7113 and not w7123;
w7125 <= not w2398 and not w7124;
w7126 <= w6704 and not w6706;
w7127 <= not w6697 and w7126;
w7128 <= not w6963 and w7127;
w7129 <= not w6697 and not w6706;
w7130 <= not w6963 and w7129;
w7131 <= not w6704 and not w7130;
w7132 <= not w7128 and not w7131;
w7133 <= w2398 and not w7113;
w7134 <= not w7123 and w7133;
w7135 <= not w7132 and not w7134;
w7136 <= not w7125 and not w7135;
w7137 <= not w2162 and not w7136;
w7138 <= not w6709 and w6716;
w7139 <= not w6718 and w7138;
w7140 <= not w6963 and w7139;
w7141 <= not w6709 and not w6718;
w7142 <= not w6963 and w7141;
w7143 <= not w6716 and not w7142;
w7144 <= not w7140 and not w7143;
w7145 <= w2162 and not w7125;
w7146 <= not w7135 and w7145;
w7147 <= not w7144 and not w7146;
w7148 <= not w7137 and not w7147;
w7149 <= not w1938 and not w7148;
w7150 <= w6728 and not w6730;
w7151 <= not w6721 and w7150;
w7152 <= not w6963 and w7151;
w7153 <= not w6721 and not w6730;
w7154 <= not w6963 and w7153;
w7155 <= not w6728 and not w7154;
w7156 <= not w7152 and not w7155;
w7157 <= w1938 and not w7137;
w7158 <= not w7147 and w7157;
w7159 <= not w7156 and not w7158;
w7160 <= not w7149 and not w7159;
w7161 <= not w1725 and not w7160;
w7162 <= not w6733 and w6740;
w7163 <= not w6742 and w7162;
w7164 <= not w6963 and w7163;
w7165 <= not w6733 and not w6742;
w7166 <= not w6963 and w7165;
w7167 <= not w6740 and not w7166;
w7168 <= not w7164 and not w7167;
w7169 <= w1725 and not w7149;
w7170 <= not w7159 and w7169;
w7171 <= not w7168 and not w7170;
w7172 <= not w7161 and not w7171;
w7173 <= not w1525 and not w7172;
w7174 <= w6752 and not w6754;
w7175 <= not w6745 and w7174;
w7176 <= not w6963 and w7175;
w7177 <= not w6745 and not w6754;
w7178 <= not w6963 and w7177;
w7179 <= not w6752 and not w7178;
w7180 <= not w7176 and not w7179;
w7181 <= w1525 and not w7161;
w7182 <= not w7171 and w7181;
w7183 <= not w7180 and not w7182;
w7184 <= not w7173 and not w7183;
w7185 <= not w1337 and not w7184;
w7186 <= not w6757 and w6764;
w7187 <= not w6766 and w7186;
w7188 <= not w6963 and w7187;
w7189 <= not w6757 and not w6766;
w7190 <= not w6963 and w7189;
w7191 <= not w6764 and not w7190;
w7192 <= not w7188 and not w7191;
w7193 <= w1337 and not w7173;
w7194 <= not w7183 and w7193;
w7195 <= not w7192 and not w7194;
w7196 <= not w7185 and not w7195;
w7197 <= not w1161 and not w7196;
w7198 <= w6776 and not w6778;
w7199 <= not w6769 and w7198;
w7200 <= not w6963 and w7199;
w7201 <= not w6769 and not w6778;
w7202 <= not w6963 and w7201;
w7203 <= not w6776 and not w7202;
w7204 <= not w7200 and not w7203;
w7205 <= w1161 and not w7185;
w7206 <= not w7195 and w7205;
w7207 <= not w7204 and not w7206;
w7208 <= not w7197 and not w7207;
w7209 <= not w997 and not w7208;
w7210 <= not w6781 and w6788;
w7211 <= not w6790 and w7210;
w7212 <= not w6963 and w7211;
w7213 <= not w6781 and not w6790;
w7214 <= not w6963 and w7213;
w7215 <= not w6788 and not w7214;
w7216 <= not w7212 and not w7215;
w7217 <= w997 and not w7197;
w7218 <= not w7207 and w7217;
w7219 <= not w7216 and not w7218;
w7220 <= not w7209 and not w7219;
w7221 <= not w845 and not w7220;
w7222 <= w6800 and not w6802;
w7223 <= not w6793 and w7222;
w7224 <= not w6963 and w7223;
w7225 <= not w6793 and not w6802;
w7226 <= not w6963 and w7225;
w7227 <= not w6800 and not w7226;
w7228 <= not w7224 and not w7227;
w7229 <= w845 and not w7209;
w7230 <= not w7219 and w7229;
w7231 <= not w7228 and not w7230;
w7232 <= not w7221 and not w7231;
w7233 <= not w705 and not w7232;
w7234 <= not w6805 and w6812;
w7235 <= not w6814 and w7234;
w7236 <= not w6963 and w7235;
w7237 <= not w6805 and not w6814;
w7238 <= not w6963 and w7237;
w7239 <= not w6812 and not w7238;
w7240 <= not w7236 and not w7239;
w7241 <= w705 and not w7221;
w7242 <= not w7231 and w7241;
w7243 <= not w7240 and not w7242;
w7244 <= not w7233 and not w7243;
w7245 <= not w577 and not w7244;
w7246 <= w6824 and not w6826;
w7247 <= not w6817 and w7246;
w7248 <= not w6963 and w7247;
w7249 <= not w6817 and not w6826;
w7250 <= not w6963 and w7249;
w7251 <= not w6824 and not w7250;
w7252 <= not w7248 and not w7251;
w7253 <= w577 and not w7233;
w7254 <= not w7243 and w7253;
w7255 <= not w7252 and not w7254;
w7256 <= not w7245 and not w7255;
w7257 <= not w460 and not w7256;
w7258 <= not w6829 and w6836;
w7259 <= not w6838 and w7258;
w7260 <= not w6963 and w7259;
w7261 <= not w6829 and not w6838;
w7262 <= not w6963 and w7261;
w7263 <= not w6836 and not w7262;
w7264 <= not w7260 and not w7263;
w7265 <= w460 and not w7245;
w7266 <= not w7255 and w7265;
w7267 <= not w7264 and not w7266;
w7268 <= not w7257 and not w7267;
w7269 <= not w356 and not w7268;
w7270 <= w6848 and not w6850;
w7271 <= not w6841 and w7270;
w7272 <= not w6963 and w7271;
w7273 <= not w6841 and not w6850;
w7274 <= not w6963 and w7273;
w7275 <= not w6848 and not w7274;
w7276 <= not w7272 and not w7275;
w7277 <= w356 and not w7257;
w7278 <= not w7267 and w7277;
w7279 <= not w7276 and not w7278;
w7280 <= not w7269 and not w7279;
w7281 <= not w264 and not w7280;
w7282 <= not w6853 and w6860;
w7283 <= not w6862 and w7282;
w7284 <= not w6963 and w7283;
w7285 <= not w6853 and not w6862;
w7286 <= not w6963 and w7285;
w7287 <= not w6860 and not w7286;
w7288 <= not w7284 and not w7287;
w7289 <= w264 and not w7269;
w7290 <= not w7279 and w7289;
w7291 <= not w7288 and not w7290;
w7292 <= not w7281 and not w7291;
w7293 <= not w184 and not w7292;
w7294 <= w6872 and not w6874;
w7295 <= not w6865 and w7294;
w7296 <= not w6963 and w7295;
w7297 <= not w6865 and not w6874;
w7298 <= not w6963 and w7297;
w7299 <= not w6872 and not w7298;
w7300 <= not w7296 and not w7299;
w7301 <= w184 and not w7281;
w7302 <= not w7291 and w7301;
w7303 <= not w7300 and not w7302;
w7304 <= not w7293 and not w7303;
w7305 <= not w115 and not w7304;
w7306 <= not w6877 and w6884;
w7307 <= not w6886 and w7306;
w7308 <= not w6963 and w7307;
w7309 <= not w6877 and not w6886;
w7310 <= not w6963 and w7309;
w7311 <= not w6884 and not w7310;
w7312 <= not w7308 and not w7311;
w7313 <= w115 and not w7293;
w7314 <= not w7303 and w7313;
w7315 <= not w7312 and not w7314;
w7316 <= not w7305 and not w7315;
w7317 <= not w60 and not w7316;
w7318 <= w6896 and not w6898;
w7319 <= not w6889 and w7318;
w7320 <= not w6963 and w7319;
w7321 <= not w6889 and not w6898;
w7322 <= not w6963 and w7321;
w7323 <= not w6896 and not w7322;
w7324 <= not w7320 and not w7323;
w7325 <= w60 and not w7305;
w7326 <= not w7315 and w7325;
w7327 <= not w7324 and not w7326;
w7328 <= not w7317 and not w7327;
w7329 <= not w22 and not w7328;
w7330 <= not w6901 and w6908;
w7331 <= not w6910 and w7330;
w7332 <= not w6963 and w7331;
w7333 <= not w6901 and not w6910;
w7334 <= not w6963 and w7333;
w7335 <= not w6908 and not w7334;
w7336 <= not w7332 and not w7335;
w7337 <= w22 and not w7317;
w7338 <= not w7327 and w7337;
w7339 <= not w7336 and not w7338;
w7340 <= not w7329 and not w7339;
w7341 <= not w5 and not w7340;
w7342 <= w6920 and not w6922;
w7343 <= not w6913 and w7342;
w7344 <= not w6963 and w7343;
w7345 <= not w6913 and not w6922;
w7346 <= not w6963 and w7345;
w7347 <= not w6920 and not w7346;
w7348 <= not w7344 and not w7347;
w7349 <= w5 and not w7329;
w7350 <= not w7339 and w7349;
w7351 <= not w7348 and not w7350;
w7352 <= not w7341 and not w7351;
w7353 <= not w6925 and w6932;
w7354 <= not w6934 and w7353;
w7355 <= not w6963 and w7354;
w7356 <= not w6925 and not w6934;
w7357 <= not w6963 and w7356;
w7358 <= not w6932 and not w7357;
w7359 <= not w7355 and not w7358;
w7360 <= not w6936 and not w6943;
w7361 <= not w6963 and w7360;
w7362 <= not w6951 and not w7361;
w7363 <= not w7359 and w7362;
w7364 <= not w7352 and w7363;
w7365 <= w0 and not w7364;
w7366 <= not w7341 and w7359;
w7367 <= not w7351 and w7366;
w7368 <= not w6943 and not w6963;
w7369 <= w6936 and not w7368;
w7370 <= not w0 and not w7360;
w7371 <= not w7369 and w7370;
w7372 <= not w6939 and not w6960;
w7373 <= not w6942 and w7372;
w7374 <= not w6955 and w7373;
w7375 <= not w6951 and w7374;
w7376 <= not w6949 and w7375;
w7377 <= not w7371 and not w7376;
w7378 <= not w7367 and w7377;
w7379 <= not w7365 and w7378;
w7380 <= a(58) and not w7379;
w7381 <= not a(56) and not a(57);
w7382 <= not a(58) and w7381;
w7383 <= not w7380 and not w7382;
w7384 <= not w6963 and not w7383;
w7385 <= not w6960 and not w7382;
w7386 <= not w6955 and w7385;
w7387 <= not w6951 and w7386;
w7388 <= not w6949 and w7387;
w7389 <= not w7380 and w7388;
w7390 <= not a(58) and not w7379;
w7391 <= a(59) and not w7390;
w7392 <= w6965 and not w7379;
w7393 <= not w7391 and not w7392;
w7394 <= not w7389 and w7393;
w7395 <= not w7384 and not w7394;
w7396 <= not w6558 and not w7395;
w7397 <= w6558 and not w7384;
w7398 <= not w7394 and w7397;
w7399 <= not w6963 and not w7376;
w7400 <= not w7371 and w7399;
w7401 <= not w7367 and w7400;
w7402 <= not w7365 and w7401;
w7403 <= not w7392 and not w7402;
w7404 <= a(60) and not w7403;
w7405 <= not a(60) and not w7402;
w7406 <= not w7392 and w7405;
w7407 <= not w7404 and not w7406;
w7408 <= not w7398 and not w7407;
w7409 <= not w7396 and not w7408;
w7410 <= not w6166 and not w7409;
w7411 <= not w6968 and not w6973;
w7412 <= not w6977 and w7411;
w7413 <= not w7379 and w7412;
w7414 <= not w7379 and w7411;
w7415 <= w6977 and not w7414;
w7416 <= not w7413 and not w7415;
w7417 <= w6166 and not w7396;
w7418 <= not w7408 and w7417;
w7419 <= not w7416 and not w7418;
w7420 <= not w7410 and not w7419;
w7421 <= not w5786 and not w7420;
w7422 <= not w6982 and w6991;
w7423 <= not w6980 and w7422;
w7424 <= not w7379 and w7423;
w7425 <= not w6980 and not w6982;
w7426 <= not w7379 and w7425;
w7427 <= not w6991 and not w7426;
w7428 <= not w7424 and not w7427;
w7429 <= w5786 and not w7410;
w7430 <= not w7419 and w7429;
w7431 <= not w7428 and not w7430;
w7432 <= not w7421 and not w7431;
w7433 <= not w5418 and not w7432;
w7434 <= not w6994 and w7000;
w7435 <= not w7002 and w7434;
w7436 <= not w7379 and w7435;
w7437 <= not w6994 and not w7002;
w7438 <= not w7379 and w7437;
w7439 <= not w7000 and not w7438;
w7440 <= not w7436 and not w7439;
w7441 <= w5418 and not w7421;
w7442 <= not w7431 and w7441;
w7443 <= not w7440 and not w7442;
w7444 <= not w7433 and not w7443;
w7445 <= not w5062 and not w7444;
w7446 <= w7012 and not w7014;
w7447 <= not w7005 and w7446;
w7448 <= not w7379 and w7447;
w7449 <= not w7005 and not w7014;
w7450 <= not w7379 and w7449;
w7451 <= not w7012 and not w7450;
w7452 <= not w7448 and not w7451;
w7453 <= w5062 and not w7433;
w7454 <= not w7443 and w7453;
w7455 <= not w7452 and not w7454;
w7456 <= not w7445 and not w7455;
w7457 <= not w4718 and not w7456;
w7458 <= w4718 and not w7445;
w7459 <= not w7455 and w7458;
w7460 <= not w7017 and w7026;
w7461 <= not w7019 and w7460;
w7462 <= not w7379 and w7461;
w7463 <= not w7017 and not w7019;
w7464 <= not w7379 and w7463;
w7465 <= not w7026 and not w7464;
w7466 <= not w7462 and not w7465;
w7467 <= not w7459 and not w7466;
w7468 <= not w7457 and not w7467;
w7469 <= not w4386 and not w7468;
w7470 <= w7036 and not w7038;
w7471 <= not w7029 and w7470;
w7472 <= not w7379 and w7471;
w7473 <= not w7029 and not w7038;
w7474 <= not w7379 and w7473;
w7475 <= not w7036 and not w7474;
w7476 <= not w7472 and not w7475;
w7477 <= w4386 and not w7457;
w7478 <= not w7467 and w7477;
w7479 <= not w7476 and not w7478;
w7480 <= not w7469 and not w7479;
w7481 <= not w4066 and not w7480;
w7482 <= not w7041 and w7048;
w7483 <= not w7050 and w7482;
w7484 <= not w7379 and w7483;
w7485 <= not w7041 and not w7050;
w7486 <= not w7379 and w7485;
w7487 <= not w7048 and not w7486;
w7488 <= not w7484 and not w7487;
w7489 <= w4066 and not w7469;
w7490 <= not w7479 and w7489;
w7491 <= not w7488 and not w7490;
w7492 <= not w7481 and not w7491;
w7493 <= not w3758 and not w7492;
w7494 <= w7060 and not w7062;
w7495 <= not w7053 and w7494;
w7496 <= not w7379 and w7495;
w7497 <= not w7053 and not w7062;
w7498 <= not w7379 and w7497;
w7499 <= not w7060 and not w7498;
w7500 <= not w7496 and not w7499;
w7501 <= w3758 and not w7481;
w7502 <= not w7491 and w7501;
w7503 <= not w7500 and not w7502;
w7504 <= not w7493 and not w7503;
w7505 <= not w3462 and not w7504;
w7506 <= not w7065 and w7072;
w7507 <= not w7074 and w7506;
w7508 <= not w7379 and w7507;
w7509 <= not w7065 and not w7074;
w7510 <= not w7379 and w7509;
w7511 <= not w7072 and not w7510;
w7512 <= not w7508 and not w7511;
w7513 <= w3462 and not w7493;
w7514 <= not w7503 and w7513;
w7515 <= not w7512 and not w7514;
w7516 <= not w7505 and not w7515;
w7517 <= not w3178 and not w7516;
w7518 <= w7084 and not w7086;
w7519 <= not w7077 and w7518;
w7520 <= not w7379 and w7519;
w7521 <= not w7077 and not w7086;
w7522 <= not w7379 and w7521;
w7523 <= not w7084 and not w7522;
w7524 <= not w7520 and not w7523;
w7525 <= w3178 and not w7505;
w7526 <= not w7515 and w7525;
w7527 <= not w7524 and not w7526;
w7528 <= not w7517 and not w7527;
w7529 <= not w2906 and not w7528;
w7530 <= not w7089 and w7096;
w7531 <= not w7098 and w7530;
w7532 <= not w7379 and w7531;
w7533 <= not w7089 and not w7098;
w7534 <= not w7379 and w7533;
w7535 <= not w7096 and not w7534;
w7536 <= not w7532 and not w7535;
w7537 <= w2906 and not w7517;
w7538 <= not w7527 and w7537;
w7539 <= not w7536 and not w7538;
w7540 <= not w7529 and not w7539;
w7541 <= not w2646 and not w7540;
w7542 <= w7108 and not w7110;
w7543 <= not w7101 and w7542;
w7544 <= not w7379 and w7543;
w7545 <= not w7101 and not w7110;
w7546 <= not w7379 and w7545;
w7547 <= not w7108 and not w7546;
w7548 <= not w7544 and not w7547;
w7549 <= w2646 and not w7529;
w7550 <= not w7539 and w7549;
w7551 <= not w7548 and not w7550;
w7552 <= not w7541 and not w7551;
w7553 <= not w2398 and not w7552;
w7554 <= not w7113 and w7120;
w7555 <= not w7122 and w7554;
w7556 <= not w7379 and w7555;
w7557 <= not w7113 and not w7122;
w7558 <= not w7379 and w7557;
w7559 <= not w7120 and not w7558;
w7560 <= not w7556 and not w7559;
w7561 <= w2398 and not w7541;
w7562 <= not w7551 and w7561;
w7563 <= not w7560 and not w7562;
w7564 <= not w7553 and not w7563;
w7565 <= not w2162 and not w7564;
w7566 <= w7132 and not w7134;
w7567 <= not w7125 and w7566;
w7568 <= not w7379 and w7567;
w7569 <= not w7125 and not w7134;
w7570 <= not w7379 and w7569;
w7571 <= not w7132 and not w7570;
w7572 <= not w7568 and not w7571;
w7573 <= w2162 and not w7553;
w7574 <= not w7563 and w7573;
w7575 <= not w7572 and not w7574;
w7576 <= not w7565 and not w7575;
w7577 <= not w1938 and not w7576;
w7578 <= not w7137 and w7144;
w7579 <= not w7146 and w7578;
w7580 <= not w7379 and w7579;
w7581 <= not w7137 and not w7146;
w7582 <= not w7379 and w7581;
w7583 <= not w7144 and not w7582;
w7584 <= not w7580 and not w7583;
w7585 <= w1938 and not w7565;
w7586 <= not w7575 and w7585;
w7587 <= not w7584 and not w7586;
w7588 <= not w7577 and not w7587;
w7589 <= not w1725 and not w7588;
w7590 <= w7156 and not w7158;
w7591 <= not w7149 and w7590;
w7592 <= not w7379 and w7591;
w7593 <= not w7149 and not w7158;
w7594 <= not w7379 and w7593;
w7595 <= not w7156 and not w7594;
w7596 <= not w7592 and not w7595;
w7597 <= w1725 and not w7577;
w7598 <= not w7587 and w7597;
w7599 <= not w7596 and not w7598;
w7600 <= not w7589 and not w7599;
w7601 <= not w1525 and not w7600;
w7602 <= not w7161 and w7168;
w7603 <= not w7170 and w7602;
w7604 <= not w7379 and w7603;
w7605 <= not w7161 and not w7170;
w7606 <= not w7379 and w7605;
w7607 <= not w7168 and not w7606;
w7608 <= not w7604 and not w7607;
w7609 <= w1525 and not w7589;
w7610 <= not w7599 and w7609;
w7611 <= not w7608 and not w7610;
w7612 <= not w7601 and not w7611;
w7613 <= not w1337 and not w7612;
w7614 <= w7180 and not w7182;
w7615 <= not w7173 and w7614;
w7616 <= not w7379 and w7615;
w7617 <= not w7173 and not w7182;
w7618 <= not w7379 and w7617;
w7619 <= not w7180 and not w7618;
w7620 <= not w7616 and not w7619;
w7621 <= w1337 and not w7601;
w7622 <= not w7611 and w7621;
w7623 <= not w7620 and not w7622;
w7624 <= not w7613 and not w7623;
w7625 <= not w1161 and not w7624;
w7626 <= not w7185 and w7192;
w7627 <= not w7194 and w7626;
w7628 <= not w7379 and w7627;
w7629 <= not w7185 and not w7194;
w7630 <= not w7379 and w7629;
w7631 <= not w7192 and not w7630;
w7632 <= not w7628 and not w7631;
w7633 <= w1161 and not w7613;
w7634 <= not w7623 and w7633;
w7635 <= not w7632 and not w7634;
w7636 <= not w7625 and not w7635;
w7637 <= not w997 and not w7636;
w7638 <= w7204 and not w7206;
w7639 <= not w7197 and w7638;
w7640 <= not w7379 and w7639;
w7641 <= not w7197 and not w7206;
w7642 <= not w7379 and w7641;
w7643 <= not w7204 and not w7642;
w7644 <= not w7640 and not w7643;
w7645 <= w997 and not w7625;
w7646 <= not w7635 and w7645;
w7647 <= not w7644 and not w7646;
w7648 <= not w7637 and not w7647;
w7649 <= not w845 and not w7648;
w7650 <= not w7209 and w7216;
w7651 <= not w7218 and w7650;
w7652 <= not w7379 and w7651;
w7653 <= not w7209 and not w7218;
w7654 <= not w7379 and w7653;
w7655 <= not w7216 and not w7654;
w7656 <= not w7652 and not w7655;
w7657 <= w845 and not w7637;
w7658 <= not w7647 and w7657;
w7659 <= not w7656 and not w7658;
w7660 <= not w7649 and not w7659;
w7661 <= not w705 and not w7660;
w7662 <= w7228 and not w7230;
w7663 <= not w7221 and w7662;
w7664 <= not w7379 and w7663;
w7665 <= not w7221 and not w7230;
w7666 <= not w7379 and w7665;
w7667 <= not w7228 and not w7666;
w7668 <= not w7664 and not w7667;
w7669 <= w705 and not w7649;
w7670 <= not w7659 and w7669;
w7671 <= not w7668 and not w7670;
w7672 <= not w7661 and not w7671;
w7673 <= not w577 and not w7672;
w7674 <= not w7233 and w7240;
w7675 <= not w7242 and w7674;
w7676 <= not w7379 and w7675;
w7677 <= not w7233 and not w7242;
w7678 <= not w7379 and w7677;
w7679 <= not w7240 and not w7678;
w7680 <= not w7676 and not w7679;
w7681 <= w577 and not w7661;
w7682 <= not w7671 and w7681;
w7683 <= not w7680 and not w7682;
w7684 <= not w7673 and not w7683;
w7685 <= not w460 and not w7684;
w7686 <= w7252 and not w7254;
w7687 <= not w7245 and w7686;
w7688 <= not w7379 and w7687;
w7689 <= not w7245 and not w7254;
w7690 <= not w7379 and w7689;
w7691 <= not w7252 and not w7690;
w7692 <= not w7688 and not w7691;
w7693 <= w460 and not w7673;
w7694 <= not w7683 and w7693;
w7695 <= not w7692 and not w7694;
w7696 <= not w7685 and not w7695;
w7697 <= not w356 and not w7696;
w7698 <= not w7257 and w7264;
w7699 <= not w7266 and w7698;
w7700 <= not w7379 and w7699;
w7701 <= not w7257 and not w7266;
w7702 <= not w7379 and w7701;
w7703 <= not w7264 and not w7702;
w7704 <= not w7700 and not w7703;
w7705 <= w356 and not w7685;
w7706 <= not w7695 and w7705;
w7707 <= not w7704 and not w7706;
w7708 <= not w7697 and not w7707;
w7709 <= not w264 and not w7708;
w7710 <= w7276 and not w7278;
w7711 <= not w7269 and w7710;
w7712 <= not w7379 and w7711;
w7713 <= not w7269 and not w7278;
w7714 <= not w7379 and w7713;
w7715 <= not w7276 and not w7714;
w7716 <= not w7712 and not w7715;
w7717 <= w264 and not w7697;
w7718 <= not w7707 and w7717;
w7719 <= not w7716 and not w7718;
w7720 <= not w7709 and not w7719;
w7721 <= not w184 and not w7720;
w7722 <= not w7281 and w7288;
w7723 <= not w7290 and w7722;
w7724 <= not w7379 and w7723;
w7725 <= not w7281 and not w7290;
w7726 <= not w7379 and w7725;
w7727 <= not w7288 and not w7726;
w7728 <= not w7724 and not w7727;
w7729 <= w184 and not w7709;
w7730 <= not w7719 and w7729;
w7731 <= not w7728 and not w7730;
w7732 <= not w7721 and not w7731;
w7733 <= not w115 and not w7732;
w7734 <= w7300 and not w7302;
w7735 <= not w7293 and w7734;
w7736 <= not w7379 and w7735;
w7737 <= not w7293 and not w7302;
w7738 <= not w7379 and w7737;
w7739 <= not w7300 and not w7738;
w7740 <= not w7736 and not w7739;
w7741 <= w115 and not w7721;
w7742 <= not w7731 and w7741;
w7743 <= not w7740 and not w7742;
w7744 <= not w7733 and not w7743;
w7745 <= not w60 and not w7744;
w7746 <= not w7305 and w7312;
w7747 <= not w7314 and w7746;
w7748 <= not w7379 and w7747;
w7749 <= not w7305 and not w7314;
w7750 <= not w7379 and w7749;
w7751 <= not w7312 and not w7750;
w7752 <= not w7748 and not w7751;
w7753 <= w60 and not w7733;
w7754 <= not w7743 and w7753;
w7755 <= not w7752 and not w7754;
w7756 <= not w7745 and not w7755;
w7757 <= not w22 and not w7756;
w7758 <= w7324 and not w7326;
w7759 <= not w7317 and w7758;
w7760 <= not w7379 and w7759;
w7761 <= not w7317 and not w7326;
w7762 <= not w7379 and w7761;
w7763 <= not w7324 and not w7762;
w7764 <= not w7760 and not w7763;
w7765 <= w22 and not w7745;
w7766 <= not w7755 and w7765;
w7767 <= not w7764 and not w7766;
w7768 <= not w7757 and not w7767;
w7769 <= not w5 and not w7768;
w7770 <= not w7329 and w7336;
w7771 <= not w7338 and w7770;
w7772 <= not w7379 and w7771;
w7773 <= not w7329 and not w7338;
w7774 <= not w7379 and w7773;
w7775 <= not w7336 and not w7774;
w7776 <= not w7772 and not w7775;
w7777 <= w5 and not w7757;
w7778 <= not w7767 and w7777;
w7779 <= not w7776 and not w7778;
w7780 <= not w7769 and not w7779;
w7781 <= w7348 and not w7350;
w7782 <= not w7341 and w7781;
w7783 <= not w7379 and w7782;
w7784 <= not w7341 and not w7350;
w7785 <= not w7379 and w7784;
w7786 <= not w7348 and not w7785;
w7787 <= not w7783 and not w7786;
w7788 <= not w7352 and not w7359;
w7789 <= not w7379 and w7788;
w7790 <= not w7367 and not w7789;
w7791 <= not w7787 and w7790;
w7792 <= not w7780 and w7791;
w7793 <= w0 and not w7792;
w7794 <= not w7769 and w7787;
w7795 <= not w7779 and w7794;
w7796 <= not w7359 and not w7379;
w7797 <= w7352 and not w7796;
w7798 <= not w0 and not w7788;
w7799 <= not w7797 and w7798;
w7800 <= not w7355 and not w7376;
w7801 <= not w7358 and w7800;
w7802 <= not w7371 and w7801;
w7803 <= not w7367 and w7802;
w7804 <= not w7365 and w7803;
w7805 <= not w7799 and not w7804;
w7806 <= not w7795 and w7805;
w7807 <= not w7793 and w7806;
w7808 <= a(56) and not w7807;
w7809 <= not a(54) and not a(55);
w7810 <= not a(56) and w7809;
w7811 <= not w7808 and not w7810;
w7812 <= not w7379 and not w7811;
w7813 <= not w7376 and not w7810;
w7814 <= not w7371 and w7813;
w7815 <= not w7367 and w7814;
w7816 <= not w7365 and w7815;
w7817 <= not w7808 and w7816;
w7818 <= not a(56) and not w7807;
w7819 <= a(57) and not w7818;
w7820 <= w7381 and not w7807;
w7821 <= not w7819 and not w7820;
w7822 <= not w7817 and w7821;
w7823 <= not w7812 and not w7822;
w7824 <= not w6963 and not w7823;
w7825 <= w6963 and not w7812;
w7826 <= not w7822 and w7825;
w7827 <= not w7379 and not w7804;
w7828 <= not w7799 and w7827;
w7829 <= not w7795 and w7828;
w7830 <= not w7793 and w7829;
w7831 <= not w7820 and not w7830;
w7832 <= a(58) and not w7831;
w7833 <= not a(58) and not w7830;
w7834 <= not w7820 and w7833;
w7835 <= not w7832 and not w7834;
w7836 <= not w7826 and not w7835;
w7837 <= not w7824 and not w7836;
w7838 <= not w6558 and not w7837;
w7839 <= not w7384 and not w7389;
w7840 <= not w7393 and w7839;
w7841 <= not w7807 and w7840;
w7842 <= not w7807 and w7839;
w7843 <= w7393 and not w7842;
w7844 <= not w7841 and not w7843;
w7845 <= w6558 and not w7824;
w7846 <= not w7836 and w7845;
w7847 <= not w7844 and not w7846;
w7848 <= not w7838 and not w7847;
w7849 <= not w6166 and not w7848;
w7850 <= not w7398 and w7407;
w7851 <= not w7396 and w7850;
w7852 <= not w7807 and w7851;
w7853 <= not w7396 and not w7398;
w7854 <= not w7807 and w7853;
w7855 <= not w7407 and not w7854;
w7856 <= not w7852 and not w7855;
w7857 <= w6166 and not w7838;
w7858 <= not w7847 and w7857;
w7859 <= not w7856 and not w7858;
w7860 <= not w7849 and not w7859;
w7861 <= not w5786 and not w7860;
w7862 <= not w7410 and w7416;
w7863 <= not w7418 and w7862;
w7864 <= not w7807 and w7863;
w7865 <= not w7410 and not w7418;
w7866 <= not w7807 and w7865;
w7867 <= not w7416 and not w7866;
w7868 <= not w7864 and not w7867;
w7869 <= w5786 and not w7849;
w7870 <= not w7859 and w7869;
w7871 <= not w7868 and not w7870;
w7872 <= not w7861 and not w7871;
w7873 <= not w5418 and not w7872;
w7874 <= w7428 and not w7430;
w7875 <= not w7421 and w7874;
w7876 <= not w7807 and w7875;
w7877 <= not w7421 and not w7430;
w7878 <= not w7807 and w7877;
w7879 <= not w7428 and not w7878;
w7880 <= not w7876 and not w7879;
w7881 <= w5418 and not w7861;
w7882 <= not w7871 and w7881;
w7883 <= not w7880 and not w7882;
w7884 <= not w7873 and not w7883;
w7885 <= not w5062 and not w7884;
w7886 <= not w7433 and w7440;
w7887 <= not w7442 and w7886;
w7888 <= not w7807 and w7887;
w7889 <= not w7433 and not w7442;
w7890 <= not w7807 and w7889;
w7891 <= not w7440 and not w7890;
w7892 <= not w7888 and not w7891;
w7893 <= w5062 and not w7873;
w7894 <= not w7883 and w7893;
w7895 <= not w7892 and not w7894;
w7896 <= not w7885 and not w7895;
w7897 <= not w4718 and not w7896;
w7898 <= w7452 and not w7454;
w7899 <= not w7445 and w7898;
w7900 <= not w7807 and w7899;
w7901 <= not w7445 and not w7454;
w7902 <= not w7807 and w7901;
w7903 <= not w7452 and not w7902;
w7904 <= not w7900 and not w7903;
w7905 <= w4718 and not w7885;
w7906 <= not w7895 and w7905;
w7907 <= not w7904 and not w7906;
w7908 <= not w7897 and not w7907;
w7909 <= not w4386 and not w7908;
w7910 <= w4386 and not w7897;
w7911 <= not w7907 and w7910;
w7912 <= not w7457 and w7466;
w7913 <= not w7459 and w7912;
w7914 <= not w7807 and w7913;
w7915 <= not w7457 and not w7459;
w7916 <= not w7807 and w7915;
w7917 <= not w7466 and not w7916;
w7918 <= not w7914 and not w7917;
w7919 <= not w7911 and not w7918;
w7920 <= not w7909 and not w7919;
w7921 <= not w4066 and not w7920;
w7922 <= w7476 and not w7478;
w7923 <= not w7469 and w7922;
w7924 <= not w7807 and w7923;
w7925 <= not w7469 and not w7478;
w7926 <= not w7807 and w7925;
w7927 <= not w7476 and not w7926;
w7928 <= not w7924 and not w7927;
w7929 <= w4066 and not w7909;
w7930 <= not w7919 and w7929;
w7931 <= not w7928 and not w7930;
w7932 <= not w7921 and not w7931;
w7933 <= not w3758 and not w7932;
w7934 <= not w7481 and w7488;
w7935 <= not w7490 and w7934;
w7936 <= not w7807 and w7935;
w7937 <= not w7481 and not w7490;
w7938 <= not w7807 and w7937;
w7939 <= not w7488 and not w7938;
w7940 <= not w7936 and not w7939;
w7941 <= w3758 and not w7921;
w7942 <= not w7931 and w7941;
w7943 <= not w7940 and not w7942;
w7944 <= not w7933 and not w7943;
w7945 <= not w3462 and not w7944;
w7946 <= w7500 and not w7502;
w7947 <= not w7493 and w7946;
w7948 <= not w7807 and w7947;
w7949 <= not w7493 and not w7502;
w7950 <= not w7807 and w7949;
w7951 <= not w7500 and not w7950;
w7952 <= not w7948 and not w7951;
w7953 <= w3462 and not w7933;
w7954 <= not w7943 and w7953;
w7955 <= not w7952 and not w7954;
w7956 <= not w7945 and not w7955;
w7957 <= not w3178 and not w7956;
w7958 <= not w7505 and w7512;
w7959 <= not w7514 and w7958;
w7960 <= not w7807 and w7959;
w7961 <= not w7505 and not w7514;
w7962 <= not w7807 and w7961;
w7963 <= not w7512 and not w7962;
w7964 <= not w7960 and not w7963;
w7965 <= w3178 and not w7945;
w7966 <= not w7955 and w7965;
w7967 <= not w7964 and not w7966;
w7968 <= not w7957 and not w7967;
w7969 <= not w2906 and not w7968;
w7970 <= w7524 and not w7526;
w7971 <= not w7517 and w7970;
w7972 <= not w7807 and w7971;
w7973 <= not w7517 and not w7526;
w7974 <= not w7807 and w7973;
w7975 <= not w7524 and not w7974;
w7976 <= not w7972 and not w7975;
w7977 <= w2906 and not w7957;
w7978 <= not w7967 and w7977;
w7979 <= not w7976 and not w7978;
w7980 <= not w7969 and not w7979;
w7981 <= not w2646 and not w7980;
w7982 <= not w7529 and w7536;
w7983 <= not w7538 and w7982;
w7984 <= not w7807 and w7983;
w7985 <= not w7529 and not w7538;
w7986 <= not w7807 and w7985;
w7987 <= not w7536 and not w7986;
w7988 <= not w7984 and not w7987;
w7989 <= w2646 and not w7969;
w7990 <= not w7979 and w7989;
w7991 <= not w7988 and not w7990;
w7992 <= not w7981 and not w7991;
w7993 <= not w2398 and not w7992;
w7994 <= w7548 and not w7550;
w7995 <= not w7541 and w7994;
w7996 <= not w7807 and w7995;
w7997 <= not w7541 and not w7550;
w7998 <= not w7807 and w7997;
w7999 <= not w7548 and not w7998;
w8000 <= not w7996 and not w7999;
w8001 <= w2398 and not w7981;
w8002 <= not w7991 and w8001;
w8003 <= not w8000 and not w8002;
w8004 <= not w7993 and not w8003;
w8005 <= not w2162 and not w8004;
w8006 <= not w7553 and w7560;
w8007 <= not w7562 and w8006;
w8008 <= not w7807 and w8007;
w8009 <= not w7553 and not w7562;
w8010 <= not w7807 and w8009;
w8011 <= not w7560 and not w8010;
w8012 <= not w8008 and not w8011;
w8013 <= w2162 and not w7993;
w8014 <= not w8003 and w8013;
w8015 <= not w8012 and not w8014;
w8016 <= not w8005 and not w8015;
w8017 <= not w1938 and not w8016;
w8018 <= w7572 and not w7574;
w8019 <= not w7565 and w8018;
w8020 <= not w7807 and w8019;
w8021 <= not w7565 and not w7574;
w8022 <= not w7807 and w8021;
w8023 <= not w7572 and not w8022;
w8024 <= not w8020 and not w8023;
w8025 <= w1938 and not w8005;
w8026 <= not w8015 and w8025;
w8027 <= not w8024 and not w8026;
w8028 <= not w8017 and not w8027;
w8029 <= not w1725 and not w8028;
w8030 <= not w7577 and w7584;
w8031 <= not w7586 and w8030;
w8032 <= not w7807 and w8031;
w8033 <= not w7577 and not w7586;
w8034 <= not w7807 and w8033;
w8035 <= not w7584 and not w8034;
w8036 <= not w8032 and not w8035;
w8037 <= w1725 and not w8017;
w8038 <= not w8027 and w8037;
w8039 <= not w8036 and not w8038;
w8040 <= not w8029 and not w8039;
w8041 <= not w1525 and not w8040;
w8042 <= w7596 and not w7598;
w8043 <= not w7589 and w8042;
w8044 <= not w7807 and w8043;
w8045 <= not w7589 and not w7598;
w8046 <= not w7807 and w8045;
w8047 <= not w7596 and not w8046;
w8048 <= not w8044 and not w8047;
w8049 <= w1525 and not w8029;
w8050 <= not w8039 and w8049;
w8051 <= not w8048 and not w8050;
w8052 <= not w8041 and not w8051;
w8053 <= not w1337 and not w8052;
w8054 <= not w7601 and w7608;
w8055 <= not w7610 and w8054;
w8056 <= not w7807 and w8055;
w8057 <= not w7601 and not w7610;
w8058 <= not w7807 and w8057;
w8059 <= not w7608 and not w8058;
w8060 <= not w8056 and not w8059;
w8061 <= w1337 and not w8041;
w8062 <= not w8051 and w8061;
w8063 <= not w8060 and not w8062;
w8064 <= not w8053 and not w8063;
w8065 <= not w1161 and not w8064;
w8066 <= w7620 and not w7622;
w8067 <= not w7613 and w8066;
w8068 <= not w7807 and w8067;
w8069 <= not w7613 and not w7622;
w8070 <= not w7807 and w8069;
w8071 <= not w7620 and not w8070;
w8072 <= not w8068 and not w8071;
w8073 <= w1161 and not w8053;
w8074 <= not w8063 and w8073;
w8075 <= not w8072 and not w8074;
w8076 <= not w8065 and not w8075;
w8077 <= not w997 and not w8076;
w8078 <= not w7625 and w7632;
w8079 <= not w7634 and w8078;
w8080 <= not w7807 and w8079;
w8081 <= not w7625 and not w7634;
w8082 <= not w7807 and w8081;
w8083 <= not w7632 and not w8082;
w8084 <= not w8080 and not w8083;
w8085 <= w997 and not w8065;
w8086 <= not w8075 and w8085;
w8087 <= not w8084 and not w8086;
w8088 <= not w8077 and not w8087;
w8089 <= not w845 and not w8088;
w8090 <= w7644 and not w7646;
w8091 <= not w7637 and w8090;
w8092 <= not w7807 and w8091;
w8093 <= not w7637 and not w7646;
w8094 <= not w7807 and w8093;
w8095 <= not w7644 and not w8094;
w8096 <= not w8092 and not w8095;
w8097 <= w845 and not w8077;
w8098 <= not w8087 and w8097;
w8099 <= not w8096 and not w8098;
w8100 <= not w8089 and not w8099;
w8101 <= not w705 and not w8100;
w8102 <= not w7649 and w7656;
w8103 <= not w7658 and w8102;
w8104 <= not w7807 and w8103;
w8105 <= not w7649 and not w7658;
w8106 <= not w7807 and w8105;
w8107 <= not w7656 and not w8106;
w8108 <= not w8104 and not w8107;
w8109 <= w705 and not w8089;
w8110 <= not w8099 and w8109;
w8111 <= not w8108 and not w8110;
w8112 <= not w8101 and not w8111;
w8113 <= not w577 and not w8112;
w8114 <= w7668 and not w7670;
w8115 <= not w7661 and w8114;
w8116 <= not w7807 and w8115;
w8117 <= not w7661 and not w7670;
w8118 <= not w7807 and w8117;
w8119 <= not w7668 and not w8118;
w8120 <= not w8116 and not w8119;
w8121 <= w577 and not w8101;
w8122 <= not w8111 and w8121;
w8123 <= not w8120 and not w8122;
w8124 <= not w8113 and not w8123;
w8125 <= not w460 and not w8124;
w8126 <= not w7673 and w7680;
w8127 <= not w7682 and w8126;
w8128 <= not w7807 and w8127;
w8129 <= not w7673 and not w7682;
w8130 <= not w7807 and w8129;
w8131 <= not w7680 and not w8130;
w8132 <= not w8128 and not w8131;
w8133 <= w460 and not w8113;
w8134 <= not w8123 and w8133;
w8135 <= not w8132 and not w8134;
w8136 <= not w8125 and not w8135;
w8137 <= not w356 and not w8136;
w8138 <= w7692 and not w7694;
w8139 <= not w7685 and w8138;
w8140 <= not w7807 and w8139;
w8141 <= not w7685 and not w7694;
w8142 <= not w7807 and w8141;
w8143 <= not w7692 and not w8142;
w8144 <= not w8140 and not w8143;
w8145 <= w356 and not w8125;
w8146 <= not w8135 and w8145;
w8147 <= not w8144 and not w8146;
w8148 <= not w8137 and not w8147;
w8149 <= not w264 and not w8148;
w8150 <= not w7697 and w7704;
w8151 <= not w7706 and w8150;
w8152 <= not w7807 and w8151;
w8153 <= not w7697 and not w7706;
w8154 <= not w7807 and w8153;
w8155 <= not w7704 and not w8154;
w8156 <= not w8152 and not w8155;
w8157 <= w264 and not w8137;
w8158 <= not w8147 and w8157;
w8159 <= not w8156 and not w8158;
w8160 <= not w8149 and not w8159;
w8161 <= not w184 and not w8160;
w8162 <= w7716 and not w7718;
w8163 <= not w7709 and w8162;
w8164 <= not w7807 and w8163;
w8165 <= not w7709 and not w7718;
w8166 <= not w7807 and w8165;
w8167 <= not w7716 and not w8166;
w8168 <= not w8164 and not w8167;
w8169 <= w184 and not w8149;
w8170 <= not w8159 and w8169;
w8171 <= not w8168 and not w8170;
w8172 <= not w8161 and not w8171;
w8173 <= not w115 and not w8172;
w8174 <= not w7721 and w7728;
w8175 <= not w7730 and w8174;
w8176 <= not w7807 and w8175;
w8177 <= not w7721 and not w7730;
w8178 <= not w7807 and w8177;
w8179 <= not w7728 and not w8178;
w8180 <= not w8176 and not w8179;
w8181 <= w115 and not w8161;
w8182 <= not w8171 and w8181;
w8183 <= not w8180 and not w8182;
w8184 <= not w8173 and not w8183;
w8185 <= not w60 and not w8184;
w8186 <= w7740 and not w7742;
w8187 <= not w7733 and w8186;
w8188 <= not w7807 and w8187;
w8189 <= not w7733 and not w7742;
w8190 <= not w7807 and w8189;
w8191 <= not w7740 and not w8190;
w8192 <= not w8188 and not w8191;
w8193 <= w60 and not w8173;
w8194 <= not w8183 and w8193;
w8195 <= not w8192 and not w8194;
w8196 <= not w8185 and not w8195;
w8197 <= not w22 and not w8196;
w8198 <= not w7745 and w7752;
w8199 <= not w7754 and w8198;
w8200 <= not w7807 and w8199;
w8201 <= not w7745 and not w7754;
w8202 <= not w7807 and w8201;
w8203 <= not w7752 and not w8202;
w8204 <= not w8200 and not w8203;
w8205 <= w22 and not w8185;
w8206 <= not w8195 and w8205;
w8207 <= not w8204 and not w8206;
w8208 <= not w8197 and not w8207;
w8209 <= not w5 and not w8208;
w8210 <= w7764 and not w7766;
w8211 <= not w7757 and w8210;
w8212 <= not w7807 and w8211;
w8213 <= not w7757 and not w7766;
w8214 <= not w7807 and w8213;
w8215 <= not w7764 and not w8214;
w8216 <= not w8212 and not w8215;
w8217 <= w5 and not w8197;
w8218 <= not w8207 and w8217;
w8219 <= not w8216 and not w8218;
w8220 <= not w8209 and not w8219;
w8221 <= not w7769 and w7776;
w8222 <= not w7778 and w8221;
w8223 <= not w7807 and w8222;
w8224 <= not w7769 and not w7778;
w8225 <= not w7807 and w8224;
w8226 <= not w7776 and not w8225;
w8227 <= not w8223 and not w8226;
w8228 <= not w7780 and not w7787;
w8229 <= not w7807 and w8228;
w8230 <= not w7795 and not w8229;
w8231 <= not w8227 and w8230;
w8232 <= not w8220 and w8231;
w8233 <= w0 and not w8232;
w8234 <= not w8209 and w8227;
w8235 <= not w8219 and w8234;
w8236 <= not w7787 and not w7807;
w8237 <= w7780 and not w8236;
w8238 <= not w0 and not w8228;
w8239 <= not w8237 and w8238;
w8240 <= not w7783 and not w7804;
w8241 <= not w7786 and w8240;
w8242 <= not w7799 and w8241;
w8243 <= not w7795 and w8242;
w8244 <= not w7793 and w8243;
w8245 <= not w8239 and not w8244;
w8246 <= not w8235 and w8245;
w8247 <= not w8233 and w8246;
w8248 <= a(54) and not w8247;
w8249 <= not a(52) and not a(53);
w8250 <= not a(54) and w8249;
w8251 <= not w8248 and not w8250;
w8252 <= not w7807 and not w8251;
w8253 <= not w7804 and not w8250;
w8254 <= not w7799 and w8253;
w8255 <= not w7795 and w8254;
w8256 <= not w7793 and w8255;
w8257 <= not w8248 and w8256;
w8258 <= not a(54) and not w8247;
w8259 <= a(55) and not w8258;
w8260 <= w7809 and not w8247;
w8261 <= not w8259 and not w8260;
w8262 <= not w8257 and w8261;
w8263 <= not w8252 and not w8262;
w8264 <= not w7379 and not w8263;
w8265 <= w7379 and not w8252;
w8266 <= not w8262 and w8265;
w8267 <= not w7807 and not w8244;
w8268 <= not w8239 and w8267;
w8269 <= not w8235 and w8268;
w8270 <= not w8233 and w8269;
w8271 <= not w8260 and not w8270;
w8272 <= a(56) and not w8271;
w8273 <= not a(56) and not w8270;
w8274 <= not w8260 and w8273;
w8275 <= not w8272 and not w8274;
w8276 <= not w8266 and not w8275;
w8277 <= not w8264 and not w8276;
w8278 <= not w6963 and not w8277;
w8279 <= not w7812 and not w7817;
w8280 <= not w7821 and w8279;
w8281 <= not w8247 and w8280;
w8282 <= not w8247 and w8279;
w8283 <= w7821 and not w8282;
w8284 <= not w8281 and not w8283;
w8285 <= w6963 and not w8264;
w8286 <= not w8276 and w8285;
w8287 <= not w8284 and not w8286;
w8288 <= not w8278 and not w8287;
w8289 <= not w6558 and not w8288;
w8290 <= not w7826 and w7835;
w8291 <= not w7824 and w8290;
w8292 <= not w8247 and w8291;
w8293 <= not w7824 and not w7826;
w8294 <= not w8247 and w8293;
w8295 <= not w7835 and not w8294;
w8296 <= not w8292 and not w8295;
w8297 <= w6558 and not w8278;
w8298 <= not w8287 and w8297;
w8299 <= not w8296 and not w8298;
w8300 <= not w8289 and not w8299;
w8301 <= not w6166 and not w8300;
w8302 <= not w7838 and w7844;
w8303 <= not w7846 and w8302;
w8304 <= not w8247 and w8303;
w8305 <= not w7838 and not w7846;
w8306 <= not w8247 and w8305;
w8307 <= not w7844 and not w8306;
w8308 <= not w8304 and not w8307;
w8309 <= w6166 and not w8289;
w8310 <= not w8299 and w8309;
w8311 <= not w8308 and not w8310;
w8312 <= not w8301 and not w8311;
w8313 <= not w5786 and not w8312;
w8314 <= w7856 and not w7858;
w8315 <= not w7849 and w8314;
w8316 <= not w8247 and w8315;
w8317 <= not w7849 and not w7858;
w8318 <= not w8247 and w8317;
w8319 <= not w7856 and not w8318;
w8320 <= not w8316 and not w8319;
w8321 <= w5786 and not w8301;
w8322 <= not w8311 and w8321;
w8323 <= not w8320 and not w8322;
w8324 <= not w8313 and not w8323;
w8325 <= not w5418 and not w8324;
w8326 <= not w7861 and w7868;
w8327 <= not w7870 and w8326;
w8328 <= not w8247 and w8327;
w8329 <= not w7861 and not w7870;
w8330 <= not w8247 and w8329;
w8331 <= not w7868 and not w8330;
w8332 <= not w8328 and not w8331;
w8333 <= w5418 and not w8313;
w8334 <= not w8323 and w8333;
w8335 <= not w8332 and not w8334;
w8336 <= not w8325 and not w8335;
w8337 <= not w5062 and not w8336;
w8338 <= w7880 and not w7882;
w8339 <= not w7873 and w8338;
w8340 <= not w8247 and w8339;
w8341 <= not w7873 and not w7882;
w8342 <= not w8247 and w8341;
w8343 <= not w7880 and not w8342;
w8344 <= not w8340 and not w8343;
w8345 <= w5062 and not w8325;
w8346 <= not w8335 and w8345;
w8347 <= not w8344 and not w8346;
w8348 <= not w8337 and not w8347;
w8349 <= not w4718 and not w8348;
w8350 <= not w7885 and w7892;
w8351 <= not w7894 and w8350;
w8352 <= not w8247 and w8351;
w8353 <= not w7885 and not w7894;
w8354 <= not w8247 and w8353;
w8355 <= not w7892 and not w8354;
w8356 <= not w8352 and not w8355;
w8357 <= w4718 and not w8337;
w8358 <= not w8347 and w8357;
w8359 <= not w8356 and not w8358;
w8360 <= not w8349 and not w8359;
w8361 <= not w4386 and not w8360;
w8362 <= w7904 and not w7906;
w8363 <= not w7897 and w8362;
w8364 <= not w8247 and w8363;
w8365 <= not w7897 and not w7906;
w8366 <= not w8247 and w8365;
w8367 <= not w7904 and not w8366;
w8368 <= not w8364 and not w8367;
w8369 <= w4386 and not w8349;
w8370 <= not w8359 and w8369;
w8371 <= not w8368 and not w8370;
w8372 <= not w8361 and not w8371;
w8373 <= not w4066 and not w8372;
w8374 <= w4066 and not w8361;
w8375 <= not w8371 and w8374;
w8376 <= not w7909 and w7918;
w8377 <= not w7911 and w8376;
w8378 <= not w8247 and w8377;
w8379 <= not w7909 and not w7911;
w8380 <= not w8247 and w8379;
w8381 <= not w7918 and not w8380;
w8382 <= not w8378 and not w8381;
w8383 <= not w8375 and not w8382;
w8384 <= not w8373 and not w8383;
w8385 <= not w3758 and not w8384;
w8386 <= w7928 and not w7930;
w8387 <= not w7921 and w8386;
w8388 <= not w8247 and w8387;
w8389 <= not w7921 and not w7930;
w8390 <= not w8247 and w8389;
w8391 <= not w7928 and not w8390;
w8392 <= not w8388 and not w8391;
w8393 <= w3758 and not w8373;
w8394 <= not w8383 and w8393;
w8395 <= not w8392 and not w8394;
w8396 <= not w8385 and not w8395;
w8397 <= not w3462 and not w8396;
w8398 <= not w7933 and w7940;
w8399 <= not w7942 and w8398;
w8400 <= not w8247 and w8399;
w8401 <= not w7933 and not w7942;
w8402 <= not w8247 and w8401;
w8403 <= not w7940 and not w8402;
w8404 <= not w8400 and not w8403;
w8405 <= w3462 and not w8385;
w8406 <= not w8395 and w8405;
w8407 <= not w8404 and not w8406;
w8408 <= not w8397 and not w8407;
w8409 <= not w3178 and not w8408;
w8410 <= w7952 and not w7954;
w8411 <= not w7945 and w8410;
w8412 <= not w8247 and w8411;
w8413 <= not w7945 and not w7954;
w8414 <= not w8247 and w8413;
w8415 <= not w7952 and not w8414;
w8416 <= not w8412 and not w8415;
w8417 <= w3178 and not w8397;
w8418 <= not w8407 and w8417;
w8419 <= not w8416 and not w8418;
w8420 <= not w8409 and not w8419;
w8421 <= not w2906 and not w8420;
w8422 <= not w7957 and w7964;
w8423 <= not w7966 and w8422;
w8424 <= not w8247 and w8423;
w8425 <= not w7957 and not w7966;
w8426 <= not w8247 and w8425;
w8427 <= not w7964 and not w8426;
w8428 <= not w8424 and not w8427;
w8429 <= w2906 and not w8409;
w8430 <= not w8419 and w8429;
w8431 <= not w8428 and not w8430;
w8432 <= not w8421 and not w8431;
w8433 <= not w2646 and not w8432;
w8434 <= w7976 and not w7978;
w8435 <= not w7969 and w8434;
w8436 <= not w8247 and w8435;
w8437 <= not w7969 and not w7978;
w8438 <= not w8247 and w8437;
w8439 <= not w7976 and not w8438;
w8440 <= not w8436 and not w8439;
w8441 <= w2646 and not w8421;
w8442 <= not w8431 and w8441;
w8443 <= not w8440 and not w8442;
w8444 <= not w8433 and not w8443;
w8445 <= not w2398 and not w8444;
w8446 <= not w7981 and w7988;
w8447 <= not w7990 and w8446;
w8448 <= not w8247 and w8447;
w8449 <= not w7981 and not w7990;
w8450 <= not w8247 and w8449;
w8451 <= not w7988 and not w8450;
w8452 <= not w8448 and not w8451;
w8453 <= w2398 and not w8433;
w8454 <= not w8443 and w8453;
w8455 <= not w8452 and not w8454;
w8456 <= not w8445 and not w8455;
w8457 <= not w2162 and not w8456;
w8458 <= w8000 and not w8002;
w8459 <= not w7993 and w8458;
w8460 <= not w8247 and w8459;
w8461 <= not w7993 and not w8002;
w8462 <= not w8247 and w8461;
w8463 <= not w8000 and not w8462;
w8464 <= not w8460 and not w8463;
w8465 <= w2162 and not w8445;
w8466 <= not w8455 and w8465;
w8467 <= not w8464 and not w8466;
w8468 <= not w8457 and not w8467;
w8469 <= not w1938 and not w8468;
w8470 <= not w8005 and w8012;
w8471 <= not w8014 and w8470;
w8472 <= not w8247 and w8471;
w8473 <= not w8005 and not w8014;
w8474 <= not w8247 and w8473;
w8475 <= not w8012 and not w8474;
w8476 <= not w8472 and not w8475;
w8477 <= w1938 and not w8457;
w8478 <= not w8467 and w8477;
w8479 <= not w8476 and not w8478;
w8480 <= not w8469 and not w8479;
w8481 <= not w1725 and not w8480;
w8482 <= w8024 and not w8026;
w8483 <= not w8017 and w8482;
w8484 <= not w8247 and w8483;
w8485 <= not w8017 and not w8026;
w8486 <= not w8247 and w8485;
w8487 <= not w8024 and not w8486;
w8488 <= not w8484 and not w8487;
w8489 <= w1725 and not w8469;
w8490 <= not w8479 and w8489;
w8491 <= not w8488 and not w8490;
w8492 <= not w8481 and not w8491;
w8493 <= not w1525 and not w8492;
w8494 <= not w8029 and w8036;
w8495 <= not w8038 and w8494;
w8496 <= not w8247 and w8495;
w8497 <= not w8029 and not w8038;
w8498 <= not w8247 and w8497;
w8499 <= not w8036 and not w8498;
w8500 <= not w8496 and not w8499;
w8501 <= w1525 and not w8481;
w8502 <= not w8491 and w8501;
w8503 <= not w8500 and not w8502;
w8504 <= not w8493 and not w8503;
w8505 <= not w1337 and not w8504;
w8506 <= w8048 and not w8050;
w8507 <= not w8041 and w8506;
w8508 <= not w8247 and w8507;
w8509 <= not w8041 and not w8050;
w8510 <= not w8247 and w8509;
w8511 <= not w8048 and not w8510;
w8512 <= not w8508 and not w8511;
w8513 <= w1337 and not w8493;
w8514 <= not w8503 and w8513;
w8515 <= not w8512 and not w8514;
w8516 <= not w8505 and not w8515;
w8517 <= not w1161 and not w8516;
w8518 <= not w8053 and w8060;
w8519 <= not w8062 and w8518;
w8520 <= not w8247 and w8519;
w8521 <= not w8053 and not w8062;
w8522 <= not w8247 and w8521;
w8523 <= not w8060 and not w8522;
w8524 <= not w8520 and not w8523;
w8525 <= w1161 and not w8505;
w8526 <= not w8515 and w8525;
w8527 <= not w8524 and not w8526;
w8528 <= not w8517 and not w8527;
w8529 <= not w997 and not w8528;
w8530 <= w8072 and not w8074;
w8531 <= not w8065 and w8530;
w8532 <= not w8247 and w8531;
w8533 <= not w8065 and not w8074;
w8534 <= not w8247 and w8533;
w8535 <= not w8072 and not w8534;
w8536 <= not w8532 and not w8535;
w8537 <= w997 and not w8517;
w8538 <= not w8527 and w8537;
w8539 <= not w8536 and not w8538;
w8540 <= not w8529 and not w8539;
w8541 <= not w845 and not w8540;
w8542 <= not w8077 and w8084;
w8543 <= not w8086 and w8542;
w8544 <= not w8247 and w8543;
w8545 <= not w8077 and not w8086;
w8546 <= not w8247 and w8545;
w8547 <= not w8084 and not w8546;
w8548 <= not w8544 and not w8547;
w8549 <= w845 and not w8529;
w8550 <= not w8539 and w8549;
w8551 <= not w8548 and not w8550;
w8552 <= not w8541 and not w8551;
w8553 <= not w705 and not w8552;
w8554 <= w8096 and not w8098;
w8555 <= not w8089 and w8554;
w8556 <= not w8247 and w8555;
w8557 <= not w8089 and not w8098;
w8558 <= not w8247 and w8557;
w8559 <= not w8096 and not w8558;
w8560 <= not w8556 and not w8559;
w8561 <= w705 and not w8541;
w8562 <= not w8551 and w8561;
w8563 <= not w8560 and not w8562;
w8564 <= not w8553 and not w8563;
w8565 <= not w577 and not w8564;
w8566 <= not w8101 and w8108;
w8567 <= not w8110 and w8566;
w8568 <= not w8247 and w8567;
w8569 <= not w8101 and not w8110;
w8570 <= not w8247 and w8569;
w8571 <= not w8108 and not w8570;
w8572 <= not w8568 and not w8571;
w8573 <= w577 and not w8553;
w8574 <= not w8563 and w8573;
w8575 <= not w8572 and not w8574;
w8576 <= not w8565 and not w8575;
w8577 <= not w460 and not w8576;
w8578 <= w8120 and not w8122;
w8579 <= not w8113 and w8578;
w8580 <= not w8247 and w8579;
w8581 <= not w8113 and not w8122;
w8582 <= not w8247 and w8581;
w8583 <= not w8120 and not w8582;
w8584 <= not w8580 and not w8583;
w8585 <= w460 and not w8565;
w8586 <= not w8575 and w8585;
w8587 <= not w8584 and not w8586;
w8588 <= not w8577 and not w8587;
w8589 <= not w356 and not w8588;
w8590 <= not w8125 and w8132;
w8591 <= not w8134 and w8590;
w8592 <= not w8247 and w8591;
w8593 <= not w8125 and not w8134;
w8594 <= not w8247 and w8593;
w8595 <= not w8132 and not w8594;
w8596 <= not w8592 and not w8595;
w8597 <= w356 and not w8577;
w8598 <= not w8587 and w8597;
w8599 <= not w8596 and not w8598;
w8600 <= not w8589 and not w8599;
w8601 <= not w264 and not w8600;
w8602 <= w8144 and not w8146;
w8603 <= not w8137 and w8602;
w8604 <= not w8247 and w8603;
w8605 <= not w8137 and not w8146;
w8606 <= not w8247 and w8605;
w8607 <= not w8144 and not w8606;
w8608 <= not w8604 and not w8607;
w8609 <= w264 and not w8589;
w8610 <= not w8599 and w8609;
w8611 <= not w8608 and not w8610;
w8612 <= not w8601 and not w8611;
w8613 <= not w184 and not w8612;
w8614 <= not w8149 and w8156;
w8615 <= not w8158 and w8614;
w8616 <= not w8247 and w8615;
w8617 <= not w8149 and not w8158;
w8618 <= not w8247 and w8617;
w8619 <= not w8156 and not w8618;
w8620 <= not w8616 and not w8619;
w8621 <= w184 and not w8601;
w8622 <= not w8611 and w8621;
w8623 <= not w8620 and not w8622;
w8624 <= not w8613 and not w8623;
w8625 <= not w115 and not w8624;
w8626 <= w8168 and not w8170;
w8627 <= not w8161 and w8626;
w8628 <= not w8247 and w8627;
w8629 <= not w8161 and not w8170;
w8630 <= not w8247 and w8629;
w8631 <= not w8168 and not w8630;
w8632 <= not w8628 and not w8631;
w8633 <= w115 and not w8613;
w8634 <= not w8623 and w8633;
w8635 <= not w8632 and not w8634;
w8636 <= not w8625 and not w8635;
w8637 <= not w60 and not w8636;
w8638 <= not w8173 and w8180;
w8639 <= not w8182 and w8638;
w8640 <= not w8247 and w8639;
w8641 <= not w8173 and not w8182;
w8642 <= not w8247 and w8641;
w8643 <= not w8180 and not w8642;
w8644 <= not w8640 and not w8643;
w8645 <= w60 and not w8625;
w8646 <= not w8635 and w8645;
w8647 <= not w8644 and not w8646;
w8648 <= not w8637 and not w8647;
w8649 <= not w22 and not w8648;
w8650 <= w8192 and not w8194;
w8651 <= not w8185 and w8650;
w8652 <= not w8247 and w8651;
w8653 <= not w8185 and not w8194;
w8654 <= not w8247 and w8653;
w8655 <= not w8192 and not w8654;
w8656 <= not w8652 and not w8655;
w8657 <= w22 and not w8637;
w8658 <= not w8647 and w8657;
w8659 <= not w8656 and not w8658;
w8660 <= not w8649 and not w8659;
w8661 <= not w5 and not w8660;
w8662 <= not w8197 and w8204;
w8663 <= not w8206 and w8662;
w8664 <= not w8247 and w8663;
w8665 <= not w8197 and not w8206;
w8666 <= not w8247 and w8665;
w8667 <= not w8204 and not w8666;
w8668 <= not w8664 and not w8667;
w8669 <= w5 and not w8649;
w8670 <= not w8659 and w8669;
w8671 <= not w8668 and not w8670;
w8672 <= not w8661 and not w8671;
w8673 <= w8216 and not w8218;
w8674 <= not w8209 and w8673;
w8675 <= not w8247 and w8674;
w8676 <= not w8209 and not w8218;
w8677 <= not w8247 and w8676;
w8678 <= not w8216 and not w8677;
w8679 <= not w8675 and not w8678;
w8680 <= not w8220 and not w8227;
w8681 <= not w8247 and w8680;
w8682 <= not w8235 and not w8681;
w8683 <= not w8679 and w8682;
w8684 <= not w8672 and w8683;
w8685 <= w0 and not w8684;
w8686 <= not w8661 and w8679;
w8687 <= not w8671 and w8686;
w8688 <= not w8227 and not w8247;
w8689 <= w8220 and not w8688;
w8690 <= not w0 and not w8680;
w8691 <= not w8689 and w8690;
w8692 <= not w8223 and not w8244;
w8693 <= not w8226 and w8692;
w8694 <= not w8239 and w8693;
w8695 <= not w8235 and w8694;
w8696 <= not w8233 and w8695;
w8697 <= not w8691 and not w8696;
w8698 <= not w8687 and w8697;
w8699 <= not w8685 and w8698;
w8700 <= a(52) and not w8699;
w8701 <= not a(50) and not a(51);
w8702 <= not a(52) and w8701;
w8703 <= not w8700 and not w8702;
w8704 <= not w8247 and not w8703;
w8705 <= not w8244 and not w8702;
w8706 <= not w8239 and w8705;
w8707 <= not w8235 and w8706;
w8708 <= not w8233 and w8707;
w8709 <= not w8700 and w8708;
w8710 <= not a(52) and not w8699;
w8711 <= a(53) and not w8710;
w8712 <= w8249 and not w8699;
w8713 <= not w8711 and not w8712;
w8714 <= not w8709 and w8713;
w8715 <= not w8704 and not w8714;
w8716 <= not w7807 and not w8715;
w8717 <= w7807 and not w8704;
w8718 <= not w8714 and w8717;
w8719 <= not w8247 and not w8696;
w8720 <= not w8691 and w8719;
w8721 <= not w8687 and w8720;
w8722 <= not w8685 and w8721;
w8723 <= not w8712 and not w8722;
w8724 <= a(54) and not w8723;
w8725 <= not a(54) and not w8722;
w8726 <= not w8712 and w8725;
w8727 <= not w8724 and not w8726;
w8728 <= not w8718 and not w8727;
w8729 <= not w8716 and not w8728;
w8730 <= not w7379 and not w8729;
w8731 <= not w8252 and not w8257;
w8732 <= not w8261 and w8731;
w8733 <= not w8699 and w8732;
w8734 <= not w8699 and w8731;
w8735 <= w8261 and not w8734;
w8736 <= not w8733 and not w8735;
w8737 <= w7379 and not w8716;
w8738 <= not w8728 and w8737;
w8739 <= not w8736 and not w8738;
w8740 <= not w8730 and not w8739;
w8741 <= not w6963 and not w8740;
w8742 <= not w8266 and w8275;
w8743 <= not w8264 and w8742;
w8744 <= not w8699 and w8743;
w8745 <= not w8264 and not w8266;
w8746 <= not w8699 and w8745;
w8747 <= not w8275 and not w8746;
w8748 <= not w8744 and not w8747;
w8749 <= w6963 and not w8730;
w8750 <= not w8739 and w8749;
w8751 <= not w8748 and not w8750;
w8752 <= not w8741 and not w8751;
w8753 <= not w6558 and not w8752;
w8754 <= not w8278 and w8284;
w8755 <= not w8286 and w8754;
w8756 <= not w8699 and w8755;
w8757 <= not w8278 and not w8286;
w8758 <= not w8699 and w8757;
w8759 <= not w8284 and not w8758;
w8760 <= not w8756 and not w8759;
w8761 <= w6558 and not w8741;
w8762 <= not w8751 and w8761;
w8763 <= not w8760 and not w8762;
w8764 <= not w8753 and not w8763;
w8765 <= not w6166 and not w8764;
w8766 <= w8296 and not w8298;
w8767 <= not w8289 and w8766;
w8768 <= not w8699 and w8767;
w8769 <= not w8289 and not w8298;
w8770 <= not w8699 and w8769;
w8771 <= not w8296 and not w8770;
w8772 <= not w8768 and not w8771;
w8773 <= w6166 and not w8753;
w8774 <= not w8763 and w8773;
w8775 <= not w8772 and not w8774;
w8776 <= not w8765 and not w8775;
w8777 <= not w5786 and not w8776;
w8778 <= not w8301 and w8308;
w8779 <= not w8310 and w8778;
w8780 <= not w8699 and w8779;
w8781 <= not w8301 and not w8310;
w8782 <= not w8699 and w8781;
w8783 <= not w8308 and not w8782;
w8784 <= not w8780 and not w8783;
w8785 <= w5786 and not w8765;
w8786 <= not w8775 and w8785;
w8787 <= not w8784 and not w8786;
w8788 <= not w8777 and not w8787;
w8789 <= not w5418 and not w8788;
w8790 <= w8320 and not w8322;
w8791 <= not w8313 and w8790;
w8792 <= not w8699 and w8791;
w8793 <= not w8313 and not w8322;
w8794 <= not w8699 and w8793;
w8795 <= not w8320 and not w8794;
w8796 <= not w8792 and not w8795;
w8797 <= w5418 and not w8777;
w8798 <= not w8787 and w8797;
w8799 <= not w8796 and not w8798;
w8800 <= not w8789 and not w8799;
w8801 <= not w5062 and not w8800;
w8802 <= not w8325 and w8332;
w8803 <= not w8334 and w8802;
w8804 <= not w8699 and w8803;
w8805 <= not w8325 and not w8334;
w8806 <= not w8699 and w8805;
w8807 <= not w8332 and not w8806;
w8808 <= not w8804 and not w8807;
w8809 <= w5062 and not w8789;
w8810 <= not w8799 and w8809;
w8811 <= not w8808 and not w8810;
w8812 <= not w8801 and not w8811;
w8813 <= not w4718 and not w8812;
w8814 <= w8344 and not w8346;
w8815 <= not w8337 and w8814;
w8816 <= not w8699 and w8815;
w8817 <= not w8337 and not w8346;
w8818 <= not w8699 and w8817;
w8819 <= not w8344 and not w8818;
w8820 <= not w8816 and not w8819;
w8821 <= w4718 and not w8801;
w8822 <= not w8811 and w8821;
w8823 <= not w8820 and not w8822;
w8824 <= not w8813 and not w8823;
w8825 <= not w4386 and not w8824;
w8826 <= not w8349 and w8356;
w8827 <= not w8358 and w8826;
w8828 <= not w8699 and w8827;
w8829 <= not w8349 and not w8358;
w8830 <= not w8699 and w8829;
w8831 <= not w8356 and not w8830;
w8832 <= not w8828 and not w8831;
w8833 <= w4386 and not w8813;
w8834 <= not w8823 and w8833;
w8835 <= not w8832 and not w8834;
w8836 <= not w8825 and not w8835;
w8837 <= not w4066 and not w8836;
w8838 <= w8368 and not w8370;
w8839 <= not w8361 and w8838;
w8840 <= not w8699 and w8839;
w8841 <= not w8361 and not w8370;
w8842 <= not w8699 and w8841;
w8843 <= not w8368 and not w8842;
w8844 <= not w8840 and not w8843;
w8845 <= w4066 and not w8825;
w8846 <= not w8835 and w8845;
w8847 <= not w8844 and not w8846;
w8848 <= not w8837 and not w8847;
w8849 <= not w3758 and not w8848;
w8850 <= w3758 and not w8837;
w8851 <= not w8847 and w8850;
w8852 <= not w8373 and w8382;
w8853 <= not w8375 and w8852;
w8854 <= not w8699 and w8853;
w8855 <= not w8373 and not w8375;
w8856 <= not w8699 and w8855;
w8857 <= not w8382 and not w8856;
w8858 <= not w8854 and not w8857;
w8859 <= not w8851 and not w8858;
w8860 <= not w8849 and not w8859;
w8861 <= not w3462 and not w8860;
w8862 <= w8392 and not w8394;
w8863 <= not w8385 and w8862;
w8864 <= not w8699 and w8863;
w8865 <= not w8385 and not w8394;
w8866 <= not w8699 and w8865;
w8867 <= not w8392 and not w8866;
w8868 <= not w8864 and not w8867;
w8869 <= w3462 and not w8849;
w8870 <= not w8859 and w8869;
w8871 <= not w8868 and not w8870;
w8872 <= not w8861 and not w8871;
w8873 <= not w3178 and not w8872;
w8874 <= not w8397 and w8404;
w8875 <= not w8406 and w8874;
w8876 <= not w8699 and w8875;
w8877 <= not w8397 and not w8406;
w8878 <= not w8699 and w8877;
w8879 <= not w8404 and not w8878;
w8880 <= not w8876 and not w8879;
w8881 <= w3178 and not w8861;
w8882 <= not w8871 and w8881;
w8883 <= not w8880 and not w8882;
w8884 <= not w8873 and not w8883;
w8885 <= not w2906 and not w8884;
w8886 <= w8416 and not w8418;
w8887 <= not w8409 and w8886;
w8888 <= not w8699 and w8887;
w8889 <= not w8409 and not w8418;
w8890 <= not w8699 and w8889;
w8891 <= not w8416 and not w8890;
w8892 <= not w8888 and not w8891;
w8893 <= w2906 and not w8873;
w8894 <= not w8883 and w8893;
w8895 <= not w8892 and not w8894;
w8896 <= not w8885 and not w8895;
w8897 <= not w2646 and not w8896;
w8898 <= not w8421 and w8428;
w8899 <= not w8430 and w8898;
w8900 <= not w8699 and w8899;
w8901 <= not w8421 and not w8430;
w8902 <= not w8699 and w8901;
w8903 <= not w8428 and not w8902;
w8904 <= not w8900 and not w8903;
w8905 <= w2646 and not w8885;
w8906 <= not w8895 and w8905;
w8907 <= not w8904 and not w8906;
w8908 <= not w8897 and not w8907;
w8909 <= not w2398 and not w8908;
w8910 <= w8440 and not w8442;
w8911 <= not w8433 and w8910;
w8912 <= not w8699 and w8911;
w8913 <= not w8433 and not w8442;
w8914 <= not w8699 and w8913;
w8915 <= not w8440 and not w8914;
w8916 <= not w8912 and not w8915;
w8917 <= w2398 and not w8897;
w8918 <= not w8907 and w8917;
w8919 <= not w8916 and not w8918;
w8920 <= not w8909 and not w8919;
w8921 <= not w2162 and not w8920;
w8922 <= not w8445 and w8452;
w8923 <= not w8454 and w8922;
w8924 <= not w8699 and w8923;
w8925 <= not w8445 and not w8454;
w8926 <= not w8699 and w8925;
w8927 <= not w8452 and not w8926;
w8928 <= not w8924 and not w8927;
w8929 <= w2162 and not w8909;
w8930 <= not w8919 and w8929;
w8931 <= not w8928 and not w8930;
w8932 <= not w8921 and not w8931;
w8933 <= not w1938 and not w8932;
w8934 <= w8464 and not w8466;
w8935 <= not w8457 and w8934;
w8936 <= not w8699 and w8935;
w8937 <= not w8457 and not w8466;
w8938 <= not w8699 and w8937;
w8939 <= not w8464 and not w8938;
w8940 <= not w8936 and not w8939;
w8941 <= w1938 and not w8921;
w8942 <= not w8931 and w8941;
w8943 <= not w8940 and not w8942;
w8944 <= not w8933 and not w8943;
w8945 <= not w1725 and not w8944;
w8946 <= not w8469 and w8476;
w8947 <= not w8478 and w8946;
w8948 <= not w8699 and w8947;
w8949 <= not w8469 and not w8478;
w8950 <= not w8699 and w8949;
w8951 <= not w8476 and not w8950;
w8952 <= not w8948 and not w8951;
w8953 <= w1725 and not w8933;
w8954 <= not w8943 and w8953;
w8955 <= not w8952 and not w8954;
w8956 <= not w8945 and not w8955;
w8957 <= not w1525 and not w8956;
w8958 <= w8488 and not w8490;
w8959 <= not w8481 and w8958;
w8960 <= not w8699 and w8959;
w8961 <= not w8481 and not w8490;
w8962 <= not w8699 and w8961;
w8963 <= not w8488 and not w8962;
w8964 <= not w8960 and not w8963;
w8965 <= w1525 and not w8945;
w8966 <= not w8955 and w8965;
w8967 <= not w8964 and not w8966;
w8968 <= not w8957 and not w8967;
w8969 <= not w1337 and not w8968;
w8970 <= not w8493 and w8500;
w8971 <= not w8502 and w8970;
w8972 <= not w8699 and w8971;
w8973 <= not w8493 and not w8502;
w8974 <= not w8699 and w8973;
w8975 <= not w8500 and not w8974;
w8976 <= not w8972 and not w8975;
w8977 <= w1337 and not w8957;
w8978 <= not w8967 and w8977;
w8979 <= not w8976 and not w8978;
w8980 <= not w8969 and not w8979;
w8981 <= not w1161 and not w8980;
w8982 <= w8512 and not w8514;
w8983 <= not w8505 and w8982;
w8984 <= not w8699 and w8983;
w8985 <= not w8505 and not w8514;
w8986 <= not w8699 and w8985;
w8987 <= not w8512 and not w8986;
w8988 <= not w8984 and not w8987;
w8989 <= w1161 and not w8969;
w8990 <= not w8979 and w8989;
w8991 <= not w8988 and not w8990;
w8992 <= not w8981 and not w8991;
w8993 <= not w997 and not w8992;
w8994 <= not w8517 and w8524;
w8995 <= not w8526 and w8994;
w8996 <= not w8699 and w8995;
w8997 <= not w8517 and not w8526;
w8998 <= not w8699 and w8997;
w8999 <= not w8524 and not w8998;
w9000 <= not w8996 and not w8999;
w9001 <= w997 and not w8981;
w9002 <= not w8991 and w9001;
w9003 <= not w9000 and not w9002;
w9004 <= not w8993 and not w9003;
w9005 <= not w845 and not w9004;
w9006 <= w8536 and not w8538;
w9007 <= not w8529 and w9006;
w9008 <= not w8699 and w9007;
w9009 <= not w8529 and not w8538;
w9010 <= not w8699 and w9009;
w9011 <= not w8536 and not w9010;
w9012 <= not w9008 and not w9011;
w9013 <= w845 and not w8993;
w9014 <= not w9003 and w9013;
w9015 <= not w9012 and not w9014;
w9016 <= not w9005 and not w9015;
w9017 <= not w705 and not w9016;
w9018 <= not w8541 and w8548;
w9019 <= not w8550 and w9018;
w9020 <= not w8699 and w9019;
w9021 <= not w8541 and not w8550;
w9022 <= not w8699 and w9021;
w9023 <= not w8548 and not w9022;
w9024 <= not w9020 and not w9023;
w9025 <= w705 and not w9005;
w9026 <= not w9015 and w9025;
w9027 <= not w9024 and not w9026;
w9028 <= not w9017 and not w9027;
w9029 <= not w577 and not w9028;
w9030 <= w8560 and not w8562;
w9031 <= not w8553 and w9030;
w9032 <= not w8699 and w9031;
w9033 <= not w8553 and not w8562;
w9034 <= not w8699 and w9033;
w9035 <= not w8560 and not w9034;
w9036 <= not w9032 and not w9035;
w9037 <= w577 and not w9017;
w9038 <= not w9027 and w9037;
w9039 <= not w9036 and not w9038;
w9040 <= not w9029 and not w9039;
w9041 <= not w460 and not w9040;
w9042 <= not w8565 and w8572;
w9043 <= not w8574 and w9042;
w9044 <= not w8699 and w9043;
w9045 <= not w8565 and not w8574;
w9046 <= not w8699 and w9045;
w9047 <= not w8572 and not w9046;
w9048 <= not w9044 and not w9047;
w9049 <= w460 and not w9029;
w9050 <= not w9039 and w9049;
w9051 <= not w9048 and not w9050;
w9052 <= not w9041 and not w9051;
w9053 <= not w356 and not w9052;
w9054 <= w8584 and not w8586;
w9055 <= not w8577 and w9054;
w9056 <= not w8699 and w9055;
w9057 <= not w8577 and not w8586;
w9058 <= not w8699 and w9057;
w9059 <= not w8584 and not w9058;
w9060 <= not w9056 and not w9059;
w9061 <= w356 and not w9041;
w9062 <= not w9051 and w9061;
w9063 <= not w9060 and not w9062;
w9064 <= not w9053 and not w9063;
w9065 <= not w264 and not w9064;
w9066 <= not w8589 and w8596;
w9067 <= not w8598 and w9066;
w9068 <= not w8699 and w9067;
w9069 <= not w8589 and not w8598;
w9070 <= not w8699 and w9069;
w9071 <= not w8596 and not w9070;
w9072 <= not w9068 and not w9071;
w9073 <= w264 and not w9053;
w9074 <= not w9063 and w9073;
w9075 <= not w9072 and not w9074;
w9076 <= not w9065 and not w9075;
w9077 <= not w184 and not w9076;
w9078 <= w8608 and not w8610;
w9079 <= not w8601 and w9078;
w9080 <= not w8699 and w9079;
w9081 <= not w8601 and not w8610;
w9082 <= not w8699 and w9081;
w9083 <= not w8608 and not w9082;
w9084 <= not w9080 and not w9083;
w9085 <= w184 and not w9065;
w9086 <= not w9075 and w9085;
w9087 <= not w9084 and not w9086;
w9088 <= not w9077 and not w9087;
w9089 <= not w115 and not w9088;
w9090 <= not w8613 and w8620;
w9091 <= not w8622 and w9090;
w9092 <= not w8699 and w9091;
w9093 <= not w8613 and not w8622;
w9094 <= not w8699 and w9093;
w9095 <= not w8620 and not w9094;
w9096 <= not w9092 and not w9095;
w9097 <= w115 and not w9077;
w9098 <= not w9087 and w9097;
w9099 <= not w9096 and not w9098;
w9100 <= not w9089 and not w9099;
w9101 <= not w60 and not w9100;
w9102 <= w8632 and not w8634;
w9103 <= not w8625 and w9102;
w9104 <= not w8699 and w9103;
w9105 <= not w8625 and not w8634;
w9106 <= not w8699 and w9105;
w9107 <= not w8632 and not w9106;
w9108 <= not w9104 and not w9107;
w9109 <= w60 and not w9089;
w9110 <= not w9099 and w9109;
w9111 <= not w9108 and not w9110;
w9112 <= not w9101 and not w9111;
w9113 <= not w22 and not w9112;
w9114 <= not w8637 and w8644;
w9115 <= not w8646 and w9114;
w9116 <= not w8699 and w9115;
w9117 <= not w8637 and not w8646;
w9118 <= not w8699 and w9117;
w9119 <= not w8644 and not w9118;
w9120 <= not w9116 and not w9119;
w9121 <= w22 and not w9101;
w9122 <= not w9111 and w9121;
w9123 <= not w9120 and not w9122;
w9124 <= not w9113 and not w9123;
w9125 <= not w5 and not w9124;
w9126 <= w8656 and not w8658;
w9127 <= not w8649 and w9126;
w9128 <= not w8699 and w9127;
w9129 <= not w8649 and not w8658;
w9130 <= not w8699 and w9129;
w9131 <= not w8656 and not w9130;
w9132 <= not w9128 and not w9131;
w9133 <= w5 and not w9113;
w9134 <= not w9123 and w9133;
w9135 <= not w9132 and not w9134;
w9136 <= not w9125 and not w9135;
w9137 <= not w8661 and w8668;
w9138 <= not w8670 and w9137;
w9139 <= not w8699 and w9138;
w9140 <= not w8661 and not w8670;
w9141 <= not w8699 and w9140;
w9142 <= not w8668 and not w9141;
w9143 <= not w9139 and not w9142;
w9144 <= not w8672 and not w8679;
w9145 <= not w8699 and w9144;
w9146 <= not w8687 and not w9145;
w9147 <= not w9143 and w9146;
w9148 <= not w9136 and w9147;
w9149 <= w0 and not w9148;
w9150 <= not w9125 and w9143;
w9151 <= not w9135 and w9150;
w9152 <= not w8679 and not w8699;
w9153 <= w8672 and not w9152;
w9154 <= not w0 and not w9144;
w9155 <= not w9153 and w9154;
w9156 <= not w8675 and not w8696;
w9157 <= not w8678 and w9156;
w9158 <= not w8691 and w9157;
w9159 <= not w8687 and w9158;
w9160 <= not w8685 and w9159;
w9161 <= not w9155 and not w9160;
w9162 <= not w9151 and w9161;
w9163 <= not w9149 and w9162;
w9164 <= a(50) and not w9163;
w9165 <= not a(48) and not a(49);
w9166 <= not a(50) and w9165;
w9167 <= not w9164 and not w9166;
w9168 <= not w8699 and not w9167;
w9169 <= not w8696 and not w9166;
w9170 <= not w8691 and w9169;
w9171 <= not w8687 and w9170;
w9172 <= not w8685 and w9171;
w9173 <= not w9164 and w9172;
w9174 <= not a(50) and not w9163;
w9175 <= a(51) and not w9174;
w9176 <= w8701 and not w9163;
w9177 <= not w9175 and not w9176;
w9178 <= not w9173 and w9177;
w9179 <= not w9168 and not w9178;
w9180 <= not w8247 and not w9179;
w9181 <= w8247 and not w9168;
w9182 <= not w9178 and w9181;
w9183 <= not w8699 and not w9160;
w9184 <= not w9155 and w9183;
w9185 <= not w9151 and w9184;
w9186 <= not w9149 and w9185;
w9187 <= not w9176 and not w9186;
w9188 <= a(52) and not w9187;
w9189 <= not a(52) and not w9186;
w9190 <= not w9176 and w9189;
w9191 <= not w9188 and not w9190;
w9192 <= not w9182 and not w9191;
w9193 <= not w9180 and not w9192;
w9194 <= not w7807 and not w9193;
w9195 <= not w8704 and not w8709;
w9196 <= not w8713 and w9195;
w9197 <= not w9163 and w9196;
w9198 <= not w9163 and w9195;
w9199 <= w8713 and not w9198;
w9200 <= not w9197 and not w9199;
w9201 <= w7807 and not w9180;
w9202 <= not w9192 and w9201;
w9203 <= not w9200 and not w9202;
w9204 <= not w9194 and not w9203;
w9205 <= not w7379 and not w9204;
w9206 <= not w8718 and w8727;
w9207 <= not w8716 and w9206;
w9208 <= not w9163 and w9207;
w9209 <= not w8716 and not w8718;
w9210 <= not w9163 and w9209;
w9211 <= not w8727 and not w9210;
w9212 <= not w9208 and not w9211;
w9213 <= w7379 and not w9194;
w9214 <= not w9203 and w9213;
w9215 <= not w9212 and not w9214;
w9216 <= not w9205 and not w9215;
w9217 <= not w6963 and not w9216;
w9218 <= not w8730 and w8736;
w9219 <= not w8738 and w9218;
w9220 <= not w9163 and w9219;
w9221 <= not w8730 and not w8738;
w9222 <= not w9163 and w9221;
w9223 <= not w8736 and not w9222;
w9224 <= not w9220 and not w9223;
w9225 <= w6963 and not w9205;
w9226 <= not w9215 and w9225;
w9227 <= not w9224 and not w9226;
w9228 <= not w9217 and not w9227;
w9229 <= not w6558 and not w9228;
w9230 <= w8748 and not w8750;
w9231 <= not w8741 and w9230;
w9232 <= not w9163 and w9231;
w9233 <= not w8741 and not w8750;
w9234 <= not w9163 and w9233;
w9235 <= not w8748 and not w9234;
w9236 <= not w9232 and not w9235;
w9237 <= w6558 and not w9217;
w9238 <= not w9227 and w9237;
w9239 <= not w9236 and not w9238;
w9240 <= not w9229 and not w9239;
w9241 <= not w6166 and not w9240;
w9242 <= not w8753 and w8760;
w9243 <= not w8762 and w9242;
w9244 <= not w9163 and w9243;
w9245 <= not w8753 and not w8762;
w9246 <= not w9163 and w9245;
w9247 <= not w8760 and not w9246;
w9248 <= not w9244 and not w9247;
w9249 <= w6166 and not w9229;
w9250 <= not w9239 and w9249;
w9251 <= not w9248 and not w9250;
w9252 <= not w9241 and not w9251;
w9253 <= not w5786 and not w9252;
w9254 <= w8772 and not w8774;
w9255 <= not w8765 and w9254;
w9256 <= not w9163 and w9255;
w9257 <= not w8765 and not w8774;
w9258 <= not w9163 and w9257;
w9259 <= not w8772 and not w9258;
w9260 <= not w9256 and not w9259;
w9261 <= w5786 and not w9241;
w9262 <= not w9251 and w9261;
w9263 <= not w9260 and not w9262;
w9264 <= not w9253 and not w9263;
w9265 <= not w5418 and not w9264;
w9266 <= not w8777 and w8784;
w9267 <= not w8786 and w9266;
w9268 <= not w9163 and w9267;
w9269 <= not w8777 and not w8786;
w9270 <= not w9163 and w9269;
w9271 <= not w8784 and not w9270;
w9272 <= not w9268 and not w9271;
w9273 <= w5418 and not w9253;
w9274 <= not w9263 and w9273;
w9275 <= not w9272 and not w9274;
w9276 <= not w9265 and not w9275;
w9277 <= not w5062 and not w9276;
w9278 <= w8796 and not w8798;
w9279 <= not w8789 and w9278;
w9280 <= not w9163 and w9279;
w9281 <= not w8789 and not w8798;
w9282 <= not w9163 and w9281;
w9283 <= not w8796 and not w9282;
w9284 <= not w9280 and not w9283;
w9285 <= w5062 and not w9265;
w9286 <= not w9275 and w9285;
w9287 <= not w9284 and not w9286;
w9288 <= not w9277 and not w9287;
w9289 <= not w4718 and not w9288;
w9290 <= not w8801 and w8808;
w9291 <= not w8810 and w9290;
w9292 <= not w9163 and w9291;
w9293 <= not w8801 and not w8810;
w9294 <= not w9163 and w9293;
w9295 <= not w8808 and not w9294;
w9296 <= not w9292 and not w9295;
w9297 <= w4718 and not w9277;
w9298 <= not w9287 and w9297;
w9299 <= not w9296 and not w9298;
w9300 <= not w9289 and not w9299;
w9301 <= not w4386 and not w9300;
w9302 <= w8820 and not w8822;
w9303 <= not w8813 and w9302;
w9304 <= not w9163 and w9303;
w9305 <= not w8813 and not w8822;
w9306 <= not w9163 and w9305;
w9307 <= not w8820 and not w9306;
w9308 <= not w9304 and not w9307;
w9309 <= w4386 and not w9289;
w9310 <= not w9299 and w9309;
w9311 <= not w9308 and not w9310;
w9312 <= not w9301 and not w9311;
w9313 <= not w4066 and not w9312;
w9314 <= not w8825 and w8832;
w9315 <= not w8834 and w9314;
w9316 <= not w9163 and w9315;
w9317 <= not w8825 and not w8834;
w9318 <= not w9163 and w9317;
w9319 <= not w8832 and not w9318;
w9320 <= not w9316 and not w9319;
w9321 <= w4066 and not w9301;
w9322 <= not w9311 and w9321;
w9323 <= not w9320 and not w9322;
w9324 <= not w9313 and not w9323;
w9325 <= not w3758 and not w9324;
w9326 <= w8844 and not w8846;
w9327 <= not w8837 and w9326;
w9328 <= not w9163 and w9327;
w9329 <= not w8837 and not w8846;
w9330 <= not w9163 and w9329;
w9331 <= not w8844 and not w9330;
w9332 <= not w9328 and not w9331;
w9333 <= w3758 and not w9313;
w9334 <= not w9323 and w9333;
w9335 <= not w9332 and not w9334;
w9336 <= not w9325 and not w9335;
w9337 <= not w3462 and not w9336;
w9338 <= w3462 and not w9325;
w9339 <= not w9335 and w9338;
w9340 <= not w8849 and w8858;
w9341 <= not w8851 and w9340;
w9342 <= not w9163 and w9341;
w9343 <= not w8849 and not w8851;
w9344 <= not w9163 and w9343;
w9345 <= not w8858 and not w9344;
w9346 <= not w9342 and not w9345;
w9347 <= not w9339 and not w9346;
w9348 <= not w9337 and not w9347;
w9349 <= not w3178 and not w9348;
w9350 <= w8868 and not w8870;
w9351 <= not w8861 and w9350;
w9352 <= not w9163 and w9351;
w9353 <= not w8861 and not w8870;
w9354 <= not w9163 and w9353;
w9355 <= not w8868 and not w9354;
w9356 <= not w9352 and not w9355;
w9357 <= w3178 and not w9337;
w9358 <= not w9347 and w9357;
w9359 <= not w9356 and not w9358;
w9360 <= not w9349 and not w9359;
w9361 <= not w2906 and not w9360;
w9362 <= not w8873 and w8880;
w9363 <= not w8882 and w9362;
w9364 <= not w9163 and w9363;
w9365 <= not w8873 and not w8882;
w9366 <= not w9163 and w9365;
w9367 <= not w8880 and not w9366;
w9368 <= not w9364 and not w9367;
w9369 <= w2906 and not w9349;
w9370 <= not w9359 and w9369;
w9371 <= not w9368 and not w9370;
w9372 <= not w9361 and not w9371;
w9373 <= not w2646 and not w9372;
w9374 <= w8892 and not w8894;
w9375 <= not w8885 and w9374;
w9376 <= not w9163 and w9375;
w9377 <= not w8885 and not w8894;
w9378 <= not w9163 and w9377;
w9379 <= not w8892 and not w9378;
w9380 <= not w9376 and not w9379;
w9381 <= w2646 and not w9361;
w9382 <= not w9371 and w9381;
w9383 <= not w9380 and not w9382;
w9384 <= not w9373 and not w9383;
w9385 <= not w2398 and not w9384;
w9386 <= not w8897 and w8904;
w9387 <= not w8906 and w9386;
w9388 <= not w9163 and w9387;
w9389 <= not w8897 and not w8906;
w9390 <= not w9163 and w9389;
w9391 <= not w8904 and not w9390;
w9392 <= not w9388 and not w9391;
w9393 <= w2398 and not w9373;
w9394 <= not w9383 and w9393;
w9395 <= not w9392 and not w9394;
w9396 <= not w9385 and not w9395;
w9397 <= not w2162 and not w9396;
w9398 <= w8916 and not w8918;
w9399 <= not w8909 and w9398;
w9400 <= not w9163 and w9399;
w9401 <= not w8909 and not w8918;
w9402 <= not w9163 and w9401;
w9403 <= not w8916 and not w9402;
w9404 <= not w9400 and not w9403;
w9405 <= w2162 and not w9385;
w9406 <= not w9395 and w9405;
w9407 <= not w9404 and not w9406;
w9408 <= not w9397 and not w9407;
w9409 <= not w1938 and not w9408;
w9410 <= not w8921 and w8928;
w9411 <= not w8930 and w9410;
w9412 <= not w9163 and w9411;
w9413 <= not w8921 and not w8930;
w9414 <= not w9163 and w9413;
w9415 <= not w8928 and not w9414;
w9416 <= not w9412 and not w9415;
w9417 <= w1938 and not w9397;
w9418 <= not w9407 and w9417;
w9419 <= not w9416 and not w9418;
w9420 <= not w9409 and not w9419;
w9421 <= not w1725 and not w9420;
w9422 <= w8940 and not w8942;
w9423 <= not w8933 and w9422;
w9424 <= not w9163 and w9423;
w9425 <= not w8933 and not w8942;
w9426 <= not w9163 and w9425;
w9427 <= not w8940 and not w9426;
w9428 <= not w9424 and not w9427;
w9429 <= w1725 and not w9409;
w9430 <= not w9419 and w9429;
w9431 <= not w9428 and not w9430;
w9432 <= not w9421 and not w9431;
w9433 <= not w1525 and not w9432;
w9434 <= not w8945 and w8952;
w9435 <= not w8954 and w9434;
w9436 <= not w9163 and w9435;
w9437 <= not w8945 and not w8954;
w9438 <= not w9163 and w9437;
w9439 <= not w8952 and not w9438;
w9440 <= not w9436 and not w9439;
w9441 <= w1525 and not w9421;
w9442 <= not w9431 and w9441;
w9443 <= not w9440 and not w9442;
w9444 <= not w9433 and not w9443;
w9445 <= not w1337 and not w9444;
w9446 <= w8964 and not w8966;
w9447 <= not w8957 and w9446;
w9448 <= not w9163 and w9447;
w9449 <= not w8957 and not w8966;
w9450 <= not w9163 and w9449;
w9451 <= not w8964 and not w9450;
w9452 <= not w9448 and not w9451;
w9453 <= w1337 and not w9433;
w9454 <= not w9443 and w9453;
w9455 <= not w9452 and not w9454;
w9456 <= not w9445 and not w9455;
w9457 <= not w1161 and not w9456;
w9458 <= not w8969 and w8976;
w9459 <= not w8978 and w9458;
w9460 <= not w9163 and w9459;
w9461 <= not w8969 and not w8978;
w9462 <= not w9163 and w9461;
w9463 <= not w8976 and not w9462;
w9464 <= not w9460 and not w9463;
w9465 <= w1161 and not w9445;
w9466 <= not w9455 and w9465;
w9467 <= not w9464 and not w9466;
w9468 <= not w9457 and not w9467;
w9469 <= not w997 and not w9468;
w9470 <= w8988 and not w8990;
w9471 <= not w8981 and w9470;
w9472 <= not w9163 and w9471;
w9473 <= not w8981 and not w8990;
w9474 <= not w9163 and w9473;
w9475 <= not w8988 and not w9474;
w9476 <= not w9472 and not w9475;
w9477 <= w997 and not w9457;
w9478 <= not w9467 and w9477;
w9479 <= not w9476 and not w9478;
w9480 <= not w9469 and not w9479;
w9481 <= not w845 and not w9480;
w9482 <= not w8993 and w9000;
w9483 <= not w9002 and w9482;
w9484 <= not w9163 and w9483;
w9485 <= not w8993 and not w9002;
w9486 <= not w9163 and w9485;
w9487 <= not w9000 and not w9486;
w9488 <= not w9484 and not w9487;
w9489 <= w845 and not w9469;
w9490 <= not w9479 and w9489;
w9491 <= not w9488 and not w9490;
w9492 <= not w9481 and not w9491;
w9493 <= not w705 and not w9492;
w9494 <= w9012 and not w9014;
w9495 <= not w9005 and w9494;
w9496 <= not w9163 and w9495;
w9497 <= not w9005 and not w9014;
w9498 <= not w9163 and w9497;
w9499 <= not w9012 and not w9498;
w9500 <= not w9496 and not w9499;
w9501 <= w705 and not w9481;
w9502 <= not w9491 and w9501;
w9503 <= not w9500 and not w9502;
w9504 <= not w9493 and not w9503;
w9505 <= not w577 and not w9504;
w9506 <= not w9017 and w9024;
w9507 <= not w9026 and w9506;
w9508 <= not w9163 and w9507;
w9509 <= not w9017 and not w9026;
w9510 <= not w9163 and w9509;
w9511 <= not w9024 and not w9510;
w9512 <= not w9508 and not w9511;
w9513 <= w577 and not w9493;
w9514 <= not w9503 and w9513;
w9515 <= not w9512 and not w9514;
w9516 <= not w9505 and not w9515;
w9517 <= not w460 and not w9516;
w9518 <= w9036 and not w9038;
w9519 <= not w9029 and w9518;
w9520 <= not w9163 and w9519;
w9521 <= not w9029 and not w9038;
w9522 <= not w9163 and w9521;
w9523 <= not w9036 and not w9522;
w9524 <= not w9520 and not w9523;
w9525 <= w460 and not w9505;
w9526 <= not w9515 and w9525;
w9527 <= not w9524 and not w9526;
w9528 <= not w9517 and not w9527;
w9529 <= not w356 and not w9528;
w9530 <= not w9041 and w9048;
w9531 <= not w9050 and w9530;
w9532 <= not w9163 and w9531;
w9533 <= not w9041 and not w9050;
w9534 <= not w9163 and w9533;
w9535 <= not w9048 and not w9534;
w9536 <= not w9532 and not w9535;
w9537 <= w356 and not w9517;
w9538 <= not w9527 and w9537;
w9539 <= not w9536 and not w9538;
w9540 <= not w9529 and not w9539;
w9541 <= not w264 and not w9540;
w9542 <= w9060 and not w9062;
w9543 <= not w9053 and w9542;
w9544 <= not w9163 and w9543;
w9545 <= not w9053 and not w9062;
w9546 <= not w9163 and w9545;
w9547 <= not w9060 and not w9546;
w9548 <= not w9544 and not w9547;
w9549 <= w264 and not w9529;
w9550 <= not w9539 and w9549;
w9551 <= not w9548 and not w9550;
w9552 <= not w9541 and not w9551;
w9553 <= not w184 and not w9552;
w9554 <= not w9065 and w9072;
w9555 <= not w9074 and w9554;
w9556 <= not w9163 and w9555;
w9557 <= not w9065 and not w9074;
w9558 <= not w9163 and w9557;
w9559 <= not w9072 and not w9558;
w9560 <= not w9556 and not w9559;
w9561 <= w184 and not w9541;
w9562 <= not w9551 and w9561;
w9563 <= not w9560 and not w9562;
w9564 <= not w9553 and not w9563;
w9565 <= not w115 and not w9564;
w9566 <= w9084 and not w9086;
w9567 <= not w9077 and w9566;
w9568 <= not w9163 and w9567;
w9569 <= not w9077 and not w9086;
w9570 <= not w9163 and w9569;
w9571 <= not w9084 and not w9570;
w9572 <= not w9568 and not w9571;
w9573 <= w115 and not w9553;
w9574 <= not w9563 and w9573;
w9575 <= not w9572 and not w9574;
w9576 <= not w9565 and not w9575;
w9577 <= not w60 and not w9576;
w9578 <= not w9089 and w9096;
w9579 <= not w9098 and w9578;
w9580 <= not w9163 and w9579;
w9581 <= not w9089 and not w9098;
w9582 <= not w9163 and w9581;
w9583 <= not w9096 and not w9582;
w9584 <= not w9580 and not w9583;
w9585 <= w60 and not w9565;
w9586 <= not w9575 and w9585;
w9587 <= not w9584 and not w9586;
w9588 <= not w9577 and not w9587;
w9589 <= not w22 and not w9588;
w9590 <= w9108 and not w9110;
w9591 <= not w9101 and w9590;
w9592 <= not w9163 and w9591;
w9593 <= not w9101 and not w9110;
w9594 <= not w9163 and w9593;
w9595 <= not w9108 and not w9594;
w9596 <= not w9592 and not w9595;
w9597 <= w22 and not w9577;
w9598 <= not w9587 and w9597;
w9599 <= not w9596 and not w9598;
w9600 <= not w9589 and not w9599;
w9601 <= not w5 and not w9600;
w9602 <= not w9113 and w9120;
w9603 <= not w9122 and w9602;
w9604 <= not w9163 and w9603;
w9605 <= not w9113 and not w9122;
w9606 <= not w9163 and w9605;
w9607 <= not w9120 and not w9606;
w9608 <= not w9604 and not w9607;
w9609 <= w5 and not w9589;
w9610 <= not w9599 and w9609;
w9611 <= not w9608 and not w9610;
w9612 <= not w9601 and not w9611;
w9613 <= w9132 and not w9134;
w9614 <= not w9125 and w9613;
w9615 <= not w9163 and w9614;
w9616 <= not w9125 and not w9134;
w9617 <= not w9163 and w9616;
w9618 <= not w9132 and not w9617;
w9619 <= not w9615 and not w9618;
w9620 <= not w9136 and not w9143;
w9621 <= not w9163 and w9620;
w9622 <= not w9151 and not w9621;
w9623 <= not w9619 and w9622;
w9624 <= not w9612 and w9623;
w9625 <= w0 and not w9624;
w9626 <= not w9601 and w9619;
w9627 <= not w9611 and w9626;
w9628 <= not w9143 and not w9163;
w9629 <= w9136 and not w9628;
w9630 <= not w0 and not w9620;
w9631 <= not w9629 and w9630;
w9632 <= not w9139 and not w9160;
w9633 <= not w9142 and w9632;
w9634 <= not w9155 and w9633;
w9635 <= not w9151 and w9634;
w9636 <= not w9149 and w9635;
w9637 <= not w9631 and not w9636;
w9638 <= not w9627 and w9637;
w9639 <= not w9625 and w9638;
w9640 <= a(48) and not w9639;
w9641 <= not a(46) and not a(47);
w9642 <= not a(48) and w9641;
w9643 <= not w9640 and not w9642;
w9644 <= not w9163 and not w9643;
w9645 <= not w9160 and not w9642;
w9646 <= not w9155 and w9645;
w9647 <= not w9151 and w9646;
w9648 <= not w9149 and w9647;
w9649 <= not w9640 and w9648;
w9650 <= not a(48) and not w9639;
w9651 <= a(49) and not w9650;
w9652 <= w9165 and not w9639;
w9653 <= not w9651 and not w9652;
w9654 <= not w9649 and w9653;
w9655 <= not w9644 and not w9654;
w9656 <= not w8699 and not w9655;
w9657 <= w8699 and not w9644;
w9658 <= not w9654 and w9657;
w9659 <= not w9163 and not w9636;
w9660 <= not w9631 and w9659;
w9661 <= not w9627 and w9660;
w9662 <= not w9625 and w9661;
w9663 <= not w9652 and not w9662;
w9664 <= a(50) and not w9663;
w9665 <= not a(50) and not w9662;
w9666 <= not w9652 and w9665;
w9667 <= not w9664 and not w9666;
w9668 <= not w9658 and not w9667;
w9669 <= not w9656 and not w9668;
w9670 <= not w8247 and not w9669;
w9671 <= not w9168 and not w9173;
w9672 <= not w9177 and w9671;
w9673 <= not w9639 and w9672;
w9674 <= not w9639 and w9671;
w9675 <= w9177 and not w9674;
w9676 <= not w9673 and not w9675;
w9677 <= w8247 and not w9656;
w9678 <= not w9668 and w9677;
w9679 <= not w9676 and not w9678;
w9680 <= not w9670 and not w9679;
w9681 <= not w7807 and not w9680;
w9682 <= not w9182 and w9191;
w9683 <= not w9180 and w9682;
w9684 <= not w9639 and w9683;
w9685 <= not w9180 and not w9182;
w9686 <= not w9639 and w9685;
w9687 <= not w9191 and not w9686;
w9688 <= not w9684 and not w9687;
w9689 <= w7807 and not w9670;
w9690 <= not w9679 and w9689;
w9691 <= not w9688 and not w9690;
w9692 <= not w9681 and not w9691;
w9693 <= not w7379 and not w9692;
w9694 <= not w9194 and w9200;
w9695 <= not w9202 and w9694;
w9696 <= not w9639 and w9695;
w9697 <= not w9194 and not w9202;
w9698 <= not w9639 and w9697;
w9699 <= not w9200 and not w9698;
w9700 <= not w9696 and not w9699;
w9701 <= w7379 and not w9681;
w9702 <= not w9691 and w9701;
w9703 <= not w9700 and not w9702;
w9704 <= not w9693 and not w9703;
w9705 <= not w6963 and not w9704;
w9706 <= w9212 and not w9214;
w9707 <= not w9205 and w9706;
w9708 <= not w9639 and w9707;
w9709 <= not w9205 and not w9214;
w9710 <= not w9639 and w9709;
w9711 <= not w9212 and not w9710;
w9712 <= not w9708 and not w9711;
w9713 <= w6963 and not w9693;
w9714 <= not w9703 and w9713;
w9715 <= not w9712 and not w9714;
w9716 <= not w9705 and not w9715;
w9717 <= not w6558 and not w9716;
w9718 <= not w9217 and w9224;
w9719 <= not w9226 and w9718;
w9720 <= not w9639 and w9719;
w9721 <= not w9217 and not w9226;
w9722 <= not w9639 and w9721;
w9723 <= not w9224 and not w9722;
w9724 <= not w9720 and not w9723;
w9725 <= w6558 and not w9705;
w9726 <= not w9715 and w9725;
w9727 <= not w9724 and not w9726;
w9728 <= not w9717 and not w9727;
w9729 <= not w6166 and not w9728;
w9730 <= w9236 and not w9238;
w9731 <= not w9229 and w9730;
w9732 <= not w9639 and w9731;
w9733 <= not w9229 and not w9238;
w9734 <= not w9639 and w9733;
w9735 <= not w9236 and not w9734;
w9736 <= not w9732 and not w9735;
w9737 <= w6166 and not w9717;
w9738 <= not w9727 and w9737;
w9739 <= not w9736 and not w9738;
w9740 <= not w9729 and not w9739;
w9741 <= not w5786 and not w9740;
w9742 <= not w9241 and w9248;
w9743 <= not w9250 and w9742;
w9744 <= not w9639 and w9743;
w9745 <= not w9241 and not w9250;
w9746 <= not w9639 and w9745;
w9747 <= not w9248 and not w9746;
w9748 <= not w9744 and not w9747;
w9749 <= w5786 and not w9729;
w9750 <= not w9739 and w9749;
w9751 <= not w9748 and not w9750;
w9752 <= not w9741 and not w9751;
w9753 <= not w5418 and not w9752;
w9754 <= w9260 and not w9262;
w9755 <= not w9253 and w9754;
w9756 <= not w9639 and w9755;
w9757 <= not w9253 and not w9262;
w9758 <= not w9639 and w9757;
w9759 <= not w9260 and not w9758;
w9760 <= not w9756 and not w9759;
w9761 <= w5418 and not w9741;
w9762 <= not w9751 and w9761;
w9763 <= not w9760 and not w9762;
w9764 <= not w9753 and not w9763;
w9765 <= not w5062 and not w9764;
w9766 <= not w9265 and w9272;
w9767 <= not w9274 and w9766;
w9768 <= not w9639 and w9767;
w9769 <= not w9265 and not w9274;
w9770 <= not w9639 and w9769;
w9771 <= not w9272 and not w9770;
w9772 <= not w9768 and not w9771;
w9773 <= w5062 and not w9753;
w9774 <= not w9763 and w9773;
w9775 <= not w9772 and not w9774;
w9776 <= not w9765 and not w9775;
w9777 <= not w4718 and not w9776;
w9778 <= w9284 and not w9286;
w9779 <= not w9277 and w9778;
w9780 <= not w9639 and w9779;
w9781 <= not w9277 and not w9286;
w9782 <= not w9639 and w9781;
w9783 <= not w9284 and not w9782;
w9784 <= not w9780 and not w9783;
w9785 <= w4718 and not w9765;
w9786 <= not w9775 and w9785;
w9787 <= not w9784 and not w9786;
w9788 <= not w9777 and not w9787;
w9789 <= not w4386 and not w9788;
w9790 <= not w9289 and w9296;
w9791 <= not w9298 and w9790;
w9792 <= not w9639 and w9791;
w9793 <= not w9289 and not w9298;
w9794 <= not w9639 and w9793;
w9795 <= not w9296 and not w9794;
w9796 <= not w9792 and not w9795;
w9797 <= w4386 and not w9777;
w9798 <= not w9787 and w9797;
w9799 <= not w9796 and not w9798;
w9800 <= not w9789 and not w9799;
w9801 <= not w4066 and not w9800;
w9802 <= w9308 and not w9310;
w9803 <= not w9301 and w9802;
w9804 <= not w9639 and w9803;
w9805 <= not w9301 and not w9310;
w9806 <= not w9639 and w9805;
w9807 <= not w9308 and not w9806;
w9808 <= not w9804 and not w9807;
w9809 <= w4066 and not w9789;
w9810 <= not w9799 and w9809;
w9811 <= not w9808 and not w9810;
w9812 <= not w9801 and not w9811;
w9813 <= not w3758 and not w9812;
w9814 <= not w9313 and w9320;
w9815 <= not w9322 and w9814;
w9816 <= not w9639 and w9815;
w9817 <= not w9313 and not w9322;
w9818 <= not w9639 and w9817;
w9819 <= not w9320 and not w9818;
w9820 <= not w9816 and not w9819;
w9821 <= w3758 and not w9801;
w9822 <= not w9811 and w9821;
w9823 <= not w9820 and not w9822;
w9824 <= not w9813 and not w9823;
w9825 <= not w3462 and not w9824;
w9826 <= w9332 and not w9334;
w9827 <= not w9325 and w9826;
w9828 <= not w9639 and w9827;
w9829 <= not w9325 and not w9334;
w9830 <= not w9639 and w9829;
w9831 <= not w9332 and not w9830;
w9832 <= not w9828 and not w9831;
w9833 <= w3462 and not w9813;
w9834 <= not w9823 and w9833;
w9835 <= not w9832 and not w9834;
w9836 <= not w9825 and not w9835;
w9837 <= not w3178 and not w9836;
w9838 <= w3178 and not w9825;
w9839 <= not w9835 and w9838;
w9840 <= not w9337 and w9346;
w9841 <= not w9339 and w9840;
w9842 <= not w9639 and w9841;
w9843 <= not w9337 and not w9339;
w9844 <= not w9639 and w9843;
w9845 <= not w9346 and not w9844;
w9846 <= not w9842 and not w9845;
w9847 <= not w9839 and not w9846;
w9848 <= not w9837 and not w9847;
w9849 <= not w2906 and not w9848;
w9850 <= w9356 and not w9358;
w9851 <= not w9349 and w9850;
w9852 <= not w9639 and w9851;
w9853 <= not w9349 and not w9358;
w9854 <= not w9639 and w9853;
w9855 <= not w9356 and not w9854;
w9856 <= not w9852 and not w9855;
w9857 <= w2906 and not w9837;
w9858 <= not w9847 and w9857;
w9859 <= not w9856 and not w9858;
w9860 <= not w9849 and not w9859;
w9861 <= not w2646 and not w9860;
w9862 <= not w9361 and w9368;
w9863 <= not w9370 and w9862;
w9864 <= not w9639 and w9863;
w9865 <= not w9361 and not w9370;
w9866 <= not w9639 and w9865;
w9867 <= not w9368 and not w9866;
w9868 <= not w9864 and not w9867;
w9869 <= w2646 and not w9849;
w9870 <= not w9859 and w9869;
w9871 <= not w9868 and not w9870;
w9872 <= not w9861 and not w9871;
w9873 <= not w2398 and not w9872;
w9874 <= w9380 and not w9382;
w9875 <= not w9373 and w9874;
w9876 <= not w9639 and w9875;
w9877 <= not w9373 and not w9382;
w9878 <= not w9639 and w9877;
w9879 <= not w9380 and not w9878;
w9880 <= not w9876 and not w9879;
w9881 <= w2398 and not w9861;
w9882 <= not w9871 and w9881;
w9883 <= not w9880 and not w9882;
w9884 <= not w9873 and not w9883;
w9885 <= not w2162 and not w9884;
w9886 <= not w9385 and w9392;
w9887 <= not w9394 and w9886;
w9888 <= not w9639 and w9887;
w9889 <= not w9385 and not w9394;
w9890 <= not w9639 and w9889;
w9891 <= not w9392 and not w9890;
w9892 <= not w9888 and not w9891;
w9893 <= w2162 and not w9873;
w9894 <= not w9883 and w9893;
w9895 <= not w9892 and not w9894;
w9896 <= not w9885 and not w9895;
w9897 <= not w1938 and not w9896;
w9898 <= w9404 and not w9406;
w9899 <= not w9397 and w9898;
w9900 <= not w9639 and w9899;
w9901 <= not w9397 and not w9406;
w9902 <= not w9639 and w9901;
w9903 <= not w9404 and not w9902;
w9904 <= not w9900 and not w9903;
w9905 <= w1938 and not w9885;
w9906 <= not w9895 and w9905;
w9907 <= not w9904 and not w9906;
w9908 <= not w9897 and not w9907;
w9909 <= not w1725 and not w9908;
w9910 <= not w9409 and w9416;
w9911 <= not w9418 and w9910;
w9912 <= not w9639 and w9911;
w9913 <= not w9409 and not w9418;
w9914 <= not w9639 and w9913;
w9915 <= not w9416 and not w9914;
w9916 <= not w9912 and not w9915;
w9917 <= w1725 and not w9897;
w9918 <= not w9907 and w9917;
w9919 <= not w9916 and not w9918;
w9920 <= not w9909 and not w9919;
w9921 <= not w1525 and not w9920;
w9922 <= w9428 and not w9430;
w9923 <= not w9421 and w9922;
w9924 <= not w9639 and w9923;
w9925 <= not w9421 and not w9430;
w9926 <= not w9639 and w9925;
w9927 <= not w9428 and not w9926;
w9928 <= not w9924 and not w9927;
w9929 <= w1525 and not w9909;
w9930 <= not w9919 and w9929;
w9931 <= not w9928 and not w9930;
w9932 <= not w9921 and not w9931;
w9933 <= not w1337 and not w9932;
w9934 <= not w9433 and w9440;
w9935 <= not w9442 and w9934;
w9936 <= not w9639 and w9935;
w9937 <= not w9433 and not w9442;
w9938 <= not w9639 and w9937;
w9939 <= not w9440 and not w9938;
w9940 <= not w9936 and not w9939;
w9941 <= w1337 and not w9921;
w9942 <= not w9931 and w9941;
w9943 <= not w9940 and not w9942;
w9944 <= not w9933 and not w9943;
w9945 <= not w1161 and not w9944;
w9946 <= w9452 and not w9454;
w9947 <= not w9445 and w9946;
w9948 <= not w9639 and w9947;
w9949 <= not w9445 and not w9454;
w9950 <= not w9639 and w9949;
w9951 <= not w9452 and not w9950;
w9952 <= not w9948 and not w9951;
w9953 <= w1161 and not w9933;
w9954 <= not w9943 and w9953;
w9955 <= not w9952 and not w9954;
w9956 <= not w9945 and not w9955;
w9957 <= not w997 and not w9956;
w9958 <= not w9457 and w9464;
w9959 <= not w9466 and w9958;
w9960 <= not w9639 and w9959;
w9961 <= not w9457 and not w9466;
w9962 <= not w9639 and w9961;
w9963 <= not w9464 and not w9962;
w9964 <= not w9960 and not w9963;
w9965 <= w997 and not w9945;
w9966 <= not w9955 and w9965;
w9967 <= not w9964 and not w9966;
w9968 <= not w9957 and not w9967;
w9969 <= not w845 and not w9968;
w9970 <= w9476 and not w9478;
w9971 <= not w9469 and w9970;
w9972 <= not w9639 and w9971;
w9973 <= not w9469 and not w9478;
w9974 <= not w9639 and w9973;
w9975 <= not w9476 and not w9974;
w9976 <= not w9972 and not w9975;
w9977 <= w845 and not w9957;
w9978 <= not w9967 and w9977;
w9979 <= not w9976 and not w9978;
w9980 <= not w9969 and not w9979;
w9981 <= not w705 and not w9980;
w9982 <= not w9481 and w9488;
w9983 <= not w9490 and w9982;
w9984 <= not w9639 and w9983;
w9985 <= not w9481 and not w9490;
w9986 <= not w9639 and w9985;
w9987 <= not w9488 and not w9986;
w9988 <= not w9984 and not w9987;
w9989 <= w705 and not w9969;
w9990 <= not w9979 and w9989;
w9991 <= not w9988 and not w9990;
w9992 <= not w9981 and not w9991;
w9993 <= not w577 and not w9992;
w9994 <= w9500 and not w9502;
w9995 <= not w9493 and w9994;
w9996 <= not w9639 and w9995;
w9997 <= not w9493 and not w9502;
w9998 <= not w9639 and w9997;
w9999 <= not w9500 and not w9998;
w10000 <= not w9996 and not w9999;
w10001 <= w577 and not w9981;
w10002 <= not w9991 and w10001;
w10003 <= not w10000 and not w10002;
w10004 <= not w9993 and not w10003;
w10005 <= not w460 and not w10004;
w10006 <= not w9505 and w9512;
w10007 <= not w9514 and w10006;
w10008 <= not w9639 and w10007;
w10009 <= not w9505 and not w9514;
w10010 <= not w9639 and w10009;
w10011 <= not w9512 and not w10010;
w10012 <= not w10008 and not w10011;
w10013 <= w460 and not w9993;
w10014 <= not w10003 and w10013;
w10015 <= not w10012 and not w10014;
w10016 <= not w10005 and not w10015;
w10017 <= not w356 and not w10016;
w10018 <= w9524 and not w9526;
w10019 <= not w9517 and w10018;
w10020 <= not w9639 and w10019;
w10021 <= not w9517 and not w9526;
w10022 <= not w9639 and w10021;
w10023 <= not w9524 and not w10022;
w10024 <= not w10020 and not w10023;
w10025 <= w356 and not w10005;
w10026 <= not w10015 and w10025;
w10027 <= not w10024 and not w10026;
w10028 <= not w10017 and not w10027;
w10029 <= not w264 and not w10028;
w10030 <= not w9529 and w9536;
w10031 <= not w9538 and w10030;
w10032 <= not w9639 and w10031;
w10033 <= not w9529 and not w9538;
w10034 <= not w9639 and w10033;
w10035 <= not w9536 and not w10034;
w10036 <= not w10032 and not w10035;
w10037 <= w264 and not w10017;
w10038 <= not w10027 and w10037;
w10039 <= not w10036 and not w10038;
w10040 <= not w10029 and not w10039;
w10041 <= not w184 and not w10040;
w10042 <= w9548 and not w9550;
w10043 <= not w9541 and w10042;
w10044 <= not w9639 and w10043;
w10045 <= not w9541 and not w9550;
w10046 <= not w9639 and w10045;
w10047 <= not w9548 and not w10046;
w10048 <= not w10044 and not w10047;
w10049 <= w184 and not w10029;
w10050 <= not w10039 and w10049;
w10051 <= not w10048 and not w10050;
w10052 <= not w10041 and not w10051;
w10053 <= not w115 and not w10052;
w10054 <= not w9553 and w9560;
w10055 <= not w9562 and w10054;
w10056 <= not w9639 and w10055;
w10057 <= not w9553 and not w9562;
w10058 <= not w9639 and w10057;
w10059 <= not w9560 and not w10058;
w10060 <= not w10056 and not w10059;
w10061 <= w115 and not w10041;
w10062 <= not w10051 and w10061;
w10063 <= not w10060 and not w10062;
w10064 <= not w10053 and not w10063;
w10065 <= not w60 and not w10064;
w10066 <= w9572 and not w9574;
w10067 <= not w9565 and w10066;
w10068 <= not w9639 and w10067;
w10069 <= not w9565 and not w9574;
w10070 <= not w9639 and w10069;
w10071 <= not w9572 and not w10070;
w10072 <= not w10068 and not w10071;
w10073 <= w60 and not w10053;
w10074 <= not w10063 and w10073;
w10075 <= not w10072 and not w10074;
w10076 <= not w10065 and not w10075;
w10077 <= not w22 and not w10076;
w10078 <= not w9577 and w9584;
w10079 <= not w9586 and w10078;
w10080 <= not w9639 and w10079;
w10081 <= not w9577 and not w9586;
w10082 <= not w9639 and w10081;
w10083 <= not w9584 and not w10082;
w10084 <= not w10080 and not w10083;
w10085 <= w22 and not w10065;
w10086 <= not w10075 and w10085;
w10087 <= not w10084 and not w10086;
w10088 <= not w10077 and not w10087;
w10089 <= not w5 and not w10088;
w10090 <= w9596 and not w9598;
w10091 <= not w9589 and w10090;
w10092 <= not w9639 and w10091;
w10093 <= not w9589 and not w9598;
w10094 <= not w9639 and w10093;
w10095 <= not w9596 and not w10094;
w10096 <= not w10092 and not w10095;
w10097 <= w5 and not w10077;
w10098 <= not w10087 and w10097;
w10099 <= not w10096 and not w10098;
w10100 <= not w10089 and not w10099;
w10101 <= not w9601 and w9608;
w10102 <= not w9610 and w10101;
w10103 <= not w9639 and w10102;
w10104 <= not w9601 and not w9610;
w10105 <= not w9639 and w10104;
w10106 <= not w9608 and not w10105;
w10107 <= not w10103 and not w10106;
w10108 <= not w9612 and not w9619;
w10109 <= not w9639 and w10108;
w10110 <= not w9627 and not w10109;
w10111 <= not w10107 and w10110;
w10112 <= not w10100 and w10111;
w10113 <= w0 and not w10112;
w10114 <= not w10089 and w10107;
w10115 <= not w10099 and w10114;
w10116 <= not w9619 and not w9639;
w10117 <= w9612 and not w10116;
w10118 <= not w0 and not w10108;
w10119 <= not w10117 and w10118;
w10120 <= not w9615 and not w9636;
w10121 <= not w9618 and w10120;
w10122 <= not w9631 and w10121;
w10123 <= not w9627 and w10122;
w10124 <= not w9625 and w10123;
w10125 <= not w10119 and not w10124;
w10126 <= not w10115 and w10125;
w10127 <= not w10113 and w10126;
w10128 <= a(46) and not w10127;
w10129 <= not a(44) and not a(45);
w10130 <= not a(46) and w10129;
w10131 <= not w10128 and not w10130;
w10132 <= not w9639 and not w10131;
w10133 <= not w9636 and not w10130;
w10134 <= not w9631 and w10133;
w10135 <= not w9627 and w10134;
w10136 <= not w9625 and w10135;
w10137 <= not w10128 and w10136;
w10138 <= not a(46) and not w10127;
w10139 <= a(47) and not w10138;
w10140 <= w9641 and not w10127;
w10141 <= not w10139 and not w10140;
w10142 <= not w10137 and w10141;
w10143 <= not w10132 and not w10142;
w10144 <= not w9163 and not w10143;
w10145 <= w9163 and not w10132;
w10146 <= not w10142 and w10145;
w10147 <= not w9639 and not w10124;
w10148 <= not w10119 and w10147;
w10149 <= not w10115 and w10148;
w10150 <= not w10113 and w10149;
w10151 <= not w10140 and not w10150;
w10152 <= a(48) and not w10151;
w10153 <= not a(48) and not w10150;
w10154 <= not w10140 and w10153;
w10155 <= not w10152 and not w10154;
w10156 <= not w10146 and not w10155;
w10157 <= not w10144 and not w10156;
w10158 <= not w8699 and not w10157;
w10159 <= not w9644 and not w9649;
w10160 <= not w9653 and w10159;
w10161 <= not w10127 and w10160;
w10162 <= not w10127 and w10159;
w10163 <= w9653 and not w10162;
w10164 <= not w10161 and not w10163;
w10165 <= w8699 and not w10144;
w10166 <= not w10156 and w10165;
w10167 <= not w10164 and not w10166;
w10168 <= not w10158 and not w10167;
w10169 <= not w8247 and not w10168;
w10170 <= not w9658 and w9667;
w10171 <= not w9656 and w10170;
w10172 <= not w10127 and w10171;
w10173 <= not w9656 and not w9658;
w10174 <= not w10127 and w10173;
w10175 <= not w9667 and not w10174;
w10176 <= not w10172 and not w10175;
w10177 <= w8247 and not w10158;
w10178 <= not w10167 and w10177;
w10179 <= not w10176 and not w10178;
w10180 <= not w10169 and not w10179;
w10181 <= not w7807 and not w10180;
w10182 <= not w9670 and w9676;
w10183 <= not w9678 and w10182;
w10184 <= not w10127 and w10183;
w10185 <= not w9670 and not w9678;
w10186 <= not w10127 and w10185;
w10187 <= not w9676 and not w10186;
w10188 <= not w10184 and not w10187;
w10189 <= w7807 and not w10169;
w10190 <= not w10179 and w10189;
w10191 <= not w10188 and not w10190;
w10192 <= not w10181 and not w10191;
w10193 <= not w7379 and not w10192;
w10194 <= w9688 and not w9690;
w10195 <= not w9681 and w10194;
w10196 <= not w10127 and w10195;
w10197 <= not w9681 and not w9690;
w10198 <= not w10127 and w10197;
w10199 <= not w9688 and not w10198;
w10200 <= not w10196 and not w10199;
w10201 <= w7379 and not w10181;
w10202 <= not w10191 and w10201;
w10203 <= not w10200 and not w10202;
w10204 <= not w10193 and not w10203;
w10205 <= not w6963 and not w10204;
w10206 <= not w9693 and w9700;
w10207 <= not w9702 and w10206;
w10208 <= not w10127 and w10207;
w10209 <= not w9693 and not w9702;
w10210 <= not w10127 and w10209;
w10211 <= not w9700 and not w10210;
w10212 <= not w10208 and not w10211;
w10213 <= w6963 and not w10193;
w10214 <= not w10203 and w10213;
w10215 <= not w10212 and not w10214;
w10216 <= not w10205 and not w10215;
w10217 <= not w6558 and not w10216;
w10218 <= w9712 and not w9714;
w10219 <= not w9705 and w10218;
w10220 <= not w10127 and w10219;
w10221 <= not w9705 and not w9714;
w10222 <= not w10127 and w10221;
w10223 <= not w9712 and not w10222;
w10224 <= not w10220 and not w10223;
w10225 <= w6558 and not w10205;
w10226 <= not w10215 and w10225;
w10227 <= not w10224 and not w10226;
w10228 <= not w10217 and not w10227;
w10229 <= not w6166 and not w10228;
w10230 <= not w9717 and w9724;
w10231 <= not w9726 and w10230;
w10232 <= not w10127 and w10231;
w10233 <= not w9717 and not w9726;
w10234 <= not w10127 and w10233;
w10235 <= not w9724 and not w10234;
w10236 <= not w10232 and not w10235;
w10237 <= w6166 and not w10217;
w10238 <= not w10227 and w10237;
w10239 <= not w10236 and not w10238;
w10240 <= not w10229 and not w10239;
w10241 <= not w5786 and not w10240;
w10242 <= w9736 and not w9738;
w10243 <= not w9729 and w10242;
w10244 <= not w10127 and w10243;
w10245 <= not w9729 and not w9738;
w10246 <= not w10127 and w10245;
w10247 <= not w9736 and not w10246;
w10248 <= not w10244 and not w10247;
w10249 <= w5786 and not w10229;
w10250 <= not w10239 and w10249;
w10251 <= not w10248 and not w10250;
w10252 <= not w10241 and not w10251;
w10253 <= not w5418 and not w10252;
w10254 <= not w9741 and w9748;
w10255 <= not w9750 and w10254;
w10256 <= not w10127 and w10255;
w10257 <= not w9741 and not w9750;
w10258 <= not w10127 and w10257;
w10259 <= not w9748 and not w10258;
w10260 <= not w10256 and not w10259;
w10261 <= w5418 and not w10241;
w10262 <= not w10251 and w10261;
w10263 <= not w10260 and not w10262;
w10264 <= not w10253 and not w10263;
w10265 <= not w5062 and not w10264;
w10266 <= w9760 and not w9762;
w10267 <= not w9753 and w10266;
w10268 <= not w10127 and w10267;
w10269 <= not w9753 and not w9762;
w10270 <= not w10127 and w10269;
w10271 <= not w9760 and not w10270;
w10272 <= not w10268 and not w10271;
w10273 <= w5062 and not w10253;
w10274 <= not w10263 and w10273;
w10275 <= not w10272 and not w10274;
w10276 <= not w10265 and not w10275;
w10277 <= not w4718 and not w10276;
w10278 <= not w9765 and w9772;
w10279 <= not w9774 and w10278;
w10280 <= not w10127 and w10279;
w10281 <= not w9765 and not w9774;
w10282 <= not w10127 and w10281;
w10283 <= not w9772 and not w10282;
w10284 <= not w10280 and not w10283;
w10285 <= w4718 and not w10265;
w10286 <= not w10275 and w10285;
w10287 <= not w10284 and not w10286;
w10288 <= not w10277 and not w10287;
w10289 <= not w4386 and not w10288;
w10290 <= w9784 and not w9786;
w10291 <= not w9777 and w10290;
w10292 <= not w10127 and w10291;
w10293 <= not w9777 and not w9786;
w10294 <= not w10127 and w10293;
w10295 <= not w9784 and not w10294;
w10296 <= not w10292 and not w10295;
w10297 <= w4386 and not w10277;
w10298 <= not w10287 and w10297;
w10299 <= not w10296 and not w10298;
w10300 <= not w10289 and not w10299;
w10301 <= not w4066 and not w10300;
w10302 <= not w9789 and w9796;
w10303 <= not w9798 and w10302;
w10304 <= not w10127 and w10303;
w10305 <= not w9789 and not w9798;
w10306 <= not w10127 and w10305;
w10307 <= not w9796 and not w10306;
w10308 <= not w10304 and not w10307;
w10309 <= w4066 and not w10289;
w10310 <= not w10299 and w10309;
w10311 <= not w10308 and not w10310;
w10312 <= not w10301 and not w10311;
w10313 <= not w3758 and not w10312;
w10314 <= w9808 and not w9810;
w10315 <= not w9801 and w10314;
w10316 <= not w10127 and w10315;
w10317 <= not w9801 and not w9810;
w10318 <= not w10127 and w10317;
w10319 <= not w9808 and not w10318;
w10320 <= not w10316 and not w10319;
w10321 <= w3758 and not w10301;
w10322 <= not w10311 and w10321;
w10323 <= not w10320 and not w10322;
w10324 <= not w10313 and not w10323;
w10325 <= not w3462 and not w10324;
w10326 <= not w9813 and w9820;
w10327 <= not w9822 and w10326;
w10328 <= not w10127 and w10327;
w10329 <= not w9813 and not w9822;
w10330 <= not w10127 and w10329;
w10331 <= not w9820 and not w10330;
w10332 <= not w10328 and not w10331;
w10333 <= w3462 and not w10313;
w10334 <= not w10323 and w10333;
w10335 <= not w10332 and not w10334;
w10336 <= not w10325 and not w10335;
w10337 <= not w3178 and not w10336;
w10338 <= w9832 and not w9834;
w10339 <= not w9825 and w10338;
w10340 <= not w10127 and w10339;
w10341 <= not w9825 and not w9834;
w10342 <= not w10127 and w10341;
w10343 <= not w9832 and not w10342;
w10344 <= not w10340 and not w10343;
w10345 <= w3178 and not w10325;
w10346 <= not w10335 and w10345;
w10347 <= not w10344 and not w10346;
w10348 <= not w10337 and not w10347;
w10349 <= not w2906 and not w10348;
w10350 <= w2906 and not w10337;
w10351 <= not w10347 and w10350;
w10352 <= not w9837 and w9846;
w10353 <= not w9839 and w10352;
w10354 <= not w10127 and w10353;
w10355 <= not w9837 and not w9839;
w10356 <= not w10127 and w10355;
w10357 <= not w9846 and not w10356;
w10358 <= not w10354 and not w10357;
w10359 <= not w10351 and not w10358;
w10360 <= not w10349 and not w10359;
w10361 <= not w2646 and not w10360;
w10362 <= w9856 and not w9858;
w10363 <= not w9849 and w10362;
w10364 <= not w10127 and w10363;
w10365 <= not w9849 and not w9858;
w10366 <= not w10127 and w10365;
w10367 <= not w9856 and not w10366;
w10368 <= not w10364 and not w10367;
w10369 <= w2646 and not w10349;
w10370 <= not w10359 and w10369;
w10371 <= not w10368 and not w10370;
w10372 <= not w10361 and not w10371;
w10373 <= not w2398 and not w10372;
w10374 <= not w9861 and w9868;
w10375 <= not w9870 and w10374;
w10376 <= not w10127 and w10375;
w10377 <= not w9861 and not w9870;
w10378 <= not w10127 and w10377;
w10379 <= not w9868 and not w10378;
w10380 <= not w10376 and not w10379;
w10381 <= w2398 and not w10361;
w10382 <= not w10371 and w10381;
w10383 <= not w10380 and not w10382;
w10384 <= not w10373 and not w10383;
w10385 <= not w2162 and not w10384;
w10386 <= w9880 and not w9882;
w10387 <= not w9873 and w10386;
w10388 <= not w10127 and w10387;
w10389 <= not w9873 and not w9882;
w10390 <= not w10127 and w10389;
w10391 <= not w9880 and not w10390;
w10392 <= not w10388 and not w10391;
w10393 <= w2162 and not w10373;
w10394 <= not w10383 and w10393;
w10395 <= not w10392 and not w10394;
w10396 <= not w10385 and not w10395;
w10397 <= not w1938 and not w10396;
w10398 <= not w9885 and w9892;
w10399 <= not w9894 and w10398;
w10400 <= not w10127 and w10399;
w10401 <= not w9885 and not w9894;
w10402 <= not w10127 and w10401;
w10403 <= not w9892 and not w10402;
w10404 <= not w10400 and not w10403;
w10405 <= w1938 and not w10385;
w10406 <= not w10395 and w10405;
w10407 <= not w10404 and not w10406;
w10408 <= not w10397 and not w10407;
w10409 <= not w1725 and not w10408;
w10410 <= w9904 and not w9906;
w10411 <= not w9897 and w10410;
w10412 <= not w10127 and w10411;
w10413 <= not w9897 and not w9906;
w10414 <= not w10127 and w10413;
w10415 <= not w9904 and not w10414;
w10416 <= not w10412 and not w10415;
w10417 <= w1725 and not w10397;
w10418 <= not w10407 and w10417;
w10419 <= not w10416 and not w10418;
w10420 <= not w10409 and not w10419;
w10421 <= not w1525 and not w10420;
w10422 <= not w9909 and w9916;
w10423 <= not w9918 and w10422;
w10424 <= not w10127 and w10423;
w10425 <= not w9909 and not w9918;
w10426 <= not w10127 and w10425;
w10427 <= not w9916 and not w10426;
w10428 <= not w10424 and not w10427;
w10429 <= w1525 and not w10409;
w10430 <= not w10419 and w10429;
w10431 <= not w10428 and not w10430;
w10432 <= not w10421 and not w10431;
w10433 <= not w1337 and not w10432;
w10434 <= w9928 and not w9930;
w10435 <= not w9921 and w10434;
w10436 <= not w10127 and w10435;
w10437 <= not w9921 and not w9930;
w10438 <= not w10127 and w10437;
w10439 <= not w9928 and not w10438;
w10440 <= not w10436 and not w10439;
w10441 <= w1337 and not w10421;
w10442 <= not w10431 and w10441;
w10443 <= not w10440 and not w10442;
w10444 <= not w10433 and not w10443;
w10445 <= not w1161 and not w10444;
w10446 <= not w9933 and w9940;
w10447 <= not w9942 and w10446;
w10448 <= not w10127 and w10447;
w10449 <= not w9933 and not w9942;
w10450 <= not w10127 and w10449;
w10451 <= not w9940 and not w10450;
w10452 <= not w10448 and not w10451;
w10453 <= w1161 and not w10433;
w10454 <= not w10443 and w10453;
w10455 <= not w10452 and not w10454;
w10456 <= not w10445 and not w10455;
w10457 <= not w997 and not w10456;
w10458 <= w9952 and not w9954;
w10459 <= not w9945 and w10458;
w10460 <= not w10127 and w10459;
w10461 <= not w9945 and not w9954;
w10462 <= not w10127 and w10461;
w10463 <= not w9952 and not w10462;
w10464 <= not w10460 and not w10463;
w10465 <= w997 and not w10445;
w10466 <= not w10455 and w10465;
w10467 <= not w10464 and not w10466;
w10468 <= not w10457 and not w10467;
w10469 <= not w845 and not w10468;
w10470 <= not w9957 and w9964;
w10471 <= not w9966 and w10470;
w10472 <= not w10127 and w10471;
w10473 <= not w9957 and not w9966;
w10474 <= not w10127 and w10473;
w10475 <= not w9964 and not w10474;
w10476 <= not w10472 and not w10475;
w10477 <= w845 and not w10457;
w10478 <= not w10467 and w10477;
w10479 <= not w10476 and not w10478;
w10480 <= not w10469 and not w10479;
w10481 <= not w705 and not w10480;
w10482 <= w9976 and not w9978;
w10483 <= not w9969 and w10482;
w10484 <= not w10127 and w10483;
w10485 <= not w9969 and not w9978;
w10486 <= not w10127 and w10485;
w10487 <= not w9976 and not w10486;
w10488 <= not w10484 and not w10487;
w10489 <= w705 and not w10469;
w10490 <= not w10479 and w10489;
w10491 <= not w10488 and not w10490;
w10492 <= not w10481 and not w10491;
w10493 <= not w577 and not w10492;
w10494 <= not w9981 and w9988;
w10495 <= not w9990 and w10494;
w10496 <= not w10127 and w10495;
w10497 <= not w9981 and not w9990;
w10498 <= not w10127 and w10497;
w10499 <= not w9988 and not w10498;
w10500 <= not w10496 and not w10499;
w10501 <= w577 and not w10481;
w10502 <= not w10491 and w10501;
w10503 <= not w10500 and not w10502;
w10504 <= not w10493 and not w10503;
w10505 <= not w460 and not w10504;
w10506 <= w10000 and not w10002;
w10507 <= not w9993 and w10506;
w10508 <= not w10127 and w10507;
w10509 <= not w9993 and not w10002;
w10510 <= not w10127 and w10509;
w10511 <= not w10000 and not w10510;
w10512 <= not w10508 and not w10511;
w10513 <= w460 and not w10493;
w10514 <= not w10503 and w10513;
w10515 <= not w10512 and not w10514;
w10516 <= not w10505 and not w10515;
w10517 <= not w356 and not w10516;
w10518 <= not w10005 and w10012;
w10519 <= not w10014 and w10518;
w10520 <= not w10127 and w10519;
w10521 <= not w10005 and not w10014;
w10522 <= not w10127 and w10521;
w10523 <= not w10012 and not w10522;
w10524 <= not w10520 and not w10523;
w10525 <= w356 and not w10505;
w10526 <= not w10515 and w10525;
w10527 <= not w10524 and not w10526;
w10528 <= not w10517 and not w10527;
w10529 <= not w264 and not w10528;
w10530 <= w10024 and not w10026;
w10531 <= not w10017 and w10530;
w10532 <= not w10127 and w10531;
w10533 <= not w10017 and not w10026;
w10534 <= not w10127 and w10533;
w10535 <= not w10024 and not w10534;
w10536 <= not w10532 and not w10535;
w10537 <= w264 and not w10517;
w10538 <= not w10527 and w10537;
w10539 <= not w10536 and not w10538;
w10540 <= not w10529 and not w10539;
w10541 <= not w184 and not w10540;
w10542 <= not w10029 and w10036;
w10543 <= not w10038 and w10542;
w10544 <= not w10127 and w10543;
w10545 <= not w10029 and not w10038;
w10546 <= not w10127 and w10545;
w10547 <= not w10036 and not w10546;
w10548 <= not w10544 and not w10547;
w10549 <= w184 and not w10529;
w10550 <= not w10539 and w10549;
w10551 <= not w10548 and not w10550;
w10552 <= not w10541 and not w10551;
w10553 <= not w115 and not w10552;
w10554 <= w10048 and not w10050;
w10555 <= not w10041 and w10554;
w10556 <= not w10127 and w10555;
w10557 <= not w10041 and not w10050;
w10558 <= not w10127 and w10557;
w10559 <= not w10048 and not w10558;
w10560 <= not w10556 and not w10559;
w10561 <= w115 and not w10541;
w10562 <= not w10551 and w10561;
w10563 <= not w10560 and not w10562;
w10564 <= not w10553 and not w10563;
w10565 <= not w60 and not w10564;
w10566 <= not w10053 and w10060;
w10567 <= not w10062 and w10566;
w10568 <= not w10127 and w10567;
w10569 <= not w10053 and not w10062;
w10570 <= not w10127 and w10569;
w10571 <= not w10060 and not w10570;
w10572 <= not w10568 and not w10571;
w10573 <= w60 and not w10553;
w10574 <= not w10563 and w10573;
w10575 <= not w10572 and not w10574;
w10576 <= not w10565 and not w10575;
w10577 <= not w22 and not w10576;
w10578 <= w10072 and not w10074;
w10579 <= not w10065 and w10578;
w10580 <= not w10127 and w10579;
w10581 <= not w10065 and not w10074;
w10582 <= not w10127 and w10581;
w10583 <= not w10072 and not w10582;
w10584 <= not w10580 and not w10583;
w10585 <= w22 and not w10565;
w10586 <= not w10575 and w10585;
w10587 <= not w10584 and not w10586;
w10588 <= not w10577 and not w10587;
w10589 <= not w5 and not w10588;
w10590 <= not w10077 and w10084;
w10591 <= not w10086 and w10590;
w10592 <= not w10127 and w10591;
w10593 <= not w10077 and not w10086;
w10594 <= not w10127 and w10593;
w10595 <= not w10084 and not w10594;
w10596 <= not w10592 and not w10595;
w10597 <= w5 and not w10577;
w10598 <= not w10587 and w10597;
w10599 <= not w10596 and not w10598;
w10600 <= not w10589 and not w10599;
w10601 <= w10096 and not w10098;
w10602 <= not w10089 and w10601;
w10603 <= not w10127 and w10602;
w10604 <= not w10089 and not w10098;
w10605 <= not w10127 and w10604;
w10606 <= not w10096 and not w10605;
w10607 <= not w10603 and not w10606;
w10608 <= not w10100 and not w10107;
w10609 <= not w10127 and w10608;
w10610 <= not w10115 and not w10609;
w10611 <= not w10607 and w10610;
w10612 <= not w10600 and w10611;
w10613 <= w0 and not w10612;
w10614 <= not w10589 and w10607;
w10615 <= not w10599 and w10614;
w10616 <= not w10107 and not w10127;
w10617 <= w10100 and not w10616;
w10618 <= not w0 and not w10608;
w10619 <= not w10617 and w10618;
w10620 <= not w10103 and not w10124;
w10621 <= not w10106 and w10620;
w10622 <= not w10119 and w10621;
w10623 <= not w10115 and w10622;
w10624 <= not w10113 and w10623;
w10625 <= not w10619 and not w10624;
w10626 <= not w10615 and w10625;
w10627 <= not w10613 and w10626;
w10628 <= a(44) and not w10627;
w10629 <= not a(42) and not a(43);
w10630 <= not a(44) and w10629;
w10631 <= not w10628 and not w10630;
w10632 <= not w10127 and not w10631;
w10633 <= not w10124 and not w10630;
w10634 <= not w10119 and w10633;
w10635 <= not w10115 and w10634;
w10636 <= not w10113 and w10635;
w10637 <= not w10628 and w10636;
w10638 <= not a(44) and not w10627;
w10639 <= a(45) and not w10638;
w10640 <= w10129 and not w10627;
w10641 <= not w10639 and not w10640;
w10642 <= not w10637 and w10641;
w10643 <= not w10632 and not w10642;
w10644 <= not w9639 and not w10643;
w10645 <= w9639 and not w10632;
w10646 <= not w10642 and w10645;
w10647 <= not w10127 and not w10624;
w10648 <= not w10619 and w10647;
w10649 <= not w10615 and w10648;
w10650 <= not w10613 and w10649;
w10651 <= not w10640 and not w10650;
w10652 <= a(46) and not w10651;
w10653 <= not a(46) and not w10650;
w10654 <= not w10640 and w10653;
w10655 <= not w10652 and not w10654;
w10656 <= not w10646 and not w10655;
w10657 <= not w10644 and not w10656;
w10658 <= not w9163 and not w10657;
w10659 <= not w10132 and not w10137;
w10660 <= not w10141 and w10659;
w10661 <= not w10627 and w10660;
w10662 <= not w10627 and w10659;
w10663 <= w10141 and not w10662;
w10664 <= not w10661 and not w10663;
w10665 <= w9163 and not w10644;
w10666 <= not w10656 and w10665;
w10667 <= not w10664 and not w10666;
w10668 <= not w10658 and not w10667;
w10669 <= not w8699 and not w10668;
w10670 <= not w10146 and w10155;
w10671 <= not w10144 and w10670;
w10672 <= not w10627 and w10671;
w10673 <= not w10144 and not w10146;
w10674 <= not w10627 and w10673;
w10675 <= not w10155 and not w10674;
w10676 <= not w10672 and not w10675;
w10677 <= w8699 and not w10658;
w10678 <= not w10667 and w10677;
w10679 <= not w10676 and not w10678;
w10680 <= not w10669 and not w10679;
w10681 <= not w8247 and not w10680;
w10682 <= not w10158 and w10164;
w10683 <= not w10166 and w10682;
w10684 <= not w10627 and w10683;
w10685 <= not w10158 and not w10166;
w10686 <= not w10627 and w10685;
w10687 <= not w10164 and not w10686;
w10688 <= not w10684 and not w10687;
w10689 <= w8247 and not w10669;
w10690 <= not w10679 and w10689;
w10691 <= not w10688 and not w10690;
w10692 <= not w10681 and not w10691;
w10693 <= not w7807 and not w10692;
w10694 <= w10176 and not w10178;
w10695 <= not w10169 and w10694;
w10696 <= not w10627 and w10695;
w10697 <= not w10169 and not w10178;
w10698 <= not w10627 and w10697;
w10699 <= not w10176 and not w10698;
w10700 <= not w10696 and not w10699;
w10701 <= w7807 and not w10681;
w10702 <= not w10691 and w10701;
w10703 <= not w10700 and not w10702;
w10704 <= not w10693 and not w10703;
w10705 <= not w7379 and not w10704;
w10706 <= not w10181 and w10188;
w10707 <= not w10190 and w10706;
w10708 <= not w10627 and w10707;
w10709 <= not w10181 and not w10190;
w10710 <= not w10627 and w10709;
w10711 <= not w10188 and not w10710;
w10712 <= not w10708 and not w10711;
w10713 <= w7379 and not w10693;
w10714 <= not w10703 and w10713;
w10715 <= not w10712 and not w10714;
w10716 <= not w10705 and not w10715;
w10717 <= not w6963 and not w10716;
w10718 <= w10200 and not w10202;
w10719 <= not w10193 and w10718;
w10720 <= not w10627 and w10719;
w10721 <= not w10193 and not w10202;
w10722 <= not w10627 and w10721;
w10723 <= not w10200 and not w10722;
w10724 <= not w10720 and not w10723;
w10725 <= w6963 and not w10705;
w10726 <= not w10715 and w10725;
w10727 <= not w10724 and not w10726;
w10728 <= not w10717 and not w10727;
w10729 <= not w6558 and not w10728;
w10730 <= not w10205 and w10212;
w10731 <= not w10214 and w10730;
w10732 <= not w10627 and w10731;
w10733 <= not w10205 and not w10214;
w10734 <= not w10627 and w10733;
w10735 <= not w10212 and not w10734;
w10736 <= not w10732 and not w10735;
w10737 <= w6558 and not w10717;
w10738 <= not w10727 and w10737;
w10739 <= not w10736 and not w10738;
w10740 <= not w10729 and not w10739;
w10741 <= not w6166 and not w10740;
w10742 <= w10224 and not w10226;
w10743 <= not w10217 and w10742;
w10744 <= not w10627 and w10743;
w10745 <= not w10217 and not w10226;
w10746 <= not w10627 and w10745;
w10747 <= not w10224 and not w10746;
w10748 <= not w10744 and not w10747;
w10749 <= w6166 and not w10729;
w10750 <= not w10739 and w10749;
w10751 <= not w10748 and not w10750;
w10752 <= not w10741 and not w10751;
w10753 <= not w5786 and not w10752;
w10754 <= not w10229 and w10236;
w10755 <= not w10238 and w10754;
w10756 <= not w10627 and w10755;
w10757 <= not w10229 and not w10238;
w10758 <= not w10627 and w10757;
w10759 <= not w10236 and not w10758;
w10760 <= not w10756 and not w10759;
w10761 <= w5786 and not w10741;
w10762 <= not w10751 and w10761;
w10763 <= not w10760 and not w10762;
w10764 <= not w10753 and not w10763;
w10765 <= not w5418 and not w10764;
w10766 <= w10248 and not w10250;
w10767 <= not w10241 and w10766;
w10768 <= not w10627 and w10767;
w10769 <= not w10241 and not w10250;
w10770 <= not w10627 and w10769;
w10771 <= not w10248 and not w10770;
w10772 <= not w10768 and not w10771;
w10773 <= w5418 and not w10753;
w10774 <= not w10763 and w10773;
w10775 <= not w10772 and not w10774;
w10776 <= not w10765 and not w10775;
w10777 <= not w5062 and not w10776;
w10778 <= not w10253 and w10260;
w10779 <= not w10262 and w10778;
w10780 <= not w10627 and w10779;
w10781 <= not w10253 and not w10262;
w10782 <= not w10627 and w10781;
w10783 <= not w10260 and not w10782;
w10784 <= not w10780 and not w10783;
w10785 <= w5062 and not w10765;
w10786 <= not w10775 and w10785;
w10787 <= not w10784 and not w10786;
w10788 <= not w10777 and not w10787;
w10789 <= not w4718 and not w10788;
w10790 <= w10272 and not w10274;
w10791 <= not w10265 and w10790;
w10792 <= not w10627 and w10791;
w10793 <= not w10265 and not w10274;
w10794 <= not w10627 and w10793;
w10795 <= not w10272 and not w10794;
w10796 <= not w10792 and not w10795;
w10797 <= w4718 and not w10777;
w10798 <= not w10787 and w10797;
w10799 <= not w10796 and not w10798;
w10800 <= not w10789 and not w10799;
w10801 <= not w4386 and not w10800;
w10802 <= not w10277 and w10284;
w10803 <= not w10286 and w10802;
w10804 <= not w10627 and w10803;
w10805 <= not w10277 and not w10286;
w10806 <= not w10627 and w10805;
w10807 <= not w10284 and not w10806;
w10808 <= not w10804 and not w10807;
w10809 <= w4386 and not w10789;
w10810 <= not w10799 and w10809;
w10811 <= not w10808 and not w10810;
w10812 <= not w10801 and not w10811;
w10813 <= not w4066 and not w10812;
w10814 <= w10296 and not w10298;
w10815 <= not w10289 and w10814;
w10816 <= not w10627 and w10815;
w10817 <= not w10289 and not w10298;
w10818 <= not w10627 and w10817;
w10819 <= not w10296 and not w10818;
w10820 <= not w10816 and not w10819;
w10821 <= w4066 and not w10801;
w10822 <= not w10811 and w10821;
w10823 <= not w10820 and not w10822;
w10824 <= not w10813 and not w10823;
w10825 <= not w3758 and not w10824;
w10826 <= not w10301 and w10308;
w10827 <= not w10310 and w10826;
w10828 <= not w10627 and w10827;
w10829 <= not w10301 and not w10310;
w10830 <= not w10627 and w10829;
w10831 <= not w10308 and not w10830;
w10832 <= not w10828 and not w10831;
w10833 <= w3758 and not w10813;
w10834 <= not w10823 and w10833;
w10835 <= not w10832 and not w10834;
w10836 <= not w10825 and not w10835;
w10837 <= not w3462 and not w10836;
w10838 <= w10320 and not w10322;
w10839 <= not w10313 and w10838;
w10840 <= not w10627 and w10839;
w10841 <= not w10313 and not w10322;
w10842 <= not w10627 and w10841;
w10843 <= not w10320 and not w10842;
w10844 <= not w10840 and not w10843;
w10845 <= w3462 and not w10825;
w10846 <= not w10835 and w10845;
w10847 <= not w10844 and not w10846;
w10848 <= not w10837 and not w10847;
w10849 <= not w3178 and not w10848;
w10850 <= not w10325 and w10332;
w10851 <= not w10334 and w10850;
w10852 <= not w10627 and w10851;
w10853 <= not w10325 and not w10334;
w10854 <= not w10627 and w10853;
w10855 <= not w10332 and not w10854;
w10856 <= not w10852 and not w10855;
w10857 <= w3178 and not w10837;
w10858 <= not w10847 and w10857;
w10859 <= not w10856 and not w10858;
w10860 <= not w10849 and not w10859;
w10861 <= not w2906 and not w10860;
w10862 <= w10344 and not w10346;
w10863 <= not w10337 and w10862;
w10864 <= not w10627 and w10863;
w10865 <= not w10337 and not w10346;
w10866 <= not w10627 and w10865;
w10867 <= not w10344 and not w10866;
w10868 <= not w10864 and not w10867;
w10869 <= w2906 and not w10849;
w10870 <= not w10859 and w10869;
w10871 <= not w10868 and not w10870;
w10872 <= not w10861 and not w10871;
w10873 <= not w2646 and not w10872;
w10874 <= w2646 and not w10861;
w10875 <= not w10871 and w10874;
w10876 <= not w10349 and w10358;
w10877 <= not w10351 and w10876;
w10878 <= not w10627 and w10877;
w10879 <= not w10349 and not w10351;
w10880 <= not w10627 and w10879;
w10881 <= not w10358 and not w10880;
w10882 <= not w10878 and not w10881;
w10883 <= not w10875 and not w10882;
w10884 <= not w10873 and not w10883;
w10885 <= not w2398 and not w10884;
w10886 <= w10368 and not w10370;
w10887 <= not w10361 and w10886;
w10888 <= not w10627 and w10887;
w10889 <= not w10361 and not w10370;
w10890 <= not w10627 and w10889;
w10891 <= not w10368 and not w10890;
w10892 <= not w10888 and not w10891;
w10893 <= w2398 and not w10873;
w10894 <= not w10883 and w10893;
w10895 <= not w10892 and not w10894;
w10896 <= not w10885 and not w10895;
w10897 <= not w2162 and not w10896;
w10898 <= not w10373 and w10380;
w10899 <= not w10382 and w10898;
w10900 <= not w10627 and w10899;
w10901 <= not w10373 and not w10382;
w10902 <= not w10627 and w10901;
w10903 <= not w10380 and not w10902;
w10904 <= not w10900 and not w10903;
w10905 <= w2162 and not w10885;
w10906 <= not w10895 and w10905;
w10907 <= not w10904 and not w10906;
w10908 <= not w10897 and not w10907;
w10909 <= not w1938 and not w10908;
w10910 <= w10392 and not w10394;
w10911 <= not w10385 and w10910;
w10912 <= not w10627 and w10911;
w10913 <= not w10385 and not w10394;
w10914 <= not w10627 and w10913;
w10915 <= not w10392 and not w10914;
w10916 <= not w10912 and not w10915;
w10917 <= w1938 and not w10897;
w10918 <= not w10907 and w10917;
w10919 <= not w10916 and not w10918;
w10920 <= not w10909 and not w10919;
w10921 <= not w1725 and not w10920;
w10922 <= not w10397 and w10404;
w10923 <= not w10406 and w10922;
w10924 <= not w10627 and w10923;
w10925 <= not w10397 and not w10406;
w10926 <= not w10627 and w10925;
w10927 <= not w10404 and not w10926;
w10928 <= not w10924 and not w10927;
w10929 <= w1725 and not w10909;
w10930 <= not w10919 and w10929;
w10931 <= not w10928 and not w10930;
w10932 <= not w10921 and not w10931;
w10933 <= not w1525 and not w10932;
w10934 <= w10416 and not w10418;
w10935 <= not w10409 and w10934;
w10936 <= not w10627 and w10935;
w10937 <= not w10409 and not w10418;
w10938 <= not w10627 and w10937;
w10939 <= not w10416 and not w10938;
w10940 <= not w10936 and not w10939;
w10941 <= w1525 and not w10921;
w10942 <= not w10931 and w10941;
w10943 <= not w10940 and not w10942;
w10944 <= not w10933 and not w10943;
w10945 <= not w1337 and not w10944;
w10946 <= not w10421 and w10428;
w10947 <= not w10430 and w10946;
w10948 <= not w10627 and w10947;
w10949 <= not w10421 and not w10430;
w10950 <= not w10627 and w10949;
w10951 <= not w10428 and not w10950;
w10952 <= not w10948 and not w10951;
w10953 <= w1337 and not w10933;
w10954 <= not w10943 and w10953;
w10955 <= not w10952 and not w10954;
w10956 <= not w10945 and not w10955;
w10957 <= not w1161 and not w10956;
w10958 <= w10440 and not w10442;
w10959 <= not w10433 and w10958;
w10960 <= not w10627 and w10959;
w10961 <= not w10433 and not w10442;
w10962 <= not w10627 and w10961;
w10963 <= not w10440 and not w10962;
w10964 <= not w10960 and not w10963;
w10965 <= w1161 and not w10945;
w10966 <= not w10955 and w10965;
w10967 <= not w10964 and not w10966;
w10968 <= not w10957 and not w10967;
w10969 <= not w997 and not w10968;
w10970 <= not w10445 and w10452;
w10971 <= not w10454 and w10970;
w10972 <= not w10627 and w10971;
w10973 <= not w10445 and not w10454;
w10974 <= not w10627 and w10973;
w10975 <= not w10452 and not w10974;
w10976 <= not w10972 and not w10975;
w10977 <= w997 and not w10957;
w10978 <= not w10967 and w10977;
w10979 <= not w10976 and not w10978;
w10980 <= not w10969 and not w10979;
w10981 <= not w845 and not w10980;
w10982 <= w10464 and not w10466;
w10983 <= not w10457 and w10982;
w10984 <= not w10627 and w10983;
w10985 <= not w10457 and not w10466;
w10986 <= not w10627 and w10985;
w10987 <= not w10464 and not w10986;
w10988 <= not w10984 and not w10987;
w10989 <= w845 and not w10969;
w10990 <= not w10979 and w10989;
w10991 <= not w10988 and not w10990;
w10992 <= not w10981 and not w10991;
w10993 <= not w705 and not w10992;
w10994 <= not w10469 and w10476;
w10995 <= not w10478 and w10994;
w10996 <= not w10627 and w10995;
w10997 <= not w10469 and not w10478;
w10998 <= not w10627 and w10997;
w10999 <= not w10476 and not w10998;
w11000 <= not w10996 and not w10999;
w11001 <= w705 and not w10981;
w11002 <= not w10991 and w11001;
w11003 <= not w11000 and not w11002;
w11004 <= not w10993 and not w11003;
w11005 <= not w577 and not w11004;
w11006 <= w10488 and not w10490;
w11007 <= not w10481 and w11006;
w11008 <= not w10627 and w11007;
w11009 <= not w10481 and not w10490;
w11010 <= not w10627 and w11009;
w11011 <= not w10488 and not w11010;
w11012 <= not w11008 and not w11011;
w11013 <= w577 and not w10993;
w11014 <= not w11003 and w11013;
w11015 <= not w11012 and not w11014;
w11016 <= not w11005 and not w11015;
w11017 <= not w460 and not w11016;
w11018 <= not w10493 and w10500;
w11019 <= not w10502 and w11018;
w11020 <= not w10627 and w11019;
w11021 <= not w10493 and not w10502;
w11022 <= not w10627 and w11021;
w11023 <= not w10500 and not w11022;
w11024 <= not w11020 and not w11023;
w11025 <= w460 and not w11005;
w11026 <= not w11015 and w11025;
w11027 <= not w11024 and not w11026;
w11028 <= not w11017 and not w11027;
w11029 <= not w356 and not w11028;
w11030 <= w10512 and not w10514;
w11031 <= not w10505 and w11030;
w11032 <= not w10627 and w11031;
w11033 <= not w10505 and not w10514;
w11034 <= not w10627 and w11033;
w11035 <= not w10512 and not w11034;
w11036 <= not w11032 and not w11035;
w11037 <= w356 and not w11017;
w11038 <= not w11027 and w11037;
w11039 <= not w11036 and not w11038;
w11040 <= not w11029 and not w11039;
w11041 <= not w264 and not w11040;
w11042 <= not w10517 and w10524;
w11043 <= not w10526 and w11042;
w11044 <= not w10627 and w11043;
w11045 <= not w10517 and not w10526;
w11046 <= not w10627 and w11045;
w11047 <= not w10524 and not w11046;
w11048 <= not w11044 and not w11047;
w11049 <= w264 and not w11029;
w11050 <= not w11039 and w11049;
w11051 <= not w11048 and not w11050;
w11052 <= not w11041 and not w11051;
w11053 <= not w184 and not w11052;
w11054 <= w10536 and not w10538;
w11055 <= not w10529 and w11054;
w11056 <= not w10627 and w11055;
w11057 <= not w10529 and not w10538;
w11058 <= not w10627 and w11057;
w11059 <= not w10536 and not w11058;
w11060 <= not w11056 and not w11059;
w11061 <= w184 and not w11041;
w11062 <= not w11051 and w11061;
w11063 <= not w11060 and not w11062;
w11064 <= not w11053 and not w11063;
w11065 <= not w115 and not w11064;
w11066 <= not w10541 and w10548;
w11067 <= not w10550 and w11066;
w11068 <= not w10627 and w11067;
w11069 <= not w10541 and not w10550;
w11070 <= not w10627 and w11069;
w11071 <= not w10548 and not w11070;
w11072 <= not w11068 and not w11071;
w11073 <= w115 and not w11053;
w11074 <= not w11063 and w11073;
w11075 <= not w11072 and not w11074;
w11076 <= not w11065 and not w11075;
w11077 <= not w60 and not w11076;
w11078 <= w10560 and not w10562;
w11079 <= not w10553 and w11078;
w11080 <= not w10627 and w11079;
w11081 <= not w10553 and not w10562;
w11082 <= not w10627 and w11081;
w11083 <= not w10560 and not w11082;
w11084 <= not w11080 and not w11083;
w11085 <= w60 and not w11065;
w11086 <= not w11075 and w11085;
w11087 <= not w11084 and not w11086;
w11088 <= not w11077 and not w11087;
w11089 <= not w22 and not w11088;
w11090 <= not w10565 and w10572;
w11091 <= not w10574 and w11090;
w11092 <= not w10627 and w11091;
w11093 <= not w10565 and not w10574;
w11094 <= not w10627 and w11093;
w11095 <= not w10572 and not w11094;
w11096 <= not w11092 and not w11095;
w11097 <= w22 and not w11077;
w11098 <= not w11087 and w11097;
w11099 <= not w11096 and not w11098;
w11100 <= not w11089 and not w11099;
w11101 <= not w5 and not w11100;
w11102 <= w10584 and not w10586;
w11103 <= not w10577 and w11102;
w11104 <= not w10627 and w11103;
w11105 <= not w10577 and not w10586;
w11106 <= not w10627 and w11105;
w11107 <= not w10584 and not w11106;
w11108 <= not w11104 and not w11107;
w11109 <= w5 and not w11089;
w11110 <= not w11099 and w11109;
w11111 <= not w11108 and not w11110;
w11112 <= not w11101 and not w11111;
w11113 <= not w10589 and w10596;
w11114 <= not w10598 and w11113;
w11115 <= not w10627 and w11114;
w11116 <= not w10589 and not w10598;
w11117 <= not w10627 and w11116;
w11118 <= not w10596 and not w11117;
w11119 <= not w11115 and not w11118;
w11120 <= not w10600 and not w10607;
w11121 <= not w10627 and w11120;
w11122 <= not w10615 and not w11121;
w11123 <= not w11119 and w11122;
w11124 <= not w11112 and w11123;
w11125 <= w0 and not w11124;
w11126 <= not w11101 and w11119;
w11127 <= not w11111 and w11126;
w11128 <= not w10607 and not w10627;
w11129 <= w10600 and not w11128;
w11130 <= not w0 and not w11120;
w11131 <= not w11129 and w11130;
w11132 <= not w10603 and not w10624;
w11133 <= not w10606 and w11132;
w11134 <= not w10619 and w11133;
w11135 <= not w10615 and w11134;
w11136 <= not w10613 and w11135;
w11137 <= not w11131 and not w11136;
w11138 <= not w11127 and w11137;
w11139 <= not w11125 and w11138;
w11140 <= a(42) and not w11139;
w11141 <= not a(40) and not a(41);
w11142 <= not a(42) and w11141;
w11143 <= not w11140 and not w11142;
w11144 <= not w10627 and not w11143;
w11145 <= not w10624 and not w11142;
w11146 <= not w10619 and w11145;
w11147 <= not w10615 and w11146;
w11148 <= not w10613 and w11147;
w11149 <= not w11140 and w11148;
w11150 <= not a(42) and not w11139;
w11151 <= a(43) and not w11150;
w11152 <= w10629 and not w11139;
w11153 <= not w11151 and not w11152;
w11154 <= not w11149 and w11153;
w11155 <= not w11144 and not w11154;
w11156 <= not w10127 and not w11155;
w11157 <= w10127 and not w11144;
w11158 <= not w11154 and w11157;
w11159 <= not w10627 and not w11136;
w11160 <= not w11131 and w11159;
w11161 <= not w11127 and w11160;
w11162 <= not w11125 and w11161;
w11163 <= not w11152 and not w11162;
w11164 <= a(44) and not w11163;
w11165 <= not a(44) and not w11162;
w11166 <= not w11152 and w11165;
w11167 <= not w11164 and not w11166;
w11168 <= not w11158 and not w11167;
w11169 <= not w11156 and not w11168;
w11170 <= not w9639 and not w11169;
w11171 <= not w10632 and not w10637;
w11172 <= not w10641 and w11171;
w11173 <= not w11139 and w11172;
w11174 <= not w11139 and w11171;
w11175 <= w10641 and not w11174;
w11176 <= not w11173 and not w11175;
w11177 <= w9639 and not w11156;
w11178 <= not w11168 and w11177;
w11179 <= not w11176 and not w11178;
w11180 <= not w11170 and not w11179;
w11181 <= not w9163 and not w11180;
w11182 <= not w10646 and w10655;
w11183 <= not w10644 and w11182;
w11184 <= not w11139 and w11183;
w11185 <= not w10644 and not w10646;
w11186 <= not w11139 and w11185;
w11187 <= not w10655 and not w11186;
w11188 <= not w11184 and not w11187;
w11189 <= w9163 and not w11170;
w11190 <= not w11179 and w11189;
w11191 <= not w11188 and not w11190;
w11192 <= not w11181 and not w11191;
w11193 <= not w8699 and not w11192;
w11194 <= not w10658 and w10664;
w11195 <= not w10666 and w11194;
w11196 <= not w11139 and w11195;
w11197 <= not w10658 and not w10666;
w11198 <= not w11139 and w11197;
w11199 <= not w10664 and not w11198;
w11200 <= not w11196 and not w11199;
w11201 <= w8699 and not w11181;
w11202 <= not w11191 and w11201;
w11203 <= not w11200 and not w11202;
w11204 <= not w11193 and not w11203;
w11205 <= not w8247 and not w11204;
w11206 <= w10676 and not w10678;
w11207 <= not w10669 and w11206;
w11208 <= not w11139 and w11207;
w11209 <= not w10669 and not w10678;
w11210 <= not w11139 and w11209;
w11211 <= not w10676 and not w11210;
w11212 <= not w11208 and not w11211;
w11213 <= w8247 and not w11193;
w11214 <= not w11203 and w11213;
w11215 <= not w11212 and not w11214;
w11216 <= not w11205 and not w11215;
w11217 <= not w7807 and not w11216;
w11218 <= not w10681 and w10688;
w11219 <= not w10690 and w11218;
w11220 <= not w11139 and w11219;
w11221 <= not w10681 and not w10690;
w11222 <= not w11139 and w11221;
w11223 <= not w10688 and not w11222;
w11224 <= not w11220 and not w11223;
w11225 <= w7807 and not w11205;
w11226 <= not w11215 and w11225;
w11227 <= not w11224 and not w11226;
w11228 <= not w11217 and not w11227;
w11229 <= not w7379 and not w11228;
w11230 <= w10700 and not w10702;
w11231 <= not w10693 and w11230;
w11232 <= not w11139 and w11231;
w11233 <= not w10693 and not w10702;
w11234 <= not w11139 and w11233;
w11235 <= not w10700 and not w11234;
w11236 <= not w11232 and not w11235;
w11237 <= w7379 and not w11217;
w11238 <= not w11227 and w11237;
w11239 <= not w11236 and not w11238;
w11240 <= not w11229 and not w11239;
w11241 <= not w6963 and not w11240;
w11242 <= not w10705 and w10712;
w11243 <= not w10714 and w11242;
w11244 <= not w11139 and w11243;
w11245 <= not w10705 and not w10714;
w11246 <= not w11139 and w11245;
w11247 <= not w10712 and not w11246;
w11248 <= not w11244 and not w11247;
w11249 <= w6963 and not w11229;
w11250 <= not w11239 and w11249;
w11251 <= not w11248 and not w11250;
w11252 <= not w11241 and not w11251;
w11253 <= not w6558 and not w11252;
w11254 <= w10724 and not w10726;
w11255 <= not w10717 and w11254;
w11256 <= not w11139 and w11255;
w11257 <= not w10717 and not w10726;
w11258 <= not w11139 and w11257;
w11259 <= not w10724 and not w11258;
w11260 <= not w11256 and not w11259;
w11261 <= w6558 and not w11241;
w11262 <= not w11251 and w11261;
w11263 <= not w11260 and not w11262;
w11264 <= not w11253 and not w11263;
w11265 <= not w6166 and not w11264;
w11266 <= not w10729 and w10736;
w11267 <= not w10738 and w11266;
w11268 <= not w11139 and w11267;
w11269 <= not w10729 and not w10738;
w11270 <= not w11139 and w11269;
w11271 <= not w10736 and not w11270;
w11272 <= not w11268 and not w11271;
w11273 <= w6166 and not w11253;
w11274 <= not w11263 and w11273;
w11275 <= not w11272 and not w11274;
w11276 <= not w11265 and not w11275;
w11277 <= not w5786 and not w11276;
w11278 <= w10748 and not w10750;
w11279 <= not w10741 and w11278;
w11280 <= not w11139 and w11279;
w11281 <= not w10741 and not w10750;
w11282 <= not w11139 and w11281;
w11283 <= not w10748 and not w11282;
w11284 <= not w11280 and not w11283;
w11285 <= w5786 and not w11265;
w11286 <= not w11275 and w11285;
w11287 <= not w11284 and not w11286;
w11288 <= not w11277 and not w11287;
w11289 <= not w5418 and not w11288;
w11290 <= not w10753 and w10760;
w11291 <= not w10762 and w11290;
w11292 <= not w11139 and w11291;
w11293 <= not w10753 and not w10762;
w11294 <= not w11139 and w11293;
w11295 <= not w10760 and not w11294;
w11296 <= not w11292 and not w11295;
w11297 <= w5418 and not w11277;
w11298 <= not w11287 and w11297;
w11299 <= not w11296 and not w11298;
w11300 <= not w11289 and not w11299;
w11301 <= not w5062 and not w11300;
w11302 <= w10772 and not w10774;
w11303 <= not w10765 and w11302;
w11304 <= not w11139 and w11303;
w11305 <= not w10765 and not w10774;
w11306 <= not w11139 and w11305;
w11307 <= not w10772 and not w11306;
w11308 <= not w11304 and not w11307;
w11309 <= w5062 and not w11289;
w11310 <= not w11299 and w11309;
w11311 <= not w11308 and not w11310;
w11312 <= not w11301 and not w11311;
w11313 <= not w4718 and not w11312;
w11314 <= not w10777 and w10784;
w11315 <= not w10786 and w11314;
w11316 <= not w11139 and w11315;
w11317 <= not w10777 and not w10786;
w11318 <= not w11139 and w11317;
w11319 <= not w10784 and not w11318;
w11320 <= not w11316 and not w11319;
w11321 <= w4718 and not w11301;
w11322 <= not w11311 and w11321;
w11323 <= not w11320 and not w11322;
w11324 <= not w11313 and not w11323;
w11325 <= not w4386 and not w11324;
w11326 <= w10796 and not w10798;
w11327 <= not w10789 and w11326;
w11328 <= not w11139 and w11327;
w11329 <= not w10789 and not w10798;
w11330 <= not w11139 and w11329;
w11331 <= not w10796 and not w11330;
w11332 <= not w11328 and not w11331;
w11333 <= w4386 and not w11313;
w11334 <= not w11323 and w11333;
w11335 <= not w11332 and not w11334;
w11336 <= not w11325 and not w11335;
w11337 <= not w4066 and not w11336;
w11338 <= not w10801 and w10808;
w11339 <= not w10810 and w11338;
w11340 <= not w11139 and w11339;
w11341 <= not w10801 and not w10810;
w11342 <= not w11139 and w11341;
w11343 <= not w10808 and not w11342;
w11344 <= not w11340 and not w11343;
w11345 <= w4066 and not w11325;
w11346 <= not w11335 and w11345;
w11347 <= not w11344 and not w11346;
w11348 <= not w11337 and not w11347;
w11349 <= not w3758 and not w11348;
w11350 <= w10820 and not w10822;
w11351 <= not w10813 and w11350;
w11352 <= not w11139 and w11351;
w11353 <= not w10813 and not w10822;
w11354 <= not w11139 and w11353;
w11355 <= not w10820 and not w11354;
w11356 <= not w11352 and not w11355;
w11357 <= w3758 and not w11337;
w11358 <= not w11347 and w11357;
w11359 <= not w11356 and not w11358;
w11360 <= not w11349 and not w11359;
w11361 <= not w3462 and not w11360;
w11362 <= not w10825 and w10832;
w11363 <= not w10834 and w11362;
w11364 <= not w11139 and w11363;
w11365 <= not w10825 and not w10834;
w11366 <= not w11139 and w11365;
w11367 <= not w10832 and not w11366;
w11368 <= not w11364 and not w11367;
w11369 <= w3462 and not w11349;
w11370 <= not w11359 and w11369;
w11371 <= not w11368 and not w11370;
w11372 <= not w11361 and not w11371;
w11373 <= not w3178 and not w11372;
w11374 <= w10844 and not w10846;
w11375 <= not w10837 and w11374;
w11376 <= not w11139 and w11375;
w11377 <= not w10837 and not w10846;
w11378 <= not w11139 and w11377;
w11379 <= not w10844 and not w11378;
w11380 <= not w11376 and not w11379;
w11381 <= w3178 and not w11361;
w11382 <= not w11371 and w11381;
w11383 <= not w11380 and not w11382;
w11384 <= not w11373 and not w11383;
w11385 <= not w2906 and not w11384;
w11386 <= not w10849 and w10856;
w11387 <= not w10858 and w11386;
w11388 <= not w11139 and w11387;
w11389 <= not w10849 and not w10858;
w11390 <= not w11139 and w11389;
w11391 <= not w10856 and not w11390;
w11392 <= not w11388 and not w11391;
w11393 <= w2906 and not w11373;
w11394 <= not w11383 and w11393;
w11395 <= not w11392 and not w11394;
w11396 <= not w11385 and not w11395;
w11397 <= not w2646 and not w11396;
w11398 <= w10868 and not w10870;
w11399 <= not w10861 and w11398;
w11400 <= not w11139 and w11399;
w11401 <= not w10861 and not w10870;
w11402 <= not w11139 and w11401;
w11403 <= not w10868 and not w11402;
w11404 <= not w11400 and not w11403;
w11405 <= w2646 and not w11385;
w11406 <= not w11395 and w11405;
w11407 <= not w11404 and not w11406;
w11408 <= not w11397 and not w11407;
w11409 <= not w2398 and not w11408;
w11410 <= w2398 and not w11397;
w11411 <= not w11407 and w11410;
w11412 <= not w10873 and w10882;
w11413 <= not w10875 and w11412;
w11414 <= not w11139 and w11413;
w11415 <= not w10873 and not w10875;
w11416 <= not w11139 and w11415;
w11417 <= not w10882 and not w11416;
w11418 <= not w11414 and not w11417;
w11419 <= not w11411 and not w11418;
w11420 <= not w11409 and not w11419;
w11421 <= not w2162 and not w11420;
w11422 <= w10892 and not w10894;
w11423 <= not w10885 and w11422;
w11424 <= not w11139 and w11423;
w11425 <= not w10885 and not w10894;
w11426 <= not w11139 and w11425;
w11427 <= not w10892 and not w11426;
w11428 <= not w11424 and not w11427;
w11429 <= w2162 and not w11409;
w11430 <= not w11419 and w11429;
w11431 <= not w11428 and not w11430;
w11432 <= not w11421 and not w11431;
w11433 <= not w1938 and not w11432;
w11434 <= not w10897 and w10904;
w11435 <= not w10906 and w11434;
w11436 <= not w11139 and w11435;
w11437 <= not w10897 and not w10906;
w11438 <= not w11139 and w11437;
w11439 <= not w10904 and not w11438;
w11440 <= not w11436 and not w11439;
w11441 <= w1938 and not w11421;
w11442 <= not w11431 and w11441;
w11443 <= not w11440 and not w11442;
w11444 <= not w11433 and not w11443;
w11445 <= not w1725 and not w11444;
w11446 <= w10916 and not w10918;
w11447 <= not w10909 and w11446;
w11448 <= not w11139 and w11447;
w11449 <= not w10909 and not w10918;
w11450 <= not w11139 and w11449;
w11451 <= not w10916 and not w11450;
w11452 <= not w11448 and not w11451;
w11453 <= w1725 and not w11433;
w11454 <= not w11443 and w11453;
w11455 <= not w11452 and not w11454;
w11456 <= not w11445 and not w11455;
w11457 <= not w1525 and not w11456;
w11458 <= not w10921 and w10928;
w11459 <= not w10930 and w11458;
w11460 <= not w11139 and w11459;
w11461 <= not w10921 and not w10930;
w11462 <= not w11139 and w11461;
w11463 <= not w10928 and not w11462;
w11464 <= not w11460 and not w11463;
w11465 <= w1525 and not w11445;
w11466 <= not w11455 and w11465;
w11467 <= not w11464 and not w11466;
w11468 <= not w11457 and not w11467;
w11469 <= not w1337 and not w11468;
w11470 <= w10940 and not w10942;
w11471 <= not w10933 and w11470;
w11472 <= not w11139 and w11471;
w11473 <= not w10933 and not w10942;
w11474 <= not w11139 and w11473;
w11475 <= not w10940 and not w11474;
w11476 <= not w11472 and not w11475;
w11477 <= w1337 and not w11457;
w11478 <= not w11467 and w11477;
w11479 <= not w11476 and not w11478;
w11480 <= not w11469 and not w11479;
w11481 <= not w1161 and not w11480;
w11482 <= not w10945 and w10952;
w11483 <= not w10954 and w11482;
w11484 <= not w11139 and w11483;
w11485 <= not w10945 and not w10954;
w11486 <= not w11139 and w11485;
w11487 <= not w10952 and not w11486;
w11488 <= not w11484 and not w11487;
w11489 <= w1161 and not w11469;
w11490 <= not w11479 and w11489;
w11491 <= not w11488 and not w11490;
w11492 <= not w11481 and not w11491;
w11493 <= not w997 and not w11492;
w11494 <= w10964 and not w10966;
w11495 <= not w10957 and w11494;
w11496 <= not w11139 and w11495;
w11497 <= not w10957 and not w10966;
w11498 <= not w11139 and w11497;
w11499 <= not w10964 and not w11498;
w11500 <= not w11496 and not w11499;
w11501 <= w997 and not w11481;
w11502 <= not w11491 and w11501;
w11503 <= not w11500 and not w11502;
w11504 <= not w11493 and not w11503;
w11505 <= not w845 and not w11504;
w11506 <= not w10969 and w10976;
w11507 <= not w10978 and w11506;
w11508 <= not w11139 and w11507;
w11509 <= not w10969 and not w10978;
w11510 <= not w11139 and w11509;
w11511 <= not w10976 and not w11510;
w11512 <= not w11508 and not w11511;
w11513 <= w845 and not w11493;
w11514 <= not w11503 and w11513;
w11515 <= not w11512 and not w11514;
w11516 <= not w11505 and not w11515;
w11517 <= not w705 and not w11516;
w11518 <= w10988 and not w10990;
w11519 <= not w10981 and w11518;
w11520 <= not w11139 and w11519;
w11521 <= not w10981 and not w10990;
w11522 <= not w11139 and w11521;
w11523 <= not w10988 and not w11522;
w11524 <= not w11520 and not w11523;
w11525 <= w705 and not w11505;
w11526 <= not w11515 and w11525;
w11527 <= not w11524 and not w11526;
w11528 <= not w11517 and not w11527;
w11529 <= not w577 and not w11528;
w11530 <= not w10993 and w11000;
w11531 <= not w11002 and w11530;
w11532 <= not w11139 and w11531;
w11533 <= not w10993 and not w11002;
w11534 <= not w11139 and w11533;
w11535 <= not w11000 and not w11534;
w11536 <= not w11532 and not w11535;
w11537 <= w577 and not w11517;
w11538 <= not w11527 and w11537;
w11539 <= not w11536 and not w11538;
w11540 <= not w11529 and not w11539;
w11541 <= not w460 and not w11540;
w11542 <= w11012 and not w11014;
w11543 <= not w11005 and w11542;
w11544 <= not w11139 and w11543;
w11545 <= not w11005 and not w11014;
w11546 <= not w11139 and w11545;
w11547 <= not w11012 and not w11546;
w11548 <= not w11544 and not w11547;
w11549 <= w460 and not w11529;
w11550 <= not w11539 and w11549;
w11551 <= not w11548 and not w11550;
w11552 <= not w11541 and not w11551;
w11553 <= not w356 and not w11552;
w11554 <= not w11017 and w11024;
w11555 <= not w11026 and w11554;
w11556 <= not w11139 and w11555;
w11557 <= not w11017 and not w11026;
w11558 <= not w11139 and w11557;
w11559 <= not w11024 and not w11558;
w11560 <= not w11556 and not w11559;
w11561 <= w356 and not w11541;
w11562 <= not w11551 and w11561;
w11563 <= not w11560 and not w11562;
w11564 <= not w11553 and not w11563;
w11565 <= not w264 and not w11564;
w11566 <= w11036 and not w11038;
w11567 <= not w11029 and w11566;
w11568 <= not w11139 and w11567;
w11569 <= not w11029 and not w11038;
w11570 <= not w11139 and w11569;
w11571 <= not w11036 and not w11570;
w11572 <= not w11568 and not w11571;
w11573 <= w264 and not w11553;
w11574 <= not w11563 and w11573;
w11575 <= not w11572 and not w11574;
w11576 <= not w11565 and not w11575;
w11577 <= not w184 and not w11576;
w11578 <= not w11041 and w11048;
w11579 <= not w11050 and w11578;
w11580 <= not w11139 and w11579;
w11581 <= not w11041 and not w11050;
w11582 <= not w11139 and w11581;
w11583 <= not w11048 and not w11582;
w11584 <= not w11580 and not w11583;
w11585 <= w184 and not w11565;
w11586 <= not w11575 and w11585;
w11587 <= not w11584 and not w11586;
w11588 <= not w11577 and not w11587;
w11589 <= not w115 and not w11588;
w11590 <= w11060 and not w11062;
w11591 <= not w11053 and w11590;
w11592 <= not w11139 and w11591;
w11593 <= not w11053 and not w11062;
w11594 <= not w11139 and w11593;
w11595 <= not w11060 and not w11594;
w11596 <= not w11592 and not w11595;
w11597 <= w115 and not w11577;
w11598 <= not w11587 and w11597;
w11599 <= not w11596 and not w11598;
w11600 <= not w11589 and not w11599;
w11601 <= not w60 and not w11600;
w11602 <= not w11065 and w11072;
w11603 <= not w11074 and w11602;
w11604 <= not w11139 and w11603;
w11605 <= not w11065 and not w11074;
w11606 <= not w11139 and w11605;
w11607 <= not w11072 and not w11606;
w11608 <= not w11604 and not w11607;
w11609 <= w60 and not w11589;
w11610 <= not w11599 and w11609;
w11611 <= not w11608 and not w11610;
w11612 <= not w11601 and not w11611;
w11613 <= not w22 and not w11612;
w11614 <= w11084 and not w11086;
w11615 <= not w11077 and w11614;
w11616 <= not w11139 and w11615;
w11617 <= not w11077 and not w11086;
w11618 <= not w11139 and w11617;
w11619 <= not w11084 and not w11618;
w11620 <= not w11616 and not w11619;
w11621 <= w22 and not w11601;
w11622 <= not w11611 and w11621;
w11623 <= not w11620 and not w11622;
w11624 <= not w11613 and not w11623;
w11625 <= not w5 and not w11624;
w11626 <= not w11089 and w11096;
w11627 <= not w11098 and w11626;
w11628 <= not w11139 and w11627;
w11629 <= not w11089 and not w11098;
w11630 <= not w11139 and w11629;
w11631 <= not w11096 and not w11630;
w11632 <= not w11628 and not w11631;
w11633 <= w5 and not w11613;
w11634 <= not w11623 and w11633;
w11635 <= not w11632 and not w11634;
w11636 <= not w11625 and not w11635;
w11637 <= w11108 and not w11110;
w11638 <= not w11101 and w11637;
w11639 <= not w11139 and w11638;
w11640 <= not w11101 and not w11110;
w11641 <= not w11139 and w11640;
w11642 <= not w11108 and not w11641;
w11643 <= not w11639 and not w11642;
w11644 <= not w11112 and not w11119;
w11645 <= not w11139 and w11644;
w11646 <= not w11127 and not w11645;
w11647 <= not w11643 and w11646;
w11648 <= not w11636 and w11647;
w11649 <= w0 and not w11648;
w11650 <= not w11625 and w11643;
w11651 <= not w11635 and w11650;
w11652 <= not w11119 and not w11139;
w11653 <= w11112 and not w11652;
w11654 <= not w0 and not w11644;
w11655 <= not w11653 and w11654;
w11656 <= not w11115 and not w11136;
w11657 <= not w11118 and w11656;
w11658 <= not w11131 and w11657;
w11659 <= not w11127 and w11658;
w11660 <= not w11125 and w11659;
w11661 <= not w11655 and not w11660;
w11662 <= not w11651 and w11661;
w11663 <= not w11649 and w11662;
w11664 <= a(40) and not w11663;
w11665 <= not a(38) and not a(39);
w11666 <= not a(40) and w11665;
w11667 <= not w11664 and not w11666;
w11668 <= not w11139 and not w11667;
w11669 <= not w11136 and not w11666;
w11670 <= not w11131 and w11669;
w11671 <= not w11127 and w11670;
w11672 <= not w11125 and w11671;
w11673 <= not w11664 and w11672;
w11674 <= not a(40) and not w11663;
w11675 <= a(41) and not w11674;
w11676 <= w11141 and not w11663;
w11677 <= not w11675 and not w11676;
w11678 <= not w11673 and w11677;
w11679 <= not w11668 and not w11678;
w11680 <= not w10627 and not w11679;
w11681 <= w10627 and not w11668;
w11682 <= not w11678 and w11681;
w11683 <= not w11139 and not w11660;
w11684 <= not w11655 and w11683;
w11685 <= not w11651 and w11684;
w11686 <= not w11649 and w11685;
w11687 <= not w11676 and not w11686;
w11688 <= a(42) and not w11687;
w11689 <= not a(42) and not w11686;
w11690 <= not w11676 and w11689;
w11691 <= not w11688 and not w11690;
w11692 <= not w11682 and not w11691;
w11693 <= not w11680 and not w11692;
w11694 <= not w10127 and not w11693;
w11695 <= not w11144 and not w11149;
w11696 <= not w11153 and w11695;
w11697 <= not w11663 and w11696;
w11698 <= not w11663 and w11695;
w11699 <= w11153 and not w11698;
w11700 <= not w11697 and not w11699;
w11701 <= w10127 and not w11680;
w11702 <= not w11692 and w11701;
w11703 <= not w11700 and not w11702;
w11704 <= not w11694 and not w11703;
w11705 <= not w9639 and not w11704;
w11706 <= not w11158 and w11167;
w11707 <= not w11156 and w11706;
w11708 <= not w11663 and w11707;
w11709 <= not w11156 and not w11158;
w11710 <= not w11663 and w11709;
w11711 <= not w11167 and not w11710;
w11712 <= not w11708 and not w11711;
w11713 <= w9639 and not w11694;
w11714 <= not w11703 and w11713;
w11715 <= not w11712 and not w11714;
w11716 <= not w11705 and not w11715;
w11717 <= not w9163 and not w11716;
w11718 <= not w11170 and w11176;
w11719 <= not w11178 and w11718;
w11720 <= not w11663 and w11719;
w11721 <= not w11170 and not w11178;
w11722 <= not w11663 and w11721;
w11723 <= not w11176 and not w11722;
w11724 <= not w11720 and not w11723;
w11725 <= w9163 and not w11705;
w11726 <= not w11715 and w11725;
w11727 <= not w11724 and not w11726;
w11728 <= not w11717 and not w11727;
w11729 <= not w8699 and not w11728;
w11730 <= w11188 and not w11190;
w11731 <= not w11181 and w11730;
w11732 <= not w11663 and w11731;
w11733 <= not w11181 and not w11190;
w11734 <= not w11663 and w11733;
w11735 <= not w11188 and not w11734;
w11736 <= not w11732 and not w11735;
w11737 <= w8699 and not w11717;
w11738 <= not w11727 and w11737;
w11739 <= not w11736 and not w11738;
w11740 <= not w11729 and not w11739;
w11741 <= not w8247 and not w11740;
w11742 <= not w11193 and w11200;
w11743 <= not w11202 and w11742;
w11744 <= not w11663 and w11743;
w11745 <= not w11193 and not w11202;
w11746 <= not w11663 and w11745;
w11747 <= not w11200 and not w11746;
w11748 <= not w11744 and not w11747;
w11749 <= w8247 and not w11729;
w11750 <= not w11739 and w11749;
w11751 <= not w11748 and not w11750;
w11752 <= not w11741 and not w11751;
w11753 <= not w7807 and not w11752;
w11754 <= w11212 and not w11214;
w11755 <= not w11205 and w11754;
w11756 <= not w11663 and w11755;
w11757 <= not w11205 and not w11214;
w11758 <= not w11663 and w11757;
w11759 <= not w11212 and not w11758;
w11760 <= not w11756 and not w11759;
w11761 <= w7807 and not w11741;
w11762 <= not w11751 and w11761;
w11763 <= not w11760 and not w11762;
w11764 <= not w11753 and not w11763;
w11765 <= not w7379 and not w11764;
w11766 <= not w11217 and w11224;
w11767 <= not w11226 and w11766;
w11768 <= not w11663 and w11767;
w11769 <= not w11217 and not w11226;
w11770 <= not w11663 and w11769;
w11771 <= not w11224 and not w11770;
w11772 <= not w11768 and not w11771;
w11773 <= w7379 and not w11753;
w11774 <= not w11763 and w11773;
w11775 <= not w11772 and not w11774;
w11776 <= not w11765 and not w11775;
w11777 <= not w6963 and not w11776;
w11778 <= w11236 and not w11238;
w11779 <= not w11229 and w11778;
w11780 <= not w11663 and w11779;
w11781 <= not w11229 and not w11238;
w11782 <= not w11663 and w11781;
w11783 <= not w11236 and not w11782;
w11784 <= not w11780 and not w11783;
w11785 <= w6963 and not w11765;
w11786 <= not w11775 and w11785;
w11787 <= not w11784 and not w11786;
w11788 <= not w11777 and not w11787;
w11789 <= not w6558 and not w11788;
w11790 <= not w11241 and w11248;
w11791 <= not w11250 and w11790;
w11792 <= not w11663 and w11791;
w11793 <= not w11241 and not w11250;
w11794 <= not w11663 and w11793;
w11795 <= not w11248 and not w11794;
w11796 <= not w11792 and not w11795;
w11797 <= w6558 and not w11777;
w11798 <= not w11787 and w11797;
w11799 <= not w11796 and not w11798;
w11800 <= not w11789 and not w11799;
w11801 <= not w6166 and not w11800;
w11802 <= w11260 and not w11262;
w11803 <= not w11253 and w11802;
w11804 <= not w11663 and w11803;
w11805 <= not w11253 and not w11262;
w11806 <= not w11663 and w11805;
w11807 <= not w11260 and not w11806;
w11808 <= not w11804 and not w11807;
w11809 <= w6166 and not w11789;
w11810 <= not w11799 and w11809;
w11811 <= not w11808 and not w11810;
w11812 <= not w11801 and not w11811;
w11813 <= not w5786 and not w11812;
w11814 <= not w11265 and w11272;
w11815 <= not w11274 and w11814;
w11816 <= not w11663 and w11815;
w11817 <= not w11265 and not w11274;
w11818 <= not w11663 and w11817;
w11819 <= not w11272 and not w11818;
w11820 <= not w11816 and not w11819;
w11821 <= w5786 and not w11801;
w11822 <= not w11811 and w11821;
w11823 <= not w11820 and not w11822;
w11824 <= not w11813 and not w11823;
w11825 <= not w5418 and not w11824;
w11826 <= w11284 and not w11286;
w11827 <= not w11277 and w11826;
w11828 <= not w11663 and w11827;
w11829 <= not w11277 and not w11286;
w11830 <= not w11663 and w11829;
w11831 <= not w11284 and not w11830;
w11832 <= not w11828 and not w11831;
w11833 <= w5418 and not w11813;
w11834 <= not w11823 and w11833;
w11835 <= not w11832 and not w11834;
w11836 <= not w11825 and not w11835;
w11837 <= not w5062 and not w11836;
w11838 <= not w11289 and w11296;
w11839 <= not w11298 and w11838;
w11840 <= not w11663 and w11839;
w11841 <= not w11289 and not w11298;
w11842 <= not w11663 and w11841;
w11843 <= not w11296 and not w11842;
w11844 <= not w11840 and not w11843;
w11845 <= w5062 and not w11825;
w11846 <= not w11835 and w11845;
w11847 <= not w11844 and not w11846;
w11848 <= not w11837 and not w11847;
w11849 <= not w4718 and not w11848;
w11850 <= w11308 and not w11310;
w11851 <= not w11301 and w11850;
w11852 <= not w11663 and w11851;
w11853 <= not w11301 and not w11310;
w11854 <= not w11663 and w11853;
w11855 <= not w11308 and not w11854;
w11856 <= not w11852 and not w11855;
w11857 <= w4718 and not w11837;
w11858 <= not w11847 and w11857;
w11859 <= not w11856 and not w11858;
w11860 <= not w11849 and not w11859;
w11861 <= not w4386 and not w11860;
w11862 <= not w11313 and w11320;
w11863 <= not w11322 and w11862;
w11864 <= not w11663 and w11863;
w11865 <= not w11313 and not w11322;
w11866 <= not w11663 and w11865;
w11867 <= not w11320 and not w11866;
w11868 <= not w11864 and not w11867;
w11869 <= w4386 and not w11849;
w11870 <= not w11859 and w11869;
w11871 <= not w11868 and not w11870;
w11872 <= not w11861 and not w11871;
w11873 <= not w4066 and not w11872;
w11874 <= w11332 and not w11334;
w11875 <= not w11325 and w11874;
w11876 <= not w11663 and w11875;
w11877 <= not w11325 and not w11334;
w11878 <= not w11663 and w11877;
w11879 <= not w11332 and not w11878;
w11880 <= not w11876 and not w11879;
w11881 <= w4066 and not w11861;
w11882 <= not w11871 and w11881;
w11883 <= not w11880 and not w11882;
w11884 <= not w11873 and not w11883;
w11885 <= not w3758 and not w11884;
w11886 <= not w11337 and w11344;
w11887 <= not w11346 and w11886;
w11888 <= not w11663 and w11887;
w11889 <= not w11337 and not w11346;
w11890 <= not w11663 and w11889;
w11891 <= not w11344 and not w11890;
w11892 <= not w11888 and not w11891;
w11893 <= w3758 and not w11873;
w11894 <= not w11883 and w11893;
w11895 <= not w11892 and not w11894;
w11896 <= not w11885 and not w11895;
w11897 <= not w3462 and not w11896;
w11898 <= w11356 and not w11358;
w11899 <= not w11349 and w11898;
w11900 <= not w11663 and w11899;
w11901 <= not w11349 and not w11358;
w11902 <= not w11663 and w11901;
w11903 <= not w11356 and not w11902;
w11904 <= not w11900 and not w11903;
w11905 <= w3462 and not w11885;
w11906 <= not w11895 and w11905;
w11907 <= not w11904 and not w11906;
w11908 <= not w11897 and not w11907;
w11909 <= not w3178 and not w11908;
w11910 <= not w11361 and w11368;
w11911 <= not w11370 and w11910;
w11912 <= not w11663 and w11911;
w11913 <= not w11361 and not w11370;
w11914 <= not w11663 and w11913;
w11915 <= not w11368 and not w11914;
w11916 <= not w11912 and not w11915;
w11917 <= w3178 and not w11897;
w11918 <= not w11907 and w11917;
w11919 <= not w11916 and not w11918;
w11920 <= not w11909 and not w11919;
w11921 <= not w2906 and not w11920;
w11922 <= w11380 and not w11382;
w11923 <= not w11373 and w11922;
w11924 <= not w11663 and w11923;
w11925 <= not w11373 and not w11382;
w11926 <= not w11663 and w11925;
w11927 <= not w11380 and not w11926;
w11928 <= not w11924 and not w11927;
w11929 <= w2906 and not w11909;
w11930 <= not w11919 and w11929;
w11931 <= not w11928 and not w11930;
w11932 <= not w11921 and not w11931;
w11933 <= not w2646 and not w11932;
w11934 <= not w11385 and w11392;
w11935 <= not w11394 and w11934;
w11936 <= not w11663 and w11935;
w11937 <= not w11385 and not w11394;
w11938 <= not w11663 and w11937;
w11939 <= not w11392 and not w11938;
w11940 <= not w11936 and not w11939;
w11941 <= w2646 and not w11921;
w11942 <= not w11931 and w11941;
w11943 <= not w11940 and not w11942;
w11944 <= not w11933 and not w11943;
w11945 <= not w2398 and not w11944;
w11946 <= w11404 and not w11406;
w11947 <= not w11397 and w11946;
w11948 <= not w11663 and w11947;
w11949 <= not w11397 and not w11406;
w11950 <= not w11663 and w11949;
w11951 <= not w11404 and not w11950;
w11952 <= not w11948 and not w11951;
w11953 <= w2398 and not w11933;
w11954 <= not w11943 and w11953;
w11955 <= not w11952 and not w11954;
w11956 <= not w11945 and not w11955;
w11957 <= not w2162 and not w11956;
w11958 <= w2162 and not w11945;
w11959 <= not w11955 and w11958;
w11960 <= not w11409 and w11418;
w11961 <= not w11411 and w11960;
w11962 <= not w11663 and w11961;
w11963 <= not w11409 and not w11411;
w11964 <= not w11663 and w11963;
w11965 <= not w11418 and not w11964;
w11966 <= not w11962 and not w11965;
w11967 <= not w11959 and not w11966;
w11968 <= not w11957 and not w11967;
w11969 <= not w1938 and not w11968;
w11970 <= w11428 and not w11430;
w11971 <= not w11421 and w11970;
w11972 <= not w11663 and w11971;
w11973 <= not w11421 and not w11430;
w11974 <= not w11663 and w11973;
w11975 <= not w11428 and not w11974;
w11976 <= not w11972 and not w11975;
w11977 <= w1938 and not w11957;
w11978 <= not w11967 and w11977;
w11979 <= not w11976 and not w11978;
w11980 <= not w11969 and not w11979;
w11981 <= not w1725 and not w11980;
w11982 <= not w11433 and w11440;
w11983 <= not w11442 and w11982;
w11984 <= not w11663 and w11983;
w11985 <= not w11433 and not w11442;
w11986 <= not w11663 and w11985;
w11987 <= not w11440 and not w11986;
w11988 <= not w11984 and not w11987;
w11989 <= w1725 and not w11969;
w11990 <= not w11979 and w11989;
w11991 <= not w11988 and not w11990;
w11992 <= not w11981 and not w11991;
w11993 <= not w1525 and not w11992;
w11994 <= w11452 and not w11454;
w11995 <= not w11445 and w11994;
w11996 <= not w11663 and w11995;
w11997 <= not w11445 and not w11454;
w11998 <= not w11663 and w11997;
w11999 <= not w11452 and not w11998;
w12000 <= not w11996 and not w11999;
w12001 <= w1525 and not w11981;
w12002 <= not w11991 and w12001;
w12003 <= not w12000 and not w12002;
w12004 <= not w11993 and not w12003;
w12005 <= not w1337 and not w12004;
w12006 <= not w11457 and w11464;
w12007 <= not w11466 and w12006;
w12008 <= not w11663 and w12007;
w12009 <= not w11457 and not w11466;
w12010 <= not w11663 and w12009;
w12011 <= not w11464 and not w12010;
w12012 <= not w12008 and not w12011;
w12013 <= w1337 and not w11993;
w12014 <= not w12003 and w12013;
w12015 <= not w12012 and not w12014;
w12016 <= not w12005 and not w12015;
w12017 <= not w1161 and not w12016;
w12018 <= w11476 and not w11478;
w12019 <= not w11469 and w12018;
w12020 <= not w11663 and w12019;
w12021 <= not w11469 and not w11478;
w12022 <= not w11663 and w12021;
w12023 <= not w11476 and not w12022;
w12024 <= not w12020 and not w12023;
w12025 <= w1161 and not w12005;
w12026 <= not w12015 and w12025;
w12027 <= not w12024 and not w12026;
w12028 <= not w12017 and not w12027;
w12029 <= not w997 and not w12028;
w12030 <= not w11481 and w11488;
w12031 <= not w11490 and w12030;
w12032 <= not w11663 and w12031;
w12033 <= not w11481 and not w11490;
w12034 <= not w11663 and w12033;
w12035 <= not w11488 and not w12034;
w12036 <= not w12032 and not w12035;
w12037 <= w997 and not w12017;
w12038 <= not w12027 and w12037;
w12039 <= not w12036 and not w12038;
w12040 <= not w12029 and not w12039;
w12041 <= not w845 and not w12040;
w12042 <= w11500 and not w11502;
w12043 <= not w11493 and w12042;
w12044 <= not w11663 and w12043;
w12045 <= not w11493 and not w11502;
w12046 <= not w11663 and w12045;
w12047 <= not w11500 and not w12046;
w12048 <= not w12044 and not w12047;
w12049 <= w845 and not w12029;
w12050 <= not w12039 and w12049;
w12051 <= not w12048 and not w12050;
w12052 <= not w12041 and not w12051;
w12053 <= not w705 and not w12052;
w12054 <= not w11505 and w11512;
w12055 <= not w11514 and w12054;
w12056 <= not w11663 and w12055;
w12057 <= not w11505 and not w11514;
w12058 <= not w11663 and w12057;
w12059 <= not w11512 and not w12058;
w12060 <= not w12056 and not w12059;
w12061 <= w705 and not w12041;
w12062 <= not w12051 and w12061;
w12063 <= not w12060 and not w12062;
w12064 <= not w12053 and not w12063;
w12065 <= not w577 and not w12064;
w12066 <= w11524 and not w11526;
w12067 <= not w11517 and w12066;
w12068 <= not w11663 and w12067;
w12069 <= not w11517 and not w11526;
w12070 <= not w11663 and w12069;
w12071 <= not w11524 and not w12070;
w12072 <= not w12068 and not w12071;
w12073 <= w577 and not w12053;
w12074 <= not w12063 and w12073;
w12075 <= not w12072 and not w12074;
w12076 <= not w12065 and not w12075;
w12077 <= not w460 and not w12076;
w12078 <= not w11529 and w11536;
w12079 <= not w11538 and w12078;
w12080 <= not w11663 and w12079;
w12081 <= not w11529 and not w11538;
w12082 <= not w11663 and w12081;
w12083 <= not w11536 and not w12082;
w12084 <= not w12080 and not w12083;
w12085 <= w460 and not w12065;
w12086 <= not w12075 and w12085;
w12087 <= not w12084 and not w12086;
w12088 <= not w12077 and not w12087;
w12089 <= not w356 and not w12088;
w12090 <= w11548 and not w11550;
w12091 <= not w11541 and w12090;
w12092 <= not w11663 and w12091;
w12093 <= not w11541 and not w11550;
w12094 <= not w11663 and w12093;
w12095 <= not w11548 and not w12094;
w12096 <= not w12092 and not w12095;
w12097 <= w356 and not w12077;
w12098 <= not w12087 and w12097;
w12099 <= not w12096 and not w12098;
w12100 <= not w12089 and not w12099;
w12101 <= not w264 and not w12100;
w12102 <= not w11553 and w11560;
w12103 <= not w11562 and w12102;
w12104 <= not w11663 and w12103;
w12105 <= not w11553 and not w11562;
w12106 <= not w11663 and w12105;
w12107 <= not w11560 and not w12106;
w12108 <= not w12104 and not w12107;
w12109 <= w264 and not w12089;
w12110 <= not w12099 and w12109;
w12111 <= not w12108 and not w12110;
w12112 <= not w12101 and not w12111;
w12113 <= not w184 and not w12112;
w12114 <= w11572 and not w11574;
w12115 <= not w11565 and w12114;
w12116 <= not w11663 and w12115;
w12117 <= not w11565 and not w11574;
w12118 <= not w11663 and w12117;
w12119 <= not w11572 and not w12118;
w12120 <= not w12116 and not w12119;
w12121 <= w184 and not w12101;
w12122 <= not w12111 and w12121;
w12123 <= not w12120 and not w12122;
w12124 <= not w12113 and not w12123;
w12125 <= not w115 and not w12124;
w12126 <= not w11577 and w11584;
w12127 <= not w11586 and w12126;
w12128 <= not w11663 and w12127;
w12129 <= not w11577 and not w11586;
w12130 <= not w11663 and w12129;
w12131 <= not w11584 and not w12130;
w12132 <= not w12128 and not w12131;
w12133 <= w115 and not w12113;
w12134 <= not w12123 and w12133;
w12135 <= not w12132 and not w12134;
w12136 <= not w12125 and not w12135;
w12137 <= not w60 and not w12136;
w12138 <= w11596 and not w11598;
w12139 <= not w11589 and w12138;
w12140 <= not w11663 and w12139;
w12141 <= not w11589 and not w11598;
w12142 <= not w11663 and w12141;
w12143 <= not w11596 and not w12142;
w12144 <= not w12140 and not w12143;
w12145 <= w60 and not w12125;
w12146 <= not w12135 and w12145;
w12147 <= not w12144 and not w12146;
w12148 <= not w12137 and not w12147;
w12149 <= not w22 and not w12148;
w12150 <= not w11601 and w11608;
w12151 <= not w11610 and w12150;
w12152 <= not w11663 and w12151;
w12153 <= not w11601 and not w11610;
w12154 <= not w11663 and w12153;
w12155 <= not w11608 and not w12154;
w12156 <= not w12152 and not w12155;
w12157 <= w22 and not w12137;
w12158 <= not w12147 and w12157;
w12159 <= not w12156 and not w12158;
w12160 <= not w12149 and not w12159;
w12161 <= not w5 and not w12160;
w12162 <= w11620 and not w11622;
w12163 <= not w11613 and w12162;
w12164 <= not w11663 and w12163;
w12165 <= not w11613 and not w11622;
w12166 <= not w11663 and w12165;
w12167 <= not w11620 and not w12166;
w12168 <= not w12164 and not w12167;
w12169 <= w5 and not w12149;
w12170 <= not w12159 and w12169;
w12171 <= not w12168 and not w12170;
w12172 <= not w12161 and not w12171;
w12173 <= not w11625 and w11632;
w12174 <= not w11634 and w12173;
w12175 <= not w11663 and w12174;
w12176 <= not w11625 and not w11634;
w12177 <= not w11663 and w12176;
w12178 <= not w11632 and not w12177;
w12179 <= not w12175 and not w12178;
w12180 <= not w11636 and not w11643;
w12181 <= not w11663 and w12180;
w12182 <= not w11651 and not w12181;
w12183 <= not w12179 and w12182;
w12184 <= not w12172 and w12183;
w12185 <= w0 and not w12184;
w12186 <= not w12161 and w12179;
w12187 <= not w12171 and w12186;
w12188 <= not w11643 and not w11663;
w12189 <= w11636 and not w12188;
w12190 <= not w0 and not w12180;
w12191 <= not w12189 and w12190;
w12192 <= not w11639 and not w11660;
w12193 <= not w11642 and w12192;
w12194 <= not w11655 and w12193;
w12195 <= not w11651 and w12194;
w12196 <= not w11649 and w12195;
w12197 <= not w12191 and not w12196;
w12198 <= not w12187 and w12197;
w12199 <= not w12185 and w12198;
w12200 <= a(38) and not w12199;
w12201 <= not a(36) and not a(37);
w12202 <= not a(38) and w12201;
w12203 <= not w12200 and not w12202;
w12204 <= not w11663 and not w12203;
w12205 <= not w11660 and not w12202;
w12206 <= not w11655 and w12205;
w12207 <= not w11651 and w12206;
w12208 <= not w11649 and w12207;
w12209 <= not w12200 and w12208;
w12210 <= not a(38) and not w12199;
w12211 <= a(39) and not w12210;
w12212 <= w11665 and not w12199;
w12213 <= not w12211 and not w12212;
w12214 <= not w12209 and w12213;
w12215 <= not w12204 and not w12214;
w12216 <= not w11139 and not w12215;
w12217 <= w11139 and not w12204;
w12218 <= not w12214 and w12217;
w12219 <= not w11663 and not w12196;
w12220 <= not w12191 and w12219;
w12221 <= not w12187 and w12220;
w12222 <= not w12185 and w12221;
w12223 <= not w12212 and not w12222;
w12224 <= a(40) and not w12223;
w12225 <= not a(40) and not w12222;
w12226 <= not w12212 and w12225;
w12227 <= not w12224 and not w12226;
w12228 <= not w12218 and not w12227;
w12229 <= not w12216 and not w12228;
w12230 <= not w10627 and not w12229;
w12231 <= not w11668 and not w11673;
w12232 <= not w11677 and w12231;
w12233 <= not w12199 and w12232;
w12234 <= not w12199 and w12231;
w12235 <= w11677 and not w12234;
w12236 <= not w12233 and not w12235;
w12237 <= w10627 and not w12216;
w12238 <= not w12228 and w12237;
w12239 <= not w12236 and not w12238;
w12240 <= not w12230 and not w12239;
w12241 <= not w10127 and not w12240;
w12242 <= not w11682 and w11691;
w12243 <= not w11680 and w12242;
w12244 <= not w12199 and w12243;
w12245 <= not w11680 and not w11682;
w12246 <= not w12199 and w12245;
w12247 <= not w11691 and not w12246;
w12248 <= not w12244 and not w12247;
w12249 <= w10127 and not w12230;
w12250 <= not w12239 and w12249;
w12251 <= not w12248 and not w12250;
w12252 <= not w12241 and not w12251;
w12253 <= not w9639 and not w12252;
w12254 <= not w11694 and w11700;
w12255 <= not w11702 and w12254;
w12256 <= not w12199 and w12255;
w12257 <= not w11694 and not w11702;
w12258 <= not w12199 and w12257;
w12259 <= not w11700 and not w12258;
w12260 <= not w12256 and not w12259;
w12261 <= w9639 and not w12241;
w12262 <= not w12251 and w12261;
w12263 <= not w12260 and not w12262;
w12264 <= not w12253 and not w12263;
w12265 <= not w9163 and not w12264;
w12266 <= w11712 and not w11714;
w12267 <= not w11705 and w12266;
w12268 <= not w12199 and w12267;
w12269 <= not w11705 and not w11714;
w12270 <= not w12199 and w12269;
w12271 <= not w11712 and not w12270;
w12272 <= not w12268 and not w12271;
w12273 <= w9163 and not w12253;
w12274 <= not w12263 and w12273;
w12275 <= not w12272 and not w12274;
w12276 <= not w12265 and not w12275;
w12277 <= not w8699 and not w12276;
w12278 <= not w11717 and w11724;
w12279 <= not w11726 and w12278;
w12280 <= not w12199 and w12279;
w12281 <= not w11717 and not w11726;
w12282 <= not w12199 and w12281;
w12283 <= not w11724 and not w12282;
w12284 <= not w12280 and not w12283;
w12285 <= w8699 and not w12265;
w12286 <= not w12275 and w12285;
w12287 <= not w12284 and not w12286;
w12288 <= not w12277 and not w12287;
w12289 <= not w8247 and not w12288;
w12290 <= w11736 and not w11738;
w12291 <= not w11729 and w12290;
w12292 <= not w12199 and w12291;
w12293 <= not w11729 and not w11738;
w12294 <= not w12199 and w12293;
w12295 <= not w11736 and not w12294;
w12296 <= not w12292 and not w12295;
w12297 <= w8247 and not w12277;
w12298 <= not w12287 and w12297;
w12299 <= not w12296 and not w12298;
w12300 <= not w12289 and not w12299;
w12301 <= not w7807 and not w12300;
w12302 <= not w11741 and w11748;
w12303 <= not w11750 and w12302;
w12304 <= not w12199 and w12303;
w12305 <= not w11741 and not w11750;
w12306 <= not w12199 and w12305;
w12307 <= not w11748 and not w12306;
w12308 <= not w12304 and not w12307;
w12309 <= w7807 and not w12289;
w12310 <= not w12299 and w12309;
w12311 <= not w12308 and not w12310;
w12312 <= not w12301 and not w12311;
w12313 <= not w7379 and not w12312;
w12314 <= w11760 and not w11762;
w12315 <= not w11753 and w12314;
w12316 <= not w12199 and w12315;
w12317 <= not w11753 and not w11762;
w12318 <= not w12199 and w12317;
w12319 <= not w11760 and not w12318;
w12320 <= not w12316 and not w12319;
w12321 <= w7379 and not w12301;
w12322 <= not w12311 and w12321;
w12323 <= not w12320 and not w12322;
w12324 <= not w12313 and not w12323;
w12325 <= not w6963 and not w12324;
w12326 <= not w11765 and w11772;
w12327 <= not w11774 and w12326;
w12328 <= not w12199 and w12327;
w12329 <= not w11765 and not w11774;
w12330 <= not w12199 and w12329;
w12331 <= not w11772 and not w12330;
w12332 <= not w12328 and not w12331;
w12333 <= w6963 and not w12313;
w12334 <= not w12323 and w12333;
w12335 <= not w12332 and not w12334;
w12336 <= not w12325 and not w12335;
w12337 <= not w6558 and not w12336;
w12338 <= w11784 and not w11786;
w12339 <= not w11777 and w12338;
w12340 <= not w12199 and w12339;
w12341 <= not w11777 and not w11786;
w12342 <= not w12199 and w12341;
w12343 <= not w11784 and not w12342;
w12344 <= not w12340 and not w12343;
w12345 <= w6558 and not w12325;
w12346 <= not w12335 and w12345;
w12347 <= not w12344 and not w12346;
w12348 <= not w12337 and not w12347;
w12349 <= not w6166 and not w12348;
w12350 <= not w11789 and w11796;
w12351 <= not w11798 and w12350;
w12352 <= not w12199 and w12351;
w12353 <= not w11789 and not w11798;
w12354 <= not w12199 and w12353;
w12355 <= not w11796 and not w12354;
w12356 <= not w12352 and not w12355;
w12357 <= w6166 and not w12337;
w12358 <= not w12347 and w12357;
w12359 <= not w12356 and not w12358;
w12360 <= not w12349 and not w12359;
w12361 <= not w5786 and not w12360;
w12362 <= w11808 and not w11810;
w12363 <= not w11801 and w12362;
w12364 <= not w12199 and w12363;
w12365 <= not w11801 and not w11810;
w12366 <= not w12199 and w12365;
w12367 <= not w11808 and not w12366;
w12368 <= not w12364 and not w12367;
w12369 <= w5786 and not w12349;
w12370 <= not w12359 and w12369;
w12371 <= not w12368 and not w12370;
w12372 <= not w12361 and not w12371;
w12373 <= not w5418 and not w12372;
w12374 <= not w11813 and w11820;
w12375 <= not w11822 and w12374;
w12376 <= not w12199 and w12375;
w12377 <= not w11813 and not w11822;
w12378 <= not w12199 and w12377;
w12379 <= not w11820 and not w12378;
w12380 <= not w12376 and not w12379;
w12381 <= w5418 and not w12361;
w12382 <= not w12371 and w12381;
w12383 <= not w12380 and not w12382;
w12384 <= not w12373 and not w12383;
w12385 <= not w5062 and not w12384;
w12386 <= w11832 and not w11834;
w12387 <= not w11825 and w12386;
w12388 <= not w12199 and w12387;
w12389 <= not w11825 and not w11834;
w12390 <= not w12199 and w12389;
w12391 <= not w11832 and not w12390;
w12392 <= not w12388 and not w12391;
w12393 <= w5062 and not w12373;
w12394 <= not w12383 and w12393;
w12395 <= not w12392 and not w12394;
w12396 <= not w12385 and not w12395;
w12397 <= not w4718 and not w12396;
w12398 <= not w11837 and w11844;
w12399 <= not w11846 and w12398;
w12400 <= not w12199 and w12399;
w12401 <= not w11837 and not w11846;
w12402 <= not w12199 and w12401;
w12403 <= not w11844 and not w12402;
w12404 <= not w12400 and not w12403;
w12405 <= w4718 and not w12385;
w12406 <= not w12395 and w12405;
w12407 <= not w12404 and not w12406;
w12408 <= not w12397 and not w12407;
w12409 <= not w4386 and not w12408;
w12410 <= w11856 and not w11858;
w12411 <= not w11849 and w12410;
w12412 <= not w12199 and w12411;
w12413 <= not w11849 and not w11858;
w12414 <= not w12199 and w12413;
w12415 <= not w11856 and not w12414;
w12416 <= not w12412 and not w12415;
w12417 <= w4386 and not w12397;
w12418 <= not w12407 and w12417;
w12419 <= not w12416 and not w12418;
w12420 <= not w12409 and not w12419;
w12421 <= not w4066 and not w12420;
w12422 <= not w11861 and w11868;
w12423 <= not w11870 and w12422;
w12424 <= not w12199 and w12423;
w12425 <= not w11861 and not w11870;
w12426 <= not w12199 and w12425;
w12427 <= not w11868 and not w12426;
w12428 <= not w12424 and not w12427;
w12429 <= w4066 and not w12409;
w12430 <= not w12419 and w12429;
w12431 <= not w12428 and not w12430;
w12432 <= not w12421 and not w12431;
w12433 <= not w3758 and not w12432;
w12434 <= w11880 and not w11882;
w12435 <= not w11873 and w12434;
w12436 <= not w12199 and w12435;
w12437 <= not w11873 and not w11882;
w12438 <= not w12199 and w12437;
w12439 <= not w11880 and not w12438;
w12440 <= not w12436 and not w12439;
w12441 <= w3758 and not w12421;
w12442 <= not w12431 and w12441;
w12443 <= not w12440 and not w12442;
w12444 <= not w12433 and not w12443;
w12445 <= not w3462 and not w12444;
w12446 <= not w11885 and w11892;
w12447 <= not w11894 and w12446;
w12448 <= not w12199 and w12447;
w12449 <= not w11885 and not w11894;
w12450 <= not w12199 and w12449;
w12451 <= not w11892 and not w12450;
w12452 <= not w12448 and not w12451;
w12453 <= w3462 and not w12433;
w12454 <= not w12443 and w12453;
w12455 <= not w12452 and not w12454;
w12456 <= not w12445 and not w12455;
w12457 <= not w3178 and not w12456;
w12458 <= w11904 and not w11906;
w12459 <= not w11897 and w12458;
w12460 <= not w12199 and w12459;
w12461 <= not w11897 and not w11906;
w12462 <= not w12199 and w12461;
w12463 <= not w11904 and not w12462;
w12464 <= not w12460 and not w12463;
w12465 <= w3178 and not w12445;
w12466 <= not w12455 and w12465;
w12467 <= not w12464 and not w12466;
w12468 <= not w12457 and not w12467;
w12469 <= not w2906 and not w12468;
w12470 <= not w11909 and w11916;
w12471 <= not w11918 and w12470;
w12472 <= not w12199 and w12471;
w12473 <= not w11909 and not w11918;
w12474 <= not w12199 and w12473;
w12475 <= not w11916 and not w12474;
w12476 <= not w12472 and not w12475;
w12477 <= w2906 and not w12457;
w12478 <= not w12467 and w12477;
w12479 <= not w12476 and not w12478;
w12480 <= not w12469 and not w12479;
w12481 <= not w2646 and not w12480;
w12482 <= w11928 and not w11930;
w12483 <= not w11921 and w12482;
w12484 <= not w12199 and w12483;
w12485 <= not w11921 and not w11930;
w12486 <= not w12199 and w12485;
w12487 <= not w11928 and not w12486;
w12488 <= not w12484 and not w12487;
w12489 <= w2646 and not w12469;
w12490 <= not w12479 and w12489;
w12491 <= not w12488 and not w12490;
w12492 <= not w12481 and not w12491;
w12493 <= not w2398 and not w12492;
w12494 <= not w11933 and w11940;
w12495 <= not w11942 and w12494;
w12496 <= not w12199 and w12495;
w12497 <= not w11933 and not w11942;
w12498 <= not w12199 and w12497;
w12499 <= not w11940 and not w12498;
w12500 <= not w12496 and not w12499;
w12501 <= w2398 and not w12481;
w12502 <= not w12491 and w12501;
w12503 <= not w12500 and not w12502;
w12504 <= not w12493 and not w12503;
w12505 <= not w2162 and not w12504;
w12506 <= w11952 and not w11954;
w12507 <= not w11945 and w12506;
w12508 <= not w12199 and w12507;
w12509 <= not w11945 and not w11954;
w12510 <= not w12199 and w12509;
w12511 <= not w11952 and not w12510;
w12512 <= not w12508 and not w12511;
w12513 <= w2162 and not w12493;
w12514 <= not w12503 and w12513;
w12515 <= not w12512 and not w12514;
w12516 <= not w12505 and not w12515;
w12517 <= not w1938 and not w12516;
w12518 <= w1938 and not w12505;
w12519 <= not w12515 and w12518;
w12520 <= not w11957 and w11966;
w12521 <= not w11959 and w12520;
w12522 <= not w12199 and w12521;
w12523 <= not w11957 and not w11959;
w12524 <= not w12199 and w12523;
w12525 <= not w11966 and not w12524;
w12526 <= not w12522 and not w12525;
w12527 <= not w12519 and not w12526;
w12528 <= not w12517 and not w12527;
w12529 <= not w1725 and not w12528;
w12530 <= w11976 and not w11978;
w12531 <= not w11969 and w12530;
w12532 <= not w12199 and w12531;
w12533 <= not w11969 and not w11978;
w12534 <= not w12199 and w12533;
w12535 <= not w11976 and not w12534;
w12536 <= not w12532 and not w12535;
w12537 <= w1725 and not w12517;
w12538 <= not w12527 and w12537;
w12539 <= not w12536 and not w12538;
w12540 <= not w12529 and not w12539;
w12541 <= not w1525 and not w12540;
w12542 <= not w11981 and w11988;
w12543 <= not w11990 and w12542;
w12544 <= not w12199 and w12543;
w12545 <= not w11981 and not w11990;
w12546 <= not w12199 and w12545;
w12547 <= not w11988 and not w12546;
w12548 <= not w12544 and not w12547;
w12549 <= w1525 and not w12529;
w12550 <= not w12539 and w12549;
w12551 <= not w12548 and not w12550;
w12552 <= not w12541 and not w12551;
w12553 <= not w1337 and not w12552;
w12554 <= w12000 and not w12002;
w12555 <= not w11993 and w12554;
w12556 <= not w12199 and w12555;
w12557 <= not w11993 and not w12002;
w12558 <= not w12199 and w12557;
w12559 <= not w12000 and not w12558;
w12560 <= not w12556 and not w12559;
w12561 <= w1337 and not w12541;
w12562 <= not w12551 and w12561;
w12563 <= not w12560 and not w12562;
w12564 <= not w12553 and not w12563;
w12565 <= not w1161 and not w12564;
w12566 <= not w12005 and w12012;
w12567 <= not w12014 and w12566;
w12568 <= not w12199 and w12567;
w12569 <= not w12005 and not w12014;
w12570 <= not w12199 and w12569;
w12571 <= not w12012 and not w12570;
w12572 <= not w12568 and not w12571;
w12573 <= w1161 and not w12553;
w12574 <= not w12563 and w12573;
w12575 <= not w12572 and not w12574;
w12576 <= not w12565 and not w12575;
w12577 <= not w997 and not w12576;
w12578 <= w12024 and not w12026;
w12579 <= not w12017 and w12578;
w12580 <= not w12199 and w12579;
w12581 <= not w12017 and not w12026;
w12582 <= not w12199 and w12581;
w12583 <= not w12024 and not w12582;
w12584 <= not w12580 and not w12583;
w12585 <= w997 and not w12565;
w12586 <= not w12575 and w12585;
w12587 <= not w12584 and not w12586;
w12588 <= not w12577 and not w12587;
w12589 <= not w845 and not w12588;
w12590 <= not w12029 and w12036;
w12591 <= not w12038 and w12590;
w12592 <= not w12199 and w12591;
w12593 <= not w12029 and not w12038;
w12594 <= not w12199 and w12593;
w12595 <= not w12036 and not w12594;
w12596 <= not w12592 and not w12595;
w12597 <= w845 and not w12577;
w12598 <= not w12587 and w12597;
w12599 <= not w12596 and not w12598;
w12600 <= not w12589 and not w12599;
w12601 <= not w705 and not w12600;
w12602 <= w12048 and not w12050;
w12603 <= not w12041 and w12602;
w12604 <= not w12199 and w12603;
w12605 <= not w12041 and not w12050;
w12606 <= not w12199 and w12605;
w12607 <= not w12048 and not w12606;
w12608 <= not w12604 and not w12607;
w12609 <= w705 and not w12589;
w12610 <= not w12599 and w12609;
w12611 <= not w12608 and not w12610;
w12612 <= not w12601 and not w12611;
w12613 <= not w577 and not w12612;
w12614 <= not w12053 and w12060;
w12615 <= not w12062 and w12614;
w12616 <= not w12199 and w12615;
w12617 <= not w12053 and not w12062;
w12618 <= not w12199 and w12617;
w12619 <= not w12060 and not w12618;
w12620 <= not w12616 and not w12619;
w12621 <= w577 and not w12601;
w12622 <= not w12611 and w12621;
w12623 <= not w12620 and not w12622;
w12624 <= not w12613 and not w12623;
w12625 <= not w460 and not w12624;
w12626 <= w12072 and not w12074;
w12627 <= not w12065 and w12626;
w12628 <= not w12199 and w12627;
w12629 <= not w12065 and not w12074;
w12630 <= not w12199 and w12629;
w12631 <= not w12072 and not w12630;
w12632 <= not w12628 and not w12631;
w12633 <= w460 and not w12613;
w12634 <= not w12623 and w12633;
w12635 <= not w12632 and not w12634;
w12636 <= not w12625 and not w12635;
w12637 <= not w356 and not w12636;
w12638 <= not w12077 and w12084;
w12639 <= not w12086 and w12638;
w12640 <= not w12199 and w12639;
w12641 <= not w12077 and not w12086;
w12642 <= not w12199 and w12641;
w12643 <= not w12084 and not w12642;
w12644 <= not w12640 and not w12643;
w12645 <= w356 and not w12625;
w12646 <= not w12635 and w12645;
w12647 <= not w12644 and not w12646;
w12648 <= not w12637 and not w12647;
w12649 <= not w264 and not w12648;
w12650 <= w12096 and not w12098;
w12651 <= not w12089 and w12650;
w12652 <= not w12199 and w12651;
w12653 <= not w12089 and not w12098;
w12654 <= not w12199 and w12653;
w12655 <= not w12096 and not w12654;
w12656 <= not w12652 and not w12655;
w12657 <= w264 and not w12637;
w12658 <= not w12647 and w12657;
w12659 <= not w12656 and not w12658;
w12660 <= not w12649 and not w12659;
w12661 <= not w184 and not w12660;
w12662 <= not w12101 and w12108;
w12663 <= not w12110 and w12662;
w12664 <= not w12199 and w12663;
w12665 <= not w12101 and not w12110;
w12666 <= not w12199 and w12665;
w12667 <= not w12108 and not w12666;
w12668 <= not w12664 and not w12667;
w12669 <= w184 and not w12649;
w12670 <= not w12659 and w12669;
w12671 <= not w12668 and not w12670;
w12672 <= not w12661 and not w12671;
w12673 <= not w115 and not w12672;
w12674 <= w12120 and not w12122;
w12675 <= not w12113 and w12674;
w12676 <= not w12199 and w12675;
w12677 <= not w12113 and not w12122;
w12678 <= not w12199 and w12677;
w12679 <= not w12120 and not w12678;
w12680 <= not w12676 and not w12679;
w12681 <= w115 and not w12661;
w12682 <= not w12671 and w12681;
w12683 <= not w12680 and not w12682;
w12684 <= not w12673 and not w12683;
w12685 <= not w60 and not w12684;
w12686 <= not w12125 and w12132;
w12687 <= not w12134 and w12686;
w12688 <= not w12199 and w12687;
w12689 <= not w12125 and not w12134;
w12690 <= not w12199 and w12689;
w12691 <= not w12132 and not w12690;
w12692 <= not w12688 and not w12691;
w12693 <= w60 and not w12673;
w12694 <= not w12683 and w12693;
w12695 <= not w12692 and not w12694;
w12696 <= not w12685 and not w12695;
w12697 <= not w22 and not w12696;
w12698 <= w12144 and not w12146;
w12699 <= not w12137 and w12698;
w12700 <= not w12199 and w12699;
w12701 <= not w12137 and not w12146;
w12702 <= not w12199 and w12701;
w12703 <= not w12144 and not w12702;
w12704 <= not w12700 and not w12703;
w12705 <= w22 and not w12685;
w12706 <= not w12695 and w12705;
w12707 <= not w12704 and not w12706;
w12708 <= not w12697 and not w12707;
w12709 <= not w5 and not w12708;
w12710 <= not w12149 and w12156;
w12711 <= not w12158 and w12710;
w12712 <= not w12199 and w12711;
w12713 <= not w12149 and not w12158;
w12714 <= not w12199 and w12713;
w12715 <= not w12156 and not w12714;
w12716 <= not w12712 and not w12715;
w12717 <= w5 and not w12697;
w12718 <= not w12707 and w12717;
w12719 <= not w12716 and not w12718;
w12720 <= not w12709 and not w12719;
w12721 <= w12168 and not w12170;
w12722 <= not w12161 and w12721;
w12723 <= not w12199 and w12722;
w12724 <= not w12161 and not w12170;
w12725 <= not w12199 and w12724;
w12726 <= not w12168 and not w12725;
w12727 <= not w12723 and not w12726;
w12728 <= not w12172 and not w12179;
w12729 <= not w12199 and w12728;
w12730 <= not w12187 and not w12729;
w12731 <= not w12727 and w12730;
w12732 <= not w12720 and w12731;
w12733 <= w0 and not w12732;
w12734 <= not w12709 and w12727;
w12735 <= not w12719 and w12734;
w12736 <= not w12179 and not w12199;
w12737 <= w12172 and not w12736;
w12738 <= not w0 and not w12728;
w12739 <= not w12737 and w12738;
w12740 <= not w12175 and not w12196;
w12741 <= not w12178 and w12740;
w12742 <= not w12191 and w12741;
w12743 <= not w12187 and w12742;
w12744 <= not w12185 and w12743;
w12745 <= not w12739 and not w12744;
w12746 <= not w12735 and w12745;
w12747 <= not w12733 and w12746;
w12748 <= a(36) and not w12747;
w12749 <= not a(34) and not a(35);
w12750 <= not a(36) and w12749;
w12751 <= not w12748 and not w12750;
w12752 <= not w12199 and not w12751;
w12753 <= not w12196 and not w12750;
w12754 <= not w12191 and w12753;
w12755 <= not w12187 and w12754;
w12756 <= not w12185 and w12755;
w12757 <= not w12748 and w12756;
w12758 <= not a(36) and not w12747;
w12759 <= a(37) and not w12758;
w12760 <= w12201 and not w12747;
w12761 <= not w12759 and not w12760;
w12762 <= not w12757 and w12761;
w12763 <= not w12752 and not w12762;
w12764 <= not w11663 and not w12763;
w12765 <= w11663 and not w12752;
w12766 <= not w12762 and w12765;
w12767 <= not w12199 and not w12744;
w12768 <= not w12739 and w12767;
w12769 <= not w12735 and w12768;
w12770 <= not w12733 and w12769;
w12771 <= not w12760 and not w12770;
w12772 <= a(38) and not w12771;
w12773 <= not a(38) and not w12770;
w12774 <= not w12760 and w12773;
w12775 <= not w12772 and not w12774;
w12776 <= not w12766 and not w12775;
w12777 <= not w12764 and not w12776;
w12778 <= not w11139 and not w12777;
w12779 <= not w12204 and not w12209;
w12780 <= not w12213 and w12779;
w12781 <= not w12747 and w12780;
w12782 <= not w12747 and w12779;
w12783 <= w12213 and not w12782;
w12784 <= not w12781 and not w12783;
w12785 <= w11139 and not w12764;
w12786 <= not w12776 and w12785;
w12787 <= not w12784 and not w12786;
w12788 <= not w12778 and not w12787;
w12789 <= not w10627 and not w12788;
w12790 <= not w12218 and w12227;
w12791 <= not w12216 and w12790;
w12792 <= not w12747 and w12791;
w12793 <= not w12216 and not w12218;
w12794 <= not w12747 and w12793;
w12795 <= not w12227 and not w12794;
w12796 <= not w12792 and not w12795;
w12797 <= w10627 and not w12778;
w12798 <= not w12787 and w12797;
w12799 <= not w12796 and not w12798;
w12800 <= not w12789 and not w12799;
w12801 <= not w10127 and not w12800;
w12802 <= not w12230 and w12236;
w12803 <= not w12238 and w12802;
w12804 <= not w12747 and w12803;
w12805 <= not w12230 and not w12238;
w12806 <= not w12747 and w12805;
w12807 <= not w12236 and not w12806;
w12808 <= not w12804 and not w12807;
w12809 <= w10127 and not w12789;
w12810 <= not w12799 and w12809;
w12811 <= not w12808 and not w12810;
w12812 <= not w12801 and not w12811;
w12813 <= not w9639 and not w12812;
w12814 <= w12248 and not w12250;
w12815 <= not w12241 and w12814;
w12816 <= not w12747 and w12815;
w12817 <= not w12241 and not w12250;
w12818 <= not w12747 and w12817;
w12819 <= not w12248 and not w12818;
w12820 <= not w12816 and not w12819;
w12821 <= w9639 and not w12801;
w12822 <= not w12811 and w12821;
w12823 <= not w12820 and not w12822;
w12824 <= not w12813 and not w12823;
w12825 <= not w9163 and not w12824;
w12826 <= not w12253 and w12260;
w12827 <= not w12262 and w12826;
w12828 <= not w12747 and w12827;
w12829 <= not w12253 and not w12262;
w12830 <= not w12747 and w12829;
w12831 <= not w12260 and not w12830;
w12832 <= not w12828 and not w12831;
w12833 <= w9163 and not w12813;
w12834 <= not w12823 and w12833;
w12835 <= not w12832 and not w12834;
w12836 <= not w12825 and not w12835;
w12837 <= not w8699 and not w12836;
w12838 <= w12272 and not w12274;
w12839 <= not w12265 and w12838;
w12840 <= not w12747 and w12839;
w12841 <= not w12265 and not w12274;
w12842 <= not w12747 and w12841;
w12843 <= not w12272 and not w12842;
w12844 <= not w12840 and not w12843;
w12845 <= w8699 and not w12825;
w12846 <= not w12835 and w12845;
w12847 <= not w12844 and not w12846;
w12848 <= not w12837 and not w12847;
w12849 <= not w8247 and not w12848;
w12850 <= not w12277 and w12284;
w12851 <= not w12286 and w12850;
w12852 <= not w12747 and w12851;
w12853 <= not w12277 and not w12286;
w12854 <= not w12747 and w12853;
w12855 <= not w12284 and not w12854;
w12856 <= not w12852 and not w12855;
w12857 <= w8247 and not w12837;
w12858 <= not w12847 and w12857;
w12859 <= not w12856 and not w12858;
w12860 <= not w12849 and not w12859;
w12861 <= not w7807 and not w12860;
w12862 <= w12296 and not w12298;
w12863 <= not w12289 and w12862;
w12864 <= not w12747 and w12863;
w12865 <= not w12289 and not w12298;
w12866 <= not w12747 and w12865;
w12867 <= not w12296 and not w12866;
w12868 <= not w12864 and not w12867;
w12869 <= w7807 and not w12849;
w12870 <= not w12859 and w12869;
w12871 <= not w12868 and not w12870;
w12872 <= not w12861 and not w12871;
w12873 <= not w7379 and not w12872;
w12874 <= not w12301 and w12308;
w12875 <= not w12310 and w12874;
w12876 <= not w12747 and w12875;
w12877 <= not w12301 and not w12310;
w12878 <= not w12747 and w12877;
w12879 <= not w12308 and not w12878;
w12880 <= not w12876 and not w12879;
w12881 <= w7379 and not w12861;
w12882 <= not w12871 and w12881;
w12883 <= not w12880 and not w12882;
w12884 <= not w12873 and not w12883;
w12885 <= not w6963 and not w12884;
w12886 <= w12320 and not w12322;
w12887 <= not w12313 and w12886;
w12888 <= not w12747 and w12887;
w12889 <= not w12313 and not w12322;
w12890 <= not w12747 and w12889;
w12891 <= not w12320 and not w12890;
w12892 <= not w12888 and not w12891;
w12893 <= w6963 and not w12873;
w12894 <= not w12883 and w12893;
w12895 <= not w12892 and not w12894;
w12896 <= not w12885 and not w12895;
w12897 <= not w6558 and not w12896;
w12898 <= not w12325 and w12332;
w12899 <= not w12334 and w12898;
w12900 <= not w12747 and w12899;
w12901 <= not w12325 and not w12334;
w12902 <= not w12747 and w12901;
w12903 <= not w12332 and not w12902;
w12904 <= not w12900 and not w12903;
w12905 <= w6558 and not w12885;
w12906 <= not w12895 and w12905;
w12907 <= not w12904 and not w12906;
w12908 <= not w12897 and not w12907;
w12909 <= not w6166 and not w12908;
w12910 <= w12344 and not w12346;
w12911 <= not w12337 and w12910;
w12912 <= not w12747 and w12911;
w12913 <= not w12337 and not w12346;
w12914 <= not w12747 and w12913;
w12915 <= not w12344 and not w12914;
w12916 <= not w12912 and not w12915;
w12917 <= w6166 and not w12897;
w12918 <= not w12907 and w12917;
w12919 <= not w12916 and not w12918;
w12920 <= not w12909 and not w12919;
w12921 <= not w5786 and not w12920;
w12922 <= not w12349 and w12356;
w12923 <= not w12358 and w12922;
w12924 <= not w12747 and w12923;
w12925 <= not w12349 and not w12358;
w12926 <= not w12747 and w12925;
w12927 <= not w12356 and not w12926;
w12928 <= not w12924 and not w12927;
w12929 <= w5786 and not w12909;
w12930 <= not w12919 and w12929;
w12931 <= not w12928 and not w12930;
w12932 <= not w12921 and not w12931;
w12933 <= not w5418 and not w12932;
w12934 <= w12368 and not w12370;
w12935 <= not w12361 and w12934;
w12936 <= not w12747 and w12935;
w12937 <= not w12361 and not w12370;
w12938 <= not w12747 and w12937;
w12939 <= not w12368 and not w12938;
w12940 <= not w12936 and not w12939;
w12941 <= w5418 and not w12921;
w12942 <= not w12931 and w12941;
w12943 <= not w12940 and not w12942;
w12944 <= not w12933 and not w12943;
w12945 <= not w5062 and not w12944;
w12946 <= not w12373 and w12380;
w12947 <= not w12382 and w12946;
w12948 <= not w12747 and w12947;
w12949 <= not w12373 and not w12382;
w12950 <= not w12747 and w12949;
w12951 <= not w12380 and not w12950;
w12952 <= not w12948 and not w12951;
w12953 <= w5062 and not w12933;
w12954 <= not w12943 and w12953;
w12955 <= not w12952 and not w12954;
w12956 <= not w12945 and not w12955;
w12957 <= not w4718 and not w12956;
w12958 <= w12392 and not w12394;
w12959 <= not w12385 and w12958;
w12960 <= not w12747 and w12959;
w12961 <= not w12385 and not w12394;
w12962 <= not w12747 and w12961;
w12963 <= not w12392 and not w12962;
w12964 <= not w12960 and not w12963;
w12965 <= w4718 and not w12945;
w12966 <= not w12955 and w12965;
w12967 <= not w12964 and not w12966;
w12968 <= not w12957 and not w12967;
w12969 <= not w4386 and not w12968;
w12970 <= not w12397 and w12404;
w12971 <= not w12406 and w12970;
w12972 <= not w12747 and w12971;
w12973 <= not w12397 and not w12406;
w12974 <= not w12747 and w12973;
w12975 <= not w12404 and not w12974;
w12976 <= not w12972 and not w12975;
w12977 <= w4386 and not w12957;
w12978 <= not w12967 and w12977;
w12979 <= not w12976 and not w12978;
w12980 <= not w12969 and not w12979;
w12981 <= not w4066 and not w12980;
w12982 <= w12416 and not w12418;
w12983 <= not w12409 and w12982;
w12984 <= not w12747 and w12983;
w12985 <= not w12409 and not w12418;
w12986 <= not w12747 and w12985;
w12987 <= not w12416 and not w12986;
w12988 <= not w12984 and not w12987;
w12989 <= w4066 and not w12969;
w12990 <= not w12979 and w12989;
w12991 <= not w12988 and not w12990;
w12992 <= not w12981 and not w12991;
w12993 <= not w3758 and not w12992;
w12994 <= not w12421 and w12428;
w12995 <= not w12430 and w12994;
w12996 <= not w12747 and w12995;
w12997 <= not w12421 and not w12430;
w12998 <= not w12747 and w12997;
w12999 <= not w12428 and not w12998;
w13000 <= not w12996 and not w12999;
w13001 <= w3758 and not w12981;
w13002 <= not w12991 and w13001;
w13003 <= not w13000 and not w13002;
w13004 <= not w12993 and not w13003;
w13005 <= not w3462 and not w13004;
w13006 <= w12440 and not w12442;
w13007 <= not w12433 and w13006;
w13008 <= not w12747 and w13007;
w13009 <= not w12433 and not w12442;
w13010 <= not w12747 and w13009;
w13011 <= not w12440 and not w13010;
w13012 <= not w13008 and not w13011;
w13013 <= w3462 and not w12993;
w13014 <= not w13003 and w13013;
w13015 <= not w13012 and not w13014;
w13016 <= not w13005 and not w13015;
w13017 <= not w3178 and not w13016;
w13018 <= not w12445 and w12452;
w13019 <= not w12454 and w13018;
w13020 <= not w12747 and w13019;
w13021 <= not w12445 and not w12454;
w13022 <= not w12747 and w13021;
w13023 <= not w12452 and not w13022;
w13024 <= not w13020 and not w13023;
w13025 <= w3178 and not w13005;
w13026 <= not w13015 and w13025;
w13027 <= not w13024 and not w13026;
w13028 <= not w13017 and not w13027;
w13029 <= not w2906 and not w13028;
w13030 <= w12464 and not w12466;
w13031 <= not w12457 and w13030;
w13032 <= not w12747 and w13031;
w13033 <= not w12457 and not w12466;
w13034 <= not w12747 and w13033;
w13035 <= not w12464 and not w13034;
w13036 <= not w13032 and not w13035;
w13037 <= w2906 and not w13017;
w13038 <= not w13027 and w13037;
w13039 <= not w13036 and not w13038;
w13040 <= not w13029 and not w13039;
w13041 <= not w2646 and not w13040;
w13042 <= not w12469 and w12476;
w13043 <= not w12478 and w13042;
w13044 <= not w12747 and w13043;
w13045 <= not w12469 and not w12478;
w13046 <= not w12747 and w13045;
w13047 <= not w12476 and not w13046;
w13048 <= not w13044 and not w13047;
w13049 <= w2646 and not w13029;
w13050 <= not w13039 and w13049;
w13051 <= not w13048 and not w13050;
w13052 <= not w13041 and not w13051;
w13053 <= not w2398 and not w13052;
w13054 <= w12488 and not w12490;
w13055 <= not w12481 and w13054;
w13056 <= not w12747 and w13055;
w13057 <= not w12481 and not w12490;
w13058 <= not w12747 and w13057;
w13059 <= not w12488 and not w13058;
w13060 <= not w13056 and not w13059;
w13061 <= w2398 and not w13041;
w13062 <= not w13051 and w13061;
w13063 <= not w13060 and not w13062;
w13064 <= not w13053 and not w13063;
w13065 <= not w2162 and not w13064;
w13066 <= not w12493 and w12500;
w13067 <= not w12502 and w13066;
w13068 <= not w12747 and w13067;
w13069 <= not w12493 and not w12502;
w13070 <= not w12747 and w13069;
w13071 <= not w12500 and not w13070;
w13072 <= not w13068 and not w13071;
w13073 <= w2162 and not w13053;
w13074 <= not w13063 and w13073;
w13075 <= not w13072 and not w13074;
w13076 <= not w13065 and not w13075;
w13077 <= not w1938 and not w13076;
w13078 <= w12512 and not w12514;
w13079 <= not w12505 and w13078;
w13080 <= not w12747 and w13079;
w13081 <= not w12505 and not w12514;
w13082 <= not w12747 and w13081;
w13083 <= not w12512 and not w13082;
w13084 <= not w13080 and not w13083;
w13085 <= w1938 and not w13065;
w13086 <= not w13075 and w13085;
w13087 <= not w13084 and not w13086;
w13088 <= not w13077 and not w13087;
w13089 <= not w1725 and not w13088;
w13090 <= w1725 and not w13077;
w13091 <= not w13087 and w13090;
w13092 <= not w12517 and w12526;
w13093 <= not w12519 and w13092;
w13094 <= not w12747 and w13093;
w13095 <= not w12517 and not w12519;
w13096 <= not w12747 and w13095;
w13097 <= not w12526 and not w13096;
w13098 <= not w13094 and not w13097;
w13099 <= not w13091 and not w13098;
w13100 <= not w13089 and not w13099;
w13101 <= not w1525 and not w13100;
w13102 <= w12536 and not w12538;
w13103 <= not w12529 and w13102;
w13104 <= not w12747 and w13103;
w13105 <= not w12529 and not w12538;
w13106 <= not w12747 and w13105;
w13107 <= not w12536 and not w13106;
w13108 <= not w13104 and not w13107;
w13109 <= w1525 and not w13089;
w13110 <= not w13099 and w13109;
w13111 <= not w13108 and not w13110;
w13112 <= not w13101 and not w13111;
w13113 <= not w1337 and not w13112;
w13114 <= not w12541 and w12548;
w13115 <= not w12550 and w13114;
w13116 <= not w12747 and w13115;
w13117 <= not w12541 and not w12550;
w13118 <= not w12747 and w13117;
w13119 <= not w12548 and not w13118;
w13120 <= not w13116 and not w13119;
w13121 <= w1337 and not w13101;
w13122 <= not w13111 and w13121;
w13123 <= not w13120 and not w13122;
w13124 <= not w13113 and not w13123;
w13125 <= not w1161 and not w13124;
w13126 <= w12560 and not w12562;
w13127 <= not w12553 and w13126;
w13128 <= not w12747 and w13127;
w13129 <= not w12553 and not w12562;
w13130 <= not w12747 and w13129;
w13131 <= not w12560 and not w13130;
w13132 <= not w13128 and not w13131;
w13133 <= w1161 and not w13113;
w13134 <= not w13123 and w13133;
w13135 <= not w13132 and not w13134;
w13136 <= not w13125 and not w13135;
w13137 <= not w997 and not w13136;
w13138 <= not w12565 and w12572;
w13139 <= not w12574 and w13138;
w13140 <= not w12747 and w13139;
w13141 <= not w12565 and not w12574;
w13142 <= not w12747 and w13141;
w13143 <= not w12572 and not w13142;
w13144 <= not w13140 and not w13143;
w13145 <= w997 and not w13125;
w13146 <= not w13135 and w13145;
w13147 <= not w13144 and not w13146;
w13148 <= not w13137 and not w13147;
w13149 <= not w845 and not w13148;
w13150 <= w12584 and not w12586;
w13151 <= not w12577 and w13150;
w13152 <= not w12747 and w13151;
w13153 <= not w12577 and not w12586;
w13154 <= not w12747 and w13153;
w13155 <= not w12584 and not w13154;
w13156 <= not w13152 and not w13155;
w13157 <= w845 and not w13137;
w13158 <= not w13147 and w13157;
w13159 <= not w13156 and not w13158;
w13160 <= not w13149 and not w13159;
w13161 <= not w705 and not w13160;
w13162 <= not w12589 and w12596;
w13163 <= not w12598 and w13162;
w13164 <= not w12747 and w13163;
w13165 <= not w12589 and not w12598;
w13166 <= not w12747 and w13165;
w13167 <= not w12596 and not w13166;
w13168 <= not w13164 and not w13167;
w13169 <= w705 and not w13149;
w13170 <= not w13159 and w13169;
w13171 <= not w13168 and not w13170;
w13172 <= not w13161 and not w13171;
w13173 <= not w577 and not w13172;
w13174 <= w12608 and not w12610;
w13175 <= not w12601 and w13174;
w13176 <= not w12747 and w13175;
w13177 <= not w12601 and not w12610;
w13178 <= not w12747 and w13177;
w13179 <= not w12608 and not w13178;
w13180 <= not w13176 and not w13179;
w13181 <= w577 and not w13161;
w13182 <= not w13171 and w13181;
w13183 <= not w13180 and not w13182;
w13184 <= not w13173 and not w13183;
w13185 <= not w460 and not w13184;
w13186 <= not w12613 and w12620;
w13187 <= not w12622 and w13186;
w13188 <= not w12747 and w13187;
w13189 <= not w12613 and not w12622;
w13190 <= not w12747 and w13189;
w13191 <= not w12620 and not w13190;
w13192 <= not w13188 and not w13191;
w13193 <= w460 and not w13173;
w13194 <= not w13183 and w13193;
w13195 <= not w13192 and not w13194;
w13196 <= not w13185 and not w13195;
w13197 <= not w356 and not w13196;
w13198 <= w12632 and not w12634;
w13199 <= not w12625 and w13198;
w13200 <= not w12747 and w13199;
w13201 <= not w12625 and not w12634;
w13202 <= not w12747 and w13201;
w13203 <= not w12632 and not w13202;
w13204 <= not w13200 and not w13203;
w13205 <= w356 and not w13185;
w13206 <= not w13195 and w13205;
w13207 <= not w13204 and not w13206;
w13208 <= not w13197 and not w13207;
w13209 <= not w264 and not w13208;
w13210 <= not w12637 and w12644;
w13211 <= not w12646 and w13210;
w13212 <= not w12747 and w13211;
w13213 <= not w12637 and not w12646;
w13214 <= not w12747 and w13213;
w13215 <= not w12644 and not w13214;
w13216 <= not w13212 and not w13215;
w13217 <= w264 and not w13197;
w13218 <= not w13207 and w13217;
w13219 <= not w13216 and not w13218;
w13220 <= not w13209 and not w13219;
w13221 <= not w184 and not w13220;
w13222 <= w12656 and not w12658;
w13223 <= not w12649 and w13222;
w13224 <= not w12747 and w13223;
w13225 <= not w12649 and not w12658;
w13226 <= not w12747 and w13225;
w13227 <= not w12656 and not w13226;
w13228 <= not w13224 and not w13227;
w13229 <= w184 and not w13209;
w13230 <= not w13219 and w13229;
w13231 <= not w13228 and not w13230;
w13232 <= not w13221 and not w13231;
w13233 <= not w115 and not w13232;
w13234 <= not w12661 and w12668;
w13235 <= not w12670 and w13234;
w13236 <= not w12747 and w13235;
w13237 <= not w12661 and not w12670;
w13238 <= not w12747 and w13237;
w13239 <= not w12668 and not w13238;
w13240 <= not w13236 and not w13239;
w13241 <= w115 and not w13221;
w13242 <= not w13231 and w13241;
w13243 <= not w13240 and not w13242;
w13244 <= not w13233 and not w13243;
w13245 <= not w60 and not w13244;
w13246 <= w12680 and not w12682;
w13247 <= not w12673 and w13246;
w13248 <= not w12747 and w13247;
w13249 <= not w12673 and not w12682;
w13250 <= not w12747 and w13249;
w13251 <= not w12680 and not w13250;
w13252 <= not w13248 and not w13251;
w13253 <= w60 and not w13233;
w13254 <= not w13243 and w13253;
w13255 <= not w13252 and not w13254;
w13256 <= not w13245 and not w13255;
w13257 <= not w22 and not w13256;
w13258 <= not w12685 and w12692;
w13259 <= not w12694 and w13258;
w13260 <= not w12747 and w13259;
w13261 <= not w12685 and not w12694;
w13262 <= not w12747 and w13261;
w13263 <= not w12692 and not w13262;
w13264 <= not w13260 and not w13263;
w13265 <= w22 and not w13245;
w13266 <= not w13255 and w13265;
w13267 <= not w13264 and not w13266;
w13268 <= not w13257 and not w13267;
w13269 <= not w5 and not w13268;
w13270 <= w12704 and not w12706;
w13271 <= not w12697 and w13270;
w13272 <= not w12747 and w13271;
w13273 <= not w12697 and not w12706;
w13274 <= not w12747 and w13273;
w13275 <= not w12704 and not w13274;
w13276 <= not w13272 and not w13275;
w13277 <= w5 and not w13257;
w13278 <= not w13267 and w13277;
w13279 <= not w13276 and not w13278;
w13280 <= not w13269 and not w13279;
w13281 <= not w12709 and w12716;
w13282 <= not w12718 and w13281;
w13283 <= not w12747 and w13282;
w13284 <= not w12709 and not w12718;
w13285 <= not w12747 and w13284;
w13286 <= not w12716 and not w13285;
w13287 <= not w13283 and not w13286;
w13288 <= not w12720 and not w12727;
w13289 <= not w12747 and w13288;
w13290 <= not w12735 and not w13289;
w13291 <= not w13287 and w13290;
w13292 <= not w13280 and w13291;
w13293 <= w0 and not w13292;
w13294 <= not w13269 and w13287;
w13295 <= not w13279 and w13294;
w13296 <= not w12727 and not w12747;
w13297 <= w12720 and not w13296;
w13298 <= not w0 and not w13288;
w13299 <= not w13297 and w13298;
w13300 <= not w12723 and not w12744;
w13301 <= not w12726 and w13300;
w13302 <= not w12739 and w13301;
w13303 <= not w12735 and w13302;
w13304 <= not w12733 and w13303;
w13305 <= not w13299 and not w13304;
w13306 <= not w13295 and w13305;
w13307 <= not w13293 and w13306;
w13308 <= a(34) and not w13307;
w13309 <= not a(32) and not a(33);
w13310 <= not a(34) and w13309;
w13311 <= not w13308 and not w13310;
w13312 <= not w12747 and not w13311;
w13313 <= not w12744 and not w13310;
w13314 <= not w12739 and w13313;
w13315 <= not w12735 and w13314;
w13316 <= not w12733 and w13315;
w13317 <= not w13308 and w13316;
w13318 <= not a(34) and not w13307;
w13319 <= a(35) and not w13318;
w13320 <= w12749 and not w13307;
w13321 <= not w13319 and not w13320;
w13322 <= not w13317 and w13321;
w13323 <= not w13312 and not w13322;
w13324 <= not w12199 and not w13323;
w13325 <= w12199 and not w13312;
w13326 <= not w13322 and w13325;
w13327 <= not w12747 and not w13304;
w13328 <= not w13299 and w13327;
w13329 <= not w13295 and w13328;
w13330 <= not w13293 and w13329;
w13331 <= not w13320 and not w13330;
w13332 <= a(36) and not w13331;
w13333 <= not a(36) and not w13330;
w13334 <= not w13320 and w13333;
w13335 <= not w13332 and not w13334;
w13336 <= not w13326 and not w13335;
w13337 <= not w13324 and not w13336;
w13338 <= not w11663 and not w13337;
w13339 <= not w12752 and not w12757;
w13340 <= not w12761 and w13339;
w13341 <= not w13307 and w13340;
w13342 <= not w13307 and w13339;
w13343 <= w12761 and not w13342;
w13344 <= not w13341 and not w13343;
w13345 <= w11663 and not w13324;
w13346 <= not w13336 and w13345;
w13347 <= not w13344 and not w13346;
w13348 <= not w13338 and not w13347;
w13349 <= not w11139 and not w13348;
w13350 <= not w12766 and w12775;
w13351 <= not w12764 and w13350;
w13352 <= not w13307 and w13351;
w13353 <= not w12764 and not w12766;
w13354 <= not w13307 and w13353;
w13355 <= not w12775 and not w13354;
w13356 <= not w13352 and not w13355;
w13357 <= w11139 and not w13338;
w13358 <= not w13347 and w13357;
w13359 <= not w13356 and not w13358;
w13360 <= not w13349 and not w13359;
w13361 <= not w10627 and not w13360;
w13362 <= not w12778 and w12784;
w13363 <= not w12786 and w13362;
w13364 <= not w13307 and w13363;
w13365 <= not w12778 and not w12786;
w13366 <= not w13307 and w13365;
w13367 <= not w12784 and not w13366;
w13368 <= not w13364 and not w13367;
w13369 <= w10627 and not w13349;
w13370 <= not w13359 and w13369;
w13371 <= not w13368 and not w13370;
w13372 <= not w13361 and not w13371;
w13373 <= not w10127 and not w13372;
w13374 <= w12796 and not w12798;
w13375 <= not w12789 and w13374;
w13376 <= not w13307 and w13375;
w13377 <= not w12789 and not w12798;
w13378 <= not w13307 and w13377;
w13379 <= not w12796 and not w13378;
w13380 <= not w13376 and not w13379;
w13381 <= w10127 and not w13361;
w13382 <= not w13371 and w13381;
w13383 <= not w13380 and not w13382;
w13384 <= not w13373 and not w13383;
w13385 <= not w9639 and not w13384;
w13386 <= not w12801 and w12808;
w13387 <= not w12810 and w13386;
w13388 <= not w13307 and w13387;
w13389 <= not w12801 and not w12810;
w13390 <= not w13307 and w13389;
w13391 <= not w12808 and not w13390;
w13392 <= not w13388 and not w13391;
w13393 <= w9639 and not w13373;
w13394 <= not w13383 and w13393;
w13395 <= not w13392 and not w13394;
w13396 <= not w13385 and not w13395;
w13397 <= not w9163 and not w13396;
w13398 <= w12820 and not w12822;
w13399 <= not w12813 and w13398;
w13400 <= not w13307 and w13399;
w13401 <= not w12813 and not w12822;
w13402 <= not w13307 and w13401;
w13403 <= not w12820 and not w13402;
w13404 <= not w13400 and not w13403;
w13405 <= w9163 and not w13385;
w13406 <= not w13395 and w13405;
w13407 <= not w13404 and not w13406;
w13408 <= not w13397 and not w13407;
w13409 <= not w8699 and not w13408;
w13410 <= not w12825 and w12832;
w13411 <= not w12834 and w13410;
w13412 <= not w13307 and w13411;
w13413 <= not w12825 and not w12834;
w13414 <= not w13307 and w13413;
w13415 <= not w12832 and not w13414;
w13416 <= not w13412 and not w13415;
w13417 <= w8699 and not w13397;
w13418 <= not w13407 and w13417;
w13419 <= not w13416 and not w13418;
w13420 <= not w13409 and not w13419;
w13421 <= not w8247 and not w13420;
w13422 <= w12844 and not w12846;
w13423 <= not w12837 and w13422;
w13424 <= not w13307 and w13423;
w13425 <= not w12837 and not w12846;
w13426 <= not w13307 and w13425;
w13427 <= not w12844 and not w13426;
w13428 <= not w13424 and not w13427;
w13429 <= w8247 and not w13409;
w13430 <= not w13419 and w13429;
w13431 <= not w13428 and not w13430;
w13432 <= not w13421 and not w13431;
w13433 <= not w7807 and not w13432;
w13434 <= not w12849 and w12856;
w13435 <= not w12858 and w13434;
w13436 <= not w13307 and w13435;
w13437 <= not w12849 and not w12858;
w13438 <= not w13307 and w13437;
w13439 <= not w12856 and not w13438;
w13440 <= not w13436 and not w13439;
w13441 <= w7807 and not w13421;
w13442 <= not w13431 and w13441;
w13443 <= not w13440 and not w13442;
w13444 <= not w13433 and not w13443;
w13445 <= not w7379 and not w13444;
w13446 <= w12868 and not w12870;
w13447 <= not w12861 and w13446;
w13448 <= not w13307 and w13447;
w13449 <= not w12861 and not w12870;
w13450 <= not w13307 and w13449;
w13451 <= not w12868 and not w13450;
w13452 <= not w13448 and not w13451;
w13453 <= w7379 and not w13433;
w13454 <= not w13443 and w13453;
w13455 <= not w13452 and not w13454;
w13456 <= not w13445 and not w13455;
w13457 <= not w6963 and not w13456;
w13458 <= not w12873 and w12880;
w13459 <= not w12882 and w13458;
w13460 <= not w13307 and w13459;
w13461 <= not w12873 and not w12882;
w13462 <= not w13307 and w13461;
w13463 <= not w12880 and not w13462;
w13464 <= not w13460 and not w13463;
w13465 <= w6963 and not w13445;
w13466 <= not w13455 and w13465;
w13467 <= not w13464 and not w13466;
w13468 <= not w13457 and not w13467;
w13469 <= not w6558 and not w13468;
w13470 <= w12892 and not w12894;
w13471 <= not w12885 and w13470;
w13472 <= not w13307 and w13471;
w13473 <= not w12885 and not w12894;
w13474 <= not w13307 and w13473;
w13475 <= not w12892 and not w13474;
w13476 <= not w13472 and not w13475;
w13477 <= w6558 and not w13457;
w13478 <= not w13467 and w13477;
w13479 <= not w13476 and not w13478;
w13480 <= not w13469 and not w13479;
w13481 <= not w6166 and not w13480;
w13482 <= not w12897 and w12904;
w13483 <= not w12906 and w13482;
w13484 <= not w13307 and w13483;
w13485 <= not w12897 and not w12906;
w13486 <= not w13307 and w13485;
w13487 <= not w12904 and not w13486;
w13488 <= not w13484 and not w13487;
w13489 <= w6166 and not w13469;
w13490 <= not w13479 and w13489;
w13491 <= not w13488 and not w13490;
w13492 <= not w13481 and not w13491;
w13493 <= not w5786 and not w13492;
w13494 <= w12916 and not w12918;
w13495 <= not w12909 and w13494;
w13496 <= not w13307 and w13495;
w13497 <= not w12909 and not w12918;
w13498 <= not w13307 and w13497;
w13499 <= not w12916 and not w13498;
w13500 <= not w13496 and not w13499;
w13501 <= w5786 and not w13481;
w13502 <= not w13491 and w13501;
w13503 <= not w13500 and not w13502;
w13504 <= not w13493 and not w13503;
w13505 <= not w5418 and not w13504;
w13506 <= not w12921 and w12928;
w13507 <= not w12930 and w13506;
w13508 <= not w13307 and w13507;
w13509 <= not w12921 and not w12930;
w13510 <= not w13307 and w13509;
w13511 <= not w12928 and not w13510;
w13512 <= not w13508 and not w13511;
w13513 <= w5418 and not w13493;
w13514 <= not w13503 and w13513;
w13515 <= not w13512 and not w13514;
w13516 <= not w13505 and not w13515;
w13517 <= not w5062 and not w13516;
w13518 <= w12940 and not w12942;
w13519 <= not w12933 and w13518;
w13520 <= not w13307 and w13519;
w13521 <= not w12933 and not w12942;
w13522 <= not w13307 and w13521;
w13523 <= not w12940 and not w13522;
w13524 <= not w13520 and not w13523;
w13525 <= w5062 and not w13505;
w13526 <= not w13515 and w13525;
w13527 <= not w13524 and not w13526;
w13528 <= not w13517 and not w13527;
w13529 <= not w4718 and not w13528;
w13530 <= not w12945 and w12952;
w13531 <= not w12954 and w13530;
w13532 <= not w13307 and w13531;
w13533 <= not w12945 and not w12954;
w13534 <= not w13307 and w13533;
w13535 <= not w12952 and not w13534;
w13536 <= not w13532 and not w13535;
w13537 <= w4718 and not w13517;
w13538 <= not w13527 and w13537;
w13539 <= not w13536 and not w13538;
w13540 <= not w13529 and not w13539;
w13541 <= not w4386 and not w13540;
w13542 <= w12964 and not w12966;
w13543 <= not w12957 and w13542;
w13544 <= not w13307 and w13543;
w13545 <= not w12957 and not w12966;
w13546 <= not w13307 and w13545;
w13547 <= not w12964 and not w13546;
w13548 <= not w13544 and not w13547;
w13549 <= w4386 and not w13529;
w13550 <= not w13539 and w13549;
w13551 <= not w13548 and not w13550;
w13552 <= not w13541 and not w13551;
w13553 <= not w4066 and not w13552;
w13554 <= not w12969 and w12976;
w13555 <= not w12978 and w13554;
w13556 <= not w13307 and w13555;
w13557 <= not w12969 and not w12978;
w13558 <= not w13307 and w13557;
w13559 <= not w12976 and not w13558;
w13560 <= not w13556 and not w13559;
w13561 <= w4066 and not w13541;
w13562 <= not w13551 and w13561;
w13563 <= not w13560 and not w13562;
w13564 <= not w13553 and not w13563;
w13565 <= not w3758 and not w13564;
w13566 <= w12988 and not w12990;
w13567 <= not w12981 and w13566;
w13568 <= not w13307 and w13567;
w13569 <= not w12981 and not w12990;
w13570 <= not w13307 and w13569;
w13571 <= not w12988 and not w13570;
w13572 <= not w13568 and not w13571;
w13573 <= w3758 and not w13553;
w13574 <= not w13563 and w13573;
w13575 <= not w13572 and not w13574;
w13576 <= not w13565 and not w13575;
w13577 <= not w3462 and not w13576;
w13578 <= not w12993 and w13000;
w13579 <= not w13002 and w13578;
w13580 <= not w13307 and w13579;
w13581 <= not w12993 and not w13002;
w13582 <= not w13307 and w13581;
w13583 <= not w13000 and not w13582;
w13584 <= not w13580 and not w13583;
w13585 <= w3462 and not w13565;
w13586 <= not w13575 and w13585;
w13587 <= not w13584 and not w13586;
w13588 <= not w13577 and not w13587;
w13589 <= not w3178 and not w13588;
w13590 <= w13012 and not w13014;
w13591 <= not w13005 and w13590;
w13592 <= not w13307 and w13591;
w13593 <= not w13005 and not w13014;
w13594 <= not w13307 and w13593;
w13595 <= not w13012 and not w13594;
w13596 <= not w13592 and not w13595;
w13597 <= w3178 and not w13577;
w13598 <= not w13587 and w13597;
w13599 <= not w13596 and not w13598;
w13600 <= not w13589 and not w13599;
w13601 <= not w2906 and not w13600;
w13602 <= not w13017 and w13024;
w13603 <= not w13026 and w13602;
w13604 <= not w13307 and w13603;
w13605 <= not w13017 and not w13026;
w13606 <= not w13307 and w13605;
w13607 <= not w13024 and not w13606;
w13608 <= not w13604 and not w13607;
w13609 <= w2906 and not w13589;
w13610 <= not w13599 and w13609;
w13611 <= not w13608 and not w13610;
w13612 <= not w13601 and not w13611;
w13613 <= not w2646 and not w13612;
w13614 <= w13036 and not w13038;
w13615 <= not w13029 and w13614;
w13616 <= not w13307 and w13615;
w13617 <= not w13029 and not w13038;
w13618 <= not w13307 and w13617;
w13619 <= not w13036 and not w13618;
w13620 <= not w13616 and not w13619;
w13621 <= w2646 and not w13601;
w13622 <= not w13611 and w13621;
w13623 <= not w13620 and not w13622;
w13624 <= not w13613 and not w13623;
w13625 <= not w2398 and not w13624;
w13626 <= not w13041 and w13048;
w13627 <= not w13050 and w13626;
w13628 <= not w13307 and w13627;
w13629 <= not w13041 and not w13050;
w13630 <= not w13307 and w13629;
w13631 <= not w13048 and not w13630;
w13632 <= not w13628 and not w13631;
w13633 <= w2398 and not w13613;
w13634 <= not w13623 and w13633;
w13635 <= not w13632 and not w13634;
w13636 <= not w13625 and not w13635;
w13637 <= not w2162 and not w13636;
w13638 <= w13060 and not w13062;
w13639 <= not w13053 and w13638;
w13640 <= not w13307 and w13639;
w13641 <= not w13053 and not w13062;
w13642 <= not w13307 and w13641;
w13643 <= not w13060 and not w13642;
w13644 <= not w13640 and not w13643;
w13645 <= w2162 and not w13625;
w13646 <= not w13635 and w13645;
w13647 <= not w13644 and not w13646;
w13648 <= not w13637 and not w13647;
w13649 <= not w1938 and not w13648;
w13650 <= not w13065 and w13072;
w13651 <= not w13074 and w13650;
w13652 <= not w13307 and w13651;
w13653 <= not w13065 and not w13074;
w13654 <= not w13307 and w13653;
w13655 <= not w13072 and not w13654;
w13656 <= not w13652 and not w13655;
w13657 <= w1938 and not w13637;
w13658 <= not w13647 and w13657;
w13659 <= not w13656 and not w13658;
w13660 <= not w13649 and not w13659;
w13661 <= not w1725 and not w13660;
w13662 <= w13084 and not w13086;
w13663 <= not w13077 and w13662;
w13664 <= not w13307 and w13663;
w13665 <= not w13077 and not w13086;
w13666 <= not w13307 and w13665;
w13667 <= not w13084 and not w13666;
w13668 <= not w13664 and not w13667;
w13669 <= w1725 and not w13649;
w13670 <= not w13659 and w13669;
w13671 <= not w13668 and not w13670;
w13672 <= not w13661 and not w13671;
w13673 <= not w1525 and not w13672;
w13674 <= w1525 and not w13661;
w13675 <= not w13671 and w13674;
w13676 <= not w13089 and w13098;
w13677 <= not w13091 and w13676;
w13678 <= not w13307 and w13677;
w13679 <= not w13089 and not w13091;
w13680 <= not w13307 and w13679;
w13681 <= not w13098 and not w13680;
w13682 <= not w13678 and not w13681;
w13683 <= not w13675 and not w13682;
w13684 <= not w13673 and not w13683;
w13685 <= not w1337 and not w13684;
w13686 <= w13108 and not w13110;
w13687 <= not w13101 and w13686;
w13688 <= not w13307 and w13687;
w13689 <= not w13101 and not w13110;
w13690 <= not w13307 and w13689;
w13691 <= not w13108 and not w13690;
w13692 <= not w13688 and not w13691;
w13693 <= w1337 and not w13673;
w13694 <= not w13683 and w13693;
w13695 <= not w13692 and not w13694;
w13696 <= not w13685 and not w13695;
w13697 <= not w1161 and not w13696;
w13698 <= not w13113 and w13120;
w13699 <= not w13122 and w13698;
w13700 <= not w13307 and w13699;
w13701 <= not w13113 and not w13122;
w13702 <= not w13307 and w13701;
w13703 <= not w13120 and not w13702;
w13704 <= not w13700 and not w13703;
w13705 <= w1161 and not w13685;
w13706 <= not w13695 and w13705;
w13707 <= not w13704 and not w13706;
w13708 <= not w13697 and not w13707;
w13709 <= not w997 and not w13708;
w13710 <= w13132 and not w13134;
w13711 <= not w13125 and w13710;
w13712 <= not w13307 and w13711;
w13713 <= not w13125 and not w13134;
w13714 <= not w13307 and w13713;
w13715 <= not w13132 and not w13714;
w13716 <= not w13712 and not w13715;
w13717 <= w997 and not w13697;
w13718 <= not w13707 and w13717;
w13719 <= not w13716 and not w13718;
w13720 <= not w13709 and not w13719;
w13721 <= not w845 and not w13720;
w13722 <= not w13137 and w13144;
w13723 <= not w13146 and w13722;
w13724 <= not w13307 and w13723;
w13725 <= not w13137 and not w13146;
w13726 <= not w13307 and w13725;
w13727 <= not w13144 and not w13726;
w13728 <= not w13724 and not w13727;
w13729 <= w845 and not w13709;
w13730 <= not w13719 and w13729;
w13731 <= not w13728 and not w13730;
w13732 <= not w13721 and not w13731;
w13733 <= not w705 and not w13732;
w13734 <= w13156 and not w13158;
w13735 <= not w13149 and w13734;
w13736 <= not w13307 and w13735;
w13737 <= not w13149 and not w13158;
w13738 <= not w13307 and w13737;
w13739 <= not w13156 and not w13738;
w13740 <= not w13736 and not w13739;
w13741 <= w705 and not w13721;
w13742 <= not w13731 and w13741;
w13743 <= not w13740 and not w13742;
w13744 <= not w13733 and not w13743;
w13745 <= not w577 and not w13744;
w13746 <= not w13161 and w13168;
w13747 <= not w13170 and w13746;
w13748 <= not w13307 and w13747;
w13749 <= not w13161 and not w13170;
w13750 <= not w13307 and w13749;
w13751 <= not w13168 and not w13750;
w13752 <= not w13748 and not w13751;
w13753 <= w577 and not w13733;
w13754 <= not w13743 and w13753;
w13755 <= not w13752 and not w13754;
w13756 <= not w13745 and not w13755;
w13757 <= not w460 and not w13756;
w13758 <= w13180 and not w13182;
w13759 <= not w13173 and w13758;
w13760 <= not w13307 and w13759;
w13761 <= not w13173 and not w13182;
w13762 <= not w13307 and w13761;
w13763 <= not w13180 and not w13762;
w13764 <= not w13760 and not w13763;
w13765 <= w460 and not w13745;
w13766 <= not w13755 and w13765;
w13767 <= not w13764 and not w13766;
w13768 <= not w13757 and not w13767;
w13769 <= not w356 and not w13768;
w13770 <= not w13185 and w13192;
w13771 <= not w13194 and w13770;
w13772 <= not w13307 and w13771;
w13773 <= not w13185 and not w13194;
w13774 <= not w13307 and w13773;
w13775 <= not w13192 and not w13774;
w13776 <= not w13772 and not w13775;
w13777 <= w356 and not w13757;
w13778 <= not w13767 and w13777;
w13779 <= not w13776 and not w13778;
w13780 <= not w13769 and not w13779;
w13781 <= not w264 and not w13780;
w13782 <= w13204 and not w13206;
w13783 <= not w13197 and w13782;
w13784 <= not w13307 and w13783;
w13785 <= not w13197 and not w13206;
w13786 <= not w13307 and w13785;
w13787 <= not w13204 and not w13786;
w13788 <= not w13784 and not w13787;
w13789 <= w264 and not w13769;
w13790 <= not w13779 and w13789;
w13791 <= not w13788 and not w13790;
w13792 <= not w13781 and not w13791;
w13793 <= not w184 and not w13792;
w13794 <= not w13209 and w13216;
w13795 <= not w13218 and w13794;
w13796 <= not w13307 and w13795;
w13797 <= not w13209 and not w13218;
w13798 <= not w13307 and w13797;
w13799 <= not w13216 and not w13798;
w13800 <= not w13796 and not w13799;
w13801 <= w184 and not w13781;
w13802 <= not w13791 and w13801;
w13803 <= not w13800 and not w13802;
w13804 <= not w13793 and not w13803;
w13805 <= not w115 and not w13804;
w13806 <= w13228 and not w13230;
w13807 <= not w13221 and w13806;
w13808 <= not w13307 and w13807;
w13809 <= not w13221 and not w13230;
w13810 <= not w13307 and w13809;
w13811 <= not w13228 and not w13810;
w13812 <= not w13808 and not w13811;
w13813 <= w115 and not w13793;
w13814 <= not w13803 and w13813;
w13815 <= not w13812 and not w13814;
w13816 <= not w13805 and not w13815;
w13817 <= not w60 and not w13816;
w13818 <= not w13233 and w13240;
w13819 <= not w13242 and w13818;
w13820 <= not w13307 and w13819;
w13821 <= not w13233 and not w13242;
w13822 <= not w13307 and w13821;
w13823 <= not w13240 and not w13822;
w13824 <= not w13820 and not w13823;
w13825 <= w60 and not w13805;
w13826 <= not w13815 and w13825;
w13827 <= not w13824 and not w13826;
w13828 <= not w13817 and not w13827;
w13829 <= not w22 and not w13828;
w13830 <= w13252 and not w13254;
w13831 <= not w13245 and w13830;
w13832 <= not w13307 and w13831;
w13833 <= not w13245 and not w13254;
w13834 <= not w13307 and w13833;
w13835 <= not w13252 and not w13834;
w13836 <= not w13832 and not w13835;
w13837 <= w22 and not w13817;
w13838 <= not w13827 and w13837;
w13839 <= not w13836 and not w13838;
w13840 <= not w13829 and not w13839;
w13841 <= not w5 and not w13840;
w13842 <= not w13257 and w13264;
w13843 <= not w13266 and w13842;
w13844 <= not w13307 and w13843;
w13845 <= not w13257 and not w13266;
w13846 <= not w13307 and w13845;
w13847 <= not w13264 and not w13846;
w13848 <= not w13844 and not w13847;
w13849 <= w5 and not w13829;
w13850 <= not w13839 and w13849;
w13851 <= not w13848 and not w13850;
w13852 <= not w13841 and not w13851;
w13853 <= w13276 and not w13278;
w13854 <= not w13269 and w13853;
w13855 <= not w13307 and w13854;
w13856 <= not w13269 and not w13278;
w13857 <= not w13307 and w13856;
w13858 <= not w13276 and not w13857;
w13859 <= not w13855 and not w13858;
w13860 <= not w13280 and not w13287;
w13861 <= not w13307 and w13860;
w13862 <= not w13295 and not w13861;
w13863 <= not w13859 and w13862;
w13864 <= not w13852 and w13863;
w13865 <= w0 and not w13864;
w13866 <= not w13841 and w13859;
w13867 <= not w13851 and w13866;
w13868 <= not w13287 and not w13307;
w13869 <= w13280 and not w13868;
w13870 <= not w0 and not w13860;
w13871 <= not w13869 and w13870;
w13872 <= not w13283 and not w13304;
w13873 <= not w13286 and w13872;
w13874 <= not w13299 and w13873;
w13875 <= not w13295 and w13874;
w13876 <= not w13293 and w13875;
w13877 <= not w13871 and not w13876;
w13878 <= not w13867 and w13877;
w13879 <= not w13865 and w13878;
w13880 <= a(32) and not w13879;
w13881 <= not a(30) and not a(31);
w13882 <= not a(32) and w13881;
w13883 <= not w13880 and not w13882;
w13884 <= not w13307 and not w13883;
w13885 <= not w13304 and not w13882;
w13886 <= not w13299 and w13885;
w13887 <= not w13295 and w13886;
w13888 <= not w13293 and w13887;
w13889 <= not w13880 and w13888;
w13890 <= not a(32) and not w13879;
w13891 <= a(33) and not w13890;
w13892 <= w13309 and not w13879;
w13893 <= not w13891 and not w13892;
w13894 <= not w13889 and w13893;
w13895 <= not w13884 and not w13894;
w13896 <= not w12747 and not w13895;
w13897 <= w12747 and not w13884;
w13898 <= not w13894 and w13897;
w13899 <= not w13307 and not w13876;
w13900 <= not w13871 and w13899;
w13901 <= not w13867 and w13900;
w13902 <= not w13865 and w13901;
w13903 <= not w13892 and not w13902;
w13904 <= a(34) and not w13903;
w13905 <= not a(34) and not w13902;
w13906 <= not w13892 and w13905;
w13907 <= not w13904 and not w13906;
w13908 <= not w13898 and not w13907;
w13909 <= not w13896 and not w13908;
w13910 <= not w12199 and not w13909;
w13911 <= not w13312 and not w13317;
w13912 <= not w13321 and w13911;
w13913 <= not w13879 and w13912;
w13914 <= not w13879 and w13911;
w13915 <= w13321 and not w13914;
w13916 <= not w13913 and not w13915;
w13917 <= w12199 and not w13896;
w13918 <= not w13908 and w13917;
w13919 <= not w13916 and not w13918;
w13920 <= not w13910 and not w13919;
w13921 <= not w11663 and not w13920;
w13922 <= not w13326 and w13335;
w13923 <= not w13324 and w13922;
w13924 <= not w13879 and w13923;
w13925 <= not w13324 and not w13326;
w13926 <= not w13879 and w13925;
w13927 <= not w13335 and not w13926;
w13928 <= not w13924 and not w13927;
w13929 <= w11663 and not w13910;
w13930 <= not w13919 and w13929;
w13931 <= not w13928 and not w13930;
w13932 <= not w13921 and not w13931;
w13933 <= not w11139 and not w13932;
w13934 <= not w13338 and w13344;
w13935 <= not w13346 and w13934;
w13936 <= not w13879 and w13935;
w13937 <= not w13338 and not w13346;
w13938 <= not w13879 and w13937;
w13939 <= not w13344 and not w13938;
w13940 <= not w13936 and not w13939;
w13941 <= w11139 and not w13921;
w13942 <= not w13931 and w13941;
w13943 <= not w13940 and not w13942;
w13944 <= not w13933 and not w13943;
w13945 <= not w10627 and not w13944;
w13946 <= w13356 and not w13358;
w13947 <= not w13349 and w13946;
w13948 <= not w13879 and w13947;
w13949 <= not w13349 and not w13358;
w13950 <= not w13879 and w13949;
w13951 <= not w13356 and not w13950;
w13952 <= not w13948 and not w13951;
w13953 <= w10627 and not w13933;
w13954 <= not w13943 and w13953;
w13955 <= not w13952 and not w13954;
w13956 <= not w13945 and not w13955;
w13957 <= not w10127 and not w13956;
w13958 <= not w13361 and w13368;
w13959 <= not w13370 and w13958;
w13960 <= not w13879 and w13959;
w13961 <= not w13361 and not w13370;
w13962 <= not w13879 and w13961;
w13963 <= not w13368 and not w13962;
w13964 <= not w13960 and not w13963;
w13965 <= w10127 and not w13945;
w13966 <= not w13955 and w13965;
w13967 <= not w13964 and not w13966;
w13968 <= not w13957 and not w13967;
w13969 <= not w9639 and not w13968;
w13970 <= w13380 and not w13382;
w13971 <= not w13373 and w13970;
w13972 <= not w13879 and w13971;
w13973 <= not w13373 and not w13382;
w13974 <= not w13879 and w13973;
w13975 <= not w13380 and not w13974;
w13976 <= not w13972 and not w13975;
w13977 <= w9639 and not w13957;
w13978 <= not w13967 and w13977;
w13979 <= not w13976 and not w13978;
w13980 <= not w13969 and not w13979;
w13981 <= not w9163 and not w13980;
w13982 <= not w13385 and w13392;
w13983 <= not w13394 and w13982;
w13984 <= not w13879 and w13983;
w13985 <= not w13385 and not w13394;
w13986 <= not w13879 and w13985;
w13987 <= not w13392 and not w13986;
w13988 <= not w13984 and not w13987;
w13989 <= w9163 and not w13969;
w13990 <= not w13979 and w13989;
w13991 <= not w13988 and not w13990;
w13992 <= not w13981 and not w13991;
w13993 <= not w8699 and not w13992;
w13994 <= w13404 and not w13406;
w13995 <= not w13397 and w13994;
w13996 <= not w13879 and w13995;
w13997 <= not w13397 and not w13406;
w13998 <= not w13879 and w13997;
w13999 <= not w13404 and not w13998;
w14000 <= not w13996 and not w13999;
w14001 <= w8699 and not w13981;
w14002 <= not w13991 and w14001;
w14003 <= not w14000 and not w14002;
w14004 <= not w13993 and not w14003;
w14005 <= not w8247 and not w14004;
w14006 <= not w13409 and w13416;
w14007 <= not w13418 and w14006;
w14008 <= not w13879 and w14007;
w14009 <= not w13409 and not w13418;
w14010 <= not w13879 and w14009;
w14011 <= not w13416 and not w14010;
w14012 <= not w14008 and not w14011;
w14013 <= w8247 and not w13993;
w14014 <= not w14003 and w14013;
w14015 <= not w14012 and not w14014;
w14016 <= not w14005 and not w14015;
w14017 <= not w7807 and not w14016;
w14018 <= w13428 and not w13430;
w14019 <= not w13421 and w14018;
w14020 <= not w13879 and w14019;
w14021 <= not w13421 and not w13430;
w14022 <= not w13879 and w14021;
w14023 <= not w13428 and not w14022;
w14024 <= not w14020 and not w14023;
w14025 <= w7807 and not w14005;
w14026 <= not w14015 and w14025;
w14027 <= not w14024 and not w14026;
w14028 <= not w14017 and not w14027;
w14029 <= not w7379 and not w14028;
w14030 <= not w13433 and w13440;
w14031 <= not w13442 and w14030;
w14032 <= not w13879 and w14031;
w14033 <= not w13433 and not w13442;
w14034 <= not w13879 and w14033;
w14035 <= not w13440 and not w14034;
w14036 <= not w14032 and not w14035;
w14037 <= w7379 and not w14017;
w14038 <= not w14027 and w14037;
w14039 <= not w14036 and not w14038;
w14040 <= not w14029 and not w14039;
w14041 <= not w6963 and not w14040;
w14042 <= w13452 and not w13454;
w14043 <= not w13445 and w14042;
w14044 <= not w13879 and w14043;
w14045 <= not w13445 and not w13454;
w14046 <= not w13879 and w14045;
w14047 <= not w13452 and not w14046;
w14048 <= not w14044 and not w14047;
w14049 <= w6963 and not w14029;
w14050 <= not w14039 and w14049;
w14051 <= not w14048 and not w14050;
w14052 <= not w14041 and not w14051;
w14053 <= not w6558 and not w14052;
w14054 <= not w13457 and w13464;
w14055 <= not w13466 and w14054;
w14056 <= not w13879 and w14055;
w14057 <= not w13457 and not w13466;
w14058 <= not w13879 and w14057;
w14059 <= not w13464 and not w14058;
w14060 <= not w14056 and not w14059;
w14061 <= w6558 and not w14041;
w14062 <= not w14051 and w14061;
w14063 <= not w14060 and not w14062;
w14064 <= not w14053 and not w14063;
w14065 <= not w6166 and not w14064;
w14066 <= w13476 and not w13478;
w14067 <= not w13469 and w14066;
w14068 <= not w13879 and w14067;
w14069 <= not w13469 and not w13478;
w14070 <= not w13879 and w14069;
w14071 <= not w13476 and not w14070;
w14072 <= not w14068 and not w14071;
w14073 <= w6166 and not w14053;
w14074 <= not w14063 and w14073;
w14075 <= not w14072 and not w14074;
w14076 <= not w14065 and not w14075;
w14077 <= not w5786 and not w14076;
w14078 <= not w13481 and w13488;
w14079 <= not w13490 and w14078;
w14080 <= not w13879 and w14079;
w14081 <= not w13481 and not w13490;
w14082 <= not w13879 and w14081;
w14083 <= not w13488 and not w14082;
w14084 <= not w14080 and not w14083;
w14085 <= w5786 and not w14065;
w14086 <= not w14075 and w14085;
w14087 <= not w14084 and not w14086;
w14088 <= not w14077 and not w14087;
w14089 <= not w5418 and not w14088;
w14090 <= w13500 and not w13502;
w14091 <= not w13493 and w14090;
w14092 <= not w13879 and w14091;
w14093 <= not w13493 and not w13502;
w14094 <= not w13879 and w14093;
w14095 <= not w13500 and not w14094;
w14096 <= not w14092 and not w14095;
w14097 <= w5418 and not w14077;
w14098 <= not w14087 and w14097;
w14099 <= not w14096 and not w14098;
w14100 <= not w14089 and not w14099;
w14101 <= not w5062 and not w14100;
w14102 <= not w13505 and w13512;
w14103 <= not w13514 and w14102;
w14104 <= not w13879 and w14103;
w14105 <= not w13505 and not w13514;
w14106 <= not w13879 and w14105;
w14107 <= not w13512 and not w14106;
w14108 <= not w14104 and not w14107;
w14109 <= w5062 and not w14089;
w14110 <= not w14099 and w14109;
w14111 <= not w14108 and not w14110;
w14112 <= not w14101 and not w14111;
w14113 <= not w4718 and not w14112;
w14114 <= w13524 and not w13526;
w14115 <= not w13517 and w14114;
w14116 <= not w13879 and w14115;
w14117 <= not w13517 and not w13526;
w14118 <= not w13879 and w14117;
w14119 <= not w13524 and not w14118;
w14120 <= not w14116 and not w14119;
w14121 <= w4718 and not w14101;
w14122 <= not w14111 and w14121;
w14123 <= not w14120 and not w14122;
w14124 <= not w14113 and not w14123;
w14125 <= not w4386 and not w14124;
w14126 <= not w13529 and w13536;
w14127 <= not w13538 and w14126;
w14128 <= not w13879 and w14127;
w14129 <= not w13529 and not w13538;
w14130 <= not w13879 and w14129;
w14131 <= not w13536 and not w14130;
w14132 <= not w14128 and not w14131;
w14133 <= w4386 and not w14113;
w14134 <= not w14123 and w14133;
w14135 <= not w14132 and not w14134;
w14136 <= not w14125 and not w14135;
w14137 <= not w4066 and not w14136;
w14138 <= w13548 and not w13550;
w14139 <= not w13541 and w14138;
w14140 <= not w13879 and w14139;
w14141 <= not w13541 and not w13550;
w14142 <= not w13879 and w14141;
w14143 <= not w13548 and not w14142;
w14144 <= not w14140 and not w14143;
w14145 <= w4066 and not w14125;
w14146 <= not w14135 and w14145;
w14147 <= not w14144 and not w14146;
w14148 <= not w14137 and not w14147;
w14149 <= not w3758 and not w14148;
w14150 <= not w13553 and w13560;
w14151 <= not w13562 and w14150;
w14152 <= not w13879 and w14151;
w14153 <= not w13553 and not w13562;
w14154 <= not w13879 and w14153;
w14155 <= not w13560 and not w14154;
w14156 <= not w14152 and not w14155;
w14157 <= w3758 and not w14137;
w14158 <= not w14147 and w14157;
w14159 <= not w14156 and not w14158;
w14160 <= not w14149 and not w14159;
w14161 <= not w3462 and not w14160;
w14162 <= w13572 and not w13574;
w14163 <= not w13565 and w14162;
w14164 <= not w13879 and w14163;
w14165 <= not w13565 and not w13574;
w14166 <= not w13879 and w14165;
w14167 <= not w13572 and not w14166;
w14168 <= not w14164 and not w14167;
w14169 <= w3462 and not w14149;
w14170 <= not w14159 and w14169;
w14171 <= not w14168 and not w14170;
w14172 <= not w14161 and not w14171;
w14173 <= not w3178 and not w14172;
w14174 <= not w13577 and w13584;
w14175 <= not w13586 and w14174;
w14176 <= not w13879 and w14175;
w14177 <= not w13577 and not w13586;
w14178 <= not w13879 and w14177;
w14179 <= not w13584 and not w14178;
w14180 <= not w14176 and not w14179;
w14181 <= w3178 and not w14161;
w14182 <= not w14171 and w14181;
w14183 <= not w14180 and not w14182;
w14184 <= not w14173 and not w14183;
w14185 <= not w2906 and not w14184;
w14186 <= w13596 and not w13598;
w14187 <= not w13589 and w14186;
w14188 <= not w13879 and w14187;
w14189 <= not w13589 and not w13598;
w14190 <= not w13879 and w14189;
w14191 <= not w13596 and not w14190;
w14192 <= not w14188 and not w14191;
w14193 <= w2906 and not w14173;
w14194 <= not w14183 and w14193;
w14195 <= not w14192 and not w14194;
w14196 <= not w14185 and not w14195;
w14197 <= not w2646 and not w14196;
w14198 <= not w13601 and w13608;
w14199 <= not w13610 and w14198;
w14200 <= not w13879 and w14199;
w14201 <= not w13601 and not w13610;
w14202 <= not w13879 and w14201;
w14203 <= not w13608 and not w14202;
w14204 <= not w14200 and not w14203;
w14205 <= w2646 and not w14185;
w14206 <= not w14195 and w14205;
w14207 <= not w14204 and not w14206;
w14208 <= not w14197 and not w14207;
w14209 <= not w2398 and not w14208;
w14210 <= w13620 and not w13622;
w14211 <= not w13613 and w14210;
w14212 <= not w13879 and w14211;
w14213 <= not w13613 and not w13622;
w14214 <= not w13879 and w14213;
w14215 <= not w13620 and not w14214;
w14216 <= not w14212 and not w14215;
w14217 <= w2398 and not w14197;
w14218 <= not w14207 and w14217;
w14219 <= not w14216 and not w14218;
w14220 <= not w14209 and not w14219;
w14221 <= not w2162 and not w14220;
w14222 <= not w13625 and w13632;
w14223 <= not w13634 and w14222;
w14224 <= not w13879 and w14223;
w14225 <= not w13625 and not w13634;
w14226 <= not w13879 and w14225;
w14227 <= not w13632 and not w14226;
w14228 <= not w14224 and not w14227;
w14229 <= w2162 and not w14209;
w14230 <= not w14219 and w14229;
w14231 <= not w14228 and not w14230;
w14232 <= not w14221 and not w14231;
w14233 <= not w1938 and not w14232;
w14234 <= w13644 and not w13646;
w14235 <= not w13637 and w14234;
w14236 <= not w13879 and w14235;
w14237 <= not w13637 and not w13646;
w14238 <= not w13879 and w14237;
w14239 <= not w13644 and not w14238;
w14240 <= not w14236 and not w14239;
w14241 <= w1938 and not w14221;
w14242 <= not w14231 and w14241;
w14243 <= not w14240 and not w14242;
w14244 <= not w14233 and not w14243;
w14245 <= not w1725 and not w14244;
w14246 <= not w13649 and w13656;
w14247 <= not w13658 and w14246;
w14248 <= not w13879 and w14247;
w14249 <= not w13649 and not w13658;
w14250 <= not w13879 and w14249;
w14251 <= not w13656 and not w14250;
w14252 <= not w14248 and not w14251;
w14253 <= w1725 and not w14233;
w14254 <= not w14243 and w14253;
w14255 <= not w14252 and not w14254;
w14256 <= not w14245 and not w14255;
w14257 <= not w1525 and not w14256;
w14258 <= w13668 and not w13670;
w14259 <= not w13661 and w14258;
w14260 <= not w13879 and w14259;
w14261 <= not w13661 and not w13670;
w14262 <= not w13879 and w14261;
w14263 <= not w13668 and not w14262;
w14264 <= not w14260 and not w14263;
w14265 <= w1525 and not w14245;
w14266 <= not w14255 and w14265;
w14267 <= not w14264 and not w14266;
w14268 <= not w14257 and not w14267;
w14269 <= not w1337 and not w14268;
w14270 <= w1337 and not w14257;
w14271 <= not w14267 and w14270;
w14272 <= not w13673 and w13682;
w14273 <= not w13675 and w14272;
w14274 <= not w13879 and w14273;
w14275 <= not w13673 and not w13675;
w14276 <= not w13879 and w14275;
w14277 <= not w13682 and not w14276;
w14278 <= not w14274 and not w14277;
w14279 <= not w14271 and not w14278;
w14280 <= not w14269 and not w14279;
w14281 <= not w1161 and not w14280;
w14282 <= w13692 and not w13694;
w14283 <= not w13685 and w14282;
w14284 <= not w13879 and w14283;
w14285 <= not w13685 and not w13694;
w14286 <= not w13879 and w14285;
w14287 <= not w13692 and not w14286;
w14288 <= not w14284 and not w14287;
w14289 <= w1161 and not w14269;
w14290 <= not w14279 and w14289;
w14291 <= not w14288 and not w14290;
w14292 <= not w14281 and not w14291;
w14293 <= not w997 and not w14292;
w14294 <= not w13697 and w13704;
w14295 <= not w13706 and w14294;
w14296 <= not w13879 and w14295;
w14297 <= not w13697 and not w13706;
w14298 <= not w13879 and w14297;
w14299 <= not w13704 and not w14298;
w14300 <= not w14296 and not w14299;
w14301 <= w997 and not w14281;
w14302 <= not w14291 and w14301;
w14303 <= not w14300 and not w14302;
w14304 <= not w14293 and not w14303;
w14305 <= not w845 and not w14304;
w14306 <= w13716 and not w13718;
w14307 <= not w13709 and w14306;
w14308 <= not w13879 and w14307;
w14309 <= not w13709 and not w13718;
w14310 <= not w13879 and w14309;
w14311 <= not w13716 and not w14310;
w14312 <= not w14308 and not w14311;
w14313 <= w845 and not w14293;
w14314 <= not w14303 and w14313;
w14315 <= not w14312 and not w14314;
w14316 <= not w14305 and not w14315;
w14317 <= not w705 and not w14316;
w14318 <= not w13721 and w13728;
w14319 <= not w13730 and w14318;
w14320 <= not w13879 and w14319;
w14321 <= not w13721 and not w13730;
w14322 <= not w13879 and w14321;
w14323 <= not w13728 and not w14322;
w14324 <= not w14320 and not w14323;
w14325 <= w705 and not w14305;
w14326 <= not w14315 and w14325;
w14327 <= not w14324 and not w14326;
w14328 <= not w14317 and not w14327;
w14329 <= not w577 and not w14328;
w14330 <= w13740 and not w13742;
w14331 <= not w13733 and w14330;
w14332 <= not w13879 and w14331;
w14333 <= not w13733 and not w13742;
w14334 <= not w13879 and w14333;
w14335 <= not w13740 and not w14334;
w14336 <= not w14332 and not w14335;
w14337 <= w577 and not w14317;
w14338 <= not w14327 and w14337;
w14339 <= not w14336 and not w14338;
w14340 <= not w14329 and not w14339;
w14341 <= not w460 and not w14340;
w14342 <= not w13745 and w13752;
w14343 <= not w13754 and w14342;
w14344 <= not w13879 and w14343;
w14345 <= not w13745 and not w13754;
w14346 <= not w13879 and w14345;
w14347 <= not w13752 and not w14346;
w14348 <= not w14344 and not w14347;
w14349 <= w460 and not w14329;
w14350 <= not w14339 and w14349;
w14351 <= not w14348 and not w14350;
w14352 <= not w14341 and not w14351;
w14353 <= not w356 and not w14352;
w14354 <= w13764 and not w13766;
w14355 <= not w13757 and w14354;
w14356 <= not w13879 and w14355;
w14357 <= not w13757 and not w13766;
w14358 <= not w13879 and w14357;
w14359 <= not w13764 and not w14358;
w14360 <= not w14356 and not w14359;
w14361 <= w356 and not w14341;
w14362 <= not w14351 and w14361;
w14363 <= not w14360 and not w14362;
w14364 <= not w14353 and not w14363;
w14365 <= not w264 and not w14364;
w14366 <= not w13769 and w13776;
w14367 <= not w13778 and w14366;
w14368 <= not w13879 and w14367;
w14369 <= not w13769 and not w13778;
w14370 <= not w13879 and w14369;
w14371 <= not w13776 and not w14370;
w14372 <= not w14368 and not w14371;
w14373 <= w264 and not w14353;
w14374 <= not w14363 and w14373;
w14375 <= not w14372 and not w14374;
w14376 <= not w14365 and not w14375;
w14377 <= not w184 and not w14376;
w14378 <= w13788 and not w13790;
w14379 <= not w13781 and w14378;
w14380 <= not w13879 and w14379;
w14381 <= not w13781 and not w13790;
w14382 <= not w13879 and w14381;
w14383 <= not w13788 and not w14382;
w14384 <= not w14380 and not w14383;
w14385 <= w184 and not w14365;
w14386 <= not w14375 and w14385;
w14387 <= not w14384 and not w14386;
w14388 <= not w14377 and not w14387;
w14389 <= not w115 and not w14388;
w14390 <= not w13793 and w13800;
w14391 <= not w13802 and w14390;
w14392 <= not w13879 and w14391;
w14393 <= not w13793 and not w13802;
w14394 <= not w13879 and w14393;
w14395 <= not w13800 and not w14394;
w14396 <= not w14392 and not w14395;
w14397 <= w115 and not w14377;
w14398 <= not w14387 and w14397;
w14399 <= not w14396 and not w14398;
w14400 <= not w14389 and not w14399;
w14401 <= not w60 and not w14400;
w14402 <= w13812 and not w13814;
w14403 <= not w13805 and w14402;
w14404 <= not w13879 and w14403;
w14405 <= not w13805 and not w13814;
w14406 <= not w13879 and w14405;
w14407 <= not w13812 and not w14406;
w14408 <= not w14404 and not w14407;
w14409 <= w60 and not w14389;
w14410 <= not w14399 and w14409;
w14411 <= not w14408 and not w14410;
w14412 <= not w14401 and not w14411;
w14413 <= not w22 and not w14412;
w14414 <= not w13817 and w13824;
w14415 <= not w13826 and w14414;
w14416 <= not w13879 and w14415;
w14417 <= not w13817 and not w13826;
w14418 <= not w13879 and w14417;
w14419 <= not w13824 and not w14418;
w14420 <= not w14416 and not w14419;
w14421 <= w22 and not w14401;
w14422 <= not w14411 and w14421;
w14423 <= not w14420 and not w14422;
w14424 <= not w14413 and not w14423;
w14425 <= not w5 and not w14424;
w14426 <= w13836 and not w13838;
w14427 <= not w13829 and w14426;
w14428 <= not w13879 and w14427;
w14429 <= not w13829 and not w13838;
w14430 <= not w13879 and w14429;
w14431 <= not w13836 and not w14430;
w14432 <= not w14428 and not w14431;
w14433 <= w5 and not w14413;
w14434 <= not w14423 and w14433;
w14435 <= not w14432 and not w14434;
w14436 <= not w14425 and not w14435;
w14437 <= not w13841 and w13848;
w14438 <= not w13850 and w14437;
w14439 <= not w13879 and w14438;
w14440 <= not w13841 and not w13850;
w14441 <= not w13879 and w14440;
w14442 <= not w13848 and not w14441;
w14443 <= not w14439 and not w14442;
w14444 <= not w13852 and not w13859;
w14445 <= not w13879 and w14444;
w14446 <= not w13867 and not w14445;
w14447 <= not w14443 and w14446;
w14448 <= not w14436 and w14447;
w14449 <= w0 and not w14448;
w14450 <= not w14425 and w14443;
w14451 <= not w14435 and w14450;
w14452 <= not w13859 and not w13879;
w14453 <= w13852 and not w14452;
w14454 <= not w0 and not w14444;
w14455 <= not w14453 and w14454;
w14456 <= not w13855 and not w13876;
w14457 <= not w13858 and w14456;
w14458 <= not w13871 and w14457;
w14459 <= not w13867 and w14458;
w14460 <= not w13865 and w14459;
w14461 <= not w14455 and not w14460;
w14462 <= not w14451 and w14461;
w14463 <= not w14449 and w14462;
w14464 <= a(30) and not w14463;
w14465 <= not a(28) and not a(29);
w14466 <= not a(30) and w14465;
w14467 <= not w14464 and not w14466;
w14468 <= not w13879 and not w14467;
w14469 <= not w13876 and not w14466;
w14470 <= not w13871 and w14469;
w14471 <= not w13867 and w14470;
w14472 <= not w13865 and w14471;
w14473 <= not w14464 and w14472;
w14474 <= not a(30) and not w14463;
w14475 <= a(31) and not w14474;
w14476 <= w13881 and not w14463;
w14477 <= not w14475 and not w14476;
w14478 <= not w14473 and w14477;
w14479 <= not w14468 and not w14478;
w14480 <= not w13307 and not w14479;
w14481 <= w13307 and not w14468;
w14482 <= not w14478 and w14481;
w14483 <= not w13879 and not w14460;
w14484 <= not w14455 and w14483;
w14485 <= not w14451 and w14484;
w14486 <= not w14449 and w14485;
w14487 <= not w14476 and not w14486;
w14488 <= a(32) and not w14487;
w14489 <= not a(32) and not w14486;
w14490 <= not w14476 and w14489;
w14491 <= not w14488 and not w14490;
w14492 <= not w14482 and not w14491;
w14493 <= not w14480 and not w14492;
w14494 <= not w12747 and not w14493;
w14495 <= not w13884 and not w13889;
w14496 <= not w13893 and w14495;
w14497 <= not w14463 and w14496;
w14498 <= not w14463 and w14495;
w14499 <= w13893 and not w14498;
w14500 <= not w14497 and not w14499;
w14501 <= w12747 and not w14480;
w14502 <= not w14492 and w14501;
w14503 <= not w14500 and not w14502;
w14504 <= not w14494 and not w14503;
w14505 <= not w12199 and not w14504;
w14506 <= not w13898 and w13907;
w14507 <= not w13896 and w14506;
w14508 <= not w14463 and w14507;
w14509 <= not w13896 and not w13898;
w14510 <= not w14463 and w14509;
w14511 <= not w13907 and not w14510;
w14512 <= not w14508 and not w14511;
w14513 <= w12199 and not w14494;
w14514 <= not w14503 and w14513;
w14515 <= not w14512 and not w14514;
w14516 <= not w14505 and not w14515;
w14517 <= not w11663 and not w14516;
w14518 <= not w13910 and w13916;
w14519 <= not w13918 and w14518;
w14520 <= not w14463 and w14519;
w14521 <= not w13910 and not w13918;
w14522 <= not w14463 and w14521;
w14523 <= not w13916 and not w14522;
w14524 <= not w14520 and not w14523;
w14525 <= w11663 and not w14505;
w14526 <= not w14515 and w14525;
w14527 <= not w14524 and not w14526;
w14528 <= not w14517 and not w14527;
w14529 <= not w11139 and not w14528;
w14530 <= w13928 and not w13930;
w14531 <= not w13921 and w14530;
w14532 <= not w14463 and w14531;
w14533 <= not w13921 and not w13930;
w14534 <= not w14463 and w14533;
w14535 <= not w13928 and not w14534;
w14536 <= not w14532 and not w14535;
w14537 <= w11139 and not w14517;
w14538 <= not w14527 and w14537;
w14539 <= not w14536 and not w14538;
w14540 <= not w14529 and not w14539;
w14541 <= not w10627 and not w14540;
w14542 <= not w13933 and w13940;
w14543 <= not w13942 and w14542;
w14544 <= not w14463 and w14543;
w14545 <= not w13933 and not w13942;
w14546 <= not w14463 and w14545;
w14547 <= not w13940 and not w14546;
w14548 <= not w14544 and not w14547;
w14549 <= w10627 and not w14529;
w14550 <= not w14539 and w14549;
w14551 <= not w14548 and not w14550;
w14552 <= not w14541 and not w14551;
w14553 <= not w10127 and not w14552;
w14554 <= w13952 and not w13954;
w14555 <= not w13945 and w14554;
w14556 <= not w14463 and w14555;
w14557 <= not w13945 and not w13954;
w14558 <= not w14463 and w14557;
w14559 <= not w13952 and not w14558;
w14560 <= not w14556 and not w14559;
w14561 <= w10127 and not w14541;
w14562 <= not w14551 and w14561;
w14563 <= not w14560 and not w14562;
w14564 <= not w14553 and not w14563;
w14565 <= not w9639 and not w14564;
w14566 <= not w13957 and w13964;
w14567 <= not w13966 and w14566;
w14568 <= not w14463 and w14567;
w14569 <= not w13957 and not w13966;
w14570 <= not w14463 and w14569;
w14571 <= not w13964 and not w14570;
w14572 <= not w14568 and not w14571;
w14573 <= w9639 and not w14553;
w14574 <= not w14563 and w14573;
w14575 <= not w14572 and not w14574;
w14576 <= not w14565 and not w14575;
w14577 <= not w9163 and not w14576;
w14578 <= w13976 and not w13978;
w14579 <= not w13969 and w14578;
w14580 <= not w14463 and w14579;
w14581 <= not w13969 and not w13978;
w14582 <= not w14463 and w14581;
w14583 <= not w13976 and not w14582;
w14584 <= not w14580 and not w14583;
w14585 <= w9163 and not w14565;
w14586 <= not w14575 and w14585;
w14587 <= not w14584 and not w14586;
w14588 <= not w14577 and not w14587;
w14589 <= not w8699 and not w14588;
w14590 <= not w13981 and w13988;
w14591 <= not w13990 and w14590;
w14592 <= not w14463 and w14591;
w14593 <= not w13981 and not w13990;
w14594 <= not w14463 and w14593;
w14595 <= not w13988 and not w14594;
w14596 <= not w14592 and not w14595;
w14597 <= w8699 and not w14577;
w14598 <= not w14587 and w14597;
w14599 <= not w14596 and not w14598;
w14600 <= not w14589 and not w14599;
w14601 <= not w8247 and not w14600;
w14602 <= w14000 and not w14002;
w14603 <= not w13993 and w14602;
w14604 <= not w14463 and w14603;
w14605 <= not w13993 and not w14002;
w14606 <= not w14463 and w14605;
w14607 <= not w14000 and not w14606;
w14608 <= not w14604 and not w14607;
w14609 <= w8247 and not w14589;
w14610 <= not w14599 and w14609;
w14611 <= not w14608 and not w14610;
w14612 <= not w14601 and not w14611;
w14613 <= not w7807 and not w14612;
w14614 <= not w14005 and w14012;
w14615 <= not w14014 and w14614;
w14616 <= not w14463 and w14615;
w14617 <= not w14005 and not w14014;
w14618 <= not w14463 and w14617;
w14619 <= not w14012 and not w14618;
w14620 <= not w14616 and not w14619;
w14621 <= w7807 and not w14601;
w14622 <= not w14611 and w14621;
w14623 <= not w14620 and not w14622;
w14624 <= not w14613 and not w14623;
w14625 <= not w7379 and not w14624;
w14626 <= w14024 and not w14026;
w14627 <= not w14017 and w14626;
w14628 <= not w14463 and w14627;
w14629 <= not w14017 and not w14026;
w14630 <= not w14463 and w14629;
w14631 <= not w14024 and not w14630;
w14632 <= not w14628 and not w14631;
w14633 <= w7379 and not w14613;
w14634 <= not w14623 and w14633;
w14635 <= not w14632 and not w14634;
w14636 <= not w14625 and not w14635;
w14637 <= not w6963 and not w14636;
w14638 <= not w14029 and w14036;
w14639 <= not w14038 and w14638;
w14640 <= not w14463 and w14639;
w14641 <= not w14029 and not w14038;
w14642 <= not w14463 and w14641;
w14643 <= not w14036 and not w14642;
w14644 <= not w14640 and not w14643;
w14645 <= w6963 and not w14625;
w14646 <= not w14635 and w14645;
w14647 <= not w14644 and not w14646;
w14648 <= not w14637 and not w14647;
w14649 <= not w6558 and not w14648;
w14650 <= w14048 and not w14050;
w14651 <= not w14041 and w14650;
w14652 <= not w14463 and w14651;
w14653 <= not w14041 and not w14050;
w14654 <= not w14463 and w14653;
w14655 <= not w14048 and not w14654;
w14656 <= not w14652 and not w14655;
w14657 <= w6558 and not w14637;
w14658 <= not w14647 and w14657;
w14659 <= not w14656 and not w14658;
w14660 <= not w14649 and not w14659;
w14661 <= not w6166 and not w14660;
w14662 <= not w14053 and w14060;
w14663 <= not w14062 and w14662;
w14664 <= not w14463 and w14663;
w14665 <= not w14053 and not w14062;
w14666 <= not w14463 and w14665;
w14667 <= not w14060 and not w14666;
w14668 <= not w14664 and not w14667;
w14669 <= w6166 and not w14649;
w14670 <= not w14659 and w14669;
w14671 <= not w14668 and not w14670;
w14672 <= not w14661 and not w14671;
w14673 <= not w5786 and not w14672;
w14674 <= w14072 and not w14074;
w14675 <= not w14065 and w14674;
w14676 <= not w14463 and w14675;
w14677 <= not w14065 and not w14074;
w14678 <= not w14463 and w14677;
w14679 <= not w14072 and not w14678;
w14680 <= not w14676 and not w14679;
w14681 <= w5786 and not w14661;
w14682 <= not w14671 and w14681;
w14683 <= not w14680 and not w14682;
w14684 <= not w14673 and not w14683;
w14685 <= not w5418 and not w14684;
w14686 <= not w14077 and w14084;
w14687 <= not w14086 and w14686;
w14688 <= not w14463 and w14687;
w14689 <= not w14077 and not w14086;
w14690 <= not w14463 and w14689;
w14691 <= not w14084 and not w14690;
w14692 <= not w14688 and not w14691;
w14693 <= w5418 and not w14673;
w14694 <= not w14683 and w14693;
w14695 <= not w14692 and not w14694;
w14696 <= not w14685 and not w14695;
w14697 <= not w5062 and not w14696;
w14698 <= w14096 and not w14098;
w14699 <= not w14089 and w14698;
w14700 <= not w14463 and w14699;
w14701 <= not w14089 and not w14098;
w14702 <= not w14463 and w14701;
w14703 <= not w14096 and not w14702;
w14704 <= not w14700 and not w14703;
w14705 <= w5062 and not w14685;
w14706 <= not w14695 and w14705;
w14707 <= not w14704 and not w14706;
w14708 <= not w14697 and not w14707;
w14709 <= not w4718 and not w14708;
w14710 <= not w14101 and w14108;
w14711 <= not w14110 and w14710;
w14712 <= not w14463 and w14711;
w14713 <= not w14101 and not w14110;
w14714 <= not w14463 and w14713;
w14715 <= not w14108 and not w14714;
w14716 <= not w14712 and not w14715;
w14717 <= w4718 and not w14697;
w14718 <= not w14707 and w14717;
w14719 <= not w14716 and not w14718;
w14720 <= not w14709 and not w14719;
w14721 <= not w4386 and not w14720;
w14722 <= w14120 and not w14122;
w14723 <= not w14113 and w14722;
w14724 <= not w14463 and w14723;
w14725 <= not w14113 and not w14122;
w14726 <= not w14463 and w14725;
w14727 <= not w14120 and not w14726;
w14728 <= not w14724 and not w14727;
w14729 <= w4386 and not w14709;
w14730 <= not w14719 and w14729;
w14731 <= not w14728 and not w14730;
w14732 <= not w14721 and not w14731;
w14733 <= not w4066 and not w14732;
w14734 <= not w14125 and w14132;
w14735 <= not w14134 and w14734;
w14736 <= not w14463 and w14735;
w14737 <= not w14125 and not w14134;
w14738 <= not w14463 and w14737;
w14739 <= not w14132 and not w14738;
w14740 <= not w14736 and not w14739;
w14741 <= w4066 and not w14721;
w14742 <= not w14731 and w14741;
w14743 <= not w14740 and not w14742;
w14744 <= not w14733 and not w14743;
w14745 <= not w3758 and not w14744;
w14746 <= w14144 and not w14146;
w14747 <= not w14137 and w14746;
w14748 <= not w14463 and w14747;
w14749 <= not w14137 and not w14146;
w14750 <= not w14463 and w14749;
w14751 <= not w14144 and not w14750;
w14752 <= not w14748 and not w14751;
w14753 <= w3758 and not w14733;
w14754 <= not w14743 and w14753;
w14755 <= not w14752 and not w14754;
w14756 <= not w14745 and not w14755;
w14757 <= not w3462 and not w14756;
w14758 <= not w14149 and w14156;
w14759 <= not w14158 and w14758;
w14760 <= not w14463 and w14759;
w14761 <= not w14149 and not w14158;
w14762 <= not w14463 and w14761;
w14763 <= not w14156 and not w14762;
w14764 <= not w14760 and not w14763;
w14765 <= w3462 and not w14745;
w14766 <= not w14755 and w14765;
w14767 <= not w14764 and not w14766;
w14768 <= not w14757 and not w14767;
w14769 <= not w3178 and not w14768;
w14770 <= w14168 and not w14170;
w14771 <= not w14161 and w14770;
w14772 <= not w14463 and w14771;
w14773 <= not w14161 and not w14170;
w14774 <= not w14463 and w14773;
w14775 <= not w14168 and not w14774;
w14776 <= not w14772 and not w14775;
w14777 <= w3178 and not w14757;
w14778 <= not w14767 and w14777;
w14779 <= not w14776 and not w14778;
w14780 <= not w14769 and not w14779;
w14781 <= not w2906 and not w14780;
w14782 <= not w14173 and w14180;
w14783 <= not w14182 and w14782;
w14784 <= not w14463 and w14783;
w14785 <= not w14173 and not w14182;
w14786 <= not w14463 and w14785;
w14787 <= not w14180 and not w14786;
w14788 <= not w14784 and not w14787;
w14789 <= w2906 and not w14769;
w14790 <= not w14779 and w14789;
w14791 <= not w14788 and not w14790;
w14792 <= not w14781 and not w14791;
w14793 <= not w2646 and not w14792;
w14794 <= w14192 and not w14194;
w14795 <= not w14185 and w14794;
w14796 <= not w14463 and w14795;
w14797 <= not w14185 and not w14194;
w14798 <= not w14463 and w14797;
w14799 <= not w14192 and not w14798;
w14800 <= not w14796 and not w14799;
w14801 <= w2646 and not w14781;
w14802 <= not w14791 and w14801;
w14803 <= not w14800 and not w14802;
w14804 <= not w14793 and not w14803;
w14805 <= not w2398 and not w14804;
w14806 <= not w14197 and w14204;
w14807 <= not w14206 and w14806;
w14808 <= not w14463 and w14807;
w14809 <= not w14197 and not w14206;
w14810 <= not w14463 and w14809;
w14811 <= not w14204 and not w14810;
w14812 <= not w14808 and not w14811;
w14813 <= w2398 and not w14793;
w14814 <= not w14803 and w14813;
w14815 <= not w14812 and not w14814;
w14816 <= not w14805 and not w14815;
w14817 <= not w2162 and not w14816;
w14818 <= w14216 and not w14218;
w14819 <= not w14209 and w14818;
w14820 <= not w14463 and w14819;
w14821 <= not w14209 and not w14218;
w14822 <= not w14463 and w14821;
w14823 <= not w14216 and not w14822;
w14824 <= not w14820 and not w14823;
w14825 <= w2162 and not w14805;
w14826 <= not w14815 and w14825;
w14827 <= not w14824 and not w14826;
w14828 <= not w14817 and not w14827;
w14829 <= not w1938 and not w14828;
w14830 <= not w14221 and w14228;
w14831 <= not w14230 and w14830;
w14832 <= not w14463 and w14831;
w14833 <= not w14221 and not w14230;
w14834 <= not w14463 and w14833;
w14835 <= not w14228 and not w14834;
w14836 <= not w14832 and not w14835;
w14837 <= w1938 and not w14817;
w14838 <= not w14827 and w14837;
w14839 <= not w14836 and not w14838;
w14840 <= not w14829 and not w14839;
w14841 <= not w1725 and not w14840;
w14842 <= w14240 and not w14242;
w14843 <= not w14233 and w14842;
w14844 <= not w14463 and w14843;
w14845 <= not w14233 and not w14242;
w14846 <= not w14463 and w14845;
w14847 <= not w14240 and not w14846;
w14848 <= not w14844 and not w14847;
w14849 <= w1725 and not w14829;
w14850 <= not w14839 and w14849;
w14851 <= not w14848 and not w14850;
w14852 <= not w14841 and not w14851;
w14853 <= not w1525 and not w14852;
w14854 <= not w14245 and w14252;
w14855 <= not w14254 and w14854;
w14856 <= not w14463 and w14855;
w14857 <= not w14245 and not w14254;
w14858 <= not w14463 and w14857;
w14859 <= not w14252 and not w14858;
w14860 <= not w14856 and not w14859;
w14861 <= w1525 and not w14841;
w14862 <= not w14851 and w14861;
w14863 <= not w14860 and not w14862;
w14864 <= not w14853 and not w14863;
w14865 <= not w1337 and not w14864;
w14866 <= w14264 and not w14266;
w14867 <= not w14257 and w14866;
w14868 <= not w14463 and w14867;
w14869 <= not w14257 and not w14266;
w14870 <= not w14463 and w14869;
w14871 <= not w14264 and not w14870;
w14872 <= not w14868 and not w14871;
w14873 <= w1337 and not w14853;
w14874 <= not w14863 and w14873;
w14875 <= not w14872 and not w14874;
w14876 <= not w14865 and not w14875;
w14877 <= not w1161 and not w14876;
w14878 <= w1161 and not w14865;
w14879 <= not w14875 and w14878;
w14880 <= not w14269 and w14278;
w14881 <= not w14271 and w14880;
w14882 <= not w14463 and w14881;
w14883 <= not w14269 and not w14271;
w14884 <= not w14463 and w14883;
w14885 <= not w14278 and not w14884;
w14886 <= not w14882 and not w14885;
w14887 <= not w14879 and not w14886;
w14888 <= not w14877 and not w14887;
w14889 <= not w997 and not w14888;
w14890 <= w14288 and not w14290;
w14891 <= not w14281 and w14890;
w14892 <= not w14463 and w14891;
w14893 <= not w14281 and not w14290;
w14894 <= not w14463 and w14893;
w14895 <= not w14288 and not w14894;
w14896 <= not w14892 and not w14895;
w14897 <= w997 and not w14877;
w14898 <= not w14887 and w14897;
w14899 <= not w14896 and not w14898;
w14900 <= not w14889 and not w14899;
w14901 <= not w845 and not w14900;
w14902 <= not w14293 and w14300;
w14903 <= not w14302 and w14902;
w14904 <= not w14463 and w14903;
w14905 <= not w14293 and not w14302;
w14906 <= not w14463 and w14905;
w14907 <= not w14300 and not w14906;
w14908 <= not w14904 and not w14907;
w14909 <= w845 and not w14889;
w14910 <= not w14899 and w14909;
w14911 <= not w14908 and not w14910;
w14912 <= not w14901 and not w14911;
w14913 <= not w705 and not w14912;
w14914 <= w14312 and not w14314;
w14915 <= not w14305 and w14914;
w14916 <= not w14463 and w14915;
w14917 <= not w14305 and not w14314;
w14918 <= not w14463 and w14917;
w14919 <= not w14312 and not w14918;
w14920 <= not w14916 and not w14919;
w14921 <= w705 and not w14901;
w14922 <= not w14911 and w14921;
w14923 <= not w14920 and not w14922;
w14924 <= not w14913 and not w14923;
w14925 <= not w577 and not w14924;
w14926 <= not w14317 and w14324;
w14927 <= not w14326 and w14926;
w14928 <= not w14463 and w14927;
w14929 <= not w14317 and not w14326;
w14930 <= not w14463 and w14929;
w14931 <= not w14324 and not w14930;
w14932 <= not w14928 and not w14931;
w14933 <= w577 and not w14913;
w14934 <= not w14923 and w14933;
w14935 <= not w14932 and not w14934;
w14936 <= not w14925 and not w14935;
w14937 <= not w460 and not w14936;
w14938 <= w14336 and not w14338;
w14939 <= not w14329 and w14938;
w14940 <= not w14463 and w14939;
w14941 <= not w14329 and not w14338;
w14942 <= not w14463 and w14941;
w14943 <= not w14336 and not w14942;
w14944 <= not w14940 and not w14943;
w14945 <= w460 and not w14925;
w14946 <= not w14935 and w14945;
w14947 <= not w14944 and not w14946;
w14948 <= not w14937 and not w14947;
w14949 <= not w356 and not w14948;
w14950 <= not w14341 and w14348;
w14951 <= not w14350 and w14950;
w14952 <= not w14463 and w14951;
w14953 <= not w14341 and not w14350;
w14954 <= not w14463 and w14953;
w14955 <= not w14348 and not w14954;
w14956 <= not w14952 and not w14955;
w14957 <= w356 and not w14937;
w14958 <= not w14947 and w14957;
w14959 <= not w14956 and not w14958;
w14960 <= not w14949 and not w14959;
w14961 <= not w264 and not w14960;
w14962 <= w14360 and not w14362;
w14963 <= not w14353 and w14962;
w14964 <= not w14463 and w14963;
w14965 <= not w14353 and not w14362;
w14966 <= not w14463 and w14965;
w14967 <= not w14360 and not w14966;
w14968 <= not w14964 and not w14967;
w14969 <= w264 and not w14949;
w14970 <= not w14959 and w14969;
w14971 <= not w14968 and not w14970;
w14972 <= not w14961 and not w14971;
w14973 <= not w184 and not w14972;
w14974 <= not w14365 and w14372;
w14975 <= not w14374 and w14974;
w14976 <= not w14463 and w14975;
w14977 <= not w14365 and not w14374;
w14978 <= not w14463 and w14977;
w14979 <= not w14372 and not w14978;
w14980 <= not w14976 and not w14979;
w14981 <= w184 and not w14961;
w14982 <= not w14971 and w14981;
w14983 <= not w14980 and not w14982;
w14984 <= not w14973 and not w14983;
w14985 <= not w115 and not w14984;
w14986 <= w14384 and not w14386;
w14987 <= not w14377 and w14986;
w14988 <= not w14463 and w14987;
w14989 <= not w14377 and not w14386;
w14990 <= not w14463 and w14989;
w14991 <= not w14384 and not w14990;
w14992 <= not w14988 and not w14991;
w14993 <= w115 and not w14973;
w14994 <= not w14983 and w14993;
w14995 <= not w14992 and not w14994;
w14996 <= not w14985 and not w14995;
w14997 <= not w60 and not w14996;
w14998 <= not w14389 and w14396;
w14999 <= not w14398 and w14998;
w15000 <= not w14463 and w14999;
w15001 <= not w14389 and not w14398;
w15002 <= not w14463 and w15001;
w15003 <= not w14396 and not w15002;
w15004 <= not w15000 and not w15003;
w15005 <= w60 and not w14985;
w15006 <= not w14995 and w15005;
w15007 <= not w15004 and not w15006;
w15008 <= not w14997 and not w15007;
w15009 <= not w22 and not w15008;
w15010 <= w14408 and not w14410;
w15011 <= not w14401 and w15010;
w15012 <= not w14463 and w15011;
w15013 <= not w14401 and not w14410;
w15014 <= not w14463 and w15013;
w15015 <= not w14408 and not w15014;
w15016 <= not w15012 and not w15015;
w15017 <= w22 and not w14997;
w15018 <= not w15007 and w15017;
w15019 <= not w15016 and not w15018;
w15020 <= not w15009 and not w15019;
w15021 <= not w5 and not w15020;
w15022 <= not w14413 and w14420;
w15023 <= not w14422 and w15022;
w15024 <= not w14463 and w15023;
w15025 <= not w14413 and not w14422;
w15026 <= not w14463 and w15025;
w15027 <= not w14420 and not w15026;
w15028 <= not w15024 and not w15027;
w15029 <= w5 and not w15009;
w15030 <= not w15019 and w15029;
w15031 <= not w15028 and not w15030;
w15032 <= not w15021 and not w15031;
w15033 <= w14432 and not w14434;
w15034 <= not w14425 and w15033;
w15035 <= not w14463 and w15034;
w15036 <= not w14425 and not w14434;
w15037 <= not w14463 and w15036;
w15038 <= not w14432 and not w15037;
w15039 <= not w15035 and not w15038;
w15040 <= not w14436 and not w14443;
w15041 <= not w14463 and w15040;
w15042 <= not w14451 and not w15041;
w15043 <= not w15039 and w15042;
w15044 <= not w15032 and w15043;
w15045 <= w0 and not w15044;
w15046 <= not w15021 and w15039;
w15047 <= not w15031 and w15046;
w15048 <= not w14443 and not w14463;
w15049 <= w14436 and not w15048;
w15050 <= not w0 and not w15040;
w15051 <= not w15049 and w15050;
w15052 <= not w14439 and not w14460;
w15053 <= not w14442 and w15052;
w15054 <= not w14455 and w15053;
w15055 <= not w14451 and w15054;
w15056 <= not w14449 and w15055;
w15057 <= not w15051 and not w15056;
w15058 <= not w15047 and w15057;
w15059 <= not w15045 and w15058;
w15060 <= a(28) and not w15059;
w15061 <= not a(26) and not a(27);
w15062 <= not a(28) and w15061;
w15063 <= not w15060 and not w15062;
w15064 <= not w14463 and not w15063;
w15065 <= not w14460 and not w15062;
w15066 <= not w14455 and w15065;
w15067 <= not w14451 and w15066;
w15068 <= not w14449 and w15067;
w15069 <= not w15060 and w15068;
w15070 <= not a(28) and not w15059;
w15071 <= a(29) and not w15070;
w15072 <= w14465 and not w15059;
w15073 <= not w15071 and not w15072;
w15074 <= not w15069 and w15073;
w15075 <= not w15064 and not w15074;
w15076 <= not w13879 and not w15075;
w15077 <= w13879 and not w15064;
w15078 <= not w15074 and w15077;
w15079 <= not w14463 and not w15056;
w15080 <= not w15051 and w15079;
w15081 <= not w15047 and w15080;
w15082 <= not w15045 and w15081;
w15083 <= not w15072 and not w15082;
w15084 <= a(30) and not w15083;
w15085 <= not a(30) and not w15082;
w15086 <= not w15072 and w15085;
w15087 <= not w15084 and not w15086;
w15088 <= not w15078 and not w15087;
w15089 <= not w15076 and not w15088;
w15090 <= not w13307 and not w15089;
w15091 <= not w14468 and not w14473;
w15092 <= not w14477 and w15091;
w15093 <= not w15059 and w15092;
w15094 <= not w15059 and w15091;
w15095 <= w14477 and not w15094;
w15096 <= not w15093 and not w15095;
w15097 <= w13307 and not w15076;
w15098 <= not w15088 and w15097;
w15099 <= not w15096 and not w15098;
w15100 <= not w15090 and not w15099;
w15101 <= not w12747 and not w15100;
w15102 <= not w14482 and w14491;
w15103 <= not w14480 and w15102;
w15104 <= not w15059 and w15103;
w15105 <= not w14480 and not w14482;
w15106 <= not w15059 and w15105;
w15107 <= not w14491 and not w15106;
w15108 <= not w15104 and not w15107;
w15109 <= w12747 and not w15090;
w15110 <= not w15099 and w15109;
w15111 <= not w15108 and not w15110;
w15112 <= not w15101 and not w15111;
w15113 <= not w12199 and not w15112;
w15114 <= not w14494 and w14500;
w15115 <= not w14502 and w15114;
w15116 <= not w15059 and w15115;
w15117 <= not w14494 and not w14502;
w15118 <= not w15059 and w15117;
w15119 <= not w14500 and not w15118;
w15120 <= not w15116 and not w15119;
w15121 <= w12199 and not w15101;
w15122 <= not w15111 and w15121;
w15123 <= not w15120 and not w15122;
w15124 <= not w15113 and not w15123;
w15125 <= not w11663 and not w15124;
w15126 <= w14512 and not w14514;
w15127 <= not w14505 and w15126;
w15128 <= not w15059 and w15127;
w15129 <= not w14505 and not w14514;
w15130 <= not w15059 and w15129;
w15131 <= not w14512 and not w15130;
w15132 <= not w15128 and not w15131;
w15133 <= w11663 and not w15113;
w15134 <= not w15123 and w15133;
w15135 <= not w15132 and not w15134;
w15136 <= not w15125 and not w15135;
w15137 <= not w11139 and not w15136;
w15138 <= not w14517 and w14524;
w15139 <= not w14526 and w15138;
w15140 <= not w15059 and w15139;
w15141 <= not w14517 and not w14526;
w15142 <= not w15059 and w15141;
w15143 <= not w14524 and not w15142;
w15144 <= not w15140 and not w15143;
w15145 <= w11139 and not w15125;
w15146 <= not w15135 and w15145;
w15147 <= not w15144 and not w15146;
w15148 <= not w15137 and not w15147;
w15149 <= not w10627 and not w15148;
w15150 <= w14536 and not w14538;
w15151 <= not w14529 and w15150;
w15152 <= not w15059 and w15151;
w15153 <= not w14529 and not w14538;
w15154 <= not w15059 and w15153;
w15155 <= not w14536 and not w15154;
w15156 <= not w15152 and not w15155;
w15157 <= w10627 and not w15137;
w15158 <= not w15147 and w15157;
w15159 <= not w15156 and not w15158;
w15160 <= not w15149 and not w15159;
w15161 <= not w10127 and not w15160;
w15162 <= not w14541 and w14548;
w15163 <= not w14550 and w15162;
w15164 <= not w15059 and w15163;
w15165 <= not w14541 and not w14550;
w15166 <= not w15059 and w15165;
w15167 <= not w14548 and not w15166;
w15168 <= not w15164 and not w15167;
w15169 <= w10127 and not w15149;
w15170 <= not w15159 and w15169;
w15171 <= not w15168 and not w15170;
w15172 <= not w15161 and not w15171;
w15173 <= not w9639 and not w15172;
w15174 <= w14560 and not w14562;
w15175 <= not w14553 and w15174;
w15176 <= not w15059 and w15175;
w15177 <= not w14553 and not w14562;
w15178 <= not w15059 and w15177;
w15179 <= not w14560 and not w15178;
w15180 <= not w15176 and not w15179;
w15181 <= w9639 and not w15161;
w15182 <= not w15171 and w15181;
w15183 <= not w15180 and not w15182;
w15184 <= not w15173 and not w15183;
w15185 <= not w9163 and not w15184;
w15186 <= not w14565 and w14572;
w15187 <= not w14574 and w15186;
w15188 <= not w15059 and w15187;
w15189 <= not w14565 and not w14574;
w15190 <= not w15059 and w15189;
w15191 <= not w14572 and not w15190;
w15192 <= not w15188 and not w15191;
w15193 <= w9163 and not w15173;
w15194 <= not w15183 and w15193;
w15195 <= not w15192 and not w15194;
w15196 <= not w15185 and not w15195;
w15197 <= not w8699 and not w15196;
w15198 <= w14584 and not w14586;
w15199 <= not w14577 and w15198;
w15200 <= not w15059 and w15199;
w15201 <= not w14577 and not w14586;
w15202 <= not w15059 and w15201;
w15203 <= not w14584 and not w15202;
w15204 <= not w15200 and not w15203;
w15205 <= w8699 and not w15185;
w15206 <= not w15195 and w15205;
w15207 <= not w15204 and not w15206;
w15208 <= not w15197 and not w15207;
w15209 <= not w8247 and not w15208;
w15210 <= not w14589 and w14596;
w15211 <= not w14598 and w15210;
w15212 <= not w15059 and w15211;
w15213 <= not w14589 and not w14598;
w15214 <= not w15059 and w15213;
w15215 <= not w14596 and not w15214;
w15216 <= not w15212 and not w15215;
w15217 <= w8247 and not w15197;
w15218 <= not w15207 and w15217;
w15219 <= not w15216 and not w15218;
w15220 <= not w15209 and not w15219;
w15221 <= not w7807 and not w15220;
w15222 <= w14608 and not w14610;
w15223 <= not w14601 and w15222;
w15224 <= not w15059 and w15223;
w15225 <= not w14601 and not w14610;
w15226 <= not w15059 and w15225;
w15227 <= not w14608 and not w15226;
w15228 <= not w15224 and not w15227;
w15229 <= w7807 and not w15209;
w15230 <= not w15219 and w15229;
w15231 <= not w15228 and not w15230;
w15232 <= not w15221 and not w15231;
w15233 <= not w7379 and not w15232;
w15234 <= not w14613 and w14620;
w15235 <= not w14622 and w15234;
w15236 <= not w15059 and w15235;
w15237 <= not w14613 and not w14622;
w15238 <= not w15059 and w15237;
w15239 <= not w14620 and not w15238;
w15240 <= not w15236 and not w15239;
w15241 <= w7379 and not w15221;
w15242 <= not w15231 and w15241;
w15243 <= not w15240 and not w15242;
w15244 <= not w15233 and not w15243;
w15245 <= not w6963 and not w15244;
w15246 <= w14632 and not w14634;
w15247 <= not w14625 and w15246;
w15248 <= not w15059 and w15247;
w15249 <= not w14625 and not w14634;
w15250 <= not w15059 and w15249;
w15251 <= not w14632 and not w15250;
w15252 <= not w15248 and not w15251;
w15253 <= w6963 and not w15233;
w15254 <= not w15243 and w15253;
w15255 <= not w15252 and not w15254;
w15256 <= not w15245 and not w15255;
w15257 <= not w6558 and not w15256;
w15258 <= not w14637 and w14644;
w15259 <= not w14646 and w15258;
w15260 <= not w15059 and w15259;
w15261 <= not w14637 and not w14646;
w15262 <= not w15059 and w15261;
w15263 <= not w14644 and not w15262;
w15264 <= not w15260 and not w15263;
w15265 <= w6558 and not w15245;
w15266 <= not w15255 and w15265;
w15267 <= not w15264 and not w15266;
w15268 <= not w15257 and not w15267;
w15269 <= not w6166 and not w15268;
w15270 <= w14656 and not w14658;
w15271 <= not w14649 and w15270;
w15272 <= not w15059 and w15271;
w15273 <= not w14649 and not w14658;
w15274 <= not w15059 and w15273;
w15275 <= not w14656 and not w15274;
w15276 <= not w15272 and not w15275;
w15277 <= w6166 and not w15257;
w15278 <= not w15267 and w15277;
w15279 <= not w15276 and not w15278;
w15280 <= not w15269 and not w15279;
w15281 <= not w5786 and not w15280;
w15282 <= not w14661 and w14668;
w15283 <= not w14670 and w15282;
w15284 <= not w15059 and w15283;
w15285 <= not w14661 and not w14670;
w15286 <= not w15059 and w15285;
w15287 <= not w14668 and not w15286;
w15288 <= not w15284 and not w15287;
w15289 <= w5786 and not w15269;
w15290 <= not w15279 and w15289;
w15291 <= not w15288 and not w15290;
w15292 <= not w15281 and not w15291;
w15293 <= not w5418 and not w15292;
w15294 <= w14680 and not w14682;
w15295 <= not w14673 and w15294;
w15296 <= not w15059 and w15295;
w15297 <= not w14673 and not w14682;
w15298 <= not w15059 and w15297;
w15299 <= not w14680 and not w15298;
w15300 <= not w15296 and not w15299;
w15301 <= w5418 and not w15281;
w15302 <= not w15291 and w15301;
w15303 <= not w15300 and not w15302;
w15304 <= not w15293 and not w15303;
w15305 <= not w5062 and not w15304;
w15306 <= not w14685 and w14692;
w15307 <= not w14694 and w15306;
w15308 <= not w15059 and w15307;
w15309 <= not w14685 and not w14694;
w15310 <= not w15059 and w15309;
w15311 <= not w14692 and not w15310;
w15312 <= not w15308 and not w15311;
w15313 <= w5062 and not w15293;
w15314 <= not w15303 and w15313;
w15315 <= not w15312 and not w15314;
w15316 <= not w15305 and not w15315;
w15317 <= not w4718 and not w15316;
w15318 <= w14704 and not w14706;
w15319 <= not w14697 and w15318;
w15320 <= not w15059 and w15319;
w15321 <= not w14697 and not w14706;
w15322 <= not w15059 and w15321;
w15323 <= not w14704 and not w15322;
w15324 <= not w15320 and not w15323;
w15325 <= w4718 and not w15305;
w15326 <= not w15315 and w15325;
w15327 <= not w15324 and not w15326;
w15328 <= not w15317 and not w15327;
w15329 <= not w4386 and not w15328;
w15330 <= not w14709 and w14716;
w15331 <= not w14718 and w15330;
w15332 <= not w15059 and w15331;
w15333 <= not w14709 and not w14718;
w15334 <= not w15059 and w15333;
w15335 <= not w14716 and not w15334;
w15336 <= not w15332 and not w15335;
w15337 <= w4386 and not w15317;
w15338 <= not w15327 and w15337;
w15339 <= not w15336 and not w15338;
w15340 <= not w15329 and not w15339;
w15341 <= not w4066 and not w15340;
w15342 <= w14728 and not w14730;
w15343 <= not w14721 and w15342;
w15344 <= not w15059 and w15343;
w15345 <= not w14721 and not w14730;
w15346 <= not w15059 and w15345;
w15347 <= not w14728 and not w15346;
w15348 <= not w15344 and not w15347;
w15349 <= w4066 and not w15329;
w15350 <= not w15339 and w15349;
w15351 <= not w15348 and not w15350;
w15352 <= not w15341 and not w15351;
w15353 <= not w3758 and not w15352;
w15354 <= not w14733 and w14740;
w15355 <= not w14742 and w15354;
w15356 <= not w15059 and w15355;
w15357 <= not w14733 and not w14742;
w15358 <= not w15059 and w15357;
w15359 <= not w14740 and not w15358;
w15360 <= not w15356 and not w15359;
w15361 <= w3758 and not w15341;
w15362 <= not w15351 and w15361;
w15363 <= not w15360 and not w15362;
w15364 <= not w15353 and not w15363;
w15365 <= not w3462 and not w15364;
w15366 <= w14752 and not w14754;
w15367 <= not w14745 and w15366;
w15368 <= not w15059 and w15367;
w15369 <= not w14745 and not w14754;
w15370 <= not w15059 and w15369;
w15371 <= not w14752 and not w15370;
w15372 <= not w15368 and not w15371;
w15373 <= w3462 and not w15353;
w15374 <= not w15363 and w15373;
w15375 <= not w15372 and not w15374;
w15376 <= not w15365 and not w15375;
w15377 <= not w3178 and not w15376;
w15378 <= not w14757 and w14764;
w15379 <= not w14766 and w15378;
w15380 <= not w15059 and w15379;
w15381 <= not w14757 and not w14766;
w15382 <= not w15059 and w15381;
w15383 <= not w14764 and not w15382;
w15384 <= not w15380 and not w15383;
w15385 <= w3178 and not w15365;
w15386 <= not w15375 and w15385;
w15387 <= not w15384 and not w15386;
w15388 <= not w15377 and not w15387;
w15389 <= not w2906 and not w15388;
w15390 <= w14776 and not w14778;
w15391 <= not w14769 and w15390;
w15392 <= not w15059 and w15391;
w15393 <= not w14769 and not w14778;
w15394 <= not w15059 and w15393;
w15395 <= not w14776 and not w15394;
w15396 <= not w15392 and not w15395;
w15397 <= w2906 and not w15377;
w15398 <= not w15387 and w15397;
w15399 <= not w15396 and not w15398;
w15400 <= not w15389 and not w15399;
w15401 <= not w2646 and not w15400;
w15402 <= not w14781 and w14788;
w15403 <= not w14790 and w15402;
w15404 <= not w15059 and w15403;
w15405 <= not w14781 and not w14790;
w15406 <= not w15059 and w15405;
w15407 <= not w14788 and not w15406;
w15408 <= not w15404 and not w15407;
w15409 <= w2646 and not w15389;
w15410 <= not w15399 and w15409;
w15411 <= not w15408 and not w15410;
w15412 <= not w15401 and not w15411;
w15413 <= not w2398 and not w15412;
w15414 <= w14800 and not w14802;
w15415 <= not w14793 and w15414;
w15416 <= not w15059 and w15415;
w15417 <= not w14793 and not w14802;
w15418 <= not w15059 and w15417;
w15419 <= not w14800 and not w15418;
w15420 <= not w15416 and not w15419;
w15421 <= w2398 and not w15401;
w15422 <= not w15411 and w15421;
w15423 <= not w15420 and not w15422;
w15424 <= not w15413 and not w15423;
w15425 <= not w2162 and not w15424;
w15426 <= not w14805 and w14812;
w15427 <= not w14814 and w15426;
w15428 <= not w15059 and w15427;
w15429 <= not w14805 and not w14814;
w15430 <= not w15059 and w15429;
w15431 <= not w14812 and not w15430;
w15432 <= not w15428 and not w15431;
w15433 <= w2162 and not w15413;
w15434 <= not w15423 and w15433;
w15435 <= not w15432 and not w15434;
w15436 <= not w15425 and not w15435;
w15437 <= not w1938 and not w15436;
w15438 <= w14824 and not w14826;
w15439 <= not w14817 and w15438;
w15440 <= not w15059 and w15439;
w15441 <= not w14817 and not w14826;
w15442 <= not w15059 and w15441;
w15443 <= not w14824 and not w15442;
w15444 <= not w15440 and not w15443;
w15445 <= w1938 and not w15425;
w15446 <= not w15435 and w15445;
w15447 <= not w15444 and not w15446;
w15448 <= not w15437 and not w15447;
w15449 <= not w1725 and not w15448;
w15450 <= not w14829 and w14836;
w15451 <= not w14838 and w15450;
w15452 <= not w15059 and w15451;
w15453 <= not w14829 and not w14838;
w15454 <= not w15059 and w15453;
w15455 <= not w14836 and not w15454;
w15456 <= not w15452 and not w15455;
w15457 <= w1725 and not w15437;
w15458 <= not w15447 and w15457;
w15459 <= not w15456 and not w15458;
w15460 <= not w15449 and not w15459;
w15461 <= not w1525 and not w15460;
w15462 <= w14848 and not w14850;
w15463 <= not w14841 and w15462;
w15464 <= not w15059 and w15463;
w15465 <= not w14841 and not w14850;
w15466 <= not w15059 and w15465;
w15467 <= not w14848 and not w15466;
w15468 <= not w15464 and not w15467;
w15469 <= w1525 and not w15449;
w15470 <= not w15459 and w15469;
w15471 <= not w15468 and not w15470;
w15472 <= not w15461 and not w15471;
w15473 <= not w1337 and not w15472;
w15474 <= not w14853 and w14860;
w15475 <= not w14862 and w15474;
w15476 <= not w15059 and w15475;
w15477 <= not w14853 and not w14862;
w15478 <= not w15059 and w15477;
w15479 <= not w14860 and not w15478;
w15480 <= not w15476 and not w15479;
w15481 <= w1337 and not w15461;
w15482 <= not w15471 and w15481;
w15483 <= not w15480 and not w15482;
w15484 <= not w15473 and not w15483;
w15485 <= not w1161 and not w15484;
w15486 <= w14872 and not w14874;
w15487 <= not w14865 and w15486;
w15488 <= not w15059 and w15487;
w15489 <= not w14865 and not w14874;
w15490 <= not w15059 and w15489;
w15491 <= not w14872 and not w15490;
w15492 <= not w15488 and not w15491;
w15493 <= w1161 and not w15473;
w15494 <= not w15483 and w15493;
w15495 <= not w15492 and not w15494;
w15496 <= not w15485 and not w15495;
w15497 <= not w997 and not w15496;
w15498 <= w997 and not w15485;
w15499 <= not w15495 and w15498;
w15500 <= not w14877 and w14886;
w15501 <= not w14879 and w15500;
w15502 <= not w15059 and w15501;
w15503 <= not w14877 and not w14879;
w15504 <= not w15059 and w15503;
w15505 <= not w14886 and not w15504;
w15506 <= not w15502 and not w15505;
w15507 <= not w15499 and not w15506;
w15508 <= not w15497 and not w15507;
w15509 <= not w845 and not w15508;
w15510 <= w14896 and not w14898;
w15511 <= not w14889 and w15510;
w15512 <= not w15059 and w15511;
w15513 <= not w14889 and not w14898;
w15514 <= not w15059 and w15513;
w15515 <= not w14896 and not w15514;
w15516 <= not w15512 and not w15515;
w15517 <= w845 and not w15497;
w15518 <= not w15507 and w15517;
w15519 <= not w15516 and not w15518;
w15520 <= not w15509 and not w15519;
w15521 <= not w705 and not w15520;
w15522 <= not w14901 and w14908;
w15523 <= not w14910 and w15522;
w15524 <= not w15059 and w15523;
w15525 <= not w14901 and not w14910;
w15526 <= not w15059 and w15525;
w15527 <= not w14908 and not w15526;
w15528 <= not w15524 and not w15527;
w15529 <= w705 and not w15509;
w15530 <= not w15519 and w15529;
w15531 <= not w15528 and not w15530;
w15532 <= not w15521 and not w15531;
w15533 <= not w577 and not w15532;
w15534 <= w14920 and not w14922;
w15535 <= not w14913 and w15534;
w15536 <= not w15059 and w15535;
w15537 <= not w14913 and not w14922;
w15538 <= not w15059 and w15537;
w15539 <= not w14920 and not w15538;
w15540 <= not w15536 and not w15539;
w15541 <= w577 and not w15521;
w15542 <= not w15531 and w15541;
w15543 <= not w15540 and not w15542;
w15544 <= not w15533 and not w15543;
w15545 <= not w460 and not w15544;
w15546 <= not w14925 and w14932;
w15547 <= not w14934 and w15546;
w15548 <= not w15059 and w15547;
w15549 <= not w14925 and not w14934;
w15550 <= not w15059 and w15549;
w15551 <= not w14932 and not w15550;
w15552 <= not w15548 and not w15551;
w15553 <= w460 and not w15533;
w15554 <= not w15543 and w15553;
w15555 <= not w15552 and not w15554;
w15556 <= not w15545 and not w15555;
w15557 <= not w356 and not w15556;
w15558 <= w14944 and not w14946;
w15559 <= not w14937 and w15558;
w15560 <= not w15059 and w15559;
w15561 <= not w14937 and not w14946;
w15562 <= not w15059 and w15561;
w15563 <= not w14944 and not w15562;
w15564 <= not w15560 and not w15563;
w15565 <= w356 and not w15545;
w15566 <= not w15555 and w15565;
w15567 <= not w15564 and not w15566;
w15568 <= not w15557 and not w15567;
w15569 <= not w264 and not w15568;
w15570 <= not w14949 and w14956;
w15571 <= not w14958 and w15570;
w15572 <= not w15059 and w15571;
w15573 <= not w14949 and not w14958;
w15574 <= not w15059 and w15573;
w15575 <= not w14956 and not w15574;
w15576 <= not w15572 and not w15575;
w15577 <= w264 and not w15557;
w15578 <= not w15567 and w15577;
w15579 <= not w15576 and not w15578;
w15580 <= not w15569 and not w15579;
w15581 <= not w184 and not w15580;
w15582 <= w14968 and not w14970;
w15583 <= not w14961 and w15582;
w15584 <= not w15059 and w15583;
w15585 <= not w14961 and not w14970;
w15586 <= not w15059 and w15585;
w15587 <= not w14968 and not w15586;
w15588 <= not w15584 and not w15587;
w15589 <= w184 and not w15569;
w15590 <= not w15579 and w15589;
w15591 <= not w15588 and not w15590;
w15592 <= not w15581 and not w15591;
w15593 <= not w115 and not w15592;
w15594 <= not w14973 and w14980;
w15595 <= not w14982 and w15594;
w15596 <= not w15059 and w15595;
w15597 <= not w14973 and not w14982;
w15598 <= not w15059 and w15597;
w15599 <= not w14980 and not w15598;
w15600 <= not w15596 and not w15599;
w15601 <= w115 and not w15581;
w15602 <= not w15591 and w15601;
w15603 <= not w15600 and not w15602;
w15604 <= not w15593 and not w15603;
w15605 <= not w60 and not w15604;
w15606 <= w14992 and not w14994;
w15607 <= not w14985 and w15606;
w15608 <= not w15059 and w15607;
w15609 <= not w14985 and not w14994;
w15610 <= not w15059 and w15609;
w15611 <= not w14992 and not w15610;
w15612 <= not w15608 and not w15611;
w15613 <= w60 and not w15593;
w15614 <= not w15603 and w15613;
w15615 <= not w15612 and not w15614;
w15616 <= not w15605 and not w15615;
w15617 <= not w22 and not w15616;
w15618 <= not w14997 and w15004;
w15619 <= not w15006 and w15618;
w15620 <= not w15059 and w15619;
w15621 <= not w14997 and not w15006;
w15622 <= not w15059 and w15621;
w15623 <= not w15004 and not w15622;
w15624 <= not w15620 and not w15623;
w15625 <= w22 and not w15605;
w15626 <= not w15615 and w15625;
w15627 <= not w15624 and not w15626;
w15628 <= not w15617 and not w15627;
w15629 <= not w5 and not w15628;
w15630 <= w15016 and not w15018;
w15631 <= not w15009 and w15630;
w15632 <= not w15059 and w15631;
w15633 <= not w15009 and not w15018;
w15634 <= not w15059 and w15633;
w15635 <= not w15016 and not w15634;
w15636 <= not w15632 and not w15635;
w15637 <= w5 and not w15617;
w15638 <= not w15627 and w15637;
w15639 <= not w15636 and not w15638;
w15640 <= not w15629 and not w15639;
w15641 <= not w15021 and w15028;
w15642 <= not w15030 and w15641;
w15643 <= not w15059 and w15642;
w15644 <= not w15021 and not w15030;
w15645 <= not w15059 and w15644;
w15646 <= not w15028 and not w15645;
w15647 <= not w15643 and not w15646;
w15648 <= not w15032 and not w15039;
w15649 <= not w15059 and w15648;
w15650 <= not w15047 and not w15649;
w15651 <= not w15647 and w15650;
w15652 <= not w15640 and w15651;
w15653 <= w0 and not w15652;
w15654 <= not w15629 and w15647;
w15655 <= not w15639 and w15654;
w15656 <= not w15039 and not w15059;
w15657 <= w15032 and not w15656;
w15658 <= not w0 and not w15648;
w15659 <= not w15657 and w15658;
w15660 <= not w15035 and not w15056;
w15661 <= not w15038 and w15660;
w15662 <= not w15051 and w15661;
w15663 <= not w15047 and w15662;
w15664 <= not w15045 and w15663;
w15665 <= not w15659 and not w15664;
w15666 <= not w15655 and w15665;
w15667 <= not w15653 and w15666;
w15668 <= a(26) and not w15667;
w15669 <= not a(24) and not a(25);
w15670 <= not a(26) and w15669;
w15671 <= not w15668 and not w15670;
w15672 <= not w15059 and not w15671;
w15673 <= not w15056 and not w15670;
w15674 <= not w15051 and w15673;
w15675 <= not w15047 and w15674;
w15676 <= not w15045 and w15675;
w15677 <= not w15668 and w15676;
w15678 <= not a(26) and not w15667;
w15679 <= a(27) and not w15678;
w15680 <= w15061 and not w15667;
w15681 <= not w15679 and not w15680;
w15682 <= not w15677 and w15681;
w15683 <= not w15672 and not w15682;
w15684 <= not w14463 and not w15683;
w15685 <= w14463 and not w15672;
w15686 <= not w15682 and w15685;
w15687 <= not w15059 and not w15664;
w15688 <= not w15659 and w15687;
w15689 <= not w15655 and w15688;
w15690 <= not w15653 and w15689;
w15691 <= not w15680 and not w15690;
w15692 <= a(28) and not w15691;
w15693 <= not a(28) and not w15690;
w15694 <= not w15680 and w15693;
w15695 <= not w15692 and not w15694;
w15696 <= not w15686 and not w15695;
w15697 <= not w15684 and not w15696;
w15698 <= not w13879 and not w15697;
w15699 <= not w15064 and not w15069;
w15700 <= not w15073 and w15699;
w15701 <= not w15667 and w15700;
w15702 <= not w15667 and w15699;
w15703 <= w15073 and not w15702;
w15704 <= not w15701 and not w15703;
w15705 <= w13879 and not w15684;
w15706 <= not w15696 and w15705;
w15707 <= not w15704 and not w15706;
w15708 <= not w15698 and not w15707;
w15709 <= not w13307 and not w15708;
w15710 <= not w15078 and w15087;
w15711 <= not w15076 and w15710;
w15712 <= not w15667 and w15711;
w15713 <= not w15076 and not w15078;
w15714 <= not w15667 and w15713;
w15715 <= not w15087 and not w15714;
w15716 <= not w15712 and not w15715;
w15717 <= w13307 and not w15698;
w15718 <= not w15707 and w15717;
w15719 <= not w15716 and not w15718;
w15720 <= not w15709 and not w15719;
w15721 <= not w12747 and not w15720;
w15722 <= not w15090 and w15096;
w15723 <= not w15098 and w15722;
w15724 <= not w15667 and w15723;
w15725 <= not w15090 and not w15098;
w15726 <= not w15667 and w15725;
w15727 <= not w15096 and not w15726;
w15728 <= not w15724 and not w15727;
w15729 <= w12747 and not w15709;
w15730 <= not w15719 and w15729;
w15731 <= not w15728 and not w15730;
w15732 <= not w15721 and not w15731;
w15733 <= not w12199 and not w15732;
w15734 <= w15108 and not w15110;
w15735 <= not w15101 and w15734;
w15736 <= not w15667 and w15735;
w15737 <= not w15101 and not w15110;
w15738 <= not w15667 and w15737;
w15739 <= not w15108 and not w15738;
w15740 <= not w15736 and not w15739;
w15741 <= w12199 and not w15721;
w15742 <= not w15731 and w15741;
w15743 <= not w15740 and not w15742;
w15744 <= not w15733 and not w15743;
w15745 <= not w11663 and not w15744;
w15746 <= not w15113 and w15120;
w15747 <= not w15122 and w15746;
w15748 <= not w15667 and w15747;
w15749 <= not w15113 and not w15122;
w15750 <= not w15667 and w15749;
w15751 <= not w15120 and not w15750;
w15752 <= not w15748 and not w15751;
w15753 <= w11663 and not w15733;
w15754 <= not w15743 and w15753;
w15755 <= not w15752 and not w15754;
w15756 <= not w15745 and not w15755;
w15757 <= not w11139 and not w15756;
w15758 <= w15132 and not w15134;
w15759 <= not w15125 and w15758;
w15760 <= not w15667 and w15759;
w15761 <= not w15125 and not w15134;
w15762 <= not w15667 and w15761;
w15763 <= not w15132 and not w15762;
w15764 <= not w15760 and not w15763;
w15765 <= w11139 and not w15745;
w15766 <= not w15755 and w15765;
w15767 <= not w15764 and not w15766;
w15768 <= not w15757 and not w15767;
w15769 <= not w10627 and not w15768;
w15770 <= not w15137 and w15144;
w15771 <= not w15146 and w15770;
w15772 <= not w15667 and w15771;
w15773 <= not w15137 and not w15146;
w15774 <= not w15667 and w15773;
w15775 <= not w15144 and not w15774;
w15776 <= not w15772 and not w15775;
w15777 <= w10627 and not w15757;
w15778 <= not w15767 and w15777;
w15779 <= not w15776 and not w15778;
w15780 <= not w15769 and not w15779;
w15781 <= not w10127 and not w15780;
w15782 <= w15156 and not w15158;
w15783 <= not w15149 and w15782;
w15784 <= not w15667 and w15783;
w15785 <= not w15149 and not w15158;
w15786 <= not w15667 and w15785;
w15787 <= not w15156 and not w15786;
w15788 <= not w15784 and not w15787;
w15789 <= w10127 and not w15769;
w15790 <= not w15779 and w15789;
w15791 <= not w15788 and not w15790;
w15792 <= not w15781 and not w15791;
w15793 <= not w9639 and not w15792;
w15794 <= not w15161 and w15168;
w15795 <= not w15170 and w15794;
w15796 <= not w15667 and w15795;
w15797 <= not w15161 and not w15170;
w15798 <= not w15667 and w15797;
w15799 <= not w15168 and not w15798;
w15800 <= not w15796 and not w15799;
w15801 <= w9639 and not w15781;
w15802 <= not w15791 and w15801;
w15803 <= not w15800 and not w15802;
w15804 <= not w15793 and not w15803;
w15805 <= not w9163 and not w15804;
w15806 <= w15180 and not w15182;
w15807 <= not w15173 and w15806;
w15808 <= not w15667 and w15807;
w15809 <= not w15173 and not w15182;
w15810 <= not w15667 and w15809;
w15811 <= not w15180 and not w15810;
w15812 <= not w15808 and not w15811;
w15813 <= w9163 and not w15793;
w15814 <= not w15803 and w15813;
w15815 <= not w15812 and not w15814;
w15816 <= not w15805 and not w15815;
w15817 <= not w8699 and not w15816;
w15818 <= not w15185 and w15192;
w15819 <= not w15194 and w15818;
w15820 <= not w15667 and w15819;
w15821 <= not w15185 and not w15194;
w15822 <= not w15667 and w15821;
w15823 <= not w15192 and not w15822;
w15824 <= not w15820 and not w15823;
w15825 <= w8699 and not w15805;
w15826 <= not w15815 and w15825;
w15827 <= not w15824 and not w15826;
w15828 <= not w15817 and not w15827;
w15829 <= not w8247 and not w15828;
w15830 <= w15204 and not w15206;
w15831 <= not w15197 and w15830;
w15832 <= not w15667 and w15831;
w15833 <= not w15197 and not w15206;
w15834 <= not w15667 and w15833;
w15835 <= not w15204 and not w15834;
w15836 <= not w15832 and not w15835;
w15837 <= w8247 and not w15817;
w15838 <= not w15827 and w15837;
w15839 <= not w15836 and not w15838;
w15840 <= not w15829 and not w15839;
w15841 <= not w7807 and not w15840;
w15842 <= not w15209 and w15216;
w15843 <= not w15218 and w15842;
w15844 <= not w15667 and w15843;
w15845 <= not w15209 and not w15218;
w15846 <= not w15667 and w15845;
w15847 <= not w15216 and not w15846;
w15848 <= not w15844 and not w15847;
w15849 <= w7807 and not w15829;
w15850 <= not w15839 and w15849;
w15851 <= not w15848 and not w15850;
w15852 <= not w15841 and not w15851;
w15853 <= not w7379 and not w15852;
w15854 <= w15228 and not w15230;
w15855 <= not w15221 and w15854;
w15856 <= not w15667 and w15855;
w15857 <= not w15221 and not w15230;
w15858 <= not w15667 and w15857;
w15859 <= not w15228 and not w15858;
w15860 <= not w15856 and not w15859;
w15861 <= w7379 and not w15841;
w15862 <= not w15851 and w15861;
w15863 <= not w15860 and not w15862;
w15864 <= not w15853 and not w15863;
w15865 <= not w6963 and not w15864;
w15866 <= not w15233 and w15240;
w15867 <= not w15242 and w15866;
w15868 <= not w15667 and w15867;
w15869 <= not w15233 and not w15242;
w15870 <= not w15667 and w15869;
w15871 <= not w15240 and not w15870;
w15872 <= not w15868 and not w15871;
w15873 <= w6963 and not w15853;
w15874 <= not w15863 and w15873;
w15875 <= not w15872 and not w15874;
w15876 <= not w15865 and not w15875;
w15877 <= not w6558 and not w15876;
w15878 <= w15252 and not w15254;
w15879 <= not w15245 and w15878;
w15880 <= not w15667 and w15879;
w15881 <= not w15245 and not w15254;
w15882 <= not w15667 and w15881;
w15883 <= not w15252 and not w15882;
w15884 <= not w15880 and not w15883;
w15885 <= w6558 and not w15865;
w15886 <= not w15875 and w15885;
w15887 <= not w15884 and not w15886;
w15888 <= not w15877 and not w15887;
w15889 <= not w6166 and not w15888;
w15890 <= not w15257 and w15264;
w15891 <= not w15266 and w15890;
w15892 <= not w15667 and w15891;
w15893 <= not w15257 and not w15266;
w15894 <= not w15667 and w15893;
w15895 <= not w15264 and not w15894;
w15896 <= not w15892 and not w15895;
w15897 <= w6166 and not w15877;
w15898 <= not w15887 and w15897;
w15899 <= not w15896 and not w15898;
w15900 <= not w15889 and not w15899;
w15901 <= not w5786 and not w15900;
w15902 <= w15276 and not w15278;
w15903 <= not w15269 and w15902;
w15904 <= not w15667 and w15903;
w15905 <= not w15269 and not w15278;
w15906 <= not w15667 and w15905;
w15907 <= not w15276 and not w15906;
w15908 <= not w15904 and not w15907;
w15909 <= w5786 and not w15889;
w15910 <= not w15899 and w15909;
w15911 <= not w15908 and not w15910;
w15912 <= not w15901 and not w15911;
w15913 <= not w5418 and not w15912;
w15914 <= not w15281 and w15288;
w15915 <= not w15290 and w15914;
w15916 <= not w15667 and w15915;
w15917 <= not w15281 and not w15290;
w15918 <= not w15667 and w15917;
w15919 <= not w15288 and not w15918;
w15920 <= not w15916 and not w15919;
w15921 <= w5418 and not w15901;
w15922 <= not w15911 and w15921;
w15923 <= not w15920 and not w15922;
w15924 <= not w15913 and not w15923;
w15925 <= not w5062 and not w15924;
w15926 <= w15300 and not w15302;
w15927 <= not w15293 and w15926;
w15928 <= not w15667 and w15927;
w15929 <= not w15293 and not w15302;
w15930 <= not w15667 and w15929;
w15931 <= not w15300 and not w15930;
w15932 <= not w15928 and not w15931;
w15933 <= w5062 and not w15913;
w15934 <= not w15923 and w15933;
w15935 <= not w15932 and not w15934;
w15936 <= not w15925 and not w15935;
w15937 <= not w4718 and not w15936;
w15938 <= not w15305 and w15312;
w15939 <= not w15314 and w15938;
w15940 <= not w15667 and w15939;
w15941 <= not w15305 and not w15314;
w15942 <= not w15667 and w15941;
w15943 <= not w15312 and not w15942;
w15944 <= not w15940 and not w15943;
w15945 <= w4718 and not w15925;
w15946 <= not w15935 and w15945;
w15947 <= not w15944 and not w15946;
w15948 <= not w15937 and not w15947;
w15949 <= not w4386 and not w15948;
w15950 <= w15324 and not w15326;
w15951 <= not w15317 and w15950;
w15952 <= not w15667 and w15951;
w15953 <= not w15317 and not w15326;
w15954 <= not w15667 and w15953;
w15955 <= not w15324 and not w15954;
w15956 <= not w15952 and not w15955;
w15957 <= w4386 and not w15937;
w15958 <= not w15947 and w15957;
w15959 <= not w15956 and not w15958;
w15960 <= not w15949 and not w15959;
w15961 <= not w4066 and not w15960;
w15962 <= not w15329 and w15336;
w15963 <= not w15338 and w15962;
w15964 <= not w15667 and w15963;
w15965 <= not w15329 and not w15338;
w15966 <= not w15667 and w15965;
w15967 <= not w15336 and not w15966;
w15968 <= not w15964 and not w15967;
w15969 <= w4066 and not w15949;
w15970 <= not w15959 and w15969;
w15971 <= not w15968 and not w15970;
w15972 <= not w15961 and not w15971;
w15973 <= not w3758 and not w15972;
w15974 <= w15348 and not w15350;
w15975 <= not w15341 and w15974;
w15976 <= not w15667 and w15975;
w15977 <= not w15341 and not w15350;
w15978 <= not w15667 and w15977;
w15979 <= not w15348 and not w15978;
w15980 <= not w15976 and not w15979;
w15981 <= w3758 and not w15961;
w15982 <= not w15971 and w15981;
w15983 <= not w15980 and not w15982;
w15984 <= not w15973 and not w15983;
w15985 <= not w3462 and not w15984;
w15986 <= not w15353 and w15360;
w15987 <= not w15362 and w15986;
w15988 <= not w15667 and w15987;
w15989 <= not w15353 and not w15362;
w15990 <= not w15667 and w15989;
w15991 <= not w15360 and not w15990;
w15992 <= not w15988 and not w15991;
w15993 <= w3462 and not w15973;
w15994 <= not w15983 and w15993;
w15995 <= not w15992 and not w15994;
w15996 <= not w15985 and not w15995;
w15997 <= not w3178 and not w15996;
w15998 <= w15372 and not w15374;
w15999 <= not w15365 and w15998;
w16000 <= not w15667 and w15999;
w16001 <= not w15365 and not w15374;
w16002 <= not w15667 and w16001;
w16003 <= not w15372 and not w16002;
w16004 <= not w16000 and not w16003;
w16005 <= w3178 and not w15985;
w16006 <= not w15995 and w16005;
w16007 <= not w16004 and not w16006;
w16008 <= not w15997 and not w16007;
w16009 <= not w2906 and not w16008;
w16010 <= not w15377 and w15384;
w16011 <= not w15386 and w16010;
w16012 <= not w15667 and w16011;
w16013 <= not w15377 and not w15386;
w16014 <= not w15667 and w16013;
w16015 <= not w15384 and not w16014;
w16016 <= not w16012 and not w16015;
w16017 <= w2906 and not w15997;
w16018 <= not w16007 and w16017;
w16019 <= not w16016 and not w16018;
w16020 <= not w16009 and not w16019;
w16021 <= not w2646 and not w16020;
w16022 <= w15396 and not w15398;
w16023 <= not w15389 and w16022;
w16024 <= not w15667 and w16023;
w16025 <= not w15389 and not w15398;
w16026 <= not w15667 and w16025;
w16027 <= not w15396 and not w16026;
w16028 <= not w16024 and not w16027;
w16029 <= w2646 and not w16009;
w16030 <= not w16019 and w16029;
w16031 <= not w16028 and not w16030;
w16032 <= not w16021 and not w16031;
w16033 <= not w2398 and not w16032;
w16034 <= not w15401 and w15408;
w16035 <= not w15410 and w16034;
w16036 <= not w15667 and w16035;
w16037 <= not w15401 and not w15410;
w16038 <= not w15667 and w16037;
w16039 <= not w15408 and not w16038;
w16040 <= not w16036 and not w16039;
w16041 <= w2398 and not w16021;
w16042 <= not w16031 and w16041;
w16043 <= not w16040 and not w16042;
w16044 <= not w16033 and not w16043;
w16045 <= not w2162 and not w16044;
w16046 <= w15420 and not w15422;
w16047 <= not w15413 and w16046;
w16048 <= not w15667 and w16047;
w16049 <= not w15413 and not w15422;
w16050 <= not w15667 and w16049;
w16051 <= not w15420 and not w16050;
w16052 <= not w16048 and not w16051;
w16053 <= w2162 and not w16033;
w16054 <= not w16043 and w16053;
w16055 <= not w16052 and not w16054;
w16056 <= not w16045 and not w16055;
w16057 <= not w1938 and not w16056;
w16058 <= not w15425 and w15432;
w16059 <= not w15434 and w16058;
w16060 <= not w15667 and w16059;
w16061 <= not w15425 and not w15434;
w16062 <= not w15667 and w16061;
w16063 <= not w15432 and not w16062;
w16064 <= not w16060 and not w16063;
w16065 <= w1938 and not w16045;
w16066 <= not w16055 and w16065;
w16067 <= not w16064 and not w16066;
w16068 <= not w16057 and not w16067;
w16069 <= not w1725 and not w16068;
w16070 <= w15444 and not w15446;
w16071 <= not w15437 and w16070;
w16072 <= not w15667 and w16071;
w16073 <= not w15437 and not w15446;
w16074 <= not w15667 and w16073;
w16075 <= not w15444 and not w16074;
w16076 <= not w16072 and not w16075;
w16077 <= w1725 and not w16057;
w16078 <= not w16067 and w16077;
w16079 <= not w16076 and not w16078;
w16080 <= not w16069 and not w16079;
w16081 <= not w1525 and not w16080;
w16082 <= not w15449 and w15456;
w16083 <= not w15458 and w16082;
w16084 <= not w15667 and w16083;
w16085 <= not w15449 and not w15458;
w16086 <= not w15667 and w16085;
w16087 <= not w15456 and not w16086;
w16088 <= not w16084 and not w16087;
w16089 <= w1525 and not w16069;
w16090 <= not w16079 and w16089;
w16091 <= not w16088 and not w16090;
w16092 <= not w16081 and not w16091;
w16093 <= not w1337 and not w16092;
w16094 <= w15468 and not w15470;
w16095 <= not w15461 and w16094;
w16096 <= not w15667 and w16095;
w16097 <= not w15461 and not w15470;
w16098 <= not w15667 and w16097;
w16099 <= not w15468 and not w16098;
w16100 <= not w16096 and not w16099;
w16101 <= w1337 and not w16081;
w16102 <= not w16091 and w16101;
w16103 <= not w16100 and not w16102;
w16104 <= not w16093 and not w16103;
w16105 <= not w1161 and not w16104;
w16106 <= not w15473 and w15480;
w16107 <= not w15482 and w16106;
w16108 <= not w15667 and w16107;
w16109 <= not w15473 and not w15482;
w16110 <= not w15667 and w16109;
w16111 <= not w15480 and not w16110;
w16112 <= not w16108 and not w16111;
w16113 <= w1161 and not w16093;
w16114 <= not w16103 and w16113;
w16115 <= not w16112 and not w16114;
w16116 <= not w16105 and not w16115;
w16117 <= not w997 and not w16116;
w16118 <= w15492 and not w15494;
w16119 <= not w15485 and w16118;
w16120 <= not w15667 and w16119;
w16121 <= not w15485 and not w15494;
w16122 <= not w15667 and w16121;
w16123 <= not w15492 and not w16122;
w16124 <= not w16120 and not w16123;
w16125 <= w997 and not w16105;
w16126 <= not w16115 and w16125;
w16127 <= not w16124 and not w16126;
w16128 <= not w16117 and not w16127;
w16129 <= not w845 and not w16128;
w16130 <= w845 and not w16117;
w16131 <= not w16127 and w16130;
w16132 <= not w15497 and w15506;
w16133 <= not w15499 and w16132;
w16134 <= not w15667 and w16133;
w16135 <= not w15497 and not w15499;
w16136 <= not w15667 and w16135;
w16137 <= not w15506 and not w16136;
w16138 <= not w16134 and not w16137;
w16139 <= not w16131 and not w16138;
w16140 <= not w16129 and not w16139;
w16141 <= not w705 and not w16140;
w16142 <= w15516 and not w15518;
w16143 <= not w15509 and w16142;
w16144 <= not w15667 and w16143;
w16145 <= not w15509 and not w15518;
w16146 <= not w15667 and w16145;
w16147 <= not w15516 and not w16146;
w16148 <= not w16144 and not w16147;
w16149 <= w705 and not w16129;
w16150 <= not w16139 and w16149;
w16151 <= not w16148 and not w16150;
w16152 <= not w16141 and not w16151;
w16153 <= not w577 and not w16152;
w16154 <= not w15521 and w15528;
w16155 <= not w15530 and w16154;
w16156 <= not w15667 and w16155;
w16157 <= not w15521 and not w15530;
w16158 <= not w15667 and w16157;
w16159 <= not w15528 and not w16158;
w16160 <= not w16156 and not w16159;
w16161 <= w577 and not w16141;
w16162 <= not w16151 and w16161;
w16163 <= not w16160 and not w16162;
w16164 <= not w16153 and not w16163;
w16165 <= not w460 and not w16164;
w16166 <= w15540 and not w15542;
w16167 <= not w15533 and w16166;
w16168 <= not w15667 and w16167;
w16169 <= not w15533 and not w15542;
w16170 <= not w15667 and w16169;
w16171 <= not w15540 and not w16170;
w16172 <= not w16168 and not w16171;
w16173 <= w460 and not w16153;
w16174 <= not w16163 and w16173;
w16175 <= not w16172 and not w16174;
w16176 <= not w16165 and not w16175;
w16177 <= not w356 and not w16176;
w16178 <= not w15545 and w15552;
w16179 <= not w15554 and w16178;
w16180 <= not w15667 and w16179;
w16181 <= not w15545 and not w15554;
w16182 <= not w15667 and w16181;
w16183 <= not w15552 and not w16182;
w16184 <= not w16180 and not w16183;
w16185 <= w356 and not w16165;
w16186 <= not w16175 and w16185;
w16187 <= not w16184 and not w16186;
w16188 <= not w16177 and not w16187;
w16189 <= not w264 and not w16188;
w16190 <= w15564 and not w15566;
w16191 <= not w15557 and w16190;
w16192 <= not w15667 and w16191;
w16193 <= not w15557 and not w15566;
w16194 <= not w15667 and w16193;
w16195 <= not w15564 and not w16194;
w16196 <= not w16192 and not w16195;
w16197 <= w264 and not w16177;
w16198 <= not w16187 and w16197;
w16199 <= not w16196 and not w16198;
w16200 <= not w16189 and not w16199;
w16201 <= not w184 and not w16200;
w16202 <= not w15569 and w15576;
w16203 <= not w15578 and w16202;
w16204 <= not w15667 and w16203;
w16205 <= not w15569 and not w15578;
w16206 <= not w15667 and w16205;
w16207 <= not w15576 and not w16206;
w16208 <= not w16204 and not w16207;
w16209 <= w184 and not w16189;
w16210 <= not w16199 and w16209;
w16211 <= not w16208 and not w16210;
w16212 <= not w16201 and not w16211;
w16213 <= not w115 and not w16212;
w16214 <= w15588 and not w15590;
w16215 <= not w15581 and w16214;
w16216 <= not w15667 and w16215;
w16217 <= not w15581 and not w15590;
w16218 <= not w15667 and w16217;
w16219 <= not w15588 and not w16218;
w16220 <= not w16216 and not w16219;
w16221 <= w115 and not w16201;
w16222 <= not w16211 and w16221;
w16223 <= not w16220 and not w16222;
w16224 <= not w16213 and not w16223;
w16225 <= not w60 and not w16224;
w16226 <= not w15593 and w15600;
w16227 <= not w15602 and w16226;
w16228 <= not w15667 and w16227;
w16229 <= not w15593 and not w15602;
w16230 <= not w15667 and w16229;
w16231 <= not w15600 and not w16230;
w16232 <= not w16228 and not w16231;
w16233 <= w60 and not w16213;
w16234 <= not w16223 and w16233;
w16235 <= not w16232 and not w16234;
w16236 <= not w16225 and not w16235;
w16237 <= not w22 and not w16236;
w16238 <= w15612 and not w15614;
w16239 <= not w15605 and w16238;
w16240 <= not w15667 and w16239;
w16241 <= not w15605 and not w15614;
w16242 <= not w15667 and w16241;
w16243 <= not w15612 and not w16242;
w16244 <= not w16240 and not w16243;
w16245 <= w22 and not w16225;
w16246 <= not w16235 and w16245;
w16247 <= not w16244 and not w16246;
w16248 <= not w16237 and not w16247;
w16249 <= not w5 and not w16248;
w16250 <= not w15617 and w15624;
w16251 <= not w15626 and w16250;
w16252 <= not w15667 and w16251;
w16253 <= not w15617 and not w15626;
w16254 <= not w15667 and w16253;
w16255 <= not w15624 and not w16254;
w16256 <= not w16252 and not w16255;
w16257 <= w5 and not w16237;
w16258 <= not w16247 and w16257;
w16259 <= not w16256 and not w16258;
w16260 <= not w16249 and not w16259;
w16261 <= w15636 and not w15638;
w16262 <= not w15629 and w16261;
w16263 <= not w15667 and w16262;
w16264 <= not w15629 and not w15638;
w16265 <= not w15667 and w16264;
w16266 <= not w15636 and not w16265;
w16267 <= not w16263 and not w16266;
w16268 <= not w15640 and not w15647;
w16269 <= not w15667 and w16268;
w16270 <= not w15655 and not w16269;
w16271 <= not w16267 and w16270;
w16272 <= not w16260 and w16271;
w16273 <= w0 and not w16272;
w16274 <= not w16249 and w16267;
w16275 <= not w16259 and w16274;
w16276 <= not w15647 and not w15667;
w16277 <= w15640 and not w16276;
w16278 <= not w0 and not w16268;
w16279 <= not w16277 and w16278;
w16280 <= not w15643 and not w15664;
w16281 <= not w15646 and w16280;
w16282 <= not w15659 and w16281;
w16283 <= not w15655 and w16282;
w16284 <= not w15653 and w16283;
w16285 <= not w16279 and not w16284;
w16286 <= not w16275 and w16285;
w16287 <= not w16273 and w16286;
w16288 <= a(24) and not w16287;
w16289 <= not a(22) and not a(23);
w16290 <= not a(24) and w16289;
w16291 <= not w16288 and not w16290;
w16292 <= not w15667 and not w16291;
w16293 <= not w15664 and not w16290;
w16294 <= not w15659 and w16293;
w16295 <= not w15655 and w16294;
w16296 <= not w15653 and w16295;
w16297 <= not w16288 and w16296;
w16298 <= not a(24) and not w16287;
w16299 <= a(25) and not w16298;
w16300 <= w15669 and not w16287;
w16301 <= not w16299 and not w16300;
w16302 <= not w16297 and w16301;
w16303 <= not w16292 and not w16302;
w16304 <= not w15059 and not w16303;
w16305 <= w15059 and not w16292;
w16306 <= not w16302 and w16305;
w16307 <= not w15667 and not w16284;
w16308 <= not w16279 and w16307;
w16309 <= not w16275 and w16308;
w16310 <= not w16273 and w16309;
w16311 <= not w16300 and not w16310;
w16312 <= a(26) and not w16311;
w16313 <= not a(26) and not w16310;
w16314 <= not w16300 and w16313;
w16315 <= not w16312 and not w16314;
w16316 <= not w16306 and not w16315;
w16317 <= not w16304 and not w16316;
w16318 <= not w14463 and not w16317;
w16319 <= not w15672 and not w15677;
w16320 <= not w15681 and w16319;
w16321 <= not w16287 and w16320;
w16322 <= not w16287 and w16319;
w16323 <= w15681 and not w16322;
w16324 <= not w16321 and not w16323;
w16325 <= w14463 and not w16304;
w16326 <= not w16316 and w16325;
w16327 <= not w16324 and not w16326;
w16328 <= not w16318 and not w16327;
w16329 <= not w13879 and not w16328;
w16330 <= not w15686 and w15695;
w16331 <= not w15684 and w16330;
w16332 <= not w16287 and w16331;
w16333 <= not w15684 and not w15686;
w16334 <= not w16287 and w16333;
w16335 <= not w15695 and not w16334;
w16336 <= not w16332 and not w16335;
w16337 <= w13879 and not w16318;
w16338 <= not w16327 and w16337;
w16339 <= not w16336 and not w16338;
w16340 <= not w16329 and not w16339;
w16341 <= not w13307 and not w16340;
w16342 <= not w15698 and w15704;
w16343 <= not w15706 and w16342;
w16344 <= not w16287 and w16343;
w16345 <= not w15698 and not w15706;
w16346 <= not w16287 and w16345;
w16347 <= not w15704 and not w16346;
w16348 <= not w16344 and not w16347;
w16349 <= w13307 and not w16329;
w16350 <= not w16339 and w16349;
w16351 <= not w16348 and not w16350;
w16352 <= not w16341 and not w16351;
w16353 <= not w12747 and not w16352;
w16354 <= w15716 and not w15718;
w16355 <= not w15709 and w16354;
w16356 <= not w16287 and w16355;
w16357 <= not w15709 and not w15718;
w16358 <= not w16287 and w16357;
w16359 <= not w15716 and not w16358;
w16360 <= not w16356 and not w16359;
w16361 <= w12747 and not w16341;
w16362 <= not w16351 and w16361;
w16363 <= not w16360 and not w16362;
w16364 <= not w16353 and not w16363;
w16365 <= not w12199 and not w16364;
w16366 <= not w15721 and w15728;
w16367 <= not w15730 and w16366;
w16368 <= not w16287 and w16367;
w16369 <= not w15721 and not w15730;
w16370 <= not w16287 and w16369;
w16371 <= not w15728 and not w16370;
w16372 <= not w16368 and not w16371;
w16373 <= w12199 and not w16353;
w16374 <= not w16363 and w16373;
w16375 <= not w16372 and not w16374;
w16376 <= not w16365 and not w16375;
w16377 <= not w11663 and not w16376;
w16378 <= w15740 and not w15742;
w16379 <= not w15733 and w16378;
w16380 <= not w16287 and w16379;
w16381 <= not w15733 and not w15742;
w16382 <= not w16287 and w16381;
w16383 <= not w15740 and not w16382;
w16384 <= not w16380 and not w16383;
w16385 <= w11663 and not w16365;
w16386 <= not w16375 and w16385;
w16387 <= not w16384 and not w16386;
w16388 <= not w16377 and not w16387;
w16389 <= not w11139 and not w16388;
w16390 <= not w15745 and w15752;
w16391 <= not w15754 and w16390;
w16392 <= not w16287 and w16391;
w16393 <= not w15745 and not w15754;
w16394 <= not w16287 and w16393;
w16395 <= not w15752 and not w16394;
w16396 <= not w16392 and not w16395;
w16397 <= w11139 and not w16377;
w16398 <= not w16387 and w16397;
w16399 <= not w16396 and not w16398;
w16400 <= not w16389 and not w16399;
w16401 <= not w10627 and not w16400;
w16402 <= w15764 and not w15766;
w16403 <= not w15757 and w16402;
w16404 <= not w16287 and w16403;
w16405 <= not w15757 and not w15766;
w16406 <= not w16287 and w16405;
w16407 <= not w15764 and not w16406;
w16408 <= not w16404 and not w16407;
w16409 <= w10627 and not w16389;
w16410 <= not w16399 and w16409;
w16411 <= not w16408 and not w16410;
w16412 <= not w16401 and not w16411;
w16413 <= not w10127 and not w16412;
w16414 <= not w15769 and w15776;
w16415 <= not w15778 and w16414;
w16416 <= not w16287 and w16415;
w16417 <= not w15769 and not w15778;
w16418 <= not w16287 and w16417;
w16419 <= not w15776 and not w16418;
w16420 <= not w16416 and not w16419;
w16421 <= w10127 and not w16401;
w16422 <= not w16411 and w16421;
w16423 <= not w16420 and not w16422;
w16424 <= not w16413 and not w16423;
w16425 <= not w9639 and not w16424;
w16426 <= w15788 and not w15790;
w16427 <= not w15781 and w16426;
w16428 <= not w16287 and w16427;
w16429 <= not w15781 and not w15790;
w16430 <= not w16287 and w16429;
w16431 <= not w15788 and not w16430;
w16432 <= not w16428 and not w16431;
w16433 <= w9639 and not w16413;
w16434 <= not w16423 and w16433;
w16435 <= not w16432 and not w16434;
w16436 <= not w16425 and not w16435;
w16437 <= not w9163 and not w16436;
w16438 <= not w15793 and w15800;
w16439 <= not w15802 and w16438;
w16440 <= not w16287 and w16439;
w16441 <= not w15793 and not w15802;
w16442 <= not w16287 and w16441;
w16443 <= not w15800 and not w16442;
w16444 <= not w16440 and not w16443;
w16445 <= w9163 and not w16425;
w16446 <= not w16435 and w16445;
w16447 <= not w16444 and not w16446;
w16448 <= not w16437 and not w16447;
w16449 <= not w8699 and not w16448;
w16450 <= w15812 and not w15814;
w16451 <= not w15805 and w16450;
w16452 <= not w16287 and w16451;
w16453 <= not w15805 and not w15814;
w16454 <= not w16287 and w16453;
w16455 <= not w15812 and not w16454;
w16456 <= not w16452 and not w16455;
w16457 <= w8699 and not w16437;
w16458 <= not w16447 and w16457;
w16459 <= not w16456 and not w16458;
w16460 <= not w16449 and not w16459;
w16461 <= not w8247 and not w16460;
w16462 <= not w15817 and w15824;
w16463 <= not w15826 and w16462;
w16464 <= not w16287 and w16463;
w16465 <= not w15817 and not w15826;
w16466 <= not w16287 and w16465;
w16467 <= not w15824 and not w16466;
w16468 <= not w16464 and not w16467;
w16469 <= w8247 and not w16449;
w16470 <= not w16459 and w16469;
w16471 <= not w16468 and not w16470;
w16472 <= not w16461 and not w16471;
w16473 <= not w7807 and not w16472;
w16474 <= w15836 and not w15838;
w16475 <= not w15829 and w16474;
w16476 <= not w16287 and w16475;
w16477 <= not w15829 and not w15838;
w16478 <= not w16287 and w16477;
w16479 <= not w15836 and not w16478;
w16480 <= not w16476 and not w16479;
w16481 <= w7807 and not w16461;
w16482 <= not w16471 and w16481;
w16483 <= not w16480 and not w16482;
w16484 <= not w16473 and not w16483;
w16485 <= not w7379 and not w16484;
w16486 <= not w15841 and w15848;
w16487 <= not w15850 and w16486;
w16488 <= not w16287 and w16487;
w16489 <= not w15841 and not w15850;
w16490 <= not w16287 and w16489;
w16491 <= not w15848 and not w16490;
w16492 <= not w16488 and not w16491;
w16493 <= w7379 and not w16473;
w16494 <= not w16483 and w16493;
w16495 <= not w16492 and not w16494;
w16496 <= not w16485 and not w16495;
w16497 <= not w6963 and not w16496;
w16498 <= w15860 and not w15862;
w16499 <= not w15853 and w16498;
w16500 <= not w16287 and w16499;
w16501 <= not w15853 and not w15862;
w16502 <= not w16287 and w16501;
w16503 <= not w15860 and not w16502;
w16504 <= not w16500 and not w16503;
w16505 <= w6963 and not w16485;
w16506 <= not w16495 and w16505;
w16507 <= not w16504 and not w16506;
w16508 <= not w16497 and not w16507;
w16509 <= not w6558 and not w16508;
w16510 <= not w15865 and w15872;
w16511 <= not w15874 and w16510;
w16512 <= not w16287 and w16511;
w16513 <= not w15865 and not w15874;
w16514 <= not w16287 and w16513;
w16515 <= not w15872 and not w16514;
w16516 <= not w16512 and not w16515;
w16517 <= w6558 and not w16497;
w16518 <= not w16507 and w16517;
w16519 <= not w16516 and not w16518;
w16520 <= not w16509 and not w16519;
w16521 <= not w6166 and not w16520;
w16522 <= w15884 and not w15886;
w16523 <= not w15877 and w16522;
w16524 <= not w16287 and w16523;
w16525 <= not w15877 and not w15886;
w16526 <= not w16287 and w16525;
w16527 <= not w15884 and not w16526;
w16528 <= not w16524 and not w16527;
w16529 <= w6166 and not w16509;
w16530 <= not w16519 and w16529;
w16531 <= not w16528 and not w16530;
w16532 <= not w16521 and not w16531;
w16533 <= not w5786 and not w16532;
w16534 <= not w15889 and w15896;
w16535 <= not w15898 and w16534;
w16536 <= not w16287 and w16535;
w16537 <= not w15889 and not w15898;
w16538 <= not w16287 and w16537;
w16539 <= not w15896 and not w16538;
w16540 <= not w16536 and not w16539;
w16541 <= w5786 and not w16521;
w16542 <= not w16531 and w16541;
w16543 <= not w16540 and not w16542;
w16544 <= not w16533 and not w16543;
w16545 <= not w5418 and not w16544;
w16546 <= w15908 and not w15910;
w16547 <= not w15901 and w16546;
w16548 <= not w16287 and w16547;
w16549 <= not w15901 and not w15910;
w16550 <= not w16287 and w16549;
w16551 <= not w15908 and not w16550;
w16552 <= not w16548 and not w16551;
w16553 <= w5418 and not w16533;
w16554 <= not w16543 and w16553;
w16555 <= not w16552 and not w16554;
w16556 <= not w16545 and not w16555;
w16557 <= not w5062 and not w16556;
w16558 <= not w15913 and w15920;
w16559 <= not w15922 and w16558;
w16560 <= not w16287 and w16559;
w16561 <= not w15913 and not w15922;
w16562 <= not w16287 and w16561;
w16563 <= not w15920 and not w16562;
w16564 <= not w16560 and not w16563;
w16565 <= w5062 and not w16545;
w16566 <= not w16555 and w16565;
w16567 <= not w16564 and not w16566;
w16568 <= not w16557 and not w16567;
w16569 <= not w4718 and not w16568;
w16570 <= w15932 and not w15934;
w16571 <= not w15925 and w16570;
w16572 <= not w16287 and w16571;
w16573 <= not w15925 and not w15934;
w16574 <= not w16287 and w16573;
w16575 <= not w15932 and not w16574;
w16576 <= not w16572 and not w16575;
w16577 <= w4718 and not w16557;
w16578 <= not w16567 and w16577;
w16579 <= not w16576 and not w16578;
w16580 <= not w16569 and not w16579;
w16581 <= not w4386 and not w16580;
w16582 <= not w15937 and w15944;
w16583 <= not w15946 and w16582;
w16584 <= not w16287 and w16583;
w16585 <= not w15937 and not w15946;
w16586 <= not w16287 and w16585;
w16587 <= not w15944 and not w16586;
w16588 <= not w16584 and not w16587;
w16589 <= w4386 and not w16569;
w16590 <= not w16579 and w16589;
w16591 <= not w16588 and not w16590;
w16592 <= not w16581 and not w16591;
w16593 <= not w4066 and not w16592;
w16594 <= w15956 and not w15958;
w16595 <= not w15949 and w16594;
w16596 <= not w16287 and w16595;
w16597 <= not w15949 and not w15958;
w16598 <= not w16287 and w16597;
w16599 <= not w15956 and not w16598;
w16600 <= not w16596 and not w16599;
w16601 <= w4066 and not w16581;
w16602 <= not w16591 and w16601;
w16603 <= not w16600 and not w16602;
w16604 <= not w16593 and not w16603;
w16605 <= not w3758 and not w16604;
w16606 <= not w15961 and w15968;
w16607 <= not w15970 and w16606;
w16608 <= not w16287 and w16607;
w16609 <= not w15961 and not w15970;
w16610 <= not w16287 and w16609;
w16611 <= not w15968 and not w16610;
w16612 <= not w16608 and not w16611;
w16613 <= w3758 and not w16593;
w16614 <= not w16603 and w16613;
w16615 <= not w16612 and not w16614;
w16616 <= not w16605 and not w16615;
w16617 <= not w3462 and not w16616;
w16618 <= w15980 and not w15982;
w16619 <= not w15973 and w16618;
w16620 <= not w16287 and w16619;
w16621 <= not w15973 and not w15982;
w16622 <= not w16287 and w16621;
w16623 <= not w15980 and not w16622;
w16624 <= not w16620 and not w16623;
w16625 <= w3462 and not w16605;
w16626 <= not w16615 and w16625;
w16627 <= not w16624 and not w16626;
w16628 <= not w16617 and not w16627;
w16629 <= not w3178 and not w16628;
w16630 <= not w15985 and w15992;
w16631 <= not w15994 and w16630;
w16632 <= not w16287 and w16631;
w16633 <= not w15985 and not w15994;
w16634 <= not w16287 and w16633;
w16635 <= not w15992 and not w16634;
w16636 <= not w16632 and not w16635;
w16637 <= w3178 and not w16617;
w16638 <= not w16627 and w16637;
w16639 <= not w16636 and not w16638;
w16640 <= not w16629 and not w16639;
w16641 <= not w2906 and not w16640;
w16642 <= w16004 and not w16006;
w16643 <= not w15997 and w16642;
w16644 <= not w16287 and w16643;
w16645 <= not w15997 and not w16006;
w16646 <= not w16287 and w16645;
w16647 <= not w16004 and not w16646;
w16648 <= not w16644 and not w16647;
w16649 <= w2906 and not w16629;
w16650 <= not w16639 and w16649;
w16651 <= not w16648 and not w16650;
w16652 <= not w16641 and not w16651;
w16653 <= not w2646 and not w16652;
w16654 <= not w16009 and w16016;
w16655 <= not w16018 and w16654;
w16656 <= not w16287 and w16655;
w16657 <= not w16009 and not w16018;
w16658 <= not w16287 and w16657;
w16659 <= not w16016 and not w16658;
w16660 <= not w16656 and not w16659;
w16661 <= w2646 and not w16641;
w16662 <= not w16651 and w16661;
w16663 <= not w16660 and not w16662;
w16664 <= not w16653 and not w16663;
w16665 <= not w2398 and not w16664;
w16666 <= w16028 and not w16030;
w16667 <= not w16021 and w16666;
w16668 <= not w16287 and w16667;
w16669 <= not w16021 and not w16030;
w16670 <= not w16287 and w16669;
w16671 <= not w16028 and not w16670;
w16672 <= not w16668 and not w16671;
w16673 <= w2398 and not w16653;
w16674 <= not w16663 and w16673;
w16675 <= not w16672 and not w16674;
w16676 <= not w16665 and not w16675;
w16677 <= not w2162 and not w16676;
w16678 <= not w16033 and w16040;
w16679 <= not w16042 and w16678;
w16680 <= not w16287 and w16679;
w16681 <= not w16033 and not w16042;
w16682 <= not w16287 and w16681;
w16683 <= not w16040 and not w16682;
w16684 <= not w16680 and not w16683;
w16685 <= w2162 and not w16665;
w16686 <= not w16675 and w16685;
w16687 <= not w16684 and not w16686;
w16688 <= not w16677 and not w16687;
w16689 <= not w1938 and not w16688;
w16690 <= w16052 and not w16054;
w16691 <= not w16045 and w16690;
w16692 <= not w16287 and w16691;
w16693 <= not w16045 and not w16054;
w16694 <= not w16287 and w16693;
w16695 <= not w16052 and not w16694;
w16696 <= not w16692 and not w16695;
w16697 <= w1938 and not w16677;
w16698 <= not w16687 and w16697;
w16699 <= not w16696 and not w16698;
w16700 <= not w16689 and not w16699;
w16701 <= not w1725 and not w16700;
w16702 <= not w16057 and w16064;
w16703 <= not w16066 and w16702;
w16704 <= not w16287 and w16703;
w16705 <= not w16057 and not w16066;
w16706 <= not w16287 and w16705;
w16707 <= not w16064 and not w16706;
w16708 <= not w16704 and not w16707;
w16709 <= w1725 and not w16689;
w16710 <= not w16699 and w16709;
w16711 <= not w16708 and not w16710;
w16712 <= not w16701 and not w16711;
w16713 <= not w1525 and not w16712;
w16714 <= w16076 and not w16078;
w16715 <= not w16069 and w16714;
w16716 <= not w16287 and w16715;
w16717 <= not w16069 and not w16078;
w16718 <= not w16287 and w16717;
w16719 <= not w16076 and not w16718;
w16720 <= not w16716 and not w16719;
w16721 <= w1525 and not w16701;
w16722 <= not w16711 and w16721;
w16723 <= not w16720 and not w16722;
w16724 <= not w16713 and not w16723;
w16725 <= not w1337 and not w16724;
w16726 <= not w16081 and w16088;
w16727 <= not w16090 and w16726;
w16728 <= not w16287 and w16727;
w16729 <= not w16081 and not w16090;
w16730 <= not w16287 and w16729;
w16731 <= not w16088 and not w16730;
w16732 <= not w16728 and not w16731;
w16733 <= w1337 and not w16713;
w16734 <= not w16723 and w16733;
w16735 <= not w16732 and not w16734;
w16736 <= not w16725 and not w16735;
w16737 <= not w1161 and not w16736;
w16738 <= w16100 and not w16102;
w16739 <= not w16093 and w16738;
w16740 <= not w16287 and w16739;
w16741 <= not w16093 and not w16102;
w16742 <= not w16287 and w16741;
w16743 <= not w16100 and not w16742;
w16744 <= not w16740 and not w16743;
w16745 <= w1161 and not w16725;
w16746 <= not w16735 and w16745;
w16747 <= not w16744 and not w16746;
w16748 <= not w16737 and not w16747;
w16749 <= not w997 and not w16748;
w16750 <= not w16105 and w16112;
w16751 <= not w16114 and w16750;
w16752 <= not w16287 and w16751;
w16753 <= not w16105 and not w16114;
w16754 <= not w16287 and w16753;
w16755 <= not w16112 and not w16754;
w16756 <= not w16752 and not w16755;
w16757 <= w997 and not w16737;
w16758 <= not w16747 and w16757;
w16759 <= not w16756 and not w16758;
w16760 <= not w16749 and not w16759;
w16761 <= not w845 and not w16760;
w16762 <= w16124 and not w16126;
w16763 <= not w16117 and w16762;
w16764 <= not w16287 and w16763;
w16765 <= not w16117 and not w16126;
w16766 <= not w16287 and w16765;
w16767 <= not w16124 and not w16766;
w16768 <= not w16764 and not w16767;
w16769 <= w845 and not w16749;
w16770 <= not w16759 and w16769;
w16771 <= not w16768 and not w16770;
w16772 <= not w16761 and not w16771;
w16773 <= not w705 and not w16772;
w16774 <= w705 and not w16761;
w16775 <= not w16771 and w16774;
w16776 <= not w16129 and w16138;
w16777 <= not w16131 and w16776;
w16778 <= not w16287 and w16777;
w16779 <= not w16129 and not w16131;
w16780 <= not w16287 and w16779;
w16781 <= not w16138 and not w16780;
w16782 <= not w16778 and not w16781;
w16783 <= not w16775 and not w16782;
w16784 <= not w16773 and not w16783;
w16785 <= not w577 and not w16784;
w16786 <= w16148 and not w16150;
w16787 <= not w16141 and w16786;
w16788 <= not w16287 and w16787;
w16789 <= not w16141 and not w16150;
w16790 <= not w16287 and w16789;
w16791 <= not w16148 and not w16790;
w16792 <= not w16788 and not w16791;
w16793 <= w577 and not w16773;
w16794 <= not w16783 and w16793;
w16795 <= not w16792 and not w16794;
w16796 <= not w16785 and not w16795;
w16797 <= not w460 and not w16796;
w16798 <= not w16153 and w16160;
w16799 <= not w16162 and w16798;
w16800 <= not w16287 and w16799;
w16801 <= not w16153 and not w16162;
w16802 <= not w16287 and w16801;
w16803 <= not w16160 and not w16802;
w16804 <= not w16800 and not w16803;
w16805 <= w460 and not w16785;
w16806 <= not w16795 and w16805;
w16807 <= not w16804 and not w16806;
w16808 <= not w16797 and not w16807;
w16809 <= not w356 and not w16808;
w16810 <= w16172 and not w16174;
w16811 <= not w16165 and w16810;
w16812 <= not w16287 and w16811;
w16813 <= not w16165 and not w16174;
w16814 <= not w16287 and w16813;
w16815 <= not w16172 and not w16814;
w16816 <= not w16812 and not w16815;
w16817 <= w356 and not w16797;
w16818 <= not w16807 and w16817;
w16819 <= not w16816 and not w16818;
w16820 <= not w16809 and not w16819;
w16821 <= not w264 and not w16820;
w16822 <= not w16177 and w16184;
w16823 <= not w16186 and w16822;
w16824 <= not w16287 and w16823;
w16825 <= not w16177 and not w16186;
w16826 <= not w16287 and w16825;
w16827 <= not w16184 and not w16826;
w16828 <= not w16824 and not w16827;
w16829 <= w264 and not w16809;
w16830 <= not w16819 and w16829;
w16831 <= not w16828 and not w16830;
w16832 <= not w16821 and not w16831;
w16833 <= not w184 and not w16832;
w16834 <= w16196 and not w16198;
w16835 <= not w16189 and w16834;
w16836 <= not w16287 and w16835;
w16837 <= not w16189 and not w16198;
w16838 <= not w16287 and w16837;
w16839 <= not w16196 and not w16838;
w16840 <= not w16836 and not w16839;
w16841 <= w184 and not w16821;
w16842 <= not w16831 and w16841;
w16843 <= not w16840 and not w16842;
w16844 <= not w16833 and not w16843;
w16845 <= not w115 and not w16844;
w16846 <= not w16201 and w16208;
w16847 <= not w16210 and w16846;
w16848 <= not w16287 and w16847;
w16849 <= not w16201 and not w16210;
w16850 <= not w16287 and w16849;
w16851 <= not w16208 and not w16850;
w16852 <= not w16848 and not w16851;
w16853 <= w115 and not w16833;
w16854 <= not w16843 and w16853;
w16855 <= not w16852 and not w16854;
w16856 <= not w16845 and not w16855;
w16857 <= not w60 and not w16856;
w16858 <= w16220 and not w16222;
w16859 <= not w16213 and w16858;
w16860 <= not w16287 and w16859;
w16861 <= not w16213 and not w16222;
w16862 <= not w16287 and w16861;
w16863 <= not w16220 and not w16862;
w16864 <= not w16860 and not w16863;
w16865 <= w60 and not w16845;
w16866 <= not w16855 and w16865;
w16867 <= not w16864 and not w16866;
w16868 <= not w16857 and not w16867;
w16869 <= not w22 and not w16868;
w16870 <= not w16225 and w16232;
w16871 <= not w16234 and w16870;
w16872 <= not w16287 and w16871;
w16873 <= not w16225 and not w16234;
w16874 <= not w16287 and w16873;
w16875 <= not w16232 and not w16874;
w16876 <= not w16872 and not w16875;
w16877 <= w22 and not w16857;
w16878 <= not w16867 and w16877;
w16879 <= not w16876 and not w16878;
w16880 <= not w16869 and not w16879;
w16881 <= not w5 and not w16880;
w16882 <= w16244 and not w16246;
w16883 <= not w16237 and w16882;
w16884 <= not w16287 and w16883;
w16885 <= not w16237 and not w16246;
w16886 <= not w16287 and w16885;
w16887 <= not w16244 and not w16886;
w16888 <= not w16884 and not w16887;
w16889 <= w5 and not w16869;
w16890 <= not w16879 and w16889;
w16891 <= not w16888 and not w16890;
w16892 <= not w16881 and not w16891;
w16893 <= not w16249 and w16256;
w16894 <= not w16258 and w16893;
w16895 <= not w16287 and w16894;
w16896 <= not w16249 and not w16258;
w16897 <= not w16287 and w16896;
w16898 <= not w16256 and not w16897;
w16899 <= not w16895 and not w16898;
w16900 <= not w16260 and not w16267;
w16901 <= not w16287 and w16900;
w16902 <= not w16275 and not w16901;
w16903 <= not w16899 and w16902;
w16904 <= not w16892 and w16903;
w16905 <= w0 and not w16904;
w16906 <= not w16881 and w16899;
w16907 <= not w16891 and w16906;
w16908 <= not w16267 and not w16287;
w16909 <= w16260 and not w16908;
w16910 <= not w0 and not w16900;
w16911 <= not w16909 and w16910;
w16912 <= not w16263 and not w16284;
w16913 <= not w16266 and w16912;
w16914 <= not w16279 and w16913;
w16915 <= not w16275 and w16914;
w16916 <= not w16273 and w16915;
w16917 <= not w16911 and not w16916;
w16918 <= not w16907 and w16917;
w16919 <= not w16905 and w16918;
w16920 <= a(22) and not w16919;
w16921 <= not a(20) and not a(21);
w16922 <= not a(22) and w16921;
w16923 <= not w16920 and not w16922;
w16924 <= not w16287 and not w16923;
w16925 <= not w16284 and not w16922;
w16926 <= not w16279 and w16925;
w16927 <= not w16275 and w16926;
w16928 <= not w16273 and w16927;
w16929 <= not w16920 and w16928;
w16930 <= not a(22) and not w16919;
w16931 <= a(23) and not w16930;
w16932 <= w16289 and not w16919;
w16933 <= not w16931 and not w16932;
w16934 <= not w16929 and w16933;
w16935 <= not w16924 and not w16934;
w16936 <= not w15667 and not w16935;
w16937 <= w15667 and not w16924;
w16938 <= not w16934 and w16937;
w16939 <= not w16287 and not w16916;
w16940 <= not w16911 and w16939;
w16941 <= not w16907 and w16940;
w16942 <= not w16905 and w16941;
w16943 <= not w16932 and not w16942;
w16944 <= a(24) and not w16943;
w16945 <= not a(24) and not w16942;
w16946 <= not w16932 and w16945;
w16947 <= not w16944 and not w16946;
w16948 <= not w16938 and not w16947;
w16949 <= not w16936 and not w16948;
w16950 <= not w15059 and not w16949;
w16951 <= not w16292 and not w16297;
w16952 <= not w16301 and w16951;
w16953 <= not w16919 and w16952;
w16954 <= not w16919 and w16951;
w16955 <= w16301 and not w16954;
w16956 <= not w16953 and not w16955;
w16957 <= w15059 and not w16936;
w16958 <= not w16948 and w16957;
w16959 <= not w16956 and not w16958;
w16960 <= not w16950 and not w16959;
w16961 <= not w14463 and not w16960;
w16962 <= not w16306 and w16315;
w16963 <= not w16304 and w16962;
w16964 <= not w16919 and w16963;
w16965 <= not w16304 and not w16306;
w16966 <= not w16919 and w16965;
w16967 <= not w16315 and not w16966;
w16968 <= not w16964 and not w16967;
w16969 <= w14463 and not w16950;
w16970 <= not w16959 and w16969;
w16971 <= not w16968 and not w16970;
w16972 <= not w16961 and not w16971;
w16973 <= not w13879 and not w16972;
w16974 <= not w16318 and w16324;
w16975 <= not w16326 and w16974;
w16976 <= not w16919 and w16975;
w16977 <= not w16318 and not w16326;
w16978 <= not w16919 and w16977;
w16979 <= not w16324 and not w16978;
w16980 <= not w16976 and not w16979;
w16981 <= w13879 and not w16961;
w16982 <= not w16971 and w16981;
w16983 <= not w16980 and not w16982;
w16984 <= not w16973 and not w16983;
w16985 <= not w13307 and not w16984;
w16986 <= w16336 and not w16338;
w16987 <= not w16329 and w16986;
w16988 <= not w16919 and w16987;
w16989 <= not w16329 and not w16338;
w16990 <= not w16919 and w16989;
w16991 <= not w16336 and not w16990;
w16992 <= not w16988 and not w16991;
w16993 <= w13307 and not w16973;
w16994 <= not w16983 and w16993;
w16995 <= not w16992 and not w16994;
w16996 <= not w16985 and not w16995;
w16997 <= not w12747 and not w16996;
w16998 <= not w16341 and w16348;
w16999 <= not w16350 and w16998;
w17000 <= not w16919 and w16999;
w17001 <= not w16341 and not w16350;
w17002 <= not w16919 and w17001;
w17003 <= not w16348 and not w17002;
w17004 <= not w17000 and not w17003;
w17005 <= w12747 and not w16985;
w17006 <= not w16995 and w17005;
w17007 <= not w17004 and not w17006;
w17008 <= not w16997 and not w17007;
w17009 <= not w12199 and not w17008;
w17010 <= w16360 and not w16362;
w17011 <= not w16353 and w17010;
w17012 <= not w16919 and w17011;
w17013 <= not w16353 and not w16362;
w17014 <= not w16919 and w17013;
w17015 <= not w16360 and not w17014;
w17016 <= not w17012 and not w17015;
w17017 <= w12199 and not w16997;
w17018 <= not w17007 and w17017;
w17019 <= not w17016 and not w17018;
w17020 <= not w17009 and not w17019;
w17021 <= not w11663 and not w17020;
w17022 <= not w16365 and w16372;
w17023 <= not w16374 and w17022;
w17024 <= not w16919 and w17023;
w17025 <= not w16365 and not w16374;
w17026 <= not w16919 and w17025;
w17027 <= not w16372 and not w17026;
w17028 <= not w17024 and not w17027;
w17029 <= w11663 and not w17009;
w17030 <= not w17019 and w17029;
w17031 <= not w17028 and not w17030;
w17032 <= not w17021 and not w17031;
w17033 <= not w11139 and not w17032;
w17034 <= w16384 and not w16386;
w17035 <= not w16377 and w17034;
w17036 <= not w16919 and w17035;
w17037 <= not w16377 and not w16386;
w17038 <= not w16919 and w17037;
w17039 <= not w16384 and not w17038;
w17040 <= not w17036 and not w17039;
w17041 <= w11139 and not w17021;
w17042 <= not w17031 and w17041;
w17043 <= not w17040 and not w17042;
w17044 <= not w17033 and not w17043;
w17045 <= not w10627 and not w17044;
w17046 <= not w16389 and w16396;
w17047 <= not w16398 and w17046;
w17048 <= not w16919 and w17047;
w17049 <= not w16389 and not w16398;
w17050 <= not w16919 and w17049;
w17051 <= not w16396 and not w17050;
w17052 <= not w17048 and not w17051;
w17053 <= w10627 and not w17033;
w17054 <= not w17043 and w17053;
w17055 <= not w17052 and not w17054;
w17056 <= not w17045 and not w17055;
w17057 <= not w10127 and not w17056;
w17058 <= w16408 and not w16410;
w17059 <= not w16401 and w17058;
w17060 <= not w16919 and w17059;
w17061 <= not w16401 and not w16410;
w17062 <= not w16919 and w17061;
w17063 <= not w16408 and not w17062;
w17064 <= not w17060 and not w17063;
w17065 <= w10127 and not w17045;
w17066 <= not w17055 and w17065;
w17067 <= not w17064 and not w17066;
w17068 <= not w17057 and not w17067;
w17069 <= not w9639 and not w17068;
w17070 <= not w16413 and w16420;
w17071 <= not w16422 and w17070;
w17072 <= not w16919 and w17071;
w17073 <= not w16413 and not w16422;
w17074 <= not w16919 and w17073;
w17075 <= not w16420 and not w17074;
w17076 <= not w17072 and not w17075;
w17077 <= w9639 and not w17057;
w17078 <= not w17067 and w17077;
w17079 <= not w17076 and not w17078;
w17080 <= not w17069 and not w17079;
w17081 <= not w9163 and not w17080;
w17082 <= w16432 and not w16434;
w17083 <= not w16425 and w17082;
w17084 <= not w16919 and w17083;
w17085 <= not w16425 and not w16434;
w17086 <= not w16919 and w17085;
w17087 <= not w16432 and not w17086;
w17088 <= not w17084 and not w17087;
w17089 <= w9163 and not w17069;
w17090 <= not w17079 and w17089;
w17091 <= not w17088 and not w17090;
w17092 <= not w17081 and not w17091;
w17093 <= not w8699 and not w17092;
w17094 <= not w16437 and w16444;
w17095 <= not w16446 and w17094;
w17096 <= not w16919 and w17095;
w17097 <= not w16437 and not w16446;
w17098 <= not w16919 and w17097;
w17099 <= not w16444 and not w17098;
w17100 <= not w17096 and not w17099;
w17101 <= w8699 and not w17081;
w17102 <= not w17091 and w17101;
w17103 <= not w17100 and not w17102;
w17104 <= not w17093 and not w17103;
w17105 <= not w8247 and not w17104;
w17106 <= w16456 and not w16458;
w17107 <= not w16449 and w17106;
w17108 <= not w16919 and w17107;
w17109 <= not w16449 and not w16458;
w17110 <= not w16919 and w17109;
w17111 <= not w16456 and not w17110;
w17112 <= not w17108 and not w17111;
w17113 <= w8247 and not w17093;
w17114 <= not w17103 and w17113;
w17115 <= not w17112 and not w17114;
w17116 <= not w17105 and not w17115;
w17117 <= not w7807 and not w17116;
w17118 <= not w16461 and w16468;
w17119 <= not w16470 and w17118;
w17120 <= not w16919 and w17119;
w17121 <= not w16461 and not w16470;
w17122 <= not w16919 and w17121;
w17123 <= not w16468 and not w17122;
w17124 <= not w17120 and not w17123;
w17125 <= w7807 and not w17105;
w17126 <= not w17115 and w17125;
w17127 <= not w17124 and not w17126;
w17128 <= not w17117 and not w17127;
w17129 <= not w7379 and not w17128;
w17130 <= w16480 and not w16482;
w17131 <= not w16473 and w17130;
w17132 <= not w16919 and w17131;
w17133 <= not w16473 and not w16482;
w17134 <= not w16919 and w17133;
w17135 <= not w16480 and not w17134;
w17136 <= not w17132 and not w17135;
w17137 <= w7379 and not w17117;
w17138 <= not w17127 and w17137;
w17139 <= not w17136 and not w17138;
w17140 <= not w17129 and not w17139;
w17141 <= not w6963 and not w17140;
w17142 <= not w16485 and w16492;
w17143 <= not w16494 and w17142;
w17144 <= not w16919 and w17143;
w17145 <= not w16485 and not w16494;
w17146 <= not w16919 and w17145;
w17147 <= not w16492 and not w17146;
w17148 <= not w17144 and not w17147;
w17149 <= w6963 and not w17129;
w17150 <= not w17139 and w17149;
w17151 <= not w17148 and not w17150;
w17152 <= not w17141 and not w17151;
w17153 <= not w6558 and not w17152;
w17154 <= w16504 and not w16506;
w17155 <= not w16497 and w17154;
w17156 <= not w16919 and w17155;
w17157 <= not w16497 and not w16506;
w17158 <= not w16919 and w17157;
w17159 <= not w16504 and not w17158;
w17160 <= not w17156 and not w17159;
w17161 <= w6558 and not w17141;
w17162 <= not w17151 and w17161;
w17163 <= not w17160 and not w17162;
w17164 <= not w17153 and not w17163;
w17165 <= not w6166 and not w17164;
w17166 <= not w16509 and w16516;
w17167 <= not w16518 and w17166;
w17168 <= not w16919 and w17167;
w17169 <= not w16509 and not w16518;
w17170 <= not w16919 and w17169;
w17171 <= not w16516 and not w17170;
w17172 <= not w17168 and not w17171;
w17173 <= w6166 and not w17153;
w17174 <= not w17163 and w17173;
w17175 <= not w17172 and not w17174;
w17176 <= not w17165 and not w17175;
w17177 <= not w5786 and not w17176;
w17178 <= w16528 and not w16530;
w17179 <= not w16521 and w17178;
w17180 <= not w16919 and w17179;
w17181 <= not w16521 and not w16530;
w17182 <= not w16919 and w17181;
w17183 <= not w16528 and not w17182;
w17184 <= not w17180 and not w17183;
w17185 <= w5786 and not w17165;
w17186 <= not w17175 and w17185;
w17187 <= not w17184 and not w17186;
w17188 <= not w17177 and not w17187;
w17189 <= not w5418 and not w17188;
w17190 <= not w16533 and w16540;
w17191 <= not w16542 and w17190;
w17192 <= not w16919 and w17191;
w17193 <= not w16533 and not w16542;
w17194 <= not w16919 and w17193;
w17195 <= not w16540 and not w17194;
w17196 <= not w17192 and not w17195;
w17197 <= w5418 and not w17177;
w17198 <= not w17187 and w17197;
w17199 <= not w17196 and not w17198;
w17200 <= not w17189 and not w17199;
w17201 <= not w5062 and not w17200;
w17202 <= w16552 and not w16554;
w17203 <= not w16545 and w17202;
w17204 <= not w16919 and w17203;
w17205 <= not w16545 and not w16554;
w17206 <= not w16919 and w17205;
w17207 <= not w16552 and not w17206;
w17208 <= not w17204 and not w17207;
w17209 <= w5062 and not w17189;
w17210 <= not w17199 and w17209;
w17211 <= not w17208 and not w17210;
w17212 <= not w17201 and not w17211;
w17213 <= not w4718 and not w17212;
w17214 <= not w16557 and w16564;
w17215 <= not w16566 and w17214;
w17216 <= not w16919 and w17215;
w17217 <= not w16557 and not w16566;
w17218 <= not w16919 and w17217;
w17219 <= not w16564 and not w17218;
w17220 <= not w17216 and not w17219;
w17221 <= w4718 and not w17201;
w17222 <= not w17211 and w17221;
w17223 <= not w17220 and not w17222;
w17224 <= not w17213 and not w17223;
w17225 <= not w4386 and not w17224;
w17226 <= w16576 and not w16578;
w17227 <= not w16569 and w17226;
w17228 <= not w16919 and w17227;
w17229 <= not w16569 and not w16578;
w17230 <= not w16919 and w17229;
w17231 <= not w16576 and not w17230;
w17232 <= not w17228 and not w17231;
w17233 <= w4386 and not w17213;
w17234 <= not w17223 and w17233;
w17235 <= not w17232 and not w17234;
w17236 <= not w17225 and not w17235;
w17237 <= not w4066 and not w17236;
w17238 <= not w16581 and w16588;
w17239 <= not w16590 and w17238;
w17240 <= not w16919 and w17239;
w17241 <= not w16581 and not w16590;
w17242 <= not w16919 and w17241;
w17243 <= not w16588 and not w17242;
w17244 <= not w17240 and not w17243;
w17245 <= w4066 and not w17225;
w17246 <= not w17235 and w17245;
w17247 <= not w17244 and not w17246;
w17248 <= not w17237 and not w17247;
w17249 <= not w3758 and not w17248;
w17250 <= w16600 and not w16602;
w17251 <= not w16593 and w17250;
w17252 <= not w16919 and w17251;
w17253 <= not w16593 and not w16602;
w17254 <= not w16919 and w17253;
w17255 <= not w16600 and not w17254;
w17256 <= not w17252 and not w17255;
w17257 <= w3758 and not w17237;
w17258 <= not w17247 and w17257;
w17259 <= not w17256 and not w17258;
w17260 <= not w17249 and not w17259;
w17261 <= not w3462 and not w17260;
w17262 <= not w16605 and w16612;
w17263 <= not w16614 and w17262;
w17264 <= not w16919 and w17263;
w17265 <= not w16605 and not w16614;
w17266 <= not w16919 and w17265;
w17267 <= not w16612 and not w17266;
w17268 <= not w17264 and not w17267;
w17269 <= w3462 and not w17249;
w17270 <= not w17259 and w17269;
w17271 <= not w17268 and not w17270;
w17272 <= not w17261 and not w17271;
w17273 <= not w3178 and not w17272;
w17274 <= w16624 and not w16626;
w17275 <= not w16617 and w17274;
w17276 <= not w16919 and w17275;
w17277 <= not w16617 and not w16626;
w17278 <= not w16919 and w17277;
w17279 <= not w16624 and not w17278;
w17280 <= not w17276 and not w17279;
w17281 <= w3178 and not w17261;
w17282 <= not w17271 and w17281;
w17283 <= not w17280 and not w17282;
w17284 <= not w17273 and not w17283;
w17285 <= not w2906 and not w17284;
w17286 <= not w16629 and w16636;
w17287 <= not w16638 and w17286;
w17288 <= not w16919 and w17287;
w17289 <= not w16629 and not w16638;
w17290 <= not w16919 and w17289;
w17291 <= not w16636 and not w17290;
w17292 <= not w17288 and not w17291;
w17293 <= w2906 and not w17273;
w17294 <= not w17283 and w17293;
w17295 <= not w17292 and not w17294;
w17296 <= not w17285 and not w17295;
w17297 <= not w2646 and not w17296;
w17298 <= w16648 and not w16650;
w17299 <= not w16641 and w17298;
w17300 <= not w16919 and w17299;
w17301 <= not w16641 and not w16650;
w17302 <= not w16919 and w17301;
w17303 <= not w16648 and not w17302;
w17304 <= not w17300 and not w17303;
w17305 <= w2646 and not w17285;
w17306 <= not w17295 and w17305;
w17307 <= not w17304 and not w17306;
w17308 <= not w17297 and not w17307;
w17309 <= not w2398 and not w17308;
w17310 <= not w16653 and w16660;
w17311 <= not w16662 and w17310;
w17312 <= not w16919 and w17311;
w17313 <= not w16653 and not w16662;
w17314 <= not w16919 and w17313;
w17315 <= not w16660 and not w17314;
w17316 <= not w17312 and not w17315;
w17317 <= w2398 and not w17297;
w17318 <= not w17307 and w17317;
w17319 <= not w17316 and not w17318;
w17320 <= not w17309 and not w17319;
w17321 <= not w2162 and not w17320;
w17322 <= w16672 and not w16674;
w17323 <= not w16665 and w17322;
w17324 <= not w16919 and w17323;
w17325 <= not w16665 and not w16674;
w17326 <= not w16919 and w17325;
w17327 <= not w16672 and not w17326;
w17328 <= not w17324 and not w17327;
w17329 <= w2162 and not w17309;
w17330 <= not w17319 and w17329;
w17331 <= not w17328 and not w17330;
w17332 <= not w17321 and not w17331;
w17333 <= not w1938 and not w17332;
w17334 <= not w16677 and w16684;
w17335 <= not w16686 and w17334;
w17336 <= not w16919 and w17335;
w17337 <= not w16677 and not w16686;
w17338 <= not w16919 and w17337;
w17339 <= not w16684 and not w17338;
w17340 <= not w17336 and not w17339;
w17341 <= w1938 and not w17321;
w17342 <= not w17331 and w17341;
w17343 <= not w17340 and not w17342;
w17344 <= not w17333 and not w17343;
w17345 <= not w1725 and not w17344;
w17346 <= w16696 and not w16698;
w17347 <= not w16689 and w17346;
w17348 <= not w16919 and w17347;
w17349 <= not w16689 and not w16698;
w17350 <= not w16919 and w17349;
w17351 <= not w16696 and not w17350;
w17352 <= not w17348 and not w17351;
w17353 <= w1725 and not w17333;
w17354 <= not w17343 and w17353;
w17355 <= not w17352 and not w17354;
w17356 <= not w17345 and not w17355;
w17357 <= not w1525 and not w17356;
w17358 <= not w16701 and w16708;
w17359 <= not w16710 and w17358;
w17360 <= not w16919 and w17359;
w17361 <= not w16701 and not w16710;
w17362 <= not w16919 and w17361;
w17363 <= not w16708 and not w17362;
w17364 <= not w17360 and not w17363;
w17365 <= w1525 and not w17345;
w17366 <= not w17355 and w17365;
w17367 <= not w17364 and not w17366;
w17368 <= not w17357 and not w17367;
w17369 <= not w1337 and not w17368;
w17370 <= w16720 and not w16722;
w17371 <= not w16713 and w17370;
w17372 <= not w16919 and w17371;
w17373 <= not w16713 and not w16722;
w17374 <= not w16919 and w17373;
w17375 <= not w16720 and not w17374;
w17376 <= not w17372 and not w17375;
w17377 <= w1337 and not w17357;
w17378 <= not w17367 and w17377;
w17379 <= not w17376 and not w17378;
w17380 <= not w17369 and not w17379;
w17381 <= not w1161 and not w17380;
w17382 <= not w16725 and w16732;
w17383 <= not w16734 and w17382;
w17384 <= not w16919 and w17383;
w17385 <= not w16725 and not w16734;
w17386 <= not w16919 and w17385;
w17387 <= not w16732 and not w17386;
w17388 <= not w17384 and not w17387;
w17389 <= w1161 and not w17369;
w17390 <= not w17379 and w17389;
w17391 <= not w17388 and not w17390;
w17392 <= not w17381 and not w17391;
w17393 <= not w997 and not w17392;
w17394 <= w16744 and not w16746;
w17395 <= not w16737 and w17394;
w17396 <= not w16919 and w17395;
w17397 <= not w16737 and not w16746;
w17398 <= not w16919 and w17397;
w17399 <= not w16744 and not w17398;
w17400 <= not w17396 and not w17399;
w17401 <= w997 and not w17381;
w17402 <= not w17391 and w17401;
w17403 <= not w17400 and not w17402;
w17404 <= not w17393 and not w17403;
w17405 <= not w845 and not w17404;
w17406 <= not w16749 and w16756;
w17407 <= not w16758 and w17406;
w17408 <= not w16919 and w17407;
w17409 <= not w16749 and not w16758;
w17410 <= not w16919 and w17409;
w17411 <= not w16756 and not w17410;
w17412 <= not w17408 and not w17411;
w17413 <= w845 and not w17393;
w17414 <= not w17403 and w17413;
w17415 <= not w17412 and not w17414;
w17416 <= not w17405 and not w17415;
w17417 <= not w705 and not w17416;
w17418 <= w16768 and not w16770;
w17419 <= not w16761 and w17418;
w17420 <= not w16919 and w17419;
w17421 <= not w16761 and not w16770;
w17422 <= not w16919 and w17421;
w17423 <= not w16768 and not w17422;
w17424 <= not w17420 and not w17423;
w17425 <= w705 and not w17405;
w17426 <= not w17415 and w17425;
w17427 <= not w17424 and not w17426;
w17428 <= not w17417 and not w17427;
w17429 <= not w577 and not w17428;
w17430 <= w577 and not w17417;
w17431 <= not w17427 and w17430;
w17432 <= not w16773 and w16782;
w17433 <= not w16775 and w17432;
w17434 <= not w16919 and w17433;
w17435 <= not w16773 and not w16775;
w17436 <= not w16919 and w17435;
w17437 <= not w16782 and not w17436;
w17438 <= not w17434 and not w17437;
w17439 <= not w17431 and not w17438;
w17440 <= not w17429 and not w17439;
w17441 <= not w460 and not w17440;
w17442 <= w16792 and not w16794;
w17443 <= not w16785 and w17442;
w17444 <= not w16919 and w17443;
w17445 <= not w16785 and not w16794;
w17446 <= not w16919 and w17445;
w17447 <= not w16792 and not w17446;
w17448 <= not w17444 and not w17447;
w17449 <= w460 and not w17429;
w17450 <= not w17439 and w17449;
w17451 <= not w17448 and not w17450;
w17452 <= not w17441 and not w17451;
w17453 <= not w356 and not w17452;
w17454 <= not w16797 and w16804;
w17455 <= not w16806 and w17454;
w17456 <= not w16919 and w17455;
w17457 <= not w16797 and not w16806;
w17458 <= not w16919 and w17457;
w17459 <= not w16804 and not w17458;
w17460 <= not w17456 and not w17459;
w17461 <= w356 and not w17441;
w17462 <= not w17451 and w17461;
w17463 <= not w17460 and not w17462;
w17464 <= not w17453 and not w17463;
w17465 <= not w264 and not w17464;
w17466 <= w16816 and not w16818;
w17467 <= not w16809 and w17466;
w17468 <= not w16919 and w17467;
w17469 <= not w16809 and not w16818;
w17470 <= not w16919 and w17469;
w17471 <= not w16816 and not w17470;
w17472 <= not w17468 and not w17471;
w17473 <= w264 and not w17453;
w17474 <= not w17463 and w17473;
w17475 <= not w17472 and not w17474;
w17476 <= not w17465 and not w17475;
w17477 <= not w184 and not w17476;
w17478 <= not w16821 and w16828;
w17479 <= not w16830 and w17478;
w17480 <= not w16919 and w17479;
w17481 <= not w16821 and not w16830;
w17482 <= not w16919 and w17481;
w17483 <= not w16828 and not w17482;
w17484 <= not w17480 and not w17483;
w17485 <= w184 and not w17465;
w17486 <= not w17475 and w17485;
w17487 <= not w17484 and not w17486;
w17488 <= not w17477 and not w17487;
w17489 <= not w115 and not w17488;
w17490 <= w16840 and not w16842;
w17491 <= not w16833 and w17490;
w17492 <= not w16919 and w17491;
w17493 <= not w16833 and not w16842;
w17494 <= not w16919 and w17493;
w17495 <= not w16840 and not w17494;
w17496 <= not w17492 and not w17495;
w17497 <= w115 and not w17477;
w17498 <= not w17487 and w17497;
w17499 <= not w17496 and not w17498;
w17500 <= not w17489 and not w17499;
w17501 <= not w60 and not w17500;
w17502 <= not w16845 and w16852;
w17503 <= not w16854 and w17502;
w17504 <= not w16919 and w17503;
w17505 <= not w16845 and not w16854;
w17506 <= not w16919 and w17505;
w17507 <= not w16852 and not w17506;
w17508 <= not w17504 and not w17507;
w17509 <= w60 and not w17489;
w17510 <= not w17499 and w17509;
w17511 <= not w17508 and not w17510;
w17512 <= not w17501 and not w17511;
w17513 <= not w22 and not w17512;
w17514 <= w16864 and not w16866;
w17515 <= not w16857 and w17514;
w17516 <= not w16919 and w17515;
w17517 <= not w16857 and not w16866;
w17518 <= not w16919 and w17517;
w17519 <= not w16864 and not w17518;
w17520 <= not w17516 and not w17519;
w17521 <= w22 and not w17501;
w17522 <= not w17511 and w17521;
w17523 <= not w17520 and not w17522;
w17524 <= not w17513 and not w17523;
w17525 <= not w5 and not w17524;
w17526 <= not w16869 and w16876;
w17527 <= not w16878 and w17526;
w17528 <= not w16919 and w17527;
w17529 <= not w16869 and not w16878;
w17530 <= not w16919 and w17529;
w17531 <= not w16876 and not w17530;
w17532 <= not w17528 and not w17531;
w17533 <= w5 and not w17513;
w17534 <= not w17523 and w17533;
w17535 <= not w17532 and not w17534;
w17536 <= not w17525 and not w17535;
w17537 <= w16888 and not w16890;
w17538 <= not w16881 and w17537;
w17539 <= not w16919 and w17538;
w17540 <= not w16881 and not w16890;
w17541 <= not w16919 and w17540;
w17542 <= not w16888 and not w17541;
w17543 <= not w17539 and not w17542;
w17544 <= not w16892 and not w16899;
w17545 <= not w16919 and w17544;
w17546 <= not w16907 and not w17545;
w17547 <= not w17543 and w17546;
w17548 <= not w17536 and w17547;
w17549 <= w0 and not w17548;
w17550 <= not w17525 and w17543;
w17551 <= not w17535 and w17550;
w17552 <= not w16899 and not w16919;
w17553 <= w16892 and not w17552;
w17554 <= not w0 and not w17544;
w17555 <= not w17553 and w17554;
w17556 <= not w16895 and not w16916;
w17557 <= not w16898 and w17556;
w17558 <= not w16911 and w17557;
w17559 <= not w16907 and w17558;
w17560 <= not w16905 and w17559;
w17561 <= not w17555 and not w17560;
w17562 <= not w17551 and w17561;
w17563 <= not w17549 and w17562;
w17564 <= a(20) and not w17563;
w17565 <= not a(18) and not a(19);
w17566 <= not a(20) and w17565;
w17567 <= not w17564 and not w17566;
w17568 <= not w16919 and not w17567;
w17569 <= not w16916 and not w17566;
w17570 <= not w16911 and w17569;
w17571 <= not w16907 and w17570;
w17572 <= not w16905 and w17571;
w17573 <= not w17564 and w17572;
w17574 <= not a(20) and not w17563;
w17575 <= a(21) and not w17574;
w17576 <= w16921 and not w17563;
w17577 <= not w17575 and not w17576;
w17578 <= not w17573 and w17577;
w17579 <= not w17568 and not w17578;
w17580 <= not w16287 and not w17579;
w17581 <= w16287 and not w17568;
w17582 <= not w17578 and w17581;
w17583 <= not w16919 and not w17560;
w17584 <= not w17555 and w17583;
w17585 <= not w17551 and w17584;
w17586 <= not w17549 and w17585;
w17587 <= not w17576 and not w17586;
w17588 <= a(22) and not w17587;
w17589 <= not a(22) and not w17586;
w17590 <= not w17576 and w17589;
w17591 <= not w17588 and not w17590;
w17592 <= not w17582 and not w17591;
w17593 <= not w17580 and not w17592;
w17594 <= not w15667 and not w17593;
w17595 <= not w16924 and not w16929;
w17596 <= not w16933 and w17595;
w17597 <= not w17563 and w17596;
w17598 <= not w17563 and w17595;
w17599 <= w16933 and not w17598;
w17600 <= not w17597 and not w17599;
w17601 <= w15667 and not w17580;
w17602 <= not w17592 and w17601;
w17603 <= not w17600 and not w17602;
w17604 <= not w17594 and not w17603;
w17605 <= not w15059 and not w17604;
w17606 <= not w16938 and w16947;
w17607 <= not w16936 and w17606;
w17608 <= not w17563 and w17607;
w17609 <= not w16936 and not w16938;
w17610 <= not w17563 and w17609;
w17611 <= not w16947 and not w17610;
w17612 <= not w17608 and not w17611;
w17613 <= w15059 and not w17594;
w17614 <= not w17603 and w17613;
w17615 <= not w17612 and not w17614;
w17616 <= not w17605 and not w17615;
w17617 <= not w14463 and not w17616;
w17618 <= not w16950 and w16956;
w17619 <= not w16958 and w17618;
w17620 <= not w17563 and w17619;
w17621 <= not w16950 and not w16958;
w17622 <= not w17563 and w17621;
w17623 <= not w16956 and not w17622;
w17624 <= not w17620 and not w17623;
w17625 <= w14463 and not w17605;
w17626 <= not w17615 and w17625;
w17627 <= not w17624 and not w17626;
w17628 <= not w17617 and not w17627;
w17629 <= not w13879 and not w17628;
w17630 <= w16968 and not w16970;
w17631 <= not w16961 and w17630;
w17632 <= not w17563 and w17631;
w17633 <= not w16961 and not w16970;
w17634 <= not w17563 and w17633;
w17635 <= not w16968 and not w17634;
w17636 <= not w17632 and not w17635;
w17637 <= w13879 and not w17617;
w17638 <= not w17627 and w17637;
w17639 <= not w17636 and not w17638;
w17640 <= not w17629 and not w17639;
w17641 <= not w13307 and not w17640;
w17642 <= not w16973 and w16980;
w17643 <= not w16982 and w17642;
w17644 <= not w17563 and w17643;
w17645 <= not w16973 and not w16982;
w17646 <= not w17563 and w17645;
w17647 <= not w16980 and not w17646;
w17648 <= not w17644 and not w17647;
w17649 <= w13307 and not w17629;
w17650 <= not w17639 and w17649;
w17651 <= not w17648 and not w17650;
w17652 <= not w17641 and not w17651;
w17653 <= not w12747 and not w17652;
w17654 <= w16992 and not w16994;
w17655 <= not w16985 and w17654;
w17656 <= not w17563 and w17655;
w17657 <= not w16985 and not w16994;
w17658 <= not w17563 and w17657;
w17659 <= not w16992 and not w17658;
w17660 <= not w17656 and not w17659;
w17661 <= w12747 and not w17641;
w17662 <= not w17651 and w17661;
w17663 <= not w17660 and not w17662;
w17664 <= not w17653 and not w17663;
w17665 <= not w12199 and not w17664;
w17666 <= not w16997 and w17004;
w17667 <= not w17006 and w17666;
w17668 <= not w17563 and w17667;
w17669 <= not w16997 and not w17006;
w17670 <= not w17563 and w17669;
w17671 <= not w17004 and not w17670;
w17672 <= not w17668 and not w17671;
w17673 <= w12199 and not w17653;
w17674 <= not w17663 and w17673;
w17675 <= not w17672 and not w17674;
w17676 <= not w17665 and not w17675;
w17677 <= not w11663 and not w17676;
w17678 <= w17016 and not w17018;
w17679 <= not w17009 and w17678;
w17680 <= not w17563 and w17679;
w17681 <= not w17009 and not w17018;
w17682 <= not w17563 and w17681;
w17683 <= not w17016 and not w17682;
w17684 <= not w17680 and not w17683;
w17685 <= w11663 and not w17665;
w17686 <= not w17675 and w17685;
w17687 <= not w17684 and not w17686;
w17688 <= not w17677 and not w17687;
w17689 <= not w11139 and not w17688;
w17690 <= not w17021 and w17028;
w17691 <= not w17030 and w17690;
w17692 <= not w17563 and w17691;
w17693 <= not w17021 and not w17030;
w17694 <= not w17563 and w17693;
w17695 <= not w17028 and not w17694;
w17696 <= not w17692 and not w17695;
w17697 <= w11139 and not w17677;
w17698 <= not w17687 and w17697;
w17699 <= not w17696 and not w17698;
w17700 <= not w17689 and not w17699;
w17701 <= not w10627 and not w17700;
w17702 <= w17040 and not w17042;
w17703 <= not w17033 and w17702;
w17704 <= not w17563 and w17703;
w17705 <= not w17033 and not w17042;
w17706 <= not w17563 and w17705;
w17707 <= not w17040 and not w17706;
w17708 <= not w17704 and not w17707;
w17709 <= w10627 and not w17689;
w17710 <= not w17699 and w17709;
w17711 <= not w17708 and not w17710;
w17712 <= not w17701 and not w17711;
w17713 <= not w10127 and not w17712;
w17714 <= not w17045 and w17052;
w17715 <= not w17054 and w17714;
w17716 <= not w17563 and w17715;
w17717 <= not w17045 and not w17054;
w17718 <= not w17563 and w17717;
w17719 <= not w17052 and not w17718;
w17720 <= not w17716 and not w17719;
w17721 <= w10127 and not w17701;
w17722 <= not w17711 and w17721;
w17723 <= not w17720 and not w17722;
w17724 <= not w17713 and not w17723;
w17725 <= not w9639 and not w17724;
w17726 <= w17064 and not w17066;
w17727 <= not w17057 and w17726;
w17728 <= not w17563 and w17727;
w17729 <= not w17057 and not w17066;
w17730 <= not w17563 and w17729;
w17731 <= not w17064 and not w17730;
w17732 <= not w17728 and not w17731;
w17733 <= w9639 and not w17713;
w17734 <= not w17723 and w17733;
w17735 <= not w17732 and not w17734;
w17736 <= not w17725 and not w17735;
w17737 <= not w9163 and not w17736;
w17738 <= not w17069 and w17076;
w17739 <= not w17078 and w17738;
w17740 <= not w17563 and w17739;
w17741 <= not w17069 and not w17078;
w17742 <= not w17563 and w17741;
w17743 <= not w17076 and not w17742;
w17744 <= not w17740 and not w17743;
w17745 <= w9163 and not w17725;
w17746 <= not w17735 and w17745;
w17747 <= not w17744 and not w17746;
w17748 <= not w17737 and not w17747;
w17749 <= not w8699 and not w17748;
w17750 <= w17088 and not w17090;
w17751 <= not w17081 and w17750;
w17752 <= not w17563 and w17751;
w17753 <= not w17081 and not w17090;
w17754 <= not w17563 and w17753;
w17755 <= not w17088 and not w17754;
w17756 <= not w17752 and not w17755;
w17757 <= w8699 and not w17737;
w17758 <= not w17747 and w17757;
w17759 <= not w17756 and not w17758;
w17760 <= not w17749 and not w17759;
w17761 <= not w8247 and not w17760;
w17762 <= not w17093 and w17100;
w17763 <= not w17102 and w17762;
w17764 <= not w17563 and w17763;
w17765 <= not w17093 and not w17102;
w17766 <= not w17563 and w17765;
w17767 <= not w17100 and not w17766;
w17768 <= not w17764 and not w17767;
w17769 <= w8247 and not w17749;
w17770 <= not w17759 and w17769;
w17771 <= not w17768 and not w17770;
w17772 <= not w17761 and not w17771;
w17773 <= not w7807 and not w17772;
w17774 <= w17112 and not w17114;
w17775 <= not w17105 and w17774;
w17776 <= not w17563 and w17775;
w17777 <= not w17105 and not w17114;
w17778 <= not w17563 and w17777;
w17779 <= not w17112 and not w17778;
w17780 <= not w17776 and not w17779;
w17781 <= w7807 and not w17761;
w17782 <= not w17771 and w17781;
w17783 <= not w17780 and not w17782;
w17784 <= not w17773 and not w17783;
w17785 <= not w7379 and not w17784;
w17786 <= not w17117 and w17124;
w17787 <= not w17126 and w17786;
w17788 <= not w17563 and w17787;
w17789 <= not w17117 and not w17126;
w17790 <= not w17563 and w17789;
w17791 <= not w17124 and not w17790;
w17792 <= not w17788 and not w17791;
w17793 <= w7379 and not w17773;
w17794 <= not w17783 and w17793;
w17795 <= not w17792 and not w17794;
w17796 <= not w17785 and not w17795;
w17797 <= not w6963 and not w17796;
w17798 <= w17136 and not w17138;
w17799 <= not w17129 and w17798;
w17800 <= not w17563 and w17799;
w17801 <= not w17129 and not w17138;
w17802 <= not w17563 and w17801;
w17803 <= not w17136 and not w17802;
w17804 <= not w17800 and not w17803;
w17805 <= w6963 and not w17785;
w17806 <= not w17795 and w17805;
w17807 <= not w17804 and not w17806;
w17808 <= not w17797 and not w17807;
w17809 <= not w6558 and not w17808;
w17810 <= not w17141 and w17148;
w17811 <= not w17150 and w17810;
w17812 <= not w17563 and w17811;
w17813 <= not w17141 and not w17150;
w17814 <= not w17563 and w17813;
w17815 <= not w17148 and not w17814;
w17816 <= not w17812 and not w17815;
w17817 <= w6558 and not w17797;
w17818 <= not w17807 and w17817;
w17819 <= not w17816 and not w17818;
w17820 <= not w17809 and not w17819;
w17821 <= not w6166 and not w17820;
w17822 <= w17160 and not w17162;
w17823 <= not w17153 and w17822;
w17824 <= not w17563 and w17823;
w17825 <= not w17153 and not w17162;
w17826 <= not w17563 and w17825;
w17827 <= not w17160 and not w17826;
w17828 <= not w17824 and not w17827;
w17829 <= w6166 and not w17809;
w17830 <= not w17819 and w17829;
w17831 <= not w17828 and not w17830;
w17832 <= not w17821 and not w17831;
w17833 <= not w5786 and not w17832;
w17834 <= not w17165 and w17172;
w17835 <= not w17174 and w17834;
w17836 <= not w17563 and w17835;
w17837 <= not w17165 and not w17174;
w17838 <= not w17563 and w17837;
w17839 <= not w17172 and not w17838;
w17840 <= not w17836 and not w17839;
w17841 <= w5786 and not w17821;
w17842 <= not w17831 and w17841;
w17843 <= not w17840 and not w17842;
w17844 <= not w17833 and not w17843;
w17845 <= not w5418 and not w17844;
w17846 <= w17184 and not w17186;
w17847 <= not w17177 and w17846;
w17848 <= not w17563 and w17847;
w17849 <= not w17177 and not w17186;
w17850 <= not w17563 and w17849;
w17851 <= not w17184 and not w17850;
w17852 <= not w17848 and not w17851;
w17853 <= w5418 and not w17833;
w17854 <= not w17843 and w17853;
w17855 <= not w17852 and not w17854;
w17856 <= not w17845 and not w17855;
w17857 <= not w5062 and not w17856;
w17858 <= not w17189 and w17196;
w17859 <= not w17198 and w17858;
w17860 <= not w17563 and w17859;
w17861 <= not w17189 and not w17198;
w17862 <= not w17563 and w17861;
w17863 <= not w17196 and not w17862;
w17864 <= not w17860 and not w17863;
w17865 <= w5062 and not w17845;
w17866 <= not w17855 and w17865;
w17867 <= not w17864 and not w17866;
w17868 <= not w17857 and not w17867;
w17869 <= not w4718 and not w17868;
w17870 <= w17208 and not w17210;
w17871 <= not w17201 and w17870;
w17872 <= not w17563 and w17871;
w17873 <= not w17201 and not w17210;
w17874 <= not w17563 and w17873;
w17875 <= not w17208 and not w17874;
w17876 <= not w17872 and not w17875;
w17877 <= w4718 and not w17857;
w17878 <= not w17867 and w17877;
w17879 <= not w17876 and not w17878;
w17880 <= not w17869 and not w17879;
w17881 <= not w4386 and not w17880;
w17882 <= not w17213 and w17220;
w17883 <= not w17222 and w17882;
w17884 <= not w17563 and w17883;
w17885 <= not w17213 and not w17222;
w17886 <= not w17563 and w17885;
w17887 <= not w17220 and not w17886;
w17888 <= not w17884 and not w17887;
w17889 <= w4386 and not w17869;
w17890 <= not w17879 and w17889;
w17891 <= not w17888 and not w17890;
w17892 <= not w17881 and not w17891;
w17893 <= not w4066 and not w17892;
w17894 <= w17232 and not w17234;
w17895 <= not w17225 and w17894;
w17896 <= not w17563 and w17895;
w17897 <= not w17225 and not w17234;
w17898 <= not w17563 and w17897;
w17899 <= not w17232 and not w17898;
w17900 <= not w17896 and not w17899;
w17901 <= w4066 and not w17881;
w17902 <= not w17891 and w17901;
w17903 <= not w17900 and not w17902;
w17904 <= not w17893 and not w17903;
w17905 <= not w3758 and not w17904;
w17906 <= not w17237 and w17244;
w17907 <= not w17246 and w17906;
w17908 <= not w17563 and w17907;
w17909 <= not w17237 and not w17246;
w17910 <= not w17563 and w17909;
w17911 <= not w17244 and not w17910;
w17912 <= not w17908 and not w17911;
w17913 <= w3758 and not w17893;
w17914 <= not w17903 and w17913;
w17915 <= not w17912 and not w17914;
w17916 <= not w17905 and not w17915;
w17917 <= not w3462 and not w17916;
w17918 <= w17256 and not w17258;
w17919 <= not w17249 and w17918;
w17920 <= not w17563 and w17919;
w17921 <= not w17249 and not w17258;
w17922 <= not w17563 and w17921;
w17923 <= not w17256 and not w17922;
w17924 <= not w17920 and not w17923;
w17925 <= w3462 and not w17905;
w17926 <= not w17915 and w17925;
w17927 <= not w17924 and not w17926;
w17928 <= not w17917 and not w17927;
w17929 <= not w3178 and not w17928;
w17930 <= not w17261 and w17268;
w17931 <= not w17270 and w17930;
w17932 <= not w17563 and w17931;
w17933 <= not w17261 and not w17270;
w17934 <= not w17563 and w17933;
w17935 <= not w17268 and not w17934;
w17936 <= not w17932 and not w17935;
w17937 <= w3178 and not w17917;
w17938 <= not w17927 and w17937;
w17939 <= not w17936 and not w17938;
w17940 <= not w17929 and not w17939;
w17941 <= not w2906 and not w17940;
w17942 <= w17280 and not w17282;
w17943 <= not w17273 and w17942;
w17944 <= not w17563 and w17943;
w17945 <= not w17273 and not w17282;
w17946 <= not w17563 and w17945;
w17947 <= not w17280 and not w17946;
w17948 <= not w17944 and not w17947;
w17949 <= w2906 and not w17929;
w17950 <= not w17939 and w17949;
w17951 <= not w17948 and not w17950;
w17952 <= not w17941 and not w17951;
w17953 <= not w2646 and not w17952;
w17954 <= not w17285 and w17292;
w17955 <= not w17294 and w17954;
w17956 <= not w17563 and w17955;
w17957 <= not w17285 and not w17294;
w17958 <= not w17563 and w17957;
w17959 <= not w17292 and not w17958;
w17960 <= not w17956 and not w17959;
w17961 <= w2646 and not w17941;
w17962 <= not w17951 and w17961;
w17963 <= not w17960 and not w17962;
w17964 <= not w17953 and not w17963;
w17965 <= not w2398 and not w17964;
w17966 <= w17304 and not w17306;
w17967 <= not w17297 and w17966;
w17968 <= not w17563 and w17967;
w17969 <= not w17297 and not w17306;
w17970 <= not w17563 and w17969;
w17971 <= not w17304 and not w17970;
w17972 <= not w17968 and not w17971;
w17973 <= w2398 and not w17953;
w17974 <= not w17963 and w17973;
w17975 <= not w17972 and not w17974;
w17976 <= not w17965 and not w17975;
w17977 <= not w2162 and not w17976;
w17978 <= not w17309 and w17316;
w17979 <= not w17318 and w17978;
w17980 <= not w17563 and w17979;
w17981 <= not w17309 and not w17318;
w17982 <= not w17563 and w17981;
w17983 <= not w17316 and not w17982;
w17984 <= not w17980 and not w17983;
w17985 <= w2162 and not w17965;
w17986 <= not w17975 and w17985;
w17987 <= not w17984 and not w17986;
w17988 <= not w17977 and not w17987;
w17989 <= not w1938 and not w17988;
w17990 <= w17328 and not w17330;
w17991 <= not w17321 and w17990;
w17992 <= not w17563 and w17991;
w17993 <= not w17321 and not w17330;
w17994 <= not w17563 and w17993;
w17995 <= not w17328 and not w17994;
w17996 <= not w17992 and not w17995;
w17997 <= w1938 and not w17977;
w17998 <= not w17987 and w17997;
w17999 <= not w17996 and not w17998;
w18000 <= not w17989 and not w17999;
w18001 <= not w1725 and not w18000;
w18002 <= not w17333 and w17340;
w18003 <= not w17342 and w18002;
w18004 <= not w17563 and w18003;
w18005 <= not w17333 and not w17342;
w18006 <= not w17563 and w18005;
w18007 <= not w17340 and not w18006;
w18008 <= not w18004 and not w18007;
w18009 <= w1725 and not w17989;
w18010 <= not w17999 and w18009;
w18011 <= not w18008 and not w18010;
w18012 <= not w18001 and not w18011;
w18013 <= not w1525 and not w18012;
w18014 <= w17352 and not w17354;
w18015 <= not w17345 and w18014;
w18016 <= not w17563 and w18015;
w18017 <= not w17345 and not w17354;
w18018 <= not w17563 and w18017;
w18019 <= not w17352 and not w18018;
w18020 <= not w18016 and not w18019;
w18021 <= w1525 and not w18001;
w18022 <= not w18011 and w18021;
w18023 <= not w18020 and not w18022;
w18024 <= not w18013 and not w18023;
w18025 <= not w1337 and not w18024;
w18026 <= not w17357 and w17364;
w18027 <= not w17366 and w18026;
w18028 <= not w17563 and w18027;
w18029 <= not w17357 and not w17366;
w18030 <= not w17563 and w18029;
w18031 <= not w17364 and not w18030;
w18032 <= not w18028 and not w18031;
w18033 <= w1337 and not w18013;
w18034 <= not w18023 and w18033;
w18035 <= not w18032 and not w18034;
w18036 <= not w18025 and not w18035;
w18037 <= not w1161 and not w18036;
w18038 <= w17376 and not w17378;
w18039 <= not w17369 and w18038;
w18040 <= not w17563 and w18039;
w18041 <= not w17369 and not w17378;
w18042 <= not w17563 and w18041;
w18043 <= not w17376 and not w18042;
w18044 <= not w18040 and not w18043;
w18045 <= w1161 and not w18025;
w18046 <= not w18035 and w18045;
w18047 <= not w18044 and not w18046;
w18048 <= not w18037 and not w18047;
w18049 <= not w997 and not w18048;
w18050 <= not w17381 and w17388;
w18051 <= not w17390 and w18050;
w18052 <= not w17563 and w18051;
w18053 <= not w17381 and not w17390;
w18054 <= not w17563 and w18053;
w18055 <= not w17388 and not w18054;
w18056 <= not w18052 and not w18055;
w18057 <= w997 and not w18037;
w18058 <= not w18047 and w18057;
w18059 <= not w18056 and not w18058;
w18060 <= not w18049 and not w18059;
w18061 <= not w845 and not w18060;
w18062 <= w17400 and not w17402;
w18063 <= not w17393 and w18062;
w18064 <= not w17563 and w18063;
w18065 <= not w17393 and not w17402;
w18066 <= not w17563 and w18065;
w18067 <= not w17400 and not w18066;
w18068 <= not w18064 and not w18067;
w18069 <= w845 and not w18049;
w18070 <= not w18059 and w18069;
w18071 <= not w18068 and not w18070;
w18072 <= not w18061 and not w18071;
w18073 <= not w705 and not w18072;
w18074 <= not w17405 and w17412;
w18075 <= not w17414 and w18074;
w18076 <= not w17563 and w18075;
w18077 <= not w17405 and not w17414;
w18078 <= not w17563 and w18077;
w18079 <= not w17412 and not w18078;
w18080 <= not w18076 and not w18079;
w18081 <= w705 and not w18061;
w18082 <= not w18071 and w18081;
w18083 <= not w18080 and not w18082;
w18084 <= not w18073 and not w18083;
w18085 <= not w577 and not w18084;
w18086 <= w17424 and not w17426;
w18087 <= not w17417 and w18086;
w18088 <= not w17563 and w18087;
w18089 <= not w17417 and not w17426;
w18090 <= not w17563 and w18089;
w18091 <= not w17424 and not w18090;
w18092 <= not w18088 and not w18091;
w18093 <= w577 and not w18073;
w18094 <= not w18083 and w18093;
w18095 <= not w18092 and not w18094;
w18096 <= not w18085 and not w18095;
w18097 <= not w460 and not w18096;
w18098 <= w460 and not w18085;
w18099 <= not w18095 and w18098;
w18100 <= not w17429 and w17438;
w18101 <= not w17431 and w18100;
w18102 <= not w17563 and w18101;
w18103 <= not w17429 and not w17431;
w18104 <= not w17563 and w18103;
w18105 <= not w17438 and not w18104;
w18106 <= not w18102 and not w18105;
w18107 <= not w18099 and not w18106;
w18108 <= not w18097 and not w18107;
w18109 <= not w356 and not w18108;
w18110 <= w17448 and not w17450;
w18111 <= not w17441 and w18110;
w18112 <= not w17563 and w18111;
w18113 <= not w17441 and not w17450;
w18114 <= not w17563 and w18113;
w18115 <= not w17448 and not w18114;
w18116 <= not w18112 and not w18115;
w18117 <= w356 and not w18097;
w18118 <= not w18107 and w18117;
w18119 <= not w18116 and not w18118;
w18120 <= not w18109 and not w18119;
w18121 <= not w264 and not w18120;
w18122 <= not w17453 and w17460;
w18123 <= not w17462 and w18122;
w18124 <= not w17563 and w18123;
w18125 <= not w17453 and not w17462;
w18126 <= not w17563 and w18125;
w18127 <= not w17460 and not w18126;
w18128 <= not w18124 and not w18127;
w18129 <= w264 and not w18109;
w18130 <= not w18119 and w18129;
w18131 <= not w18128 and not w18130;
w18132 <= not w18121 and not w18131;
w18133 <= not w184 and not w18132;
w18134 <= w17472 and not w17474;
w18135 <= not w17465 and w18134;
w18136 <= not w17563 and w18135;
w18137 <= not w17465 and not w17474;
w18138 <= not w17563 and w18137;
w18139 <= not w17472 and not w18138;
w18140 <= not w18136 and not w18139;
w18141 <= w184 and not w18121;
w18142 <= not w18131 and w18141;
w18143 <= not w18140 and not w18142;
w18144 <= not w18133 and not w18143;
w18145 <= not w115 and not w18144;
w18146 <= not w17477 and w17484;
w18147 <= not w17486 and w18146;
w18148 <= not w17563 and w18147;
w18149 <= not w17477 and not w17486;
w18150 <= not w17563 and w18149;
w18151 <= not w17484 and not w18150;
w18152 <= not w18148 and not w18151;
w18153 <= w115 and not w18133;
w18154 <= not w18143 and w18153;
w18155 <= not w18152 and not w18154;
w18156 <= not w18145 and not w18155;
w18157 <= not w60 and not w18156;
w18158 <= w17496 and not w17498;
w18159 <= not w17489 and w18158;
w18160 <= not w17563 and w18159;
w18161 <= not w17489 and not w17498;
w18162 <= not w17563 and w18161;
w18163 <= not w17496 and not w18162;
w18164 <= not w18160 and not w18163;
w18165 <= w60 and not w18145;
w18166 <= not w18155 and w18165;
w18167 <= not w18164 and not w18166;
w18168 <= not w18157 and not w18167;
w18169 <= not w22 and not w18168;
w18170 <= not w17501 and w17508;
w18171 <= not w17510 and w18170;
w18172 <= not w17563 and w18171;
w18173 <= not w17501 and not w17510;
w18174 <= not w17563 and w18173;
w18175 <= not w17508 and not w18174;
w18176 <= not w18172 and not w18175;
w18177 <= w22 and not w18157;
w18178 <= not w18167 and w18177;
w18179 <= not w18176 and not w18178;
w18180 <= not w18169 and not w18179;
w18181 <= not w5 and not w18180;
w18182 <= w17520 and not w17522;
w18183 <= not w17513 and w18182;
w18184 <= not w17563 and w18183;
w18185 <= not w17513 and not w17522;
w18186 <= not w17563 and w18185;
w18187 <= not w17520 and not w18186;
w18188 <= not w18184 and not w18187;
w18189 <= w5 and not w18169;
w18190 <= not w18179 and w18189;
w18191 <= not w18188 and not w18190;
w18192 <= not w18181 and not w18191;
w18193 <= not w17525 and w17532;
w18194 <= not w17534 and w18193;
w18195 <= not w17563 and w18194;
w18196 <= not w17525 and not w17534;
w18197 <= not w17563 and w18196;
w18198 <= not w17532 and not w18197;
w18199 <= not w18195 and not w18198;
w18200 <= not w17536 and not w17543;
w18201 <= not w17563 and w18200;
w18202 <= not w17551 and not w18201;
w18203 <= not w18199 and w18202;
w18204 <= not w18192 and w18203;
w18205 <= w0 and not w18204;
w18206 <= not w18181 and w18199;
w18207 <= not w18191 and w18206;
w18208 <= not w17543 and not w17563;
w18209 <= w17536 and not w18208;
w18210 <= not w0 and not w18200;
w18211 <= not w18209 and w18210;
w18212 <= not w17539 and not w17560;
w18213 <= not w17542 and w18212;
w18214 <= not w17555 and w18213;
w18215 <= not w17551 and w18214;
w18216 <= not w17549 and w18215;
w18217 <= not w18211 and not w18216;
w18218 <= not w18207 and w18217;
w18219 <= not w18205 and w18218;
w18220 <= a(18) and not w18219;
w18221 <= not a(16) and not a(17);
w18222 <= not a(18) and w18221;
w18223 <= not w18220 and not w18222;
w18224 <= not w17563 and not w18223;
w18225 <= not w17560 and not w18222;
w18226 <= not w17555 and w18225;
w18227 <= not w17551 and w18226;
w18228 <= not w17549 and w18227;
w18229 <= not w18220 and w18228;
w18230 <= not a(18) and not w18219;
w18231 <= a(19) and not w18230;
w18232 <= w17565 and not w18219;
w18233 <= not w18231 and not w18232;
w18234 <= not w18229 and w18233;
w18235 <= not w18224 and not w18234;
w18236 <= not w16919 and not w18235;
w18237 <= w16919 and not w18224;
w18238 <= not w18234 and w18237;
w18239 <= not w17563 and not w18216;
w18240 <= not w18211 and w18239;
w18241 <= not w18207 and w18240;
w18242 <= not w18205 and w18241;
w18243 <= not w18232 and not w18242;
w18244 <= a(20) and not w18243;
w18245 <= not a(20) and not w18242;
w18246 <= not w18232 and w18245;
w18247 <= not w18244 and not w18246;
w18248 <= not w18238 and not w18247;
w18249 <= not w18236 and not w18248;
w18250 <= not w16287 and not w18249;
w18251 <= not w17568 and not w17573;
w18252 <= not w17577 and w18251;
w18253 <= not w18219 and w18252;
w18254 <= not w18219 and w18251;
w18255 <= w17577 and not w18254;
w18256 <= not w18253 and not w18255;
w18257 <= w16287 and not w18236;
w18258 <= not w18248 and w18257;
w18259 <= not w18256 and not w18258;
w18260 <= not w18250 and not w18259;
w18261 <= not w15667 and not w18260;
w18262 <= not w17582 and w17591;
w18263 <= not w17580 and w18262;
w18264 <= not w18219 and w18263;
w18265 <= not w17580 and not w17582;
w18266 <= not w18219 and w18265;
w18267 <= not w17591 and not w18266;
w18268 <= not w18264 and not w18267;
w18269 <= w15667 and not w18250;
w18270 <= not w18259 and w18269;
w18271 <= not w18268 and not w18270;
w18272 <= not w18261 and not w18271;
w18273 <= not w15059 and not w18272;
w18274 <= not w17594 and w17600;
w18275 <= not w17602 and w18274;
w18276 <= not w18219 and w18275;
w18277 <= not w17594 and not w17602;
w18278 <= not w18219 and w18277;
w18279 <= not w17600 and not w18278;
w18280 <= not w18276 and not w18279;
w18281 <= w15059 and not w18261;
w18282 <= not w18271 and w18281;
w18283 <= not w18280 and not w18282;
w18284 <= not w18273 and not w18283;
w18285 <= not w14463 and not w18284;
w18286 <= w17612 and not w17614;
w18287 <= not w17605 and w18286;
w18288 <= not w18219 and w18287;
w18289 <= not w17605 and not w17614;
w18290 <= not w18219 and w18289;
w18291 <= not w17612 and not w18290;
w18292 <= not w18288 and not w18291;
w18293 <= w14463 and not w18273;
w18294 <= not w18283 and w18293;
w18295 <= not w18292 and not w18294;
w18296 <= not w18285 and not w18295;
w18297 <= not w13879 and not w18296;
w18298 <= not w17617 and w17624;
w18299 <= not w17626 and w18298;
w18300 <= not w18219 and w18299;
w18301 <= not w17617 and not w17626;
w18302 <= not w18219 and w18301;
w18303 <= not w17624 and not w18302;
w18304 <= not w18300 and not w18303;
w18305 <= w13879 and not w18285;
w18306 <= not w18295 and w18305;
w18307 <= not w18304 and not w18306;
w18308 <= not w18297 and not w18307;
w18309 <= not w13307 and not w18308;
w18310 <= w17636 and not w17638;
w18311 <= not w17629 and w18310;
w18312 <= not w18219 and w18311;
w18313 <= not w17629 and not w17638;
w18314 <= not w18219 and w18313;
w18315 <= not w17636 and not w18314;
w18316 <= not w18312 and not w18315;
w18317 <= w13307 and not w18297;
w18318 <= not w18307 and w18317;
w18319 <= not w18316 and not w18318;
w18320 <= not w18309 and not w18319;
w18321 <= not w12747 and not w18320;
w18322 <= not w17641 and w17648;
w18323 <= not w17650 and w18322;
w18324 <= not w18219 and w18323;
w18325 <= not w17641 and not w17650;
w18326 <= not w18219 and w18325;
w18327 <= not w17648 and not w18326;
w18328 <= not w18324 and not w18327;
w18329 <= w12747 and not w18309;
w18330 <= not w18319 and w18329;
w18331 <= not w18328 and not w18330;
w18332 <= not w18321 and not w18331;
w18333 <= not w12199 and not w18332;
w18334 <= w17660 and not w17662;
w18335 <= not w17653 and w18334;
w18336 <= not w18219 and w18335;
w18337 <= not w17653 and not w17662;
w18338 <= not w18219 and w18337;
w18339 <= not w17660 and not w18338;
w18340 <= not w18336 and not w18339;
w18341 <= w12199 and not w18321;
w18342 <= not w18331 and w18341;
w18343 <= not w18340 and not w18342;
w18344 <= not w18333 and not w18343;
w18345 <= not w11663 and not w18344;
w18346 <= not w17665 and w17672;
w18347 <= not w17674 and w18346;
w18348 <= not w18219 and w18347;
w18349 <= not w17665 and not w17674;
w18350 <= not w18219 and w18349;
w18351 <= not w17672 and not w18350;
w18352 <= not w18348 and not w18351;
w18353 <= w11663 and not w18333;
w18354 <= not w18343 and w18353;
w18355 <= not w18352 and not w18354;
w18356 <= not w18345 and not w18355;
w18357 <= not w11139 and not w18356;
w18358 <= w17684 and not w17686;
w18359 <= not w17677 and w18358;
w18360 <= not w18219 and w18359;
w18361 <= not w17677 and not w17686;
w18362 <= not w18219 and w18361;
w18363 <= not w17684 and not w18362;
w18364 <= not w18360 and not w18363;
w18365 <= w11139 and not w18345;
w18366 <= not w18355 and w18365;
w18367 <= not w18364 and not w18366;
w18368 <= not w18357 and not w18367;
w18369 <= not w10627 and not w18368;
w18370 <= not w17689 and w17696;
w18371 <= not w17698 and w18370;
w18372 <= not w18219 and w18371;
w18373 <= not w17689 and not w17698;
w18374 <= not w18219 and w18373;
w18375 <= not w17696 and not w18374;
w18376 <= not w18372 and not w18375;
w18377 <= w10627 and not w18357;
w18378 <= not w18367 and w18377;
w18379 <= not w18376 and not w18378;
w18380 <= not w18369 and not w18379;
w18381 <= not w10127 and not w18380;
w18382 <= w17708 and not w17710;
w18383 <= not w17701 and w18382;
w18384 <= not w18219 and w18383;
w18385 <= not w17701 and not w17710;
w18386 <= not w18219 and w18385;
w18387 <= not w17708 and not w18386;
w18388 <= not w18384 and not w18387;
w18389 <= w10127 and not w18369;
w18390 <= not w18379 and w18389;
w18391 <= not w18388 and not w18390;
w18392 <= not w18381 and not w18391;
w18393 <= not w9639 and not w18392;
w18394 <= not w17713 and w17720;
w18395 <= not w17722 and w18394;
w18396 <= not w18219 and w18395;
w18397 <= not w17713 and not w17722;
w18398 <= not w18219 and w18397;
w18399 <= not w17720 and not w18398;
w18400 <= not w18396 and not w18399;
w18401 <= w9639 and not w18381;
w18402 <= not w18391 and w18401;
w18403 <= not w18400 and not w18402;
w18404 <= not w18393 and not w18403;
w18405 <= not w9163 and not w18404;
w18406 <= w17732 and not w17734;
w18407 <= not w17725 and w18406;
w18408 <= not w18219 and w18407;
w18409 <= not w17725 and not w17734;
w18410 <= not w18219 and w18409;
w18411 <= not w17732 and not w18410;
w18412 <= not w18408 and not w18411;
w18413 <= w9163 and not w18393;
w18414 <= not w18403 and w18413;
w18415 <= not w18412 and not w18414;
w18416 <= not w18405 and not w18415;
w18417 <= not w8699 and not w18416;
w18418 <= not w17737 and w17744;
w18419 <= not w17746 and w18418;
w18420 <= not w18219 and w18419;
w18421 <= not w17737 and not w17746;
w18422 <= not w18219 and w18421;
w18423 <= not w17744 and not w18422;
w18424 <= not w18420 and not w18423;
w18425 <= w8699 and not w18405;
w18426 <= not w18415 and w18425;
w18427 <= not w18424 and not w18426;
w18428 <= not w18417 and not w18427;
w18429 <= not w8247 and not w18428;
w18430 <= w17756 and not w17758;
w18431 <= not w17749 and w18430;
w18432 <= not w18219 and w18431;
w18433 <= not w17749 and not w17758;
w18434 <= not w18219 and w18433;
w18435 <= not w17756 and not w18434;
w18436 <= not w18432 and not w18435;
w18437 <= w8247 and not w18417;
w18438 <= not w18427 and w18437;
w18439 <= not w18436 and not w18438;
w18440 <= not w18429 and not w18439;
w18441 <= not w7807 and not w18440;
w18442 <= not w17761 and w17768;
w18443 <= not w17770 and w18442;
w18444 <= not w18219 and w18443;
w18445 <= not w17761 and not w17770;
w18446 <= not w18219 and w18445;
w18447 <= not w17768 and not w18446;
w18448 <= not w18444 and not w18447;
w18449 <= w7807 and not w18429;
w18450 <= not w18439 and w18449;
w18451 <= not w18448 and not w18450;
w18452 <= not w18441 and not w18451;
w18453 <= not w7379 and not w18452;
w18454 <= w17780 and not w17782;
w18455 <= not w17773 and w18454;
w18456 <= not w18219 and w18455;
w18457 <= not w17773 and not w17782;
w18458 <= not w18219 and w18457;
w18459 <= not w17780 and not w18458;
w18460 <= not w18456 and not w18459;
w18461 <= w7379 and not w18441;
w18462 <= not w18451 and w18461;
w18463 <= not w18460 and not w18462;
w18464 <= not w18453 and not w18463;
w18465 <= not w6963 and not w18464;
w18466 <= not w17785 and w17792;
w18467 <= not w17794 and w18466;
w18468 <= not w18219 and w18467;
w18469 <= not w17785 and not w17794;
w18470 <= not w18219 and w18469;
w18471 <= not w17792 and not w18470;
w18472 <= not w18468 and not w18471;
w18473 <= w6963 and not w18453;
w18474 <= not w18463 and w18473;
w18475 <= not w18472 and not w18474;
w18476 <= not w18465 and not w18475;
w18477 <= not w6558 and not w18476;
w18478 <= w17804 and not w17806;
w18479 <= not w17797 and w18478;
w18480 <= not w18219 and w18479;
w18481 <= not w17797 and not w17806;
w18482 <= not w18219 and w18481;
w18483 <= not w17804 and not w18482;
w18484 <= not w18480 and not w18483;
w18485 <= w6558 and not w18465;
w18486 <= not w18475 and w18485;
w18487 <= not w18484 and not w18486;
w18488 <= not w18477 and not w18487;
w18489 <= not w6166 and not w18488;
w18490 <= not w17809 and w17816;
w18491 <= not w17818 and w18490;
w18492 <= not w18219 and w18491;
w18493 <= not w17809 and not w17818;
w18494 <= not w18219 and w18493;
w18495 <= not w17816 and not w18494;
w18496 <= not w18492 and not w18495;
w18497 <= w6166 and not w18477;
w18498 <= not w18487 and w18497;
w18499 <= not w18496 and not w18498;
w18500 <= not w18489 and not w18499;
w18501 <= not w5786 and not w18500;
w18502 <= w17828 and not w17830;
w18503 <= not w17821 and w18502;
w18504 <= not w18219 and w18503;
w18505 <= not w17821 and not w17830;
w18506 <= not w18219 and w18505;
w18507 <= not w17828 and not w18506;
w18508 <= not w18504 and not w18507;
w18509 <= w5786 and not w18489;
w18510 <= not w18499 and w18509;
w18511 <= not w18508 and not w18510;
w18512 <= not w18501 and not w18511;
w18513 <= not w5418 and not w18512;
w18514 <= not w17833 and w17840;
w18515 <= not w17842 and w18514;
w18516 <= not w18219 and w18515;
w18517 <= not w17833 and not w17842;
w18518 <= not w18219 and w18517;
w18519 <= not w17840 and not w18518;
w18520 <= not w18516 and not w18519;
w18521 <= w5418 and not w18501;
w18522 <= not w18511 and w18521;
w18523 <= not w18520 and not w18522;
w18524 <= not w18513 and not w18523;
w18525 <= not w5062 and not w18524;
w18526 <= w17852 and not w17854;
w18527 <= not w17845 and w18526;
w18528 <= not w18219 and w18527;
w18529 <= not w17845 and not w17854;
w18530 <= not w18219 and w18529;
w18531 <= not w17852 and not w18530;
w18532 <= not w18528 and not w18531;
w18533 <= w5062 and not w18513;
w18534 <= not w18523 and w18533;
w18535 <= not w18532 and not w18534;
w18536 <= not w18525 and not w18535;
w18537 <= not w4718 and not w18536;
w18538 <= not w17857 and w17864;
w18539 <= not w17866 and w18538;
w18540 <= not w18219 and w18539;
w18541 <= not w17857 and not w17866;
w18542 <= not w18219 and w18541;
w18543 <= not w17864 and not w18542;
w18544 <= not w18540 and not w18543;
w18545 <= w4718 and not w18525;
w18546 <= not w18535 and w18545;
w18547 <= not w18544 and not w18546;
w18548 <= not w18537 and not w18547;
w18549 <= not w4386 and not w18548;
w18550 <= w17876 and not w17878;
w18551 <= not w17869 and w18550;
w18552 <= not w18219 and w18551;
w18553 <= not w17869 and not w17878;
w18554 <= not w18219 and w18553;
w18555 <= not w17876 and not w18554;
w18556 <= not w18552 and not w18555;
w18557 <= w4386 and not w18537;
w18558 <= not w18547 and w18557;
w18559 <= not w18556 and not w18558;
w18560 <= not w18549 and not w18559;
w18561 <= not w4066 and not w18560;
w18562 <= not w17881 and w17888;
w18563 <= not w17890 and w18562;
w18564 <= not w18219 and w18563;
w18565 <= not w17881 and not w17890;
w18566 <= not w18219 and w18565;
w18567 <= not w17888 and not w18566;
w18568 <= not w18564 and not w18567;
w18569 <= w4066 and not w18549;
w18570 <= not w18559 and w18569;
w18571 <= not w18568 and not w18570;
w18572 <= not w18561 and not w18571;
w18573 <= not w3758 and not w18572;
w18574 <= w17900 and not w17902;
w18575 <= not w17893 and w18574;
w18576 <= not w18219 and w18575;
w18577 <= not w17893 and not w17902;
w18578 <= not w18219 and w18577;
w18579 <= not w17900 and not w18578;
w18580 <= not w18576 and not w18579;
w18581 <= w3758 and not w18561;
w18582 <= not w18571 and w18581;
w18583 <= not w18580 and not w18582;
w18584 <= not w18573 and not w18583;
w18585 <= not w3462 and not w18584;
w18586 <= not w17905 and w17912;
w18587 <= not w17914 and w18586;
w18588 <= not w18219 and w18587;
w18589 <= not w17905 and not w17914;
w18590 <= not w18219 and w18589;
w18591 <= not w17912 and not w18590;
w18592 <= not w18588 and not w18591;
w18593 <= w3462 and not w18573;
w18594 <= not w18583 and w18593;
w18595 <= not w18592 and not w18594;
w18596 <= not w18585 and not w18595;
w18597 <= not w3178 and not w18596;
w18598 <= w17924 and not w17926;
w18599 <= not w17917 and w18598;
w18600 <= not w18219 and w18599;
w18601 <= not w17917 and not w17926;
w18602 <= not w18219 and w18601;
w18603 <= not w17924 and not w18602;
w18604 <= not w18600 and not w18603;
w18605 <= w3178 and not w18585;
w18606 <= not w18595 and w18605;
w18607 <= not w18604 and not w18606;
w18608 <= not w18597 and not w18607;
w18609 <= not w2906 and not w18608;
w18610 <= not w17929 and w17936;
w18611 <= not w17938 and w18610;
w18612 <= not w18219 and w18611;
w18613 <= not w17929 and not w17938;
w18614 <= not w18219 and w18613;
w18615 <= not w17936 and not w18614;
w18616 <= not w18612 and not w18615;
w18617 <= w2906 and not w18597;
w18618 <= not w18607 and w18617;
w18619 <= not w18616 and not w18618;
w18620 <= not w18609 and not w18619;
w18621 <= not w2646 and not w18620;
w18622 <= w17948 and not w17950;
w18623 <= not w17941 and w18622;
w18624 <= not w18219 and w18623;
w18625 <= not w17941 and not w17950;
w18626 <= not w18219 and w18625;
w18627 <= not w17948 and not w18626;
w18628 <= not w18624 and not w18627;
w18629 <= w2646 and not w18609;
w18630 <= not w18619 and w18629;
w18631 <= not w18628 and not w18630;
w18632 <= not w18621 and not w18631;
w18633 <= not w2398 and not w18632;
w18634 <= not w17953 and w17960;
w18635 <= not w17962 and w18634;
w18636 <= not w18219 and w18635;
w18637 <= not w17953 and not w17962;
w18638 <= not w18219 and w18637;
w18639 <= not w17960 and not w18638;
w18640 <= not w18636 and not w18639;
w18641 <= w2398 and not w18621;
w18642 <= not w18631 and w18641;
w18643 <= not w18640 and not w18642;
w18644 <= not w18633 and not w18643;
w18645 <= not w2162 and not w18644;
w18646 <= w17972 and not w17974;
w18647 <= not w17965 and w18646;
w18648 <= not w18219 and w18647;
w18649 <= not w17965 and not w17974;
w18650 <= not w18219 and w18649;
w18651 <= not w17972 and not w18650;
w18652 <= not w18648 and not w18651;
w18653 <= w2162 and not w18633;
w18654 <= not w18643 and w18653;
w18655 <= not w18652 and not w18654;
w18656 <= not w18645 and not w18655;
w18657 <= not w1938 and not w18656;
w18658 <= not w17977 and w17984;
w18659 <= not w17986 and w18658;
w18660 <= not w18219 and w18659;
w18661 <= not w17977 and not w17986;
w18662 <= not w18219 and w18661;
w18663 <= not w17984 and not w18662;
w18664 <= not w18660 and not w18663;
w18665 <= w1938 and not w18645;
w18666 <= not w18655 and w18665;
w18667 <= not w18664 and not w18666;
w18668 <= not w18657 and not w18667;
w18669 <= not w1725 and not w18668;
w18670 <= w17996 and not w17998;
w18671 <= not w17989 and w18670;
w18672 <= not w18219 and w18671;
w18673 <= not w17989 and not w17998;
w18674 <= not w18219 and w18673;
w18675 <= not w17996 and not w18674;
w18676 <= not w18672 and not w18675;
w18677 <= w1725 and not w18657;
w18678 <= not w18667 and w18677;
w18679 <= not w18676 and not w18678;
w18680 <= not w18669 and not w18679;
w18681 <= not w1525 and not w18680;
w18682 <= not w18001 and w18008;
w18683 <= not w18010 and w18682;
w18684 <= not w18219 and w18683;
w18685 <= not w18001 and not w18010;
w18686 <= not w18219 and w18685;
w18687 <= not w18008 and not w18686;
w18688 <= not w18684 and not w18687;
w18689 <= w1525 and not w18669;
w18690 <= not w18679 and w18689;
w18691 <= not w18688 and not w18690;
w18692 <= not w18681 and not w18691;
w18693 <= not w1337 and not w18692;
w18694 <= w18020 and not w18022;
w18695 <= not w18013 and w18694;
w18696 <= not w18219 and w18695;
w18697 <= not w18013 and not w18022;
w18698 <= not w18219 and w18697;
w18699 <= not w18020 and not w18698;
w18700 <= not w18696 and not w18699;
w18701 <= w1337 and not w18681;
w18702 <= not w18691 and w18701;
w18703 <= not w18700 and not w18702;
w18704 <= not w18693 and not w18703;
w18705 <= not w1161 and not w18704;
w18706 <= not w18025 and w18032;
w18707 <= not w18034 and w18706;
w18708 <= not w18219 and w18707;
w18709 <= not w18025 and not w18034;
w18710 <= not w18219 and w18709;
w18711 <= not w18032 and not w18710;
w18712 <= not w18708 and not w18711;
w18713 <= w1161 and not w18693;
w18714 <= not w18703 and w18713;
w18715 <= not w18712 and not w18714;
w18716 <= not w18705 and not w18715;
w18717 <= not w997 and not w18716;
w18718 <= w18044 and not w18046;
w18719 <= not w18037 and w18718;
w18720 <= not w18219 and w18719;
w18721 <= not w18037 and not w18046;
w18722 <= not w18219 and w18721;
w18723 <= not w18044 and not w18722;
w18724 <= not w18720 and not w18723;
w18725 <= w997 and not w18705;
w18726 <= not w18715 and w18725;
w18727 <= not w18724 and not w18726;
w18728 <= not w18717 and not w18727;
w18729 <= not w845 and not w18728;
w18730 <= not w18049 and w18056;
w18731 <= not w18058 and w18730;
w18732 <= not w18219 and w18731;
w18733 <= not w18049 and not w18058;
w18734 <= not w18219 and w18733;
w18735 <= not w18056 and not w18734;
w18736 <= not w18732 and not w18735;
w18737 <= w845 and not w18717;
w18738 <= not w18727 and w18737;
w18739 <= not w18736 and not w18738;
w18740 <= not w18729 and not w18739;
w18741 <= not w705 and not w18740;
w18742 <= w18068 and not w18070;
w18743 <= not w18061 and w18742;
w18744 <= not w18219 and w18743;
w18745 <= not w18061 and not w18070;
w18746 <= not w18219 and w18745;
w18747 <= not w18068 and not w18746;
w18748 <= not w18744 and not w18747;
w18749 <= w705 and not w18729;
w18750 <= not w18739 and w18749;
w18751 <= not w18748 and not w18750;
w18752 <= not w18741 and not w18751;
w18753 <= not w577 and not w18752;
w18754 <= not w18073 and w18080;
w18755 <= not w18082 and w18754;
w18756 <= not w18219 and w18755;
w18757 <= not w18073 and not w18082;
w18758 <= not w18219 and w18757;
w18759 <= not w18080 and not w18758;
w18760 <= not w18756 and not w18759;
w18761 <= w577 and not w18741;
w18762 <= not w18751 and w18761;
w18763 <= not w18760 and not w18762;
w18764 <= not w18753 and not w18763;
w18765 <= not w460 and not w18764;
w18766 <= w18092 and not w18094;
w18767 <= not w18085 and w18766;
w18768 <= not w18219 and w18767;
w18769 <= not w18085 and not w18094;
w18770 <= not w18219 and w18769;
w18771 <= not w18092 and not w18770;
w18772 <= not w18768 and not w18771;
w18773 <= w460 and not w18753;
w18774 <= not w18763 and w18773;
w18775 <= not w18772 and not w18774;
w18776 <= not w18765 and not w18775;
w18777 <= not w356 and not w18776;
w18778 <= w356 and not w18765;
w18779 <= not w18775 and w18778;
w18780 <= not w18097 and w18106;
w18781 <= not w18099 and w18780;
w18782 <= not w18219 and w18781;
w18783 <= not w18097 and not w18099;
w18784 <= not w18219 and w18783;
w18785 <= not w18106 and not w18784;
w18786 <= not w18782 and not w18785;
w18787 <= not w18779 and not w18786;
w18788 <= not w18777 and not w18787;
w18789 <= not w264 and not w18788;
w18790 <= w18116 and not w18118;
w18791 <= not w18109 and w18790;
w18792 <= not w18219 and w18791;
w18793 <= not w18109 and not w18118;
w18794 <= not w18219 and w18793;
w18795 <= not w18116 and not w18794;
w18796 <= not w18792 and not w18795;
w18797 <= w264 and not w18777;
w18798 <= not w18787 and w18797;
w18799 <= not w18796 and not w18798;
w18800 <= not w18789 and not w18799;
w18801 <= not w184 and not w18800;
w18802 <= not w18121 and w18128;
w18803 <= not w18130 and w18802;
w18804 <= not w18219 and w18803;
w18805 <= not w18121 and not w18130;
w18806 <= not w18219 and w18805;
w18807 <= not w18128 and not w18806;
w18808 <= not w18804 and not w18807;
w18809 <= w184 and not w18789;
w18810 <= not w18799 and w18809;
w18811 <= not w18808 and not w18810;
w18812 <= not w18801 and not w18811;
w18813 <= not w115 and not w18812;
w18814 <= w18140 and not w18142;
w18815 <= not w18133 and w18814;
w18816 <= not w18219 and w18815;
w18817 <= not w18133 and not w18142;
w18818 <= not w18219 and w18817;
w18819 <= not w18140 and not w18818;
w18820 <= not w18816 and not w18819;
w18821 <= w115 and not w18801;
w18822 <= not w18811 and w18821;
w18823 <= not w18820 and not w18822;
w18824 <= not w18813 and not w18823;
w18825 <= not w60 and not w18824;
w18826 <= not w18145 and w18152;
w18827 <= not w18154 and w18826;
w18828 <= not w18219 and w18827;
w18829 <= not w18145 and not w18154;
w18830 <= not w18219 and w18829;
w18831 <= not w18152 and not w18830;
w18832 <= not w18828 and not w18831;
w18833 <= w60 and not w18813;
w18834 <= not w18823 and w18833;
w18835 <= not w18832 and not w18834;
w18836 <= not w18825 and not w18835;
w18837 <= not w22 and not w18836;
w18838 <= w18164 and not w18166;
w18839 <= not w18157 and w18838;
w18840 <= not w18219 and w18839;
w18841 <= not w18157 and not w18166;
w18842 <= not w18219 and w18841;
w18843 <= not w18164 and not w18842;
w18844 <= not w18840 and not w18843;
w18845 <= w22 and not w18825;
w18846 <= not w18835 and w18845;
w18847 <= not w18844 and not w18846;
w18848 <= not w18837 and not w18847;
w18849 <= not w5 and not w18848;
w18850 <= not w18169 and w18176;
w18851 <= not w18178 and w18850;
w18852 <= not w18219 and w18851;
w18853 <= not w18169 and not w18178;
w18854 <= not w18219 and w18853;
w18855 <= not w18176 and not w18854;
w18856 <= not w18852 and not w18855;
w18857 <= w5 and not w18837;
w18858 <= not w18847 and w18857;
w18859 <= not w18856 and not w18858;
w18860 <= not w18849 and not w18859;
w18861 <= w18188 and not w18190;
w18862 <= not w18181 and w18861;
w18863 <= not w18219 and w18862;
w18864 <= not w18181 and not w18190;
w18865 <= not w18219 and w18864;
w18866 <= not w18188 and not w18865;
w18867 <= not w18863 and not w18866;
w18868 <= not w18192 and not w18199;
w18869 <= not w18219 and w18868;
w18870 <= not w18207 and not w18869;
w18871 <= not w18867 and w18870;
w18872 <= not w18860 and w18871;
w18873 <= w0 and not w18872;
w18874 <= not w18849 and w18867;
w18875 <= not w18859 and w18874;
w18876 <= not w18199 and not w18219;
w18877 <= w18192 and not w18876;
w18878 <= not w0 and not w18868;
w18879 <= not w18877 and w18878;
w18880 <= not w18195 and not w18216;
w18881 <= not w18198 and w18880;
w18882 <= not w18211 and w18881;
w18883 <= not w18207 and w18882;
w18884 <= not w18205 and w18883;
w18885 <= not w18879 and not w18884;
w18886 <= not w18875 and w18885;
w18887 <= not w18873 and w18886;
w18888 <= a(16) and not w18887;
w18889 <= not a(14) and not a(15);
w18890 <= not a(16) and w18889;
w18891 <= not w18888 and not w18890;
w18892 <= not w18219 and not w18891;
w18893 <= not w18216 and not w18890;
w18894 <= not w18211 and w18893;
w18895 <= not w18207 and w18894;
w18896 <= not w18205 and w18895;
w18897 <= not w18888 and w18896;
w18898 <= not a(16) and not w18887;
w18899 <= a(17) and not w18898;
w18900 <= w18221 and not w18887;
w18901 <= not w18899 and not w18900;
w18902 <= not w18897 and w18901;
w18903 <= not w18892 and not w18902;
w18904 <= not w17563 and not w18903;
w18905 <= w17563 and not w18892;
w18906 <= not w18902 and w18905;
w18907 <= not w18219 and not w18884;
w18908 <= not w18879 and w18907;
w18909 <= not w18875 and w18908;
w18910 <= not w18873 and w18909;
w18911 <= not w18900 and not w18910;
w18912 <= a(18) and not w18911;
w18913 <= not a(18) and not w18910;
w18914 <= not w18900 and w18913;
w18915 <= not w18912 and not w18914;
w18916 <= not w18906 and not w18915;
w18917 <= not w18904 and not w18916;
w18918 <= not w16919 and not w18917;
w18919 <= not w18224 and not w18229;
w18920 <= not w18233 and w18919;
w18921 <= not w18887 and w18920;
w18922 <= not w18887 and w18919;
w18923 <= w18233 and not w18922;
w18924 <= not w18921 and not w18923;
w18925 <= w16919 and not w18904;
w18926 <= not w18916 and w18925;
w18927 <= not w18924 and not w18926;
w18928 <= not w18918 and not w18927;
w18929 <= not w16287 and not w18928;
w18930 <= not w18238 and w18247;
w18931 <= not w18236 and w18930;
w18932 <= not w18887 and w18931;
w18933 <= not w18236 and not w18238;
w18934 <= not w18887 and w18933;
w18935 <= not w18247 and not w18934;
w18936 <= not w18932 and not w18935;
w18937 <= w16287 and not w18918;
w18938 <= not w18927 and w18937;
w18939 <= not w18936 and not w18938;
w18940 <= not w18929 and not w18939;
w18941 <= not w15667 and not w18940;
w18942 <= not w18250 and w18256;
w18943 <= not w18258 and w18942;
w18944 <= not w18887 and w18943;
w18945 <= not w18250 and not w18258;
w18946 <= not w18887 and w18945;
w18947 <= not w18256 and not w18946;
w18948 <= not w18944 and not w18947;
w18949 <= w15667 and not w18929;
w18950 <= not w18939 and w18949;
w18951 <= not w18948 and not w18950;
w18952 <= not w18941 and not w18951;
w18953 <= not w15059 and not w18952;
w18954 <= w18268 and not w18270;
w18955 <= not w18261 and w18954;
w18956 <= not w18887 and w18955;
w18957 <= not w18261 and not w18270;
w18958 <= not w18887 and w18957;
w18959 <= not w18268 and not w18958;
w18960 <= not w18956 and not w18959;
w18961 <= w15059 and not w18941;
w18962 <= not w18951 and w18961;
w18963 <= not w18960 and not w18962;
w18964 <= not w18953 and not w18963;
w18965 <= not w14463 and not w18964;
w18966 <= not w18273 and w18280;
w18967 <= not w18282 and w18966;
w18968 <= not w18887 and w18967;
w18969 <= not w18273 and not w18282;
w18970 <= not w18887 and w18969;
w18971 <= not w18280 and not w18970;
w18972 <= not w18968 and not w18971;
w18973 <= w14463 and not w18953;
w18974 <= not w18963 and w18973;
w18975 <= not w18972 and not w18974;
w18976 <= not w18965 and not w18975;
w18977 <= not w13879 and not w18976;
w18978 <= w18292 and not w18294;
w18979 <= not w18285 and w18978;
w18980 <= not w18887 and w18979;
w18981 <= not w18285 and not w18294;
w18982 <= not w18887 and w18981;
w18983 <= not w18292 and not w18982;
w18984 <= not w18980 and not w18983;
w18985 <= w13879 and not w18965;
w18986 <= not w18975 and w18985;
w18987 <= not w18984 and not w18986;
w18988 <= not w18977 and not w18987;
w18989 <= not w13307 and not w18988;
w18990 <= not w18297 and w18304;
w18991 <= not w18306 and w18990;
w18992 <= not w18887 and w18991;
w18993 <= not w18297 and not w18306;
w18994 <= not w18887 and w18993;
w18995 <= not w18304 and not w18994;
w18996 <= not w18992 and not w18995;
w18997 <= w13307 and not w18977;
w18998 <= not w18987 and w18997;
w18999 <= not w18996 and not w18998;
w19000 <= not w18989 and not w18999;
w19001 <= not w12747 and not w19000;
w19002 <= w18316 and not w18318;
w19003 <= not w18309 and w19002;
w19004 <= not w18887 and w19003;
w19005 <= not w18309 and not w18318;
w19006 <= not w18887 and w19005;
w19007 <= not w18316 and not w19006;
w19008 <= not w19004 and not w19007;
w19009 <= w12747 and not w18989;
w19010 <= not w18999 and w19009;
w19011 <= not w19008 and not w19010;
w19012 <= not w19001 and not w19011;
w19013 <= not w12199 and not w19012;
w19014 <= not w18321 and w18328;
w19015 <= not w18330 and w19014;
w19016 <= not w18887 and w19015;
w19017 <= not w18321 and not w18330;
w19018 <= not w18887 and w19017;
w19019 <= not w18328 and not w19018;
w19020 <= not w19016 and not w19019;
w19021 <= w12199 and not w19001;
w19022 <= not w19011 and w19021;
w19023 <= not w19020 and not w19022;
w19024 <= not w19013 and not w19023;
w19025 <= not w11663 and not w19024;
w19026 <= w18340 and not w18342;
w19027 <= not w18333 and w19026;
w19028 <= not w18887 and w19027;
w19029 <= not w18333 and not w18342;
w19030 <= not w18887 and w19029;
w19031 <= not w18340 and not w19030;
w19032 <= not w19028 and not w19031;
w19033 <= w11663 and not w19013;
w19034 <= not w19023 and w19033;
w19035 <= not w19032 and not w19034;
w19036 <= not w19025 and not w19035;
w19037 <= not w11139 and not w19036;
w19038 <= not w18345 and w18352;
w19039 <= not w18354 and w19038;
w19040 <= not w18887 and w19039;
w19041 <= not w18345 and not w18354;
w19042 <= not w18887 and w19041;
w19043 <= not w18352 and not w19042;
w19044 <= not w19040 and not w19043;
w19045 <= w11139 and not w19025;
w19046 <= not w19035 and w19045;
w19047 <= not w19044 and not w19046;
w19048 <= not w19037 and not w19047;
w19049 <= not w10627 and not w19048;
w19050 <= w18364 and not w18366;
w19051 <= not w18357 and w19050;
w19052 <= not w18887 and w19051;
w19053 <= not w18357 and not w18366;
w19054 <= not w18887 and w19053;
w19055 <= not w18364 and not w19054;
w19056 <= not w19052 and not w19055;
w19057 <= w10627 and not w19037;
w19058 <= not w19047 and w19057;
w19059 <= not w19056 and not w19058;
w19060 <= not w19049 and not w19059;
w19061 <= not w10127 and not w19060;
w19062 <= not w18369 and w18376;
w19063 <= not w18378 and w19062;
w19064 <= not w18887 and w19063;
w19065 <= not w18369 and not w18378;
w19066 <= not w18887 and w19065;
w19067 <= not w18376 and not w19066;
w19068 <= not w19064 and not w19067;
w19069 <= w10127 and not w19049;
w19070 <= not w19059 and w19069;
w19071 <= not w19068 and not w19070;
w19072 <= not w19061 and not w19071;
w19073 <= not w9639 and not w19072;
w19074 <= w18388 and not w18390;
w19075 <= not w18381 and w19074;
w19076 <= not w18887 and w19075;
w19077 <= not w18381 and not w18390;
w19078 <= not w18887 and w19077;
w19079 <= not w18388 and not w19078;
w19080 <= not w19076 and not w19079;
w19081 <= w9639 and not w19061;
w19082 <= not w19071 and w19081;
w19083 <= not w19080 and not w19082;
w19084 <= not w19073 and not w19083;
w19085 <= not w9163 and not w19084;
w19086 <= not w18393 and w18400;
w19087 <= not w18402 and w19086;
w19088 <= not w18887 and w19087;
w19089 <= not w18393 and not w18402;
w19090 <= not w18887 and w19089;
w19091 <= not w18400 and not w19090;
w19092 <= not w19088 and not w19091;
w19093 <= w9163 and not w19073;
w19094 <= not w19083 and w19093;
w19095 <= not w19092 and not w19094;
w19096 <= not w19085 and not w19095;
w19097 <= not w8699 and not w19096;
w19098 <= w18412 and not w18414;
w19099 <= not w18405 and w19098;
w19100 <= not w18887 and w19099;
w19101 <= not w18405 and not w18414;
w19102 <= not w18887 and w19101;
w19103 <= not w18412 and not w19102;
w19104 <= not w19100 and not w19103;
w19105 <= w8699 and not w19085;
w19106 <= not w19095 and w19105;
w19107 <= not w19104 and not w19106;
w19108 <= not w19097 and not w19107;
w19109 <= not w8247 and not w19108;
w19110 <= not w18417 and w18424;
w19111 <= not w18426 and w19110;
w19112 <= not w18887 and w19111;
w19113 <= not w18417 and not w18426;
w19114 <= not w18887 and w19113;
w19115 <= not w18424 and not w19114;
w19116 <= not w19112 and not w19115;
w19117 <= w8247 and not w19097;
w19118 <= not w19107 and w19117;
w19119 <= not w19116 and not w19118;
w19120 <= not w19109 and not w19119;
w19121 <= not w7807 and not w19120;
w19122 <= w18436 and not w18438;
w19123 <= not w18429 and w19122;
w19124 <= not w18887 and w19123;
w19125 <= not w18429 and not w18438;
w19126 <= not w18887 and w19125;
w19127 <= not w18436 and not w19126;
w19128 <= not w19124 and not w19127;
w19129 <= w7807 and not w19109;
w19130 <= not w19119 and w19129;
w19131 <= not w19128 and not w19130;
w19132 <= not w19121 and not w19131;
w19133 <= not w7379 and not w19132;
w19134 <= not w18441 and w18448;
w19135 <= not w18450 and w19134;
w19136 <= not w18887 and w19135;
w19137 <= not w18441 and not w18450;
w19138 <= not w18887 and w19137;
w19139 <= not w18448 and not w19138;
w19140 <= not w19136 and not w19139;
w19141 <= w7379 and not w19121;
w19142 <= not w19131 and w19141;
w19143 <= not w19140 and not w19142;
w19144 <= not w19133 and not w19143;
w19145 <= not w6963 and not w19144;
w19146 <= w18460 and not w18462;
w19147 <= not w18453 and w19146;
w19148 <= not w18887 and w19147;
w19149 <= not w18453 and not w18462;
w19150 <= not w18887 and w19149;
w19151 <= not w18460 and not w19150;
w19152 <= not w19148 and not w19151;
w19153 <= w6963 and not w19133;
w19154 <= not w19143 and w19153;
w19155 <= not w19152 and not w19154;
w19156 <= not w19145 and not w19155;
w19157 <= not w6558 and not w19156;
w19158 <= not w18465 and w18472;
w19159 <= not w18474 and w19158;
w19160 <= not w18887 and w19159;
w19161 <= not w18465 and not w18474;
w19162 <= not w18887 and w19161;
w19163 <= not w18472 and not w19162;
w19164 <= not w19160 and not w19163;
w19165 <= w6558 and not w19145;
w19166 <= not w19155 and w19165;
w19167 <= not w19164 and not w19166;
w19168 <= not w19157 and not w19167;
w19169 <= not w6166 and not w19168;
w19170 <= w18484 and not w18486;
w19171 <= not w18477 and w19170;
w19172 <= not w18887 and w19171;
w19173 <= not w18477 and not w18486;
w19174 <= not w18887 and w19173;
w19175 <= not w18484 and not w19174;
w19176 <= not w19172 and not w19175;
w19177 <= w6166 and not w19157;
w19178 <= not w19167 and w19177;
w19179 <= not w19176 and not w19178;
w19180 <= not w19169 and not w19179;
w19181 <= not w5786 and not w19180;
w19182 <= not w18489 and w18496;
w19183 <= not w18498 and w19182;
w19184 <= not w18887 and w19183;
w19185 <= not w18489 and not w18498;
w19186 <= not w18887 and w19185;
w19187 <= not w18496 and not w19186;
w19188 <= not w19184 and not w19187;
w19189 <= w5786 and not w19169;
w19190 <= not w19179 and w19189;
w19191 <= not w19188 and not w19190;
w19192 <= not w19181 and not w19191;
w19193 <= not w5418 and not w19192;
w19194 <= w18508 and not w18510;
w19195 <= not w18501 and w19194;
w19196 <= not w18887 and w19195;
w19197 <= not w18501 and not w18510;
w19198 <= not w18887 and w19197;
w19199 <= not w18508 and not w19198;
w19200 <= not w19196 and not w19199;
w19201 <= w5418 and not w19181;
w19202 <= not w19191 and w19201;
w19203 <= not w19200 and not w19202;
w19204 <= not w19193 and not w19203;
w19205 <= not w5062 and not w19204;
w19206 <= not w18513 and w18520;
w19207 <= not w18522 and w19206;
w19208 <= not w18887 and w19207;
w19209 <= not w18513 and not w18522;
w19210 <= not w18887 and w19209;
w19211 <= not w18520 and not w19210;
w19212 <= not w19208 and not w19211;
w19213 <= w5062 and not w19193;
w19214 <= not w19203 and w19213;
w19215 <= not w19212 and not w19214;
w19216 <= not w19205 and not w19215;
w19217 <= not w4718 and not w19216;
w19218 <= w18532 and not w18534;
w19219 <= not w18525 and w19218;
w19220 <= not w18887 and w19219;
w19221 <= not w18525 and not w18534;
w19222 <= not w18887 and w19221;
w19223 <= not w18532 and not w19222;
w19224 <= not w19220 and not w19223;
w19225 <= w4718 and not w19205;
w19226 <= not w19215 and w19225;
w19227 <= not w19224 and not w19226;
w19228 <= not w19217 and not w19227;
w19229 <= not w4386 and not w19228;
w19230 <= not w18537 and w18544;
w19231 <= not w18546 and w19230;
w19232 <= not w18887 and w19231;
w19233 <= not w18537 and not w18546;
w19234 <= not w18887 and w19233;
w19235 <= not w18544 and not w19234;
w19236 <= not w19232 and not w19235;
w19237 <= w4386 and not w19217;
w19238 <= not w19227 and w19237;
w19239 <= not w19236 and not w19238;
w19240 <= not w19229 and not w19239;
w19241 <= not w4066 and not w19240;
w19242 <= w18556 and not w18558;
w19243 <= not w18549 and w19242;
w19244 <= not w18887 and w19243;
w19245 <= not w18549 and not w18558;
w19246 <= not w18887 and w19245;
w19247 <= not w18556 and not w19246;
w19248 <= not w19244 and not w19247;
w19249 <= w4066 and not w19229;
w19250 <= not w19239 and w19249;
w19251 <= not w19248 and not w19250;
w19252 <= not w19241 and not w19251;
w19253 <= not w3758 and not w19252;
w19254 <= not w18561 and w18568;
w19255 <= not w18570 and w19254;
w19256 <= not w18887 and w19255;
w19257 <= not w18561 and not w18570;
w19258 <= not w18887 and w19257;
w19259 <= not w18568 and not w19258;
w19260 <= not w19256 and not w19259;
w19261 <= w3758 and not w19241;
w19262 <= not w19251 and w19261;
w19263 <= not w19260 and not w19262;
w19264 <= not w19253 and not w19263;
w19265 <= not w3462 and not w19264;
w19266 <= w18580 and not w18582;
w19267 <= not w18573 and w19266;
w19268 <= not w18887 and w19267;
w19269 <= not w18573 and not w18582;
w19270 <= not w18887 and w19269;
w19271 <= not w18580 and not w19270;
w19272 <= not w19268 and not w19271;
w19273 <= w3462 and not w19253;
w19274 <= not w19263 and w19273;
w19275 <= not w19272 and not w19274;
w19276 <= not w19265 and not w19275;
w19277 <= not w3178 and not w19276;
w19278 <= not w18585 and w18592;
w19279 <= not w18594 and w19278;
w19280 <= not w18887 and w19279;
w19281 <= not w18585 and not w18594;
w19282 <= not w18887 and w19281;
w19283 <= not w18592 and not w19282;
w19284 <= not w19280 and not w19283;
w19285 <= w3178 and not w19265;
w19286 <= not w19275 and w19285;
w19287 <= not w19284 and not w19286;
w19288 <= not w19277 and not w19287;
w19289 <= not w2906 and not w19288;
w19290 <= w18604 and not w18606;
w19291 <= not w18597 and w19290;
w19292 <= not w18887 and w19291;
w19293 <= not w18597 and not w18606;
w19294 <= not w18887 and w19293;
w19295 <= not w18604 and not w19294;
w19296 <= not w19292 and not w19295;
w19297 <= w2906 and not w19277;
w19298 <= not w19287 and w19297;
w19299 <= not w19296 and not w19298;
w19300 <= not w19289 and not w19299;
w19301 <= not w2646 and not w19300;
w19302 <= not w18609 and w18616;
w19303 <= not w18618 and w19302;
w19304 <= not w18887 and w19303;
w19305 <= not w18609 and not w18618;
w19306 <= not w18887 and w19305;
w19307 <= not w18616 and not w19306;
w19308 <= not w19304 and not w19307;
w19309 <= w2646 and not w19289;
w19310 <= not w19299 and w19309;
w19311 <= not w19308 and not w19310;
w19312 <= not w19301 and not w19311;
w19313 <= not w2398 and not w19312;
w19314 <= w18628 and not w18630;
w19315 <= not w18621 and w19314;
w19316 <= not w18887 and w19315;
w19317 <= not w18621 and not w18630;
w19318 <= not w18887 and w19317;
w19319 <= not w18628 and not w19318;
w19320 <= not w19316 and not w19319;
w19321 <= w2398 and not w19301;
w19322 <= not w19311 and w19321;
w19323 <= not w19320 and not w19322;
w19324 <= not w19313 and not w19323;
w19325 <= not w2162 and not w19324;
w19326 <= not w18633 and w18640;
w19327 <= not w18642 and w19326;
w19328 <= not w18887 and w19327;
w19329 <= not w18633 and not w18642;
w19330 <= not w18887 and w19329;
w19331 <= not w18640 and not w19330;
w19332 <= not w19328 and not w19331;
w19333 <= w2162 and not w19313;
w19334 <= not w19323 and w19333;
w19335 <= not w19332 and not w19334;
w19336 <= not w19325 and not w19335;
w19337 <= not w1938 and not w19336;
w19338 <= w18652 and not w18654;
w19339 <= not w18645 and w19338;
w19340 <= not w18887 and w19339;
w19341 <= not w18645 and not w18654;
w19342 <= not w18887 and w19341;
w19343 <= not w18652 and not w19342;
w19344 <= not w19340 and not w19343;
w19345 <= w1938 and not w19325;
w19346 <= not w19335 and w19345;
w19347 <= not w19344 and not w19346;
w19348 <= not w19337 and not w19347;
w19349 <= not w1725 and not w19348;
w19350 <= not w18657 and w18664;
w19351 <= not w18666 and w19350;
w19352 <= not w18887 and w19351;
w19353 <= not w18657 and not w18666;
w19354 <= not w18887 and w19353;
w19355 <= not w18664 and not w19354;
w19356 <= not w19352 and not w19355;
w19357 <= w1725 and not w19337;
w19358 <= not w19347 and w19357;
w19359 <= not w19356 and not w19358;
w19360 <= not w19349 and not w19359;
w19361 <= not w1525 and not w19360;
w19362 <= w18676 and not w18678;
w19363 <= not w18669 and w19362;
w19364 <= not w18887 and w19363;
w19365 <= not w18669 and not w18678;
w19366 <= not w18887 and w19365;
w19367 <= not w18676 and not w19366;
w19368 <= not w19364 and not w19367;
w19369 <= w1525 and not w19349;
w19370 <= not w19359 and w19369;
w19371 <= not w19368 and not w19370;
w19372 <= not w19361 and not w19371;
w19373 <= not w1337 and not w19372;
w19374 <= not w18681 and w18688;
w19375 <= not w18690 and w19374;
w19376 <= not w18887 and w19375;
w19377 <= not w18681 and not w18690;
w19378 <= not w18887 and w19377;
w19379 <= not w18688 and not w19378;
w19380 <= not w19376 and not w19379;
w19381 <= w1337 and not w19361;
w19382 <= not w19371 and w19381;
w19383 <= not w19380 and not w19382;
w19384 <= not w19373 and not w19383;
w19385 <= not w1161 and not w19384;
w19386 <= w18700 and not w18702;
w19387 <= not w18693 and w19386;
w19388 <= not w18887 and w19387;
w19389 <= not w18693 and not w18702;
w19390 <= not w18887 and w19389;
w19391 <= not w18700 and not w19390;
w19392 <= not w19388 and not w19391;
w19393 <= w1161 and not w19373;
w19394 <= not w19383 and w19393;
w19395 <= not w19392 and not w19394;
w19396 <= not w19385 and not w19395;
w19397 <= not w997 and not w19396;
w19398 <= not w18705 and w18712;
w19399 <= not w18714 and w19398;
w19400 <= not w18887 and w19399;
w19401 <= not w18705 and not w18714;
w19402 <= not w18887 and w19401;
w19403 <= not w18712 and not w19402;
w19404 <= not w19400 and not w19403;
w19405 <= w997 and not w19385;
w19406 <= not w19395 and w19405;
w19407 <= not w19404 and not w19406;
w19408 <= not w19397 and not w19407;
w19409 <= not w845 and not w19408;
w19410 <= w18724 and not w18726;
w19411 <= not w18717 and w19410;
w19412 <= not w18887 and w19411;
w19413 <= not w18717 and not w18726;
w19414 <= not w18887 and w19413;
w19415 <= not w18724 and not w19414;
w19416 <= not w19412 and not w19415;
w19417 <= w845 and not w19397;
w19418 <= not w19407 and w19417;
w19419 <= not w19416 and not w19418;
w19420 <= not w19409 and not w19419;
w19421 <= not w705 and not w19420;
w19422 <= not w18729 and w18736;
w19423 <= not w18738 and w19422;
w19424 <= not w18887 and w19423;
w19425 <= not w18729 and not w18738;
w19426 <= not w18887 and w19425;
w19427 <= not w18736 and not w19426;
w19428 <= not w19424 and not w19427;
w19429 <= w705 and not w19409;
w19430 <= not w19419 and w19429;
w19431 <= not w19428 and not w19430;
w19432 <= not w19421 and not w19431;
w19433 <= not w577 and not w19432;
w19434 <= w18748 and not w18750;
w19435 <= not w18741 and w19434;
w19436 <= not w18887 and w19435;
w19437 <= not w18741 and not w18750;
w19438 <= not w18887 and w19437;
w19439 <= not w18748 and not w19438;
w19440 <= not w19436 and not w19439;
w19441 <= w577 and not w19421;
w19442 <= not w19431 and w19441;
w19443 <= not w19440 and not w19442;
w19444 <= not w19433 and not w19443;
w19445 <= not w460 and not w19444;
w19446 <= not w18753 and w18760;
w19447 <= not w18762 and w19446;
w19448 <= not w18887 and w19447;
w19449 <= not w18753 and not w18762;
w19450 <= not w18887 and w19449;
w19451 <= not w18760 and not w19450;
w19452 <= not w19448 and not w19451;
w19453 <= w460 and not w19433;
w19454 <= not w19443 and w19453;
w19455 <= not w19452 and not w19454;
w19456 <= not w19445 and not w19455;
w19457 <= not w356 and not w19456;
w19458 <= w18772 and not w18774;
w19459 <= not w18765 and w19458;
w19460 <= not w18887 and w19459;
w19461 <= not w18765 and not w18774;
w19462 <= not w18887 and w19461;
w19463 <= not w18772 and not w19462;
w19464 <= not w19460 and not w19463;
w19465 <= w356 and not w19445;
w19466 <= not w19455 and w19465;
w19467 <= not w19464 and not w19466;
w19468 <= not w19457 and not w19467;
w19469 <= not w264 and not w19468;
w19470 <= w264 and not w19457;
w19471 <= not w19467 and w19470;
w19472 <= not w18777 and w18786;
w19473 <= not w18779 and w19472;
w19474 <= not w18887 and w19473;
w19475 <= not w18777 and not w18779;
w19476 <= not w18887 and w19475;
w19477 <= not w18786 and not w19476;
w19478 <= not w19474 and not w19477;
w19479 <= not w19471 and not w19478;
w19480 <= not w19469 and not w19479;
w19481 <= not w184 and not w19480;
w19482 <= w18796 and not w18798;
w19483 <= not w18789 and w19482;
w19484 <= not w18887 and w19483;
w19485 <= not w18789 and not w18798;
w19486 <= not w18887 and w19485;
w19487 <= not w18796 and not w19486;
w19488 <= not w19484 and not w19487;
w19489 <= w184 and not w19469;
w19490 <= not w19479 and w19489;
w19491 <= not w19488 and not w19490;
w19492 <= not w19481 and not w19491;
w19493 <= not w115 and not w19492;
w19494 <= not w18801 and w18808;
w19495 <= not w18810 and w19494;
w19496 <= not w18887 and w19495;
w19497 <= not w18801 and not w18810;
w19498 <= not w18887 and w19497;
w19499 <= not w18808 and not w19498;
w19500 <= not w19496 and not w19499;
w19501 <= w115 and not w19481;
w19502 <= not w19491 and w19501;
w19503 <= not w19500 and not w19502;
w19504 <= not w19493 and not w19503;
w19505 <= not w60 and not w19504;
w19506 <= w18820 and not w18822;
w19507 <= not w18813 and w19506;
w19508 <= not w18887 and w19507;
w19509 <= not w18813 and not w18822;
w19510 <= not w18887 and w19509;
w19511 <= not w18820 and not w19510;
w19512 <= not w19508 and not w19511;
w19513 <= w60 and not w19493;
w19514 <= not w19503 and w19513;
w19515 <= not w19512 and not w19514;
w19516 <= not w19505 and not w19515;
w19517 <= not w22 and not w19516;
w19518 <= not w18825 and w18832;
w19519 <= not w18834 and w19518;
w19520 <= not w18887 and w19519;
w19521 <= not w18825 and not w18834;
w19522 <= not w18887 and w19521;
w19523 <= not w18832 and not w19522;
w19524 <= not w19520 and not w19523;
w19525 <= w22 and not w19505;
w19526 <= not w19515 and w19525;
w19527 <= not w19524 and not w19526;
w19528 <= not w19517 and not w19527;
w19529 <= not w5 and not w19528;
w19530 <= w18844 and not w18846;
w19531 <= not w18837 and w19530;
w19532 <= not w18887 and w19531;
w19533 <= not w18837 and not w18846;
w19534 <= not w18887 and w19533;
w19535 <= not w18844 and not w19534;
w19536 <= not w19532 and not w19535;
w19537 <= w5 and not w19517;
w19538 <= not w19527 and w19537;
w19539 <= not w19536 and not w19538;
w19540 <= not w19529 and not w19539;
w19541 <= not w18849 and w18856;
w19542 <= not w18858 and w19541;
w19543 <= not w18887 and w19542;
w19544 <= not w18849 and not w18858;
w19545 <= not w18887 and w19544;
w19546 <= not w18856 and not w19545;
w19547 <= not w19543 and not w19546;
w19548 <= not w18860 and not w18867;
w19549 <= not w18887 and w19548;
w19550 <= not w18875 and not w19549;
w19551 <= not w19547 and w19550;
w19552 <= not w19540 and w19551;
w19553 <= w0 and not w19552;
w19554 <= not w19529 and w19547;
w19555 <= not w19539 and w19554;
w19556 <= not w18867 and not w18887;
w19557 <= w18860 and not w19556;
w19558 <= not w0 and not w19548;
w19559 <= not w19557 and w19558;
w19560 <= not w18863 and not w18884;
w19561 <= not w18866 and w19560;
w19562 <= not w18879 and w19561;
w19563 <= not w18875 and w19562;
w19564 <= not w18873 and w19563;
w19565 <= not w19559 and not w19564;
w19566 <= not w19555 and w19565;
w19567 <= not w19553 and w19566;
w19568 <= a(14) and not w19567;
w19569 <= not a(12) and not a(13);
w19570 <= not a(14) and w19569;
w19571 <= not w19568 and not w19570;
w19572 <= not w18887 and not w19571;
w19573 <= not w18884 and not w19570;
w19574 <= not w18879 and w19573;
w19575 <= not w18875 and w19574;
w19576 <= not w18873 and w19575;
w19577 <= not w19568 and w19576;
w19578 <= not a(14) and not w19567;
w19579 <= a(15) and not w19578;
w19580 <= w18889 and not w19567;
w19581 <= not w19579 and not w19580;
w19582 <= not w19577 and w19581;
w19583 <= not w19572 and not w19582;
w19584 <= not w18219 and not w19583;
w19585 <= w18219 and not w19572;
w19586 <= not w19582 and w19585;
w19587 <= not w18887 and not w19564;
w19588 <= not w19559 and w19587;
w19589 <= not w19555 and w19588;
w19590 <= not w19553 and w19589;
w19591 <= not w19580 and not w19590;
w19592 <= a(16) and not w19591;
w19593 <= not a(16) and not w19590;
w19594 <= not w19580 and w19593;
w19595 <= not w19592 and not w19594;
w19596 <= not w19586 and not w19595;
w19597 <= not w19584 and not w19596;
w19598 <= not w17563 and not w19597;
w19599 <= not w18892 and not w18897;
w19600 <= not w18901 and w19599;
w19601 <= not w19567 and w19600;
w19602 <= not w19567 and w19599;
w19603 <= w18901 and not w19602;
w19604 <= not w19601 and not w19603;
w19605 <= w17563 and not w19584;
w19606 <= not w19596 and w19605;
w19607 <= not w19604 and not w19606;
w19608 <= not w19598 and not w19607;
w19609 <= not w16919 and not w19608;
w19610 <= not w18906 and w18915;
w19611 <= not w18904 and w19610;
w19612 <= not w19567 and w19611;
w19613 <= not w18904 and not w18906;
w19614 <= not w19567 and w19613;
w19615 <= not w18915 and not w19614;
w19616 <= not w19612 and not w19615;
w19617 <= w16919 and not w19598;
w19618 <= not w19607 and w19617;
w19619 <= not w19616 and not w19618;
w19620 <= not w19609 and not w19619;
w19621 <= not w16287 and not w19620;
w19622 <= not w18918 and w18924;
w19623 <= not w18926 and w19622;
w19624 <= not w19567 and w19623;
w19625 <= not w18918 and not w18926;
w19626 <= not w19567 and w19625;
w19627 <= not w18924 and not w19626;
w19628 <= not w19624 and not w19627;
w19629 <= w16287 and not w19609;
w19630 <= not w19619 and w19629;
w19631 <= not w19628 and not w19630;
w19632 <= not w19621 and not w19631;
w19633 <= not w15667 and not w19632;
w19634 <= w18936 and not w18938;
w19635 <= not w18929 and w19634;
w19636 <= not w19567 and w19635;
w19637 <= not w18929 and not w18938;
w19638 <= not w19567 and w19637;
w19639 <= not w18936 and not w19638;
w19640 <= not w19636 and not w19639;
w19641 <= w15667 and not w19621;
w19642 <= not w19631 and w19641;
w19643 <= not w19640 and not w19642;
w19644 <= not w19633 and not w19643;
w19645 <= not w15059 and not w19644;
w19646 <= not w18941 and w18948;
w19647 <= not w18950 and w19646;
w19648 <= not w19567 and w19647;
w19649 <= not w18941 and not w18950;
w19650 <= not w19567 and w19649;
w19651 <= not w18948 and not w19650;
w19652 <= not w19648 and not w19651;
w19653 <= w15059 and not w19633;
w19654 <= not w19643 and w19653;
w19655 <= not w19652 and not w19654;
w19656 <= not w19645 and not w19655;
w19657 <= not w14463 and not w19656;
w19658 <= w18960 and not w18962;
w19659 <= not w18953 and w19658;
w19660 <= not w19567 and w19659;
w19661 <= not w18953 and not w18962;
w19662 <= not w19567 and w19661;
w19663 <= not w18960 and not w19662;
w19664 <= not w19660 and not w19663;
w19665 <= w14463 and not w19645;
w19666 <= not w19655 and w19665;
w19667 <= not w19664 and not w19666;
w19668 <= not w19657 and not w19667;
w19669 <= not w13879 and not w19668;
w19670 <= not w18965 and w18972;
w19671 <= not w18974 and w19670;
w19672 <= not w19567 and w19671;
w19673 <= not w18965 and not w18974;
w19674 <= not w19567 and w19673;
w19675 <= not w18972 and not w19674;
w19676 <= not w19672 and not w19675;
w19677 <= w13879 and not w19657;
w19678 <= not w19667 and w19677;
w19679 <= not w19676 and not w19678;
w19680 <= not w19669 and not w19679;
w19681 <= not w13307 and not w19680;
w19682 <= w18984 and not w18986;
w19683 <= not w18977 and w19682;
w19684 <= not w19567 and w19683;
w19685 <= not w18977 and not w18986;
w19686 <= not w19567 and w19685;
w19687 <= not w18984 and not w19686;
w19688 <= not w19684 and not w19687;
w19689 <= w13307 and not w19669;
w19690 <= not w19679 and w19689;
w19691 <= not w19688 and not w19690;
w19692 <= not w19681 and not w19691;
w19693 <= not w12747 and not w19692;
w19694 <= not w18989 and w18996;
w19695 <= not w18998 and w19694;
w19696 <= not w19567 and w19695;
w19697 <= not w18989 and not w18998;
w19698 <= not w19567 and w19697;
w19699 <= not w18996 and not w19698;
w19700 <= not w19696 and not w19699;
w19701 <= w12747 and not w19681;
w19702 <= not w19691 and w19701;
w19703 <= not w19700 and not w19702;
w19704 <= not w19693 and not w19703;
w19705 <= not w12199 and not w19704;
w19706 <= w19008 and not w19010;
w19707 <= not w19001 and w19706;
w19708 <= not w19567 and w19707;
w19709 <= not w19001 and not w19010;
w19710 <= not w19567 and w19709;
w19711 <= not w19008 and not w19710;
w19712 <= not w19708 and not w19711;
w19713 <= w12199 and not w19693;
w19714 <= not w19703 and w19713;
w19715 <= not w19712 and not w19714;
w19716 <= not w19705 and not w19715;
w19717 <= not w11663 and not w19716;
w19718 <= not w19013 and w19020;
w19719 <= not w19022 and w19718;
w19720 <= not w19567 and w19719;
w19721 <= not w19013 and not w19022;
w19722 <= not w19567 and w19721;
w19723 <= not w19020 and not w19722;
w19724 <= not w19720 and not w19723;
w19725 <= w11663 and not w19705;
w19726 <= not w19715 and w19725;
w19727 <= not w19724 and not w19726;
w19728 <= not w19717 and not w19727;
w19729 <= not w11139 and not w19728;
w19730 <= w19032 and not w19034;
w19731 <= not w19025 and w19730;
w19732 <= not w19567 and w19731;
w19733 <= not w19025 and not w19034;
w19734 <= not w19567 and w19733;
w19735 <= not w19032 and not w19734;
w19736 <= not w19732 and not w19735;
w19737 <= w11139 and not w19717;
w19738 <= not w19727 and w19737;
w19739 <= not w19736 and not w19738;
w19740 <= not w19729 and not w19739;
w19741 <= not w10627 and not w19740;
w19742 <= not w19037 and w19044;
w19743 <= not w19046 and w19742;
w19744 <= not w19567 and w19743;
w19745 <= not w19037 and not w19046;
w19746 <= not w19567 and w19745;
w19747 <= not w19044 and not w19746;
w19748 <= not w19744 and not w19747;
w19749 <= w10627 and not w19729;
w19750 <= not w19739 and w19749;
w19751 <= not w19748 and not w19750;
w19752 <= not w19741 and not w19751;
w19753 <= not w10127 and not w19752;
w19754 <= w19056 and not w19058;
w19755 <= not w19049 and w19754;
w19756 <= not w19567 and w19755;
w19757 <= not w19049 and not w19058;
w19758 <= not w19567 and w19757;
w19759 <= not w19056 and not w19758;
w19760 <= not w19756 and not w19759;
w19761 <= w10127 and not w19741;
w19762 <= not w19751 and w19761;
w19763 <= not w19760 and not w19762;
w19764 <= not w19753 and not w19763;
w19765 <= not w9639 and not w19764;
w19766 <= not w19061 and w19068;
w19767 <= not w19070 and w19766;
w19768 <= not w19567 and w19767;
w19769 <= not w19061 and not w19070;
w19770 <= not w19567 and w19769;
w19771 <= not w19068 and not w19770;
w19772 <= not w19768 and not w19771;
w19773 <= w9639 and not w19753;
w19774 <= not w19763 and w19773;
w19775 <= not w19772 and not w19774;
w19776 <= not w19765 and not w19775;
w19777 <= not w9163 and not w19776;
w19778 <= w19080 and not w19082;
w19779 <= not w19073 and w19778;
w19780 <= not w19567 and w19779;
w19781 <= not w19073 and not w19082;
w19782 <= not w19567 and w19781;
w19783 <= not w19080 and not w19782;
w19784 <= not w19780 and not w19783;
w19785 <= w9163 and not w19765;
w19786 <= not w19775 and w19785;
w19787 <= not w19784 and not w19786;
w19788 <= not w19777 and not w19787;
w19789 <= not w8699 and not w19788;
w19790 <= not w19085 and w19092;
w19791 <= not w19094 and w19790;
w19792 <= not w19567 and w19791;
w19793 <= not w19085 and not w19094;
w19794 <= not w19567 and w19793;
w19795 <= not w19092 and not w19794;
w19796 <= not w19792 and not w19795;
w19797 <= w8699 and not w19777;
w19798 <= not w19787 and w19797;
w19799 <= not w19796 and not w19798;
w19800 <= not w19789 and not w19799;
w19801 <= not w8247 and not w19800;
w19802 <= w19104 and not w19106;
w19803 <= not w19097 and w19802;
w19804 <= not w19567 and w19803;
w19805 <= not w19097 and not w19106;
w19806 <= not w19567 and w19805;
w19807 <= not w19104 and not w19806;
w19808 <= not w19804 and not w19807;
w19809 <= w8247 and not w19789;
w19810 <= not w19799 and w19809;
w19811 <= not w19808 and not w19810;
w19812 <= not w19801 and not w19811;
w19813 <= not w7807 and not w19812;
w19814 <= not w19109 and w19116;
w19815 <= not w19118 and w19814;
w19816 <= not w19567 and w19815;
w19817 <= not w19109 and not w19118;
w19818 <= not w19567 and w19817;
w19819 <= not w19116 and not w19818;
w19820 <= not w19816 and not w19819;
w19821 <= w7807 and not w19801;
w19822 <= not w19811 and w19821;
w19823 <= not w19820 and not w19822;
w19824 <= not w19813 and not w19823;
w19825 <= not w7379 and not w19824;
w19826 <= w19128 and not w19130;
w19827 <= not w19121 and w19826;
w19828 <= not w19567 and w19827;
w19829 <= not w19121 and not w19130;
w19830 <= not w19567 and w19829;
w19831 <= not w19128 and not w19830;
w19832 <= not w19828 and not w19831;
w19833 <= w7379 and not w19813;
w19834 <= not w19823 and w19833;
w19835 <= not w19832 and not w19834;
w19836 <= not w19825 and not w19835;
w19837 <= not w6963 and not w19836;
w19838 <= not w19133 and w19140;
w19839 <= not w19142 and w19838;
w19840 <= not w19567 and w19839;
w19841 <= not w19133 and not w19142;
w19842 <= not w19567 and w19841;
w19843 <= not w19140 and not w19842;
w19844 <= not w19840 and not w19843;
w19845 <= w6963 and not w19825;
w19846 <= not w19835 and w19845;
w19847 <= not w19844 and not w19846;
w19848 <= not w19837 and not w19847;
w19849 <= not w6558 and not w19848;
w19850 <= w19152 and not w19154;
w19851 <= not w19145 and w19850;
w19852 <= not w19567 and w19851;
w19853 <= not w19145 and not w19154;
w19854 <= not w19567 and w19853;
w19855 <= not w19152 and not w19854;
w19856 <= not w19852 and not w19855;
w19857 <= w6558 and not w19837;
w19858 <= not w19847 and w19857;
w19859 <= not w19856 and not w19858;
w19860 <= not w19849 and not w19859;
w19861 <= not w6166 and not w19860;
w19862 <= not w19157 and w19164;
w19863 <= not w19166 and w19862;
w19864 <= not w19567 and w19863;
w19865 <= not w19157 and not w19166;
w19866 <= not w19567 and w19865;
w19867 <= not w19164 and not w19866;
w19868 <= not w19864 and not w19867;
w19869 <= w6166 and not w19849;
w19870 <= not w19859 and w19869;
w19871 <= not w19868 and not w19870;
w19872 <= not w19861 and not w19871;
w19873 <= not w5786 and not w19872;
w19874 <= w19176 and not w19178;
w19875 <= not w19169 and w19874;
w19876 <= not w19567 and w19875;
w19877 <= not w19169 and not w19178;
w19878 <= not w19567 and w19877;
w19879 <= not w19176 and not w19878;
w19880 <= not w19876 and not w19879;
w19881 <= w5786 and not w19861;
w19882 <= not w19871 and w19881;
w19883 <= not w19880 and not w19882;
w19884 <= not w19873 and not w19883;
w19885 <= not w5418 and not w19884;
w19886 <= not w19181 and w19188;
w19887 <= not w19190 and w19886;
w19888 <= not w19567 and w19887;
w19889 <= not w19181 and not w19190;
w19890 <= not w19567 and w19889;
w19891 <= not w19188 and not w19890;
w19892 <= not w19888 and not w19891;
w19893 <= w5418 and not w19873;
w19894 <= not w19883 and w19893;
w19895 <= not w19892 and not w19894;
w19896 <= not w19885 and not w19895;
w19897 <= not w5062 and not w19896;
w19898 <= w19200 and not w19202;
w19899 <= not w19193 and w19898;
w19900 <= not w19567 and w19899;
w19901 <= not w19193 and not w19202;
w19902 <= not w19567 and w19901;
w19903 <= not w19200 and not w19902;
w19904 <= not w19900 and not w19903;
w19905 <= w5062 and not w19885;
w19906 <= not w19895 and w19905;
w19907 <= not w19904 and not w19906;
w19908 <= not w19897 and not w19907;
w19909 <= not w4718 and not w19908;
w19910 <= not w19205 and w19212;
w19911 <= not w19214 and w19910;
w19912 <= not w19567 and w19911;
w19913 <= not w19205 and not w19214;
w19914 <= not w19567 and w19913;
w19915 <= not w19212 and not w19914;
w19916 <= not w19912 and not w19915;
w19917 <= w4718 and not w19897;
w19918 <= not w19907 and w19917;
w19919 <= not w19916 and not w19918;
w19920 <= not w19909 and not w19919;
w19921 <= not w4386 and not w19920;
w19922 <= w19224 and not w19226;
w19923 <= not w19217 and w19922;
w19924 <= not w19567 and w19923;
w19925 <= not w19217 and not w19226;
w19926 <= not w19567 and w19925;
w19927 <= not w19224 and not w19926;
w19928 <= not w19924 and not w19927;
w19929 <= w4386 and not w19909;
w19930 <= not w19919 and w19929;
w19931 <= not w19928 and not w19930;
w19932 <= not w19921 and not w19931;
w19933 <= not w4066 and not w19932;
w19934 <= not w19229 and w19236;
w19935 <= not w19238 and w19934;
w19936 <= not w19567 and w19935;
w19937 <= not w19229 and not w19238;
w19938 <= not w19567 and w19937;
w19939 <= not w19236 and not w19938;
w19940 <= not w19936 and not w19939;
w19941 <= w4066 and not w19921;
w19942 <= not w19931 and w19941;
w19943 <= not w19940 and not w19942;
w19944 <= not w19933 and not w19943;
w19945 <= not w3758 and not w19944;
w19946 <= w19248 and not w19250;
w19947 <= not w19241 and w19946;
w19948 <= not w19567 and w19947;
w19949 <= not w19241 and not w19250;
w19950 <= not w19567 and w19949;
w19951 <= not w19248 and not w19950;
w19952 <= not w19948 and not w19951;
w19953 <= w3758 and not w19933;
w19954 <= not w19943 and w19953;
w19955 <= not w19952 and not w19954;
w19956 <= not w19945 and not w19955;
w19957 <= not w3462 and not w19956;
w19958 <= not w19253 and w19260;
w19959 <= not w19262 and w19958;
w19960 <= not w19567 and w19959;
w19961 <= not w19253 and not w19262;
w19962 <= not w19567 and w19961;
w19963 <= not w19260 and not w19962;
w19964 <= not w19960 and not w19963;
w19965 <= w3462 and not w19945;
w19966 <= not w19955 and w19965;
w19967 <= not w19964 and not w19966;
w19968 <= not w19957 and not w19967;
w19969 <= not w3178 and not w19968;
w19970 <= w19272 and not w19274;
w19971 <= not w19265 and w19970;
w19972 <= not w19567 and w19971;
w19973 <= not w19265 and not w19274;
w19974 <= not w19567 and w19973;
w19975 <= not w19272 and not w19974;
w19976 <= not w19972 and not w19975;
w19977 <= w3178 and not w19957;
w19978 <= not w19967 and w19977;
w19979 <= not w19976 and not w19978;
w19980 <= not w19969 and not w19979;
w19981 <= not w2906 and not w19980;
w19982 <= not w19277 and w19284;
w19983 <= not w19286 and w19982;
w19984 <= not w19567 and w19983;
w19985 <= not w19277 and not w19286;
w19986 <= not w19567 and w19985;
w19987 <= not w19284 and not w19986;
w19988 <= not w19984 and not w19987;
w19989 <= w2906 and not w19969;
w19990 <= not w19979 and w19989;
w19991 <= not w19988 and not w19990;
w19992 <= not w19981 and not w19991;
w19993 <= not w2646 and not w19992;
w19994 <= w19296 and not w19298;
w19995 <= not w19289 and w19994;
w19996 <= not w19567 and w19995;
w19997 <= not w19289 and not w19298;
w19998 <= not w19567 and w19997;
w19999 <= not w19296 and not w19998;
w20000 <= not w19996 and not w19999;
w20001 <= w2646 and not w19981;
w20002 <= not w19991 and w20001;
w20003 <= not w20000 and not w20002;
w20004 <= not w19993 and not w20003;
w20005 <= not w2398 and not w20004;
w20006 <= not w19301 and w19308;
w20007 <= not w19310 and w20006;
w20008 <= not w19567 and w20007;
w20009 <= not w19301 and not w19310;
w20010 <= not w19567 and w20009;
w20011 <= not w19308 and not w20010;
w20012 <= not w20008 and not w20011;
w20013 <= w2398 and not w19993;
w20014 <= not w20003 and w20013;
w20015 <= not w20012 and not w20014;
w20016 <= not w20005 and not w20015;
w20017 <= not w2162 and not w20016;
w20018 <= w19320 and not w19322;
w20019 <= not w19313 and w20018;
w20020 <= not w19567 and w20019;
w20021 <= not w19313 and not w19322;
w20022 <= not w19567 and w20021;
w20023 <= not w19320 and not w20022;
w20024 <= not w20020 and not w20023;
w20025 <= w2162 and not w20005;
w20026 <= not w20015 and w20025;
w20027 <= not w20024 and not w20026;
w20028 <= not w20017 and not w20027;
w20029 <= not w1938 and not w20028;
w20030 <= not w19325 and w19332;
w20031 <= not w19334 and w20030;
w20032 <= not w19567 and w20031;
w20033 <= not w19325 and not w19334;
w20034 <= not w19567 and w20033;
w20035 <= not w19332 and not w20034;
w20036 <= not w20032 and not w20035;
w20037 <= w1938 and not w20017;
w20038 <= not w20027 and w20037;
w20039 <= not w20036 and not w20038;
w20040 <= not w20029 and not w20039;
w20041 <= not w1725 and not w20040;
w20042 <= w19344 and not w19346;
w20043 <= not w19337 and w20042;
w20044 <= not w19567 and w20043;
w20045 <= not w19337 and not w19346;
w20046 <= not w19567 and w20045;
w20047 <= not w19344 and not w20046;
w20048 <= not w20044 and not w20047;
w20049 <= w1725 and not w20029;
w20050 <= not w20039 and w20049;
w20051 <= not w20048 and not w20050;
w20052 <= not w20041 and not w20051;
w20053 <= not w1525 and not w20052;
w20054 <= not w19349 and w19356;
w20055 <= not w19358 and w20054;
w20056 <= not w19567 and w20055;
w20057 <= not w19349 and not w19358;
w20058 <= not w19567 and w20057;
w20059 <= not w19356 and not w20058;
w20060 <= not w20056 and not w20059;
w20061 <= w1525 and not w20041;
w20062 <= not w20051 and w20061;
w20063 <= not w20060 and not w20062;
w20064 <= not w20053 and not w20063;
w20065 <= not w1337 and not w20064;
w20066 <= w19368 and not w19370;
w20067 <= not w19361 and w20066;
w20068 <= not w19567 and w20067;
w20069 <= not w19361 and not w19370;
w20070 <= not w19567 and w20069;
w20071 <= not w19368 and not w20070;
w20072 <= not w20068 and not w20071;
w20073 <= w1337 and not w20053;
w20074 <= not w20063 and w20073;
w20075 <= not w20072 and not w20074;
w20076 <= not w20065 and not w20075;
w20077 <= not w1161 and not w20076;
w20078 <= not w19373 and w19380;
w20079 <= not w19382 and w20078;
w20080 <= not w19567 and w20079;
w20081 <= not w19373 and not w19382;
w20082 <= not w19567 and w20081;
w20083 <= not w19380 and not w20082;
w20084 <= not w20080 and not w20083;
w20085 <= w1161 and not w20065;
w20086 <= not w20075 and w20085;
w20087 <= not w20084 and not w20086;
w20088 <= not w20077 and not w20087;
w20089 <= not w997 and not w20088;
w20090 <= w19392 and not w19394;
w20091 <= not w19385 and w20090;
w20092 <= not w19567 and w20091;
w20093 <= not w19385 and not w19394;
w20094 <= not w19567 and w20093;
w20095 <= not w19392 and not w20094;
w20096 <= not w20092 and not w20095;
w20097 <= w997 and not w20077;
w20098 <= not w20087 and w20097;
w20099 <= not w20096 and not w20098;
w20100 <= not w20089 and not w20099;
w20101 <= not w845 and not w20100;
w20102 <= not w19397 and w19404;
w20103 <= not w19406 and w20102;
w20104 <= not w19567 and w20103;
w20105 <= not w19397 and not w19406;
w20106 <= not w19567 and w20105;
w20107 <= not w19404 and not w20106;
w20108 <= not w20104 and not w20107;
w20109 <= w845 and not w20089;
w20110 <= not w20099 and w20109;
w20111 <= not w20108 and not w20110;
w20112 <= not w20101 and not w20111;
w20113 <= not w705 and not w20112;
w20114 <= w19416 and not w19418;
w20115 <= not w19409 and w20114;
w20116 <= not w19567 and w20115;
w20117 <= not w19409 and not w19418;
w20118 <= not w19567 and w20117;
w20119 <= not w19416 and not w20118;
w20120 <= not w20116 and not w20119;
w20121 <= w705 and not w20101;
w20122 <= not w20111 and w20121;
w20123 <= not w20120 and not w20122;
w20124 <= not w20113 and not w20123;
w20125 <= not w577 and not w20124;
w20126 <= not w19421 and w19428;
w20127 <= not w19430 and w20126;
w20128 <= not w19567 and w20127;
w20129 <= not w19421 and not w19430;
w20130 <= not w19567 and w20129;
w20131 <= not w19428 and not w20130;
w20132 <= not w20128 and not w20131;
w20133 <= w577 and not w20113;
w20134 <= not w20123 and w20133;
w20135 <= not w20132 and not w20134;
w20136 <= not w20125 and not w20135;
w20137 <= not w460 and not w20136;
w20138 <= w19440 and not w19442;
w20139 <= not w19433 and w20138;
w20140 <= not w19567 and w20139;
w20141 <= not w19433 and not w19442;
w20142 <= not w19567 and w20141;
w20143 <= not w19440 and not w20142;
w20144 <= not w20140 and not w20143;
w20145 <= w460 and not w20125;
w20146 <= not w20135 and w20145;
w20147 <= not w20144 and not w20146;
w20148 <= not w20137 and not w20147;
w20149 <= not w356 and not w20148;
w20150 <= not w19445 and w19452;
w20151 <= not w19454 and w20150;
w20152 <= not w19567 and w20151;
w20153 <= not w19445 and not w19454;
w20154 <= not w19567 and w20153;
w20155 <= not w19452 and not w20154;
w20156 <= not w20152 and not w20155;
w20157 <= w356 and not w20137;
w20158 <= not w20147 and w20157;
w20159 <= not w20156 and not w20158;
w20160 <= not w20149 and not w20159;
w20161 <= not w264 and not w20160;
w20162 <= w19464 and not w19466;
w20163 <= not w19457 and w20162;
w20164 <= not w19567 and w20163;
w20165 <= not w19457 and not w19466;
w20166 <= not w19567 and w20165;
w20167 <= not w19464 and not w20166;
w20168 <= not w20164 and not w20167;
w20169 <= w264 and not w20149;
w20170 <= not w20159 and w20169;
w20171 <= not w20168 and not w20170;
w20172 <= not w20161 and not w20171;
w20173 <= not w184 and not w20172;
w20174 <= w184 and not w20161;
w20175 <= not w20171 and w20174;
w20176 <= not w19469 and w19478;
w20177 <= not w19471 and w20176;
w20178 <= not w19567 and w20177;
w20179 <= not w19469 and not w19471;
w20180 <= not w19567 and w20179;
w20181 <= not w19478 and not w20180;
w20182 <= not w20178 and not w20181;
w20183 <= not w20175 and not w20182;
w20184 <= not w20173 and not w20183;
w20185 <= not w115 and not w20184;
w20186 <= w19488 and not w19490;
w20187 <= not w19481 and w20186;
w20188 <= not w19567 and w20187;
w20189 <= not w19481 and not w19490;
w20190 <= not w19567 and w20189;
w20191 <= not w19488 and not w20190;
w20192 <= not w20188 and not w20191;
w20193 <= w115 and not w20173;
w20194 <= not w20183 and w20193;
w20195 <= not w20192 and not w20194;
w20196 <= not w20185 and not w20195;
w20197 <= not w60 and not w20196;
w20198 <= not w19493 and w19500;
w20199 <= not w19502 and w20198;
w20200 <= not w19567 and w20199;
w20201 <= not w19493 and not w19502;
w20202 <= not w19567 and w20201;
w20203 <= not w19500 and not w20202;
w20204 <= not w20200 and not w20203;
w20205 <= w60 and not w20185;
w20206 <= not w20195 and w20205;
w20207 <= not w20204 and not w20206;
w20208 <= not w20197 and not w20207;
w20209 <= not w22 and not w20208;
w20210 <= w19512 and not w19514;
w20211 <= not w19505 and w20210;
w20212 <= not w19567 and w20211;
w20213 <= not w19505 and not w19514;
w20214 <= not w19567 and w20213;
w20215 <= not w19512 and not w20214;
w20216 <= not w20212 and not w20215;
w20217 <= w22 and not w20197;
w20218 <= not w20207 and w20217;
w20219 <= not w20216 and not w20218;
w20220 <= not w20209 and not w20219;
w20221 <= not w5 and not w20220;
w20222 <= not w19517 and w19524;
w20223 <= not w19526 and w20222;
w20224 <= not w19567 and w20223;
w20225 <= not w19517 and not w19526;
w20226 <= not w19567 and w20225;
w20227 <= not w19524 and not w20226;
w20228 <= not w20224 and not w20227;
w20229 <= w5 and not w20209;
w20230 <= not w20219 and w20229;
w20231 <= not w20228 and not w20230;
w20232 <= not w20221 and not w20231;
w20233 <= w19536 and not w19538;
w20234 <= not w19529 and w20233;
w20235 <= not w19567 and w20234;
w20236 <= not w19529 and not w19538;
w20237 <= not w19567 and w20236;
w20238 <= not w19536 and not w20237;
w20239 <= not w20235 and not w20238;
w20240 <= not w19540 and not w19547;
w20241 <= not w19567 and w20240;
w20242 <= not w19555 and not w20241;
w20243 <= not w20239 and w20242;
w20244 <= not w20232 and w20243;
w20245 <= w0 and not w20244;
w20246 <= not w20221 and w20239;
w20247 <= not w20231 and w20246;
w20248 <= not w19547 and not w19567;
w20249 <= w19540 and not w20248;
w20250 <= not w0 and not w20240;
w20251 <= not w20249 and w20250;
w20252 <= not w19543 and not w19564;
w20253 <= not w19546 and w20252;
w20254 <= not w19559 and w20253;
w20255 <= not w19555 and w20254;
w20256 <= not w19553 and w20255;
w20257 <= not w20251 and not w20256;
w20258 <= not w20247 and w20257;
w20259 <= not w20245 and w20258;
w20260 <= a(12) and not w20259;
w20261 <= not a(10) and not a(11);
w20262 <= not a(12) and w20261;
w20263 <= not w20260 and not w20262;
w20264 <= not w19567 and not w20263;
w20265 <= not w19564 and not w20262;
w20266 <= not w19559 and w20265;
w20267 <= not w19555 and w20266;
w20268 <= not w19553 and w20267;
w20269 <= not w20260 and w20268;
w20270 <= not a(12) and not w20259;
w20271 <= a(13) and not w20270;
w20272 <= w19569 and not w20259;
w20273 <= not w20271 and not w20272;
w20274 <= not w20269 and w20273;
w20275 <= not w20264 and not w20274;
w20276 <= not w18887 and not w20275;
w20277 <= w18887 and not w20264;
w20278 <= not w20274 and w20277;
w20279 <= not w19567 and not w20256;
w20280 <= not w20251 and w20279;
w20281 <= not w20247 and w20280;
w20282 <= not w20245 and w20281;
w20283 <= not w20272 and not w20282;
w20284 <= a(14) and not w20283;
w20285 <= not a(14) and not w20282;
w20286 <= not w20272 and w20285;
w20287 <= not w20284 and not w20286;
w20288 <= not w20278 and not w20287;
w20289 <= not w20276 and not w20288;
w20290 <= not w18219 and not w20289;
w20291 <= not w19572 and not w19577;
w20292 <= not w19581 and w20291;
w20293 <= not w20259 and w20292;
w20294 <= not w20259 and w20291;
w20295 <= w19581 and not w20294;
w20296 <= not w20293 and not w20295;
w20297 <= w18219 and not w20276;
w20298 <= not w20288 and w20297;
w20299 <= not w20296 and not w20298;
w20300 <= not w20290 and not w20299;
w20301 <= not w17563 and not w20300;
w20302 <= not w19586 and w19595;
w20303 <= not w19584 and w20302;
w20304 <= not w20259 and w20303;
w20305 <= not w19584 and not w19586;
w20306 <= not w20259 and w20305;
w20307 <= not w19595 and not w20306;
w20308 <= not w20304 and not w20307;
w20309 <= w17563 and not w20290;
w20310 <= not w20299 and w20309;
w20311 <= not w20308 and not w20310;
w20312 <= not w20301 and not w20311;
w20313 <= not w16919 and not w20312;
w20314 <= not w19598 and w19604;
w20315 <= not w19606 and w20314;
w20316 <= not w20259 and w20315;
w20317 <= not w19598 and not w19606;
w20318 <= not w20259 and w20317;
w20319 <= not w19604 and not w20318;
w20320 <= not w20316 and not w20319;
w20321 <= w16919 and not w20301;
w20322 <= not w20311 and w20321;
w20323 <= not w20320 and not w20322;
w20324 <= not w20313 and not w20323;
w20325 <= not w16287 and not w20324;
w20326 <= w19616 and not w19618;
w20327 <= not w19609 and w20326;
w20328 <= not w20259 and w20327;
w20329 <= not w19609 and not w19618;
w20330 <= not w20259 and w20329;
w20331 <= not w19616 and not w20330;
w20332 <= not w20328 and not w20331;
w20333 <= w16287 and not w20313;
w20334 <= not w20323 and w20333;
w20335 <= not w20332 and not w20334;
w20336 <= not w20325 and not w20335;
w20337 <= not w15667 and not w20336;
w20338 <= not w19621 and w19628;
w20339 <= not w19630 and w20338;
w20340 <= not w20259 and w20339;
w20341 <= not w19621 and not w19630;
w20342 <= not w20259 and w20341;
w20343 <= not w19628 and not w20342;
w20344 <= not w20340 and not w20343;
w20345 <= w15667 and not w20325;
w20346 <= not w20335 and w20345;
w20347 <= not w20344 and not w20346;
w20348 <= not w20337 and not w20347;
w20349 <= not w15059 and not w20348;
w20350 <= w19640 and not w19642;
w20351 <= not w19633 and w20350;
w20352 <= not w20259 and w20351;
w20353 <= not w19633 and not w19642;
w20354 <= not w20259 and w20353;
w20355 <= not w19640 and not w20354;
w20356 <= not w20352 and not w20355;
w20357 <= w15059 and not w20337;
w20358 <= not w20347 and w20357;
w20359 <= not w20356 and not w20358;
w20360 <= not w20349 and not w20359;
w20361 <= not w14463 and not w20360;
w20362 <= not w19645 and w19652;
w20363 <= not w19654 and w20362;
w20364 <= not w20259 and w20363;
w20365 <= not w19645 and not w19654;
w20366 <= not w20259 and w20365;
w20367 <= not w19652 and not w20366;
w20368 <= not w20364 and not w20367;
w20369 <= w14463 and not w20349;
w20370 <= not w20359 and w20369;
w20371 <= not w20368 and not w20370;
w20372 <= not w20361 and not w20371;
w20373 <= not w13879 and not w20372;
w20374 <= w19664 and not w19666;
w20375 <= not w19657 and w20374;
w20376 <= not w20259 and w20375;
w20377 <= not w19657 and not w19666;
w20378 <= not w20259 and w20377;
w20379 <= not w19664 and not w20378;
w20380 <= not w20376 and not w20379;
w20381 <= w13879 and not w20361;
w20382 <= not w20371 and w20381;
w20383 <= not w20380 and not w20382;
w20384 <= not w20373 and not w20383;
w20385 <= not w13307 and not w20384;
w20386 <= not w19669 and w19676;
w20387 <= not w19678 and w20386;
w20388 <= not w20259 and w20387;
w20389 <= not w19669 and not w19678;
w20390 <= not w20259 and w20389;
w20391 <= not w19676 and not w20390;
w20392 <= not w20388 and not w20391;
w20393 <= w13307 and not w20373;
w20394 <= not w20383 and w20393;
w20395 <= not w20392 and not w20394;
w20396 <= not w20385 and not w20395;
w20397 <= not w12747 and not w20396;
w20398 <= w19688 and not w19690;
w20399 <= not w19681 and w20398;
w20400 <= not w20259 and w20399;
w20401 <= not w19681 and not w19690;
w20402 <= not w20259 and w20401;
w20403 <= not w19688 and not w20402;
w20404 <= not w20400 and not w20403;
w20405 <= w12747 and not w20385;
w20406 <= not w20395 and w20405;
w20407 <= not w20404 and not w20406;
w20408 <= not w20397 and not w20407;
w20409 <= not w12199 and not w20408;
w20410 <= not w19693 and w19700;
w20411 <= not w19702 and w20410;
w20412 <= not w20259 and w20411;
w20413 <= not w19693 and not w19702;
w20414 <= not w20259 and w20413;
w20415 <= not w19700 and not w20414;
w20416 <= not w20412 and not w20415;
w20417 <= w12199 and not w20397;
w20418 <= not w20407 and w20417;
w20419 <= not w20416 and not w20418;
w20420 <= not w20409 and not w20419;
w20421 <= not w11663 and not w20420;
w20422 <= w19712 and not w19714;
w20423 <= not w19705 and w20422;
w20424 <= not w20259 and w20423;
w20425 <= not w19705 and not w19714;
w20426 <= not w20259 and w20425;
w20427 <= not w19712 and not w20426;
w20428 <= not w20424 and not w20427;
w20429 <= w11663 and not w20409;
w20430 <= not w20419 and w20429;
w20431 <= not w20428 and not w20430;
w20432 <= not w20421 and not w20431;
w20433 <= not w11139 and not w20432;
w20434 <= not w19717 and w19724;
w20435 <= not w19726 and w20434;
w20436 <= not w20259 and w20435;
w20437 <= not w19717 and not w19726;
w20438 <= not w20259 and w20437;
w20439 <= not w19724 and not w20438;
w20440 <= not w20436 and not w20439;
w20441 <= w11139 and not w20421;
w20442 <= not w20431 and w20441;
w20443 <= not w20440 and not w20442;
w20444 <= not w20433 and not w20443;
w20445 <= not w10627 and not w20444;
w20446 <= w19736 and not w19738;
w20447 <= not w19729 and w20446;
w20448 <= not w20259 and w20447;
w20449 <= not w19729 and not w19738;
w20450 <= not w20259 and w20449;
w20451 <= not w19736 and not w20450;
w20452 <= not w20448 and not w20451;
w20453 <= w10627 and not w20433;
w20454 <= not w20443 and w20453;
w20455 <= not w20452 and not w20454;
w20456 <= not w20445 and not w20455;
w20457 <= not w10127 and not w20456;
w20458 <= not w19741 and w19748;
w20459 <= not w19750 and w20458;
w20460 <= not w20259 and w20459;
w20461 <= not w19741 and not w19750;
w20462 <= not w20259 and w20461;
w20463 <= not w19748 and not w20462;
w20464 <= not w20460 and not w20463;
w20465 <= w10127 and not w20445;
w20466 <= not w20455 and w20465;
w20467 <= not w20464 and not w20466;
w20468 <= not w20457 and not w20467;
w20469 <= not w9639 and not w20468;
w20470 <= w19760 and not w19762;
w20471 <= not w19753 and w20470;
w20472 <= not w20259 and w20471;
w20473 <= not w19753 and not w19762;
w20474 <= not w20259 and w20473;
w20475 <= not w19760 and not w20474;
w20476 <= not w20472 and not w20475;
w20477 <= w9639 and not w20457;
w20478 <= not w20467 and w20477;
w20479 <= not w20476 and not w20478;
w20480 <= not w20469 and not w20479;
w20481 <= not w9163 and not w20480;
w20482 <= not w19765 and w19772;
w20483 <= not w19774 and w20482;
w20484 <= not w20259 and w20483;
w20485 <= not w19765 and not w19774;
w20486 <= not w20259 and w20485;
w20487 <= not w19772 and not w20486;
w20488 <= not w20484 and not w20487;
w20489 <= w9163 and not w20469;
w20490 <= not w20479 and w20489;
w20491 <= not w20488 and not w20490;
w20492 <= not w20481 and not w20491;
w20493 <= not w8699 and not w20492;
w20494 <= w19784 and not w19786;
w20495 <= not w19777 and w20494;
w20496 <= not w20259 and w20495;
w20497 <= not w19777 and not w19786;
w20498 <= not w20259 and w20497;
w20499 <= not w19784 and not w20498;
w20500 <= not w20496 and not w20499;
w20501 <= w8699 and not w20481;
w20502 <= not w20491 and w20501;
w20503 <= not w20500 and not w20502;
w20504 <= not w20493 and not w20503;
w20505 <= not w8247 and not w20504;
w20506 <= not w19789 and w19796;
w20507 <= not w19798 and w20506;
w20508 <= not w20259 and w20507;
w20509 <= not w19789 and not w19798;
w20510 <= not w20259 and w20509;
w20511 <= not w19796 and not w20510;
w20512 <= not w20508 and not w20511;
w20513 <= w8247 and not w20493;
w20514 <= not w20503 and w20513;
w20515 <= not w20512 and not w20514;
w20516 <= not w20505 and not w20515;
w20517 <= not w7807 and not w20516;
w20518 <= w19808 and not w19810;
w20519 <= not w19801 and w20518;
w20520 <= not w20259 and w20519;
w20521 <= not w19801 and not w19810;
w20522 <= not w20259 and w20521;
w20523 <= not w19808 and not w20522;
w20524 <= not w20520 and not w20523;
w20525 <= w7807 and not w20505;
w20526 <= not w20515 and w20525;
w20527 <= not w20524 and not w20526;
w20528 <= not w20517 and not w20527;
w20529 <= not w7379 and not w20528;
w20530 <= not w19813 and w19820;
w20531 <= not w19822 and w20530;
w20532 <= not w20259 and w20531;
w20533 <= not w19813 and not w19822;
w20534 <= not w20259 and w20533;
w20535 <= not w19820 and not w20534;
w20536 <= not w20532 and not w20535;
w20537 <= w7379 and not w20517;
w20538 <= not w20527 and w20537;
w20539 <= not w20536 and not w20538;
w20540 <= not w20529 and not w20539;
w20541 <= not w6963 and not w20540;
w20542 <= w19832 and not w19834;
w20543 <= not w19825 and w20542;
w20544 <= not w20259 and w20543;
w20545 <= not w19825 and not w19834;
w20546 <= not w20259 and w20545;
w20547 <= not w19832 and not w20546;
w20548 <= not w20544 and not w20547;
w20549 <= w6963 and not w20529;
w20550 <= not w20539 and w20549;
w20551 <= not w20548 and not w20550;
w20552 <= not w20541 and not w20551;
w20553 <= not w6558 and not w20552;
w20554 <= not w19837 and w19844;
w20555 <= not w19846 and w20554;
w20556 <= not w20259 and w20555;
w20557 <= not w19837 and not w19846;
w20558 <= not w20259 and w20557;
w20559 <= not w19844 and not w20558;
w20560 <= not w20556 and not w20559;
w20561 <= w6558 and not w20541;
w20562 <= not w20551 and w20561;
w20563 <= not w20560 and not w20562;
w20564 <= not w20553 and not w20563;
w20565 <= not w6166 and not w20564;
w20566 <= w19856 and not w19858;
w20567 <= not w19849 and w20566;
w20568 <= not w20259 and w20567;
w20569 <= not w19849 and not w19858;
w20570 <= not w20259 and w20569;
w20571 <= not w19856 and not w20570;
w20572 <= not w20568 and not w20571;
w20573 <= w6166 and not w20553;
w20574 <= not w20563 and w20573;
w20575 <= not w20572 and not w20574;
w20576 <= not w20565 and not w20575;
w20577 <= not w5786 and not w20576;
w20578 <= not w19861 and w19868;
w20579 <= not w19870 and w20578;
w20580 <= not w20259 and w20579;
w20581 <= not w19861 and not w19870;
w20582 <= not w20259 and w20581;
w20583 <= not w19868 and not w20582;
w20584 <= not w20580 and not w20583;
w20585 <= w5786 and not w20565;
w20586 <= not w20575 and w20585;
w20587 <= not w20584 and not w20586;
w20588 <= not w20577 and not w20587;
w20589 <= not w5418 and not w20588;
w20590 <= w19880 and not w19882;
w20591 <= not w19873 and w20590;
w20592 <= not w20259 and w20591;
w20593 <= not w19873 and not w19882;
w20594 <= not w20259 and w20593;
w20595 <= not w19880 and not w20594;
w20596 <= not w20592 and not w20595;
w20597 <= w5418 and not w20577;
w20598 <= not w20587 and w20597;
w20599 <= not w20596 and not w20598;
w20600 <= not w20589 and not w20599;
w20601 <= not w5062 and not w20600;
w20602 <= not w19885 and w19892;
w20603 <= not w19894 and w20602;
w20604 <= not w20259 and w20603;
w20605 <= not w19885 and not w19894;
w20606 <= not w20259 and w20605;
w20607 <= not w19892 and not w20606;
w20608 <= not w20604 and not w20607;
w20609 <= w5062 and not w20589;
w20610 <= not w20599 and w20609;
w20611 <= not w20608 and not w20610;
w20612 <= not w20601 and not w20611;
w20613 <= not w4718 and not w20612;
w20614 <= w19904 and not w19906;
w20615 <= not w19897 and w20614;
w20616 <= not w20259 and w20615;
w20617 <= not w19897 and not w19906;
w20618 <= not w20259 and w20617;
w20619 <= not w19904 and not w20618;
w20620 <= not w20616 and not w20619;
w20621 <= w4718 and not w20601;
w20622 <= not w20611 and w20621;
w20623 <= not w20620 and not w20622;
w20624 <= not w20613 and not w20623;
w20625 <= not w4386 and not w20624;
w20626 <= not w19909 and w19916;
w20627 <= not w19918 and w20626;
w20628 <= not w20259 and w20627;
w20629 <= not w19909 and not w19918;
w20630 <= not w20259 and w20629;
w20631 <= not w19916 and not w20630;
w20632 <= not w20628 and not w20631;
w20633 <= w4386 and not w20613;
w20634 <= not w20623 and w20633;
w20635 <= not w20632 and not w20634;
w20636 <= not w20625 and not w20635;
w20637 <= not w4066 and not w20636;
w20638 <= w19928 and not w19930;
w20639 <= not w19921 and w20638;
w20640 <= not w20259 and w20639;
w20641 <= not w19921 and not w19930;
w20642 <= not w20259 and w20641;
w20643 <= not w19928 and not w20642;
w20644 <= not w20640 and not w20643;
w20645 <= w4066 and not w20625;
w20646 <= not w20635 and w20645;
w20647 <= not w20644 and not w20646;
w20648 <= not w20637 and not w20647;
w20649 <= not w3758 and not w20648;
w20650 <= not w19933 and w19940;
w20651 <= not w19942 and w20650;
w20652 <= not w20259 and w20651;
w20653 <= not w19933 and not w19942;
w20654 <= not w20259 and w20653;
w20655 <= not w19940 and not w20654;
w20656 <= not w20652 and not w20655;
w20657 <= w3758 and not w20637;
w20658 <= not w20647 and w20657;
w20659 <= not w20656 and not w20658;
w20660 <= not w20649 and not w20659;
w20661 <= not w3462 and not w20660;
w20662 <= w19952 and not w19954;
w20663 <= not w19945 and w20662;
w20664 <= not w20259 and w20663;
w20665 <= not w19945 and not w19954;
w20666 <= not w20259 and w20665;
w20667 <= not w19952 and not w20666;
w20668 <= not w20664 and not w20667;
w20669 <= w3462 and not w20649;
w20670 <= not w20659 and w20669;
w20671 <= not w20668 and not w20670;
w20672 <= not w20661 and not w20671;
w20673 <= not w3178 and not w20672;
w20674 <= not w19957 and w19964;
w20675 <= not w19966 and w20674;
w20676 <= not w20259 and w20675;
w20677 <= not w19957 and not w19966;
w20678 <= not w20259 and w20677;
w20679 <= not w19964 and not w20678;
w20680 <= not w20676 and not w20679;
w20681 <= w3178 and not w20661;
w20682 <= not w20671 and w20681;
w20683 <= not w20680 and not w20682;
w20684 <= not w20673 and not w20683;
w20685 <= not w2906 and not w20684;
w20686 <= w19976 and not w19978;
w20687 <= not w19969 and w20686;
w20688 <= not w20259 and w20687;
w20689 <= not w19969 and not w19978;
w20690 <= not w20259 and w20689;
w20691 <= not w19976 and not w20690;
w20692 <= not w20688 and not w20691;
w20693 <= w2906 and not w20673;
w20694 <= not w20683 and w20693;
w20695 <= not w20692 and not w20694;
w20696 <= not w20685 and not w20695;
w20697 <= not w2646 and not w20696;
w20698 <= not w19981 and w19988;
w20699 <= not w19990 and w20698;
w20700 <= not w20259 and w20699;
w20701 <= not w19981 and not w19990;
w20702 <= not w20259 and w20701;
w20703 <= not w19988 and not w20702;
w20704 <= not w20700 and not w20703;
w20705 <= w2646 and not w20685;
w20706 <= not w20695 and w20705;
w20707 <= not w20704 and not w20706;
w20708 <= not w20697 and not w20707;
w20709 <= not w2398 and not w20708;
w20710 <= w20000 and not w20002;
w20711 <= not w19993 and w20710;
w20712 <= not w20259 and w20711;
w20713 <= not w19993 and not w20002;
w20714 <= not w20259 and w20713;
w20715 <= not w20000 and not w20714;
w20716 <= not w20712 and not w20715;
w20717 <= w2398 and not w20697;
w20718 <= not w20707 and w20717;
w20719 <= not w20716 and not w20718;
w20720 <= not w20709 and not w20719;
w20721 <= not w2162 and not w20720;
w20722 <= not w20005 and w20012;
w20723 <= not w20014 and w20722;
w20724 <= not w20259 and w20723;
w20725 <= not w20005 and not w20014;
w20726 <= not w20259 and w20725;
w20727 <= not w20012 and not w20726;
w20728 <= not w20724 and not w20727;
w20729 <= w2162 and not w20709;
w20730 <= not w20719 and w20729;
w20731 <= not w20728 and not w20730;
w20732 <= not w20721 and not w20731;
w20733 <= not w1938 and not w20732;
w20734 <= w20024 and not w20026;
w20735 <= not w20017 and w20734;
w20736 <= not w20259 and w20735;
w20737 <= not w20017 and not w20026;
w20738 <= not w20259 and w20737;
w20739 <= not w20024 and not w20738;
w20740 <= not w20736 and not w20739;
w20741 <= w1938 and not w20721;
w20742 <= not w20731 and w20741;
w20743 <= not w20740 and not w20742;
w20744 <= not w20733 and not w20743;
w20745 <= not w1725 and not w20744;
w20746 <= not w20029 and w20036;
w20747 <= not w20038 and w20746;
w20748 <= not w20259 and w20747;
w20749 <= not w20029 and not w20038;
w20750 <= not w20259 and w20749;
w20751 <= not w20036 and not w20750;
w20752 <= not w20748 and not w20751;
w20753 <= w1725 and not w20733;
w20754 <= not w20743 and w20753;
w20755 <= not w20752 and not w20754;
w20756 <= not w20745 and not w20755;
w20757 <= not w1525 and not w20756;
w20758 <= w20048 and not w20050;
w20759 <= not w20041 and w20758;
w20760 <= not w20259 and w20759;
w20761 <= not w20041 and not w20050;
w20762 <= not w20259 and w20761;
w20763 <= not w20048 and not w20762;
w20764 <= not w20760 and not w20763;
w20765 <= w1525 and not w20745;
w20766 <= not w20755 and w20765;
w20767 <= not w20764 and not w20766;
w20768 <= not w20757 and not w20767;
w20769 <= not w1337 and not w20768;
w20770 <= not w20053 and w20060;
w20771 <= not w20062 and w20770;
w20772 <= not w20259 and w20771;
w20773 <= not w20053 and not w20062;
w20774 <= not w20259 and w20773;
w20775 <= not w20060 and not w20774;
w20776 <= not w20772 and not w20775;
w20777 <= w1337 and not w20757;
w20778 <= not w20767 and w20777;
w20779 <= not w20776 and not w20778;
w20780 <= not w20769 and not w20779;
w20781 <= not w1161 and not w20780;
w20782 <= w20072 and not w20074;
w20783 <= not w20065 and w20782;
w20784 <= not w20259 and w20783;
w20785 <= not w20065 and not w20074;
w20786 <= not w20259 and w20785;
w20787 <= not w20072 and not w20786;
w20788 <= not w20784 and not w20787;
w20789 <= w1161 and not w20769;
w20790 <= not w20779 and w20789;
w20791 <= not w20788 and not w20790;
w20792 <= not w20781 and not w20791;
w20793 <= not w997 and not w20792;
w20794 <= not w20077 and w20084;
w20795 <= not w20086 and w20794;
w20796 <= not w20259 and w20795;
w20797 <= not w20077 and not w20086;
w20798 <= not w20259 and w20797;
w20799 <= not w20084 and not w20798;
w20800 <= not w20796 and not w20799;
w20801 <= w997 and not w20781;
w20802 <= not w20791 and w20801;
w20803 <= not w20800 and not w20802;
w20804 <= not w20793 and not w20803;
w20805 <= not w845 and not w20804;
w20806 <= w20096 and not w20098;
w20807 <= not w20089 and w20806;
w20808 <= not w20259 and w20807;
w20809 <= not w20089 and not w20098;
w20810 <= not w20259 and w20809;
w20811 <= not w20096 and not w20810;
w20812 <= not w20808 and not w20811;
w20813 <= w845 and not w20793;
w20814 <= not w20803 and w20813;
w20815 <= not w20812 and not w20814;
w20816 <= not w20805 and not w20815;
w20817 <= not w705 and not w20816;
w20818 <= not w20101 and w20108;
w20819 <= not w20110 and w20818;
w20820 <= not w20259 and w20819;
w20821 <= not w20101 and not w20110;
w20822 <= not w20259 and w20821;
w20823 <= not w20108 and not w20822;
w20824 <= not w20820 and not w20823;
w20825 <= w705 and not w20805;
w20826 <= not w20815 and w20825;
w20827 <= not w20824 and not w20826;
w20828 <= not w20817 and not w20827;
w20829 <= not w577 and not w20828;
w20830 <= w20120 and not w20122;
w20831 <= not w20113 and w20830;
w20832 <= not w20259 and w20831;
w20833 <= not w20113 and not w20122;
w20834 <= not w20259 and w20833;
w20835 <= not w20120 and not w20834;
w20836 <= not w20832 and not w20835;
w20837 <= w577 and not w20817;
w20838 <= not w20827 and w20837;
w20839 <= not w20836 and not w20838;
w20840 <= not w20829 and not w20839;
w20841 <= not w460 and not w20840;
w20842 <= not w20125 and w20132;
w20843 <= not w20134 and w20842;
w20844 <= not w20259 and w20843;
w20845 <= not w20125 and not w20134;
w20846 <= not w20259 and w20845;
w20847 <= not w20132 and not w20846;
w20848 <= not w20844 and not w20847;
w20849 <= w460 and not w20829;
w20850 <= not w20839 and w20849;
w20851 <= not w20848 and not w20850;
w20852 <= not w20841 and not w20851;
w20853 <= not w356 and not w20852;
w20854 <= w20144 and not w20146;
w20855 <= not w20137 and w20854;
w20856 <= not w20259 and w20855;
w20857 <= not w20137 and not w20146;
w20858 <= not w20259 and w20857;
w20859 <= not w20144 and not w20858;
w20860 <= not w20856 and not w20859;
w20861 <= w356 and not w20841;
w20862 <= not w20851 and w20861;
w20863 <= not w20860 and not w20862;
w20864 <= not w20853 and not w20863;
w20865 <= not w264 and not w20864;
w20866 <= not w20149 and w20156;
w20867 <= not w20158 and w20866;
w20868 <= not w20259 and w20867;
w20869 <= not w20149 and not w20158;
w20870 <= not w20259 and w20869;
w20871 <= not w20156 and not w20870;
w20872 <= not w20868 and not w20871;
w20873 <= w264 and not w20853;
w20874 <= not w20863 and w20873;
w20875 <= not w20872 and not w20874;
w20876 <= not w20865 and not w20875;
w20877 <= not w184 and not w20876;
w20878 <= w20168 and not w20170;
w20879 <= not w20161 and w20878;
w20880 <= not w20259 and w20879;
w20881 <= not w20161 and not w20170;
w20882 <= not w20259 and w20881;
w20883 <= not w20168 and not w20882;
w20884 <= not w20880 and not w20883;
w20885 <= w184 and not w20865;
w20886 <= not w20875 and w20885;
w20887 <= not w20884 and not w20886;
w20888 <= not w20877 and not w20887;
w20889 <= not w115 and not w20888;
w20890 <= w115 and not w20877;
w20891 <= not w20887 and w20890;
w20892 <= not w20173 and w20182;
w20893 <= not w20175 and w20892;
w20894 <= not w20259 and w20893;
w20895 <= not w20173 and not w20175;
w20896 <= not w20259 and w20895;
w20897 <= not w20182 and not w20896;
w20898 <= not w20894 and not w20897;
w20899 <= not w20891 and not w20898;
w20900 <= not w20889 and not w20899;
w20901 <= not w60 and not w20900;
w20902 <= w20192 and not w20194;
w20903 <= not w20185 and w20902;
w20904 <= not w20259 and w20903;
w20905 <= not w20185 and not w20194;
w20906 <= not w20259 and w20905;
w20907 <= not w20192 and not w20906;
w20908 <= not w20904 and not w20907;
w20909 <= w60 and not w20889;
w20910 <= not w20899 and w20909;
w20911 <= not w20908 and not w20910;
w20912 <= not w20901 and not w20911;
w20913 <= not w22 and not w20912;
w20914 <= not w20197 and w20204;
w20915 <= not w20206 and w20914;
w20916 <= not w20259 and w20915;
w20917 <= not w20197 and not w20206;
w20918 <= not w20259 and w20917;
w20919 <= not w20204 and not w20918;
w20920 <= not w20916 and not w20919;
w20921 <= w22 and not w20901;
w20922 <= not w20911 and w20921;
w20923 <= not w20920 and not w20922;
w20924 <= not w20913 and not w20923;
w20925 <= not w5 and not w20924;
w20926 <= w20216 and not w20218;
w20927 <= not w20209 and w20926;
w20928 <= not w20259 and w20927;
w20929 <= not w20209 and not w20218;
w20930 <= not w20259 and w20929;
w20931 <= not w20216 and not w20930;
w20932 <= not w20928 and not w20931;
w20933 <= w5 and not w20913;
w20934 <= not w20923 and w20933;
w20935 <= not w20932 and not w20934;
w20936 <= not w20925 and not w20935;
w20937 <= not w20221 and w20228;
w20938 <= not w20230 and w20937;
w20939 <= not w20259 and w20938;
w20940 <= not w20221 and not w20230;
w20941 <= not w20259 and w20940;
w20942 <= not w20228 and not w20941;
w20943 <= not w20939 and not w20942;
w20944 <= not w20232 and not w20239;
w20945 <= not w20259 and w20944;
w20946 <= not w20247 and not w20945;
w20947 <= not w20943 and w20946;
w20948 <= not w20936 and w20947;
w20949 <= w0 and not w20948;
w20950 <= not w20925 and w20943;
w20951 <= not w20935 and w20950;
w20952 <= not w20239 and not w20259;
w20953 <= w20232 and not w20952;
w20954 <= not w0 and not w20944;
w20955 <= not w20953 and w20954;
w20956 <= not w20951 and not w20955;
w20957 <= not w20949 and w20956;
w20958 <= a(10) and not w20957;
w20959 <= not a(8) and not a(9);
w20960 <= not a(10) and w20959;
w20961 <= not w20958 and not w20960;
w20962 <= not w20259 and not w20961;
w20963 <= not w20256 and not w20960;
w20964 <= not w20251 and w20963;
w20965 <= not w20247 and w20964;
w20966 <= not w20245 and w20965;
w20967 <= not w20958 and w20966;
w20968 <= not a(10) and not w20957;
w20969 <= a(11) and not w20968;
w20970 <= w20261 and not w20957;
w20971 <= not w20969 and not w20970;
w20972 <= not w20967 and w20971;
w20973 <= not w20962 and not w20972;
w20974 <= not w19567 and not w20973;
w20975 <= w19567 and not w20962;
w20976 <= not w20972 and w20975;
w20977 <= not w20259 and not w20955;
w20978 <= not w20951 and w20977;
w20979 <= not w20949 and w20978;
w20980 <= not w20970 and not w20979;
w20981 <= a(12) and not w20980;
w20982 <= not a(12) and not w20979;
w20983 <= not w20970 and w20982;
w20984 <= not w20981 and not w20983;
w20985 <= not w20976 and not w20984;
w20986 <= not w20974 and not w20985;
w20987 <= not w18887 and not w20986;
w20988 <= not w20264 and not w20269;
w20989 <= not w20273 and w20988;
w20990 <= not w20957 and w20989;
w20991 <= not w20957 and w20988;
w20992 <= w20273 and not w20991;
w20993 <= not w20990 and not w20992;
w20994 <= w18887 and not w20974;
w20995 <= not w20985 and w20994;
w20996 <= not w20993 and not w20995;
w20997 <= not w20987 and not w20996;
w20998 <= not w18219 and not w20997;
w20999 <= not w20278 and w20287;
w21000 <= not w20276 and w20999;
w21001 <= not w20957 and w21000;
w21002 <= not w20276 and not w20278;
w21003 <= not w20957 and w21002;
w21004 <= not w20287 and not w21003;
w21005 <= not w21001 and not w21004;
w21006 <= w18219 and not w20987;
w21007 <= not w20996 and w21006;
w21008 <= not w21005 and not w21007;
w21009 <= not w20998 and not w21008;
w21010 <= not w17563 and not w21009;
w21011 <= not w20290 and w20296;
w21012 <= not w20298 and w21011;
w21013 <= not w20957 and w21012;
w21014 <= not w20290 and not w20298;
w21015 <= not w20957 and w21014;
w21016 <= not w20296 and not w21015;
w21017 <= not w21013 and not w21016;
w21018 <= w17563 and not w20998;
w21019 <= not w21008 and w21018;
w21020 <= not w21017 and not w21019;
w21021 <= not w21010 and not w21020;
w21022 <= not w16919 and not w21021;
w21023 <= w20308 and not w20310;
w21024 <= not w20301 and w21023;
w21025 <= not w20957 and w21024;
w21026 <= not w20301 and not w20310;
w21027 <= not w20957 and w21026;
w21028 <= not w20308 and not w21027;
w21029 <= not w21025 and not w21028;
w21030 <= w16919 and not w21010;
w21031 <= not w21020 and w21030;
w21032 <= not w21029 and not w21031;
w21033 <= not w21022 and not w21032;
w21034 <= not w16287 and not w21033;
w21035 <= not w20313 and w20320;
w21036 <= not w20322 and w21035;
w21037 <= not w20957 and w21036;
w21038 <= not w20313 and not w20322;
w21039 <= not w20957 and w21038;
w21040 <= not w20320 and not w21039;
w21041 <= not w21037 and not w21040;
w21042 <= w16287 and not w21022;
w21043 <= not w21032 and w21042;
w21044 <= not w21041 and not w21043;
w21045 <= not w21034 and not w21044;
w21046 <= not w15667 and not w21045;
w21047 <= w20332 and not w20334;
w21048 <= not w20325 and w21047;
w21049 <= not w20957 and w21048;
w21050 <= not w20325 and not w20334;
w21051 <= not w20957 and w21050;
w21052 <= not w20332 and not w21051;
w21053 <= not w21049 and not w21052;
w21054 <= w15667 and not w21034;
w21055 <= not w21044 and w21054;
w21056 <= not w21053 and not w21055;
w21057 <= not w21046 and not w21056;
w21058 <= not w15059 and not w21057;
w21059 <= not w20337 and w20344;
w21060 <= not w20346 and w21059;
w21061 <= not w20957 and w21060;
w21062 <= not w20337 and not w20346;
w21063 <= not w20957 and w21062;
w21064 <= not w20344 and not w21063;
w21065 <= not w21061 and not w21064;
w21066 <= w15059 and not w21046;
w21067 <= not w21056 and w21066;
w21068 <= not w21065 and not w21067;
w21069 <= not w21058 and not w21068;
w21070 <= not w14463 and not w21069;
w21071 <= w20356 and not w20358;
w21072 <= not w20349 and w21071;
w21073 <= not w20957 and w21072;
w21074 <= not w20349 and not w20358;
w21075 <= not w20957 and w21074;
w21076 <= not w20356 and not w21075;
w21077 <= not w21073 and not w21076;
w21078 <= w14463 and not w21058;
w21079 <= not w21068 and w21078;
w21080 <= not w21077 and not w21079;
w21081 <= not w21070 and not w21080;
w21082 <= not w13879 and not w21081;
w21083 <= not w20361 and w20368;
w21084 <= not w20370 and w21083;
w21085 <= not w20957 and w21084;
w21086 <= not w20361 and not w20370;
w21087 <= not w20957 and w21086;
w21088 <= not w20368 and not w21087;
w21089 <= not w21085 and not w21088;
w21090 <= w13879 and not w21070;
w21091 <= not w21080 and w21090;
w21092 <= not w21089 and not w21091;
w21093 <= not w21082 and not w21092;
w21094 <= not w13307 and not w21093;
w21095 <= w20380 and not w20382;
w21096 <= not w20373 and w21095;
w21097 <= not w20957 and w21096;
w21098 <= not w20373 and not w20382;
w21099 <= not w20957 and w21098;
w21100 <= not w20380 and not w21099;
w21101 <= not w21097 and not w21100;
w21102 <= w13307 and not w21082;
w21103 <= not w21092 and w21102;
w21104 <= not w21101 and not w21103;
w21105 <= not w21094 and not w21104;
w21106 <= not w12747 and not w21105;
w21107 <= not w20385 and w20392;
w21108 <= not w20394 and w21107;
w21109 <= not w20957 and w21108;
w21110 <= not w20385 and not w20394;
w21111 <= not w20957 and w21110;
w21112 <= not w20392 and not w21111;
w21113 <= not w21109 and not w21112;
w21114 <= w12747 and not w21094;
w21115 <= not w21104 and w21114;
w21116 <= not w21113 and not w21115;
w21117 <= not w21106 and not w21116;
w21118 <= not w12199 and not w21117;
w21119 <= w20404 and not w20406;
w21120 <= not w20397 and w21119;
w21121 <= not w20957 and w21120;
w21122 <= not w20397 and not w20406;
w21123 <= not w20957 and w21122;
w21124 <= not w20404 and not w21123;
w21125 <= not w21121 and not w21124;
w21126 <= w12199 and not w21106;
w21127 <= not w21116 and w21126;
w21128 <= not w21125 and not w21127;
w21129 <= not w21118 and not w21128;
w21130 <= not w11663 and not w21129;
w21131 <= not w20409 and w20416;
w21132 <= not w20418 and w21131;
w21133 <= not w20957 and w21132;
w21134 <= not w20409 and not w20418;
w21135 <= not w20957 and w21134;
w21136 <= not w20416 and not w21135;
w21137 <= not w21133 and not w21136;
w21138 <= w11663 and not w21118;
w21139 <= not w21128 and w21138;
w21140 <= not w21137 and not w21139;
w21141 <= not w21130 and not w21140;
w21142 <= not w11139 and not w21141;
w21143 <= w20428 and not w20430;
w21144 <= not w20421 and w21143;
w21145 <= not w20957 and w21144;
w21146 <= not w20421 and not w20430;
w21147 <= not w20957 and w21146;
w21148 <= not w20428 and not w21147;
w21149 <= not w21145 and not w21148;
w21150 <= w11139 and not w21130;
w21151 <= not w21140 and w21150;
w21152 <= not w21149 and not w21151;
w21153 <= not w21142 and not w21152;
w21154 <= not w10627 and not w21153;
w21155 <= not w20433 and w20440;
w21156 <= not w20442 and w21155;
w21157 <= not w20957 and w21156;
w21158 <= not w20433 and not w20442;
w21159 <= not w20957 and w21158;
w21160 <= not w20440 and not w21159;
w21161 <= not w21157 and not w21160;
w21162 <= w10627 and not w21142;
w21163 <= not w21152 and w21162;
w21164 <= not w21161 and not w21163;
w21165 <= not w21154 and not w21164;
w21166 <= not w10127 and not w21165;
w21167 <= w20452 and not w20454;
w21168 <= not w20445 and w21167;
w21169 <= not w20957 and w21168;
w21170 <= not w20445 and not w20454;
w21171 <= not w20957 and w21170;
w21172 <= not w20452 and not w21171;
w21173 <= not w21169 and not w21172;
w21174 <= w10127 and not w21154;
w21175 <= not w21164 and w21174;
w21176 <= not w21173 and not w21175;
w21177 <= not w21166 and not w21176;
w21178 <= not w9639 and not w21177;
w21179 <= not w20457 and w20464;
w21180 <= not w20466 and w21179;
w21181 <= not w20957 and w21180;
w21182 <= not w20457 and not w20466;
w21183 <= not w20957 and w21182;
w21184 <= not w20464 and not w21183;
w21185 <= not w21181 and not w21184;
w21186 <= w9639 and not w21166;
w21187 <= not w21176 and w21186;
w21188 <= not w21185 and not w21187;
w21189 <= not w21178 and not w21188;
w21190 <= not w9163 and not w21189;
w21191 <= w20476 and not w20478;
w21192 <= not w20469 and w21191;
w21193 <= not w20957 and w21192;
w21194 <= not w20469 and not w20478;
w21195 <= not w20957 and w21194;
w21196 <= not w20476 and not w21195;
w21197 <= not w21193 and not w21196;
w21198 <= w9163 and not w21178;
w21199 <= not w21188 and w21198;
w21200 <= not w21197 and not w21199;
w21201 <= not w21190 and not w21200;
w21202 <= not w8699 and not w21201;
w21203 <= not w20481 and w20488;
w21204 <= not w20490 and w21203;
w21205 <= not w20957 and w21204;
w21206 <= not w20481 and not w20490;
w21207 <= not w20957 and w21206;
w21208 <= not w20488 and not w21207;
w21209 <= not w21205 and not w21208;
w21210 <= w8699 and not w21190;
w21211 <= not w21200 and w21210;
w21212 <= not w21209 and not w21211;
w21213 <= not w21202 and not w21212;
w21214 <= not w8247 and not w21213;
w21215 <= w20500 and not w20502;
w21216 <= not w20493 and w21215;
w21217 <= not w20957 and w21216;
w21218 <= not w20493 and not w20502;
w21219 <= not w20957 and w21218;
w21220 <= not w20500 and not w21219;
w21221 <= not w21217 and not w21220;
w21222 <= w8247 and not w21202;
w21223 <= not w21212 and w21222;
w21224 <= not w21221 and not w21223;
w21225 <= not w21214 and not w21224;
w21226 <= not w7807 and not w21225;
w21227 <= not w20505 and w20512;
w21228 <= not w20514 and w21227;
w21229 <= not w20957 and w21228;
w21230 <= not w20505 and not w20514;
w21231 <= not w20957 and w21230;
w21232 <= not w20512 and not w21231;
w21233 <= not w21229 and not w21232;
w21234 <= w7807 and not w21214;
w21235 <= not w21224 and w21234;
w21236 <= not w21233 and not w21235;
w21237 <= not w21226 and not w21236;
w21238 <= not w7379 and not w21237;
w21239 <= w20524 and not w20526;
w21240 <= not w20517 and w21239;
w21241 <= not w20957 and w21240;
w21242 <= not w20517 and not w20526;
w21243 <= not w20957 and w21242;
w21244 <= not w20524 and not w21243;
w21245 <= not w21241 and not w21244;
w21246 <= w7379 and not w21226;
w21247 <= not w21236 and w21246;
w21248 <= not w21245 and not w21247;
w21249 <= not w21238 and not w21248;
w21250 <= not w6963 and not w21249;
w21251 <= not w20529 and w20536;
w21252 <= not w20538 and w21251;
w21253 <= not w20957 and w21252;
w21254 <= not w20529 and not w20538;
w21255 <= not w20957 and w21254;
w21256 <= not w20536 and not w21255;
w21257 <= not w21253 and not w21256;
w21258 <= w6963 and not w21238;
w21259 <= not w21248 and w21258;
w21260 <= not w21257 and not w21259;
w21261 <= not w21250 and not w21260;
w21262 <= not w6558 and not w21261;
w21263 <= w20548 and not w20550;
w21264 <= not w20541 and w21263;
w21265 <= not w20957 and w21264;
w21266 <= not w20541 and not w20550;
w21267 <= not w20957 and w21266;
w21268 <= not w20548 and not w21267;
w21269 <= not w21265 and not w21268;
w21270 <= w6558 and not w21250;
w21271 <= not w21260 and w21270;
w21272 <= not w21269 and not w21271;
w21273 <= not w21262 and not w21272;
w21274 <= not w6166 and not w21273;
w21275 <= not w20553 and w20560;
w21276 <= not w20562 and w21275;
w21277 <= not w20957 and w21276;
w21278 <= not w20553 and not w20562;
w21279 <= not w20957 and w21278;
w21280 <= not w20560 and not w21279;
w21281 <= not w21277 and not w21280;
w21282 <= w6166 and not w21262;
w21283 <= not w21272 and w21282;
w21284 <= not w21281 and not w21283;
w21285 <= not w21274 and not w21284;
w21286 <= not w5786 and not w21285;
w21287 <= w20572 and not w20574;
w21288 <= not w20565 and w21287;
w21289 <= not w20957 and w21288;
w21290 <= not w20565 and not w20574;
w21291 <= not w20957 and w21290;
w21292 <= not w20572 and not w21291;
w21293 <= not w21289 and not w21292;
w21294 <= w5786 and not w21274;
w21295 <= not w21284 and w21294;
w21296 <= not w21293 and not w21295;
w21297 <= not w21286 and not w21296;
w21298 <= not w5418 and not w21297;
w21299 <= not w20577 and w20584;
w21300 <= not w20586 and w21299;
w21301 <= not w20957 and w21300;
w21302 <= not w20577 and not w20586;
w21303 <= not w20957 and w21302;
w21304 <= not w20584 and not w21303;
w21305 <= not w21301 and not w21304;
w21306 <= w5418 and not w21286;
w21307 <= not w21296 and w21306;
w21308 <= not w21305 and not w21307;
w21309 <= not w21298 and not w21308;
w21310 <= not w5062 and not w21309;
w21311 <= w20596 and not w20598;
w21312 <= not w20589 and w21311;
w21313 <= not w20957 and w21312;
w21314 <= not w20589 and not w20598;
w21315 <= not w20957 and w21314;
w21316 <= not w20596 and not w21315;
w21317 <= not w21313 and not w21316;
w21318 <= w5062 and not w21298;
w21319 <= not w21308 and w21318;
w21320 <= not w21317 and not w21319;
w21321 <= not w21310 and not w21320;
w21322 <= not w4718 and not w21321;
w21323 <= not w20601 and w20608;
w21324 <= not w20610 and w21323;
w21325 <= not w20957 and w21324;
w21326 <= not w20601 and not w20610;
w21327 <= not w20957 and w21326;
w21328 <= not w20608 and not w21327;
w21329 <= not w21325 and not w21328;
w21330 <= w4718 and not w21310;
w21331 <= not w21320 and w21330;
w21332 <= not w21329 and not w21331;
w21333 <= not w21322 and not w21332;
w21334 <= not w4386 and not w21333;
w21335 <= w20620 and not w20622;
w21336 <= not w20613 and w21335;
w21337 <= not w20957 and w21336;
w21338 <= not w20613 and not w20622;
w21339 <= not w20957 and w21338;
w21340 <= not w20620 and not w21339;
w21341 <= not w21337 and not w21340;
w21342 <= w4386 and not w21322;
w21343 <= not w21332 and w21342;
w21344 <= not w21341 and not w21343;
w21345 <= not w21334 and not w21344;
w21346 <= not w4066 and not w21345;
w21347 <= not w20625 and w20632;
w21348 <= not w20634 and w21347;
w21349 <= not w20957 and w21348;
w21350 <= not w20625 and not w20634;
w21351 <= not w20957 and w21350;
w21352 <= not w20632 and not w21351;
w21353 <= not w21349 and not w21352;
w21354 <= w4066 and not w21334;
w21355 <= not w21344 and w21354;
w21356 <= not w21353 and not w21355;
w21357 <= not w21346 and not w21356;
w21358 <= not w3758 and not w21357;
w21359 <= w20644 and not w20646;
w21360 <= not w20637 and w21359;
w21361 <= not w20957 and w21360;
w21362 <= not w20637 and not w20646;
w21363 <= not w20957 and w21362;
w21364 <= not w20644 and not w21363;
w21365 <= not w21361 and not w21364;
w21366 <= w3758 and not w21346;
w21367 <= not w21356 and w21366;
w21368 <= not w21365 and not w21367;
w21369 <= not w21358 and not w21368;
w21370 <= not w3462 and not w21369;
w21371 <= not w20649 and w20656;
w21372 <= not w20658 and w21371;
w21373 <= not w20957 and w21372;
w21374 <= not w20649 and not w20658;
w21375 <= not w20957 and w21374;
w21376 <= not w20656 and not w21375;
w21377 <= not w21373 and not w21376;
w21378 <= w3462 and not w21358;
w21379 <= not w21368 and w21378;
w21380 <= not w21377 and not w21379;
w21381 <= not w21370 and not w21380;
w21382 <= not w3178 and not w21381;
w21383 <= w20668 and not w20670;
w21384 <= not w20661 and w21383;
w21385 <= not w20957 and w21384;
w21386 <= not w20661 and not w20670;
w21387 <= not w20957 and w21386;
w21388 <= not w20668 and not w21387;
w21389 <= not w21385 and not w21388;
w21390 <= w3178 and not w21370;
w21391 <= not w21380 and w21390;
w21392 <= not w21389 and not w21391;
w21393 <= not w21382 and not w21392;
w21394 <= not w2906 and not w21393;
w21395 <= not w20673 and w20680;
w21396 <= not w20682 and w21395;
w21397 <= not w20957 and w21396;
w21398 <= not w20673 and not w20682;
w21399 <= not w20957 and w21398;
w21400 <= not w20680 and not w21399;
w21401 <= not w21397 and not w21400;
w21402 <= w2906 and not w21382;
w21403 <= not w21392 and w21402;
w21404 <= not w21401 and not w21403;
w21405 <= not w21394 and not w21404;
w21406 <= not w2646 and not w21405;
w21407 <= w20692 and not w20694;
w21408 <= not w20685 and w21407;
w21409 <= not w20957 and w21408;
w21410 <= not w20685 and not w20694;
w21411 <= not w20957 and w21410;
w21412 <= not w20692 and not w21411;
w21413 <= not w21409 and not w21412;
w21414 <= w2646 and not w21394;
w21415 <= not w21404 and w21414;
w21416 <= not w21413 and not w21415;
w21417 <= not w21406 and not w21416;
w21418 <= not w2398 and not w21417;
w21419 <= not w20697 and w20704;
w21420 <= not w20706 and w21419;
w21421 <= not w20957 and w21420;
w21422 <= not w20697 and not w20706;
w21423 <= not w20957 and w21422;
w21424 <= not w20704 and not w21423;
w21425 <= not w21421 and not w21424;
w21426 <= w2398 and not w21406;
w21427 <= not w21416 and w21426;
w21428 <= not w21425 and not w21427;
w21429 <= not w21418 and not w21428;
w21430 <= not w2162 and not w21429;
w21431 <= w20716 and not w20718;
w21432 <= not w20709 and w21431;
w21433 <= not w20957 and w21432;
w21434 <= not w20709 and not w20718;
w21435 <= not w20957 and w21434;
w21436 <= not w20716 and not w21435;
w21437 <= not w21433 and not w21436;
w21438 <= w2162 and not w21418;
w21439 <= not w21428 and w21438;
w21440 <= not w21437 and not w21439;
w21441 <= not w21430 and not w21440;
w21442 <= not w1938 and not w21441;
w21443 <= not w20721 and w20728;
w21444 <= not w20730 and w21443;
w21445 <= not w20957 and w21444;
w21446 <= not w20721 and not w20730;
w21447 <= not w20957 and w21446;
w21448 <= not w20728 and not w21447;
w21449 <= not w21445 and not w21448;
w21450 <= w1938 and not w21430;
w21451 <= not w21440 and w21450;
w21452 <= not w21449 and not w21451;
w21453 <= not w21442 and not w21452;
w21454 <= not w1725 and not w21453;
w21455 <= w20740 and not w20742;
w21456 <= not w20733 and w21455;
w21457 <= not w20957 and w21456;
w21458 <= not w20733 and not w20742;
w21459 <= not w20957 and w21458;
w21460 <= not w20740 and not w21459;
w21461 <= not w21457 and not w21460;
w21462 <= w1725 and not w21442;
w21463 <= not w21452 and w21462;
w21464 <= not w21461 and not w21463;
w21465 <= not w21454 and not w21464;
w21466 <= not w1525 and not w21465;
w21467 <= not w20745 and w20752;
w21468 <= not w20754 and w21467;
w21469 <= not w20957 and w21468;
w21470 <= not w20745 and not w20754;
w21471 <= not w20957 and w21470;
w21472 <= not w20752 and not w21471;
w21473 <= not w21469 and not w21472;
w21474 <= w1525 and not w21454;
w21475 <= not w21464 and w21474;
w21476 <= not w21473 and not w21475;
w21477 <= not w21466 and not w21476;
w21478 <= not w1337 and not w21477;
w21479 <= w20764 and not w20766;
w21480 <= not w20757 and w21479;
w21481 <= not w20957 and w21480;
w21482 <= not w20757 and not w20766;
w21483 <= not w20957 and w21482;
w21484 <= not w20764 and not w21483;
w21485 <= not w21481 and not w21484;
w21486 <= w1337 and not w21466;
w21487 <= not w21476 and w21486;
w21488 <= not w21485 and not w21487;
w21489 <= not w21478 and not w21488;
w21490 <= not w1161 and not w21489;
w21491 <= not w20769 and w20776;
w21492 <= not w20778 and w21491;
w21493 <= not w20957 and w21492;
w21494 <= not w20769 and not w20778;
w21495 <= not w20957 and w21494;
w21496 <= not w20776 and not w21495;
w21497 <= not w21493 and not w21496;
w21498 <= w1161 and not w21478;
w21499 <= not w21488 and w21498;
w21500 <= not w21497 and not w21499;
w21501 <= not w21490 and not w21500;
w21502 <= not w997 and not w21501;
w21503 <= w20788 and not w20790;
w21504 <= not w20781 and w21503;
w21505 <= not w20957 and w21504;
w21506 <= not w20781 and not w20790;
w21507 <= not w20957 and w21506;
w21508 <= not w20788 and not w21507;
w21509 <= not w21505 and not w21508;
w21510 <= w997 and not w21490;
w21511 <= not w21500 and w21510;
w21512 <= not w21509 and not w21511;
w21513 <= not w21502 and not w21512;
w21514 <= not w845 and not w21513;
w21515 <= not w20793 and w20800;
w21516 <= not w20802 and w21515;
w21517 <= not w20957 and w21516;
w21518 <= not w20793 and not w20802;
w21519 <= not w20957 and w21518;
w21520 <= not w20800 and not w21519;
w21521 <= not w21517 and not w21520;
w21522 <= w845 and not w21502;
w21523 <= not w21512 and w21522;
w21524 <= not w21521 and not w21523;
w21525 <= not w21514 and not w21524;
w21526 <= not w705 and not w21525;
w21527 <= w20812 and not w20814;
w21528 <= not w20805 and w21527;
w21529 <= not w20957 and w21528;
w21530 <= not w20805 and not w20814;
w21531 <= not w20957 and w21530;
w21532 <= not w20812 and not w21531;
w21533 <= not w21529 and not w21532;
w21534 <= w705 and not w21514;
w21535 <= not w21524 and w21534;
w21536 <= not w21533 and not w21535;
w21537 <= not w21526 and not w21536;
w21538 <= not w577 and not w21537;
w21539 <= not w20817 and w20824;
w21540 <= not w20826 and w21539;
w21541 <= not w20957 and w21540;
w21542 <= not w20817 and not w20826;
w21543 <= not w20957 and w21542;
w21544 <= not w20824 and not w21543;
w21545 <= not w21541 and not w21544;
w21546 <= w577 and not w21526;
w21547 <= not w21536 and w21546;
w21548 <= not w21545 and not w21547;
w21549 <= not w21538 and not w21548;
w21550 <= not w460 and not w21549;
w21551 <= w20836 and not w20838;
w21552 <= not w20829 and w21551;
w21553 <= not w20957 and w21552;
w21554 <= not w20829 and not w20838;
w21555 <= not w20957 and w21554;
w21556 <= not w20836 and not w21555;
w21557 <= not w21553 and not w21556;
w21558 <= w460 and not w21538;
w21559 <= not w21548 and w21558;
w21560 <= not w21557 and not w21559;
w21561 <= not w21550 and not w21560;
w21562 <= not w356 and not w21561;
w21563 <= not w20841 and w20848;
w21564 <= not w20850 and w21563;
w21565 <= not w20957 and w21564;
w21566 <= not w20841 and not w20850;
w21567 <= not w20957 and w21566;
w21568 <= not w20848 and not w21567;
w21569 <= not w21565 and not w21568;
w21570 <= w356 and not w21550;
w21571 <= not w21560 and w21570;
w21572 <= not w21569 and not w21571;
w21573 <= not w21562 and not w21572;
w21574 <= not w264 and not w21573;
w21575 <= w20860 and not w20862;
w21576 <= not w20853 and w21575;
w21577 <= not w20957 and w21576;
w21578 <= not w20853 and not w20862;
w21579 <= not w20957 and w21578;
w21580 <= not w20860 and not w21579;
w21581 <= not w21577 and not w21580;
w21582 <= w264 and not w21562;
w21583 <= not w21572 and w21582;
w21584 <= not w21581 and not w21583;
w21585 <= not w21574 and not w21584;
w21586 <= not w184 and not w21585;
w21587 <= not w20865 and w20872;
w21588 <= not w20874 and w21587;
w21589 <= not w20957 and w21588;
w21590 <= not w20865 and not w20874;
w21591 <= not w20957 and w21590;
w21592 <= not w20872 and not w21591;
w21593 <= not w21589 and not w21592;
w21594 <= w184 and not w21574;
w21595 <= not w21584 and w21594;
w21596 <= not w21593 and not w21595;
w21597 <= not w21586 and not w21596;
w21598 <= not w115 and not w21597;
w21599 <= w20884 and not w20886;
w21600 <= not w20877 and w21599;
w21601 <= not w20957 and w21600;
w21602 <= not w20877 and not w20886;
w21603 <= not w20957 and w21602;
w21604 <= not w20884 and not w21603;
w21605 <= not w21601 and not w21604;
w21606 <= w115 and not w21586;
w21607 <= not w21596 and w21606;
w21608 <= not w21605 and not w21607;
w21609 <= not w21598 and not w21608;
w21610 <= not w60 and not w21609;
w21611 <= w60 and not w21598;
w21612 <= not w21608 and w21611;
w21613 <= not w20889 and w20898;
w21614 <= not w20891 and w21613;
w21615 <= not w20957 and w21614;
w21616 <= not w20889 and not w20891;
w21617 <= not w20957 and w21616;
w21618 <= not w20898 and not w21617;
w21619 <= not w21615 and not w21618;
w21620 <= not w21612 and not w21619;
w21621 <= not w21610 and not w21620;
w21622 <= not w22 and not w21621;
w21623 <= w20908 and not w20910;
w21624 <= not w20901 and w21623;
w21625 <= not w20957 and w21624;
w21626 <= not w20901 and not w20910;
w21627 <= not w20957 and w21626;
w21628 <= not w20908 and not w21627;
w21629 <= not w21625 and not w21628;
w21630 <= w22 and not w21610;
w21631 <= not w21620 and w21630;
w21632 <= not w21629 and not w21631;
w21633 <= not w21622 and not w21632;
w21634 <= not w5 and not w21633;
w21635 <= not w20913 and w20920;
w21636 <= not w20922 and w21635;
w21637 <= not w20957 and w21636;
w21638 <= not w20913 and not w20922;
w21639 <= not w20957 and w21638;
w21640 <= not w20920 and not w21639;
w21641 <= not w21637 and not w21640;
w21642 <= w5 and not w21622;
w21643 <= not w21632 and w21642;
w21644 <= not w21641 and not w21643;
w21645 <= not w21634 and not w21644;
w21646 <= w20932 and not w20934;
w21647 <= not w20925 and w21646;
w21648 <= not w20957 and w21647;
w21649 <= not w20925 and not w20934;
w21650 <= not w20957 and w21649;
w21651 <= not w20932 and not w21650;
w21652 <= not w21648 and not w21651;
w21653 <= not w20936 and not w20943;
w21654 <= not w20957 and w21653;
w21655 <= not w20951 and not w21654;
w21656 <= not w21652 and w21655;
w21657 <= not w21645 and w21656;
w21658 <= w0 and not w21657;
w21659 <= not w21634 and w21652;
w21660 <= not w21644 and w21659;
w21661 <= not w20943 and not w20957;
w21662 <= w20936 and not w21661;
w21663 <= not w0 and not w21653;
w21664 <= not w21662 and w21663;
w21665 <= not w21660 and not w21664;
w21666 <= not w21658 and w21665;
w21667 <= a(8) and not w21666;
w21668 <= not a(6) and not a(7);
w21669 <= not a(8) and w21668;
w21670 <= not w21667 and not w21669;
w21671 <= not w20957 and not w21670;
w21672 <= not w20955 and not w21669;
w21673 <= not w20951 and w21672;
w21674 <= not w20949 and w21673;
w21675 <= not w21667 and w21674;
w21676 <= not a(8) and not w21666;
w21677 <= a(9) and not w21676;
w21678 <= w20959 and not w21666;
w21679 <= not w21677 and not w21678;
w21680 <= not w21675 and w21679;
w21681 <= not w21671 and not w21680;
w21682 <= not w20259 and not w21681;
w21683 <= w20259 and not w21671;
w21684 <= not w21680 and w21683;
w21685 <= not w20957 and not w21664;
w21686 <= not w21660 and w21685;
w21687 <= not w21658 and w21686;
w21688 <= not w21678 and not w21687;
w21689 <= a(10) and not w21688;
w21690 <= not a(10) and not w21687;
w21691 <= not w21678 and w21690;
w21692 <= not w21689 and not w21691;
w21693 <= not w21684 and not w21692;
w21694 <= not w21682 and not w21693;
w21695 <= not w19567 and not w21694;
w21696 <= not w20962 and not w20967;
w21697 <= not w20971 and w21696;
w21698 <= not w21666 and w21697;
w21699 <= not w21666 and w21696;
w21700 <= w20971 and not w21699;
w21701 <= not w21698 and not w21700;
w21702 <= w19567 and not w21682;
w21703 <= not w21693 and w21702;
w21704 <= not w21701 and not w21703;
w21705 <= not w21695 and not w21704;
w21706 <= not w18887 and not w21705;
w21707 <= not w20976 and w20984;
w21708 <= not w20974 and w21707;
w21709 <= not w21666 and w21708;
w21710 <= not w20974 and not w20976;
w21711 <= not w21666 and w21710;
w21712 <= not w20984 and not w21711;
w21713 <= not w21709 and not w21712;
w21714 <= w18887 and not w21695;
w21715 <= not w21704 and w21714;
w21716 <= not w21713 and not w21715;
w21717 <= not w21706 and not w21716;
w21718 <= not w18219 and not w21717;
w21719 <= not w20987 and w20993;
w21720 <= not w20995 and w21719;
w21721 <= not w21666 and w21720;
w21722 <= not w20987 and not w20995;
w21723 <= not w21666 and w21722;
w21724 <= not w20993 and not w21723;
w21725 <= not w21721 and not w21724;
w21726 <= w18219 and not w21706;
w21727 <= not w21716 and w21726;
w21728 <= not w21725 and not w21727;
w21729 <= not w21718 and not w21728;
w21730 <= not w17563 and not w21729;
w21731 <= w21005 and not w21007;
w21732 <= not w20998 and w21731;
w21733 <= not w21666 and w21732;
w21734 <= not w20998 and not w21007;
w21735 <= not w21666 and w21734;
w21736 <= not w21005 and not w21735;
w21737 <= not w21733 and not w21736;
w21738 <= w17563 and not w21718;
w21739 <= not w21728 and w21738;
w21740 <= not w21737 and not w21739;
w21741 <= not w21730 and not w21740;
w21742 <= not w16919 and not w21741;
w21743 <= not w21010 and w21017;
w21744 <= not w21019 and w21743;
w21745 <= not w21666 and w21744;
w21746 <= not w21010 and not w21019;
w21747 <= not w21666 and w21746;
w21748 <= not w21017 and not w21747;
w21749 <= not w21745 and not w21748;
w21750 <= w16919 and not w21730;
w21751 <= not w21740 and w21750;
w21752 <= not w21749 and not w21751;
w21753 <= not w21742 and not w21752;
w21754 <= not w16287 and not w21753;
w21755 <= w21029 and not w21031;
w21756 <= not w21022 and w21755;
w21757 <= not w21666 and w21756;
w21758 <= not w21022 and not w21031;
w21759 <= not w21666 and w21758;
w21760 <= not w21029 and not w21759;
w21761 <= not w21757 and not w21760;
w21762 <= w16287 and not w21742;
w21763 <= not w21752 and w21762;
w21764 <= not w21761 and not w21763;
w21765 <= not w21754 and not w21764;
w21766 <= not w15667 and not w21765;
w21767 <= not w21034 and w21041;
w21768 <= not w21043 and w21767;
w21769 <= not w21666 and w21768;
w21770 <= not w21034 and not w21043;
w21771 <= not w21666 and w21770;
w21772 <= not w21041 and not w21771;
w21773 <= not w21769 and not w21772;
w21774 <= w15667 and not w21754;
w21775 <= not w21764 and w21774;
w21776 <= not w21773 and not w21775;
w21777 <= not w21766 and not w21776;
w21778 <= not w15059 and not w21777;
w21779 <= w21053 and not w21055;
w21780 <= not w21046 and w21779;
w21781 <= not w21666 and w21780;
w21782 <= not w21046 and not w21055;
w21783 <= not w21666 and w21782;
w21784 <= not w21053 and not w21783;
w21785 <= not w21781 and not w21784;
w21786 <= w15059 and not w21766;
w21787 <= not w21776 and w21786;
w21788 <= not w21785 and not w21787;
w21789 <= not w21778 and not w21788;
w21790 <= not w14463 and not w21789;
w21791 <= not w21058 and w21065;
w21792 <= not w21067 and w21791;
w21793 <= not w21666 and w21792;
w21794 <= not w21058 and not w21067;
w21795 <= not w21666 and w21794;
w21796 <= not w21065 and not w21795;
w21797 <= not w21793 and not w21796;
w21798 <= w14463 and not w21778;
w21799 <= not w21788 and w21798;
w21800 <= not w21797 and not w21799;
w21801 <= not w21790 and not w21800;
w21802 <= not w13879 and not w21801;
w21803 <= w21077 and not w21079;
w21804 <= not w21070 and w21803;
w21805 <= not w21666 and w21804;
w21806 <= not w21070 and not w21079;
w21807 <= not w21666 and w21806;
w21808 <= not w21077 and not w21807;
w21809 <= not w21805 and not w21808;
w21810 <= w13879 and not w21790;
w21811 <= not w21800 and w21810;
w21812 <= not w21809 and not w21811;
w21813 <= not w21802 and not w21812;
w21814 <= not w13307 and not w21813;
w21815 <= not w21082 and w21089;
w21816 <= not w21091 and w21815;
w21817 <= not w21666 and w21816;
w21818 <= not w21082 and not w21091;
w21819 <= not w21666 and w21818;
w21820 <= not w21089 and not w21819;
w21821 <= not w21817 and not w21820;
w21822 <= w13307 and not w21802;
w21823 <= not w21812 and w21822;
w21824 <= not w21821 and not w21823;
w21825 <= not w21814 and not w21824;
w21826 <= not w12747 and not w21825;
w21827 <= w21101 and not w21103;
w21828 <= not w21094 and w21827;
w21829 <= not w21666 and w21828;
w21830 <= not w21094 and not w21103;
w21831 <= not w21666 and w21830;
w21832 <= not w21101 and not w21831;
w21833 <= not w21829 and not w21832;
w21834 <= w12747 and not w21814;
w21835 <= not w21824 and w21834;
w21836 <= not w21833 and not w21835;
w21837 <= not w21826 and not w21836;
w21838 <= not w12199 and not w21837;
w21839 <= not w21106 and w21113;
w21840 <= not w21115 and w21839;
w21841 <= not w21666 and w21840;
w21842 <= not w21106 and not w21115;
w21843 <= not w21666 and w21842;
w21844 <= not w21113 and not w21843;
w21845 <= not w21841 and not w21844;
w21846 <= w12199 and not w21826;
w21847 <= not w21836 and w21846;
w21848 <= not w21845 and not w21847;
w21849 <= not w21838 and not w21848;
w21850 <= not w11663 and not w21849;
w21851 <= w21125 and not w21127;
w21852 <= not w21118 and w21851;
w21853 <= not w21666 and w21852;
w21854 <= not w21118 and not w21127;
w21855 <= not w21666 and w21854;
w21856 <= not w21125 and not w21855;
w21857 <= not w21853 and not w21856;
w21858 <= w11663 and not w21838;
w21859 <= not w21848 and w21858;
w21860 <= not w21857 and not w21859;
w21861 <= not w21850 and not w21860;
w21862 <= not w11139 and not w21861;
w21863 <= not w21130 and w21137;
w21864 <= not w21139 and w21863;
w21865 <= not w21666 and w21864;
w21866 <= not w21130 and not w21139;
w21867 <= not w21666 and w21866;
w21868 <= not w21137 and not w21867;
w21869 <= not w21865 and not w21868;
w21870 <= w11139 and not w21850;
w21871 <= not w21860 and w21870;
w21872 <= not w21869 and not w21871;
w21873 <= not w21862 and not w21872;
w21874 <= not w10627 and not w21873;
w21875 <= w21149 and not w21151;
w21876 <= not w21142 and w21875;
w21877 <= not w21666 and w21876;
w21878 <= not w21142 and not w21151;
w21879 <= not w21666 and w21878;
w21880 <= not w21149 and not w21879;
w21881 <= not w21877 and not w21880;
w21882 <= w10627 and not w21862;
w21883 <= not w21872 and w21882;
w21884 <= not w21881 and not w21883;
w21885 <= not w21874 and not w21884;
w21886 <= not w10127 and not w21885;
w21887 <= not w21154 and w21161;
w21888 <= not w21163 and w21887;
w21889 <= not w21666 and w21888;
w21890 <= not w21154 and not w21163;
w21891 <= not w21666 and w21890;
w21892 <= not w21161 and not w21891;
w21893 <= not w21889 and not w21892;
w21894 <= w10127 and not w21874;
w21895 <= not w21884 and w21894;
w21896 <= not w21893 and not w21895;
w21897 <= not w21886 and not w21896;
w21898 <= not w9639 and not w21897;
w21899 <= w21173 and not w21175;
w21900 <= not w21166 and w21899;
w21901 <= not w21666 and w21900;
w21902 <= not w21166 and not w21175;
w21903 <= not w21666 and w21902;
w21904 <= not w21173 and not w21903;
w21905 <= not w21901 and not w21904;
w21906 <= w9639 and not w21886;
w21907 <= not w21896 and w21906;
w21908 <= not w21905 and not w21907;
w21909 <= not w21898 and not w21908;
w21910 <= not w9163 and not w21909;
w21911 <= not w21178 and w21185;
w21912 <= not w21187 and w21911;
w21913 <= not w21666 and w21912;
w21914 <= not w21178 and not w21187;
w21915 <= not w21666 and w21914;
w21916 <= not w21185 and not w21915;
w21917 <= not w21913 and not w21916;
w21918 <= w9163 and not w21898;
w21919 <= not w21908 and w21918;
w21920 <= not w21917 and not w21919;
w21921 <= not w21910 and not w21920;
w21922 <= not w8699 and not w21921;
w21923 <= w21197 and not w21199;
w21924 <= not w21190 and w21923;
w21925 <= not w21666 and w21924;
w21926 <= not w21190 and not w21199;
w21927 <= not w21666 and w21926;
w21928 <= not w21197 and not w21927;
w21929 <= not w21925 and not w21928;
w21930 <= w8699 and not w21910;
w21931 <= not w21920 and w21930;
w21932 <= not w21929 and not w21931;
w21933 <= not w21922 and not w21932;
w21934 <= not w8247 and not w21933;
w21935 <= not w21202 and w21209;
w21936 <= not w21211 and w21935;
w21937 <= not w21666 and w21936;
w21938 <= not w21202 and not w21211;
w21939 <= not w21666 and w21938;
w21940 <= not w21209 and not w21939;
w21941 <= not w21937 and not w21940;
w21942 <= w8247 and not w21922;
w21943 <= not w21932 and w21942;
w21944 <= not w21941 and not w21943;
w21945 <= not w21934 and not w21944;
w21946 <= not w7807 and not w21945;
w21947 <= w21221 and not w21223;
w21948 <= not w21214 and w21947;
w21949 <= not w21666 and w21948;
w21950 <= not w21214 and not w21223;
w21951 <= not w21666 and w21950;
w21952 <= not w21221 and not w21951;
w21953 <= not w21949 and not w21952;
w21954 <= w7807 and not w21934;
w21955 <= not w21944 and w21954;
w21956 <= not w21953 and not w21955;
w21957 <= not w21946 and not w21956;
w21958 <= not w7379 and not w21957;
w21959 <= not w21226 and w21233;
w21960 <= not w21235 and w21959;
w21961 <= not w21666 and w21960;
w21962 <= not w21226 and not w21235;
w21963 <= not w21666 and w21962;
w21964 <= not w21233 and not w21963;
w21965 <= not w21961 and not w21964;
w21966 <= w7379 and not w21946;
w21967 <= not w21956 and w21966;
w21968 <= not w21965 and not w21967;
w21969 <= not w21958 and not w21968;
w21970 <= not w6963 and not w21969;
w21971 <= w21245 and not w21247;
w21972 <= not w21238 and w21971;
w21973 <= not w21666 and w21972;
w21974 <= not w21238 and not w21247;
w21975 <= not w21666 and w21974;
w21976 <= not w21245 and not w21975;
w21977 <= not w21973 and not w21976;
w21978 <= w6963 and not w21958;
w21979 <= not w21968 and w21978;
w21980 <= not w21977 and not w21979;
w21981 <= not w21970 and not w21980;
w21982 <= not w6558 and not w21981;
w21983 <= not w21250 and w21257;
w21984 <= not w21259 and w21983;
w21985 <= not w21666 and w21984;
w21986 <= not w21250 and not w21259;
w21987 <= not w21666 and w21986;
w21988 <= not w21257 and not w21987;
w21989 <= not w21985 and not w21988;
w21990 <= w6558 and not w21970;
w21991 <= not w21980 and w21990;
w21992 <= not w21989 and not w21991;
w21993 <= not w21982 and not w21992;
w21994 <= not w6166 and not w21993;
w21995 <= w21269 and not w21271;
w21996 <= not w21262 and w21995;
w21997 <= not w21666 and w21996;
w21998 <= not w21262 and not w21271;
w21999 <= not w21666 and w21998;
w22000 <= not w21269 and not w21999;
w22001 <= not w21997 and not w22000;
w22002 <= w6166 and not w21982;
w22003 <= not w21992 and w22002;
w22004 <= not w22001 and not w22003;
w22005 <= not w21994 and not w22004;
w22006 <= not w5786 and not w22005;
w22007 <= not w21274 and w21281;
w22008 <= not w21283 and w22007;
w22009 <= not w21666 and w22008;
w22010 <= not w21274 and not w21283;
w22011 <= not w21666 and w22010;
w22012 <= not w21281 and not w22011;
w22013 <= not w22009 and not w22012;
w22014 <= w5786 and not w21994;
w22015 <= not w22004 and w22014;
w22016 <= not w22013 and not w22015;
w22017 <= not w22006 and not w22016;
w22018 <= not w5418 and not w22017;
w22019 <= w21293 and not w21295;
w22020 <= not w21286 and w22019;
w22021 <= not w21666 and w22020;
w22022 <= not w21286 and not w21295;
w22023 <= not w21666 and w22022;
w22024 <= not w21293 and not w22023;
w22025 <= not w22021 and not w22024;
w22026 <= w5418 and not w22006;
w22027 <= not w22016 and w22026;
w22028 <= not w22025 and not w22027;
w22029 <= not w22018 and not w22028;
w22030 <= not w5062 and not w22029;
w22031 <= not w21298 and w21305;
w22032 <= not w21307 and w22031;
w22033 <= not w21666 and w22032;
w22034 <= not w21298 and not w21307;
w22035 <= not w21666 and w22034;
w22036 <= not w21305 and not w22035;
w22037 <= not w22033 and not w22036;
w22038 <= w5062 and not w22018;
w22039 <= not w22028 and w22038;
w22040 <= not w22037 and not w22039;
w22041 <= not w22030 and not w22040;
w22042 <= not w4718 and not w22041;
w22043 <= w21317 and not w21319;
w22044 <= not w21310 and w22043;
w22045 <= not w21666 and w22044;
w22046 <= not w21310 and not w21319;
w22047 <= not w21666 and w22046;
w22048 <= not w21317 and not w22047;
w22049 <= not w22045 and not w22048;
w22050 <= w4718 and not w22030;
w22051 <= not w22040 and w22050;
w22052 <= not w22049 and not w22051;
w22053 <= not w22042 and not w22052;
w22054 <= not w4386 and not w22053;
w22055 <= not w21322 and w21329;
w22056 <= not w21331 and w22055;
w22057 <= not w21666 and w22056;
w22058 <= not w21322 and not w21331;
w22059 <= not w21666 and w22058;
w22060 <= not w21329 and not w22059;
w22061 <= not w22057 and not w22060;
w22062 <= w4386 and not w22042;
w22063 <= not w22052 and w22062;
w22064 <= not w22061 and not w22063;
w22065 <= not w22054 and not w22064;
w22066 <= not w4066 and not w22065;
w22067 <= w21341 and not w21343;
w22068 <= not w21334 and w22067;
w22069 <= not w21666 and w22068;
w22070 <= not w21334 and not w21343;
w22071 <= not w21666 and w22070;
w22072 <= not w21341 and not w22071;
w22073 <= not w22069 and not w22072;
w22074 <= w4066 and not w22054;
w22075 <= not w22064 and w22074;
w22076 <= not w22073 and not w22075;
w22077 <= not w22066 and not w22076;
w22078 <= not w3758 and not w22077;
w22079 <= not w21346 and w21353;
w22080 <= not w21355 and w22079;
w22081 <= not w21666 and w22080;
w22082 <= not w21346 and not w21355;
w22083 <= not w21666 and w22082;
w22084 <= not w21353 and not w22083;
w22085 <= not w22081 and not w22084;
w22086 <= w3758 and not w22066;
w22087 <= not w22076 and w22086;
w22088 <= not w22085 and not w22087;
w22089 <= not w22078 and not w22088;
w22090 <= not w3462 and not w22089;
w22091 <= w21365 and not w21367;
w22092 <= not w21358 and w22091;
w22093 <= not w21666 and w22092;
w22094 <= not w21358 and not w21367;
w22095 <= not w21666 and w22094;
w22096 <= not w21365 and not w22095;
w22097 <= not w22093 and not w22096;
w22098 <= w3462 and not w22078;
w22099 <= not w22088 and w22098;
w22100 <= not w22097 and not w22099;
w22101 <= not w22090 and not w22100;
w22102 <= not w3178 and not w22101;
w22103 <= not w21370 and w21377;
w22104 <= not w21379 and w22103;
w22105 <= not w21666 and w22104;
w22106 <= not w21370 and not w21379;
w22107 <= not w21666 and w22106;
w22108 <= not w21377 and not w22107;
w22109 <= not w22105 and not w22108;
w22110 <= w3178 and not w22090;
w22111 <= not w22100 and w22110;
w22112 <= not w22109 and not w22111;
w22113 <= not w22102 and not w22112;
w22114 <= not w2906 and not w22113;
w22115 <= w21389 and not w21391;
w22116 <= not w21382 and w22115;
w22117 <= not w21666 and w22116;
w22118 <= not w21382 and not w21391;
w22119 <= not w21666 and w22118;
w22120 <= not w21389 and not w22119;
w22121 <= not w22117 and not w22120;
w22122 <= w2906 and not w22102;
w22123 <= not w22112 and w22122;
w22124 <= not w22121 and not w22123;
w22125 <= not w22114 and not w22124;
w22126 <= not w2646 and not w22125;
w22127 <= not w21394 and w21401;
w22128 <= not w21403 and w22127;
w22129 <= not w21666 and w22128;
w22130 <= not w21394 and not w21403;
w22131 <= not w21666 and w22130;
w22132 <= not w21401 and not w22131;
w22133 <= not w22129 and not w22132;
w22134 <= w2646 and not w22114;
w22135 <= not w22124 and w22134;
w22136 <= not w22133 and not w22135;
w22137 <= not w22126 and not w22136;
w22138 <= not w2398 and not w22137;
w22139 <= w21413 and not w21415;
w22140 <= not w21406 and w22139;
w22141 <= not w21666 and w22140;
w22142 <= not w21406 and not w21415;
w22143 <= not w21666 and w22142;
w22144 <= not w21413 and not w22143;
w22145 <= not w22141 and not w22144;
w22146 <= w2398 and not w22126;
w22147 <= not w22136 and w22146;
w22148 <= not w22145 and not w22147;
w22149 <= not w22138 and not w22148;
w22150 <= not w2162 and not w22149;
w22151 <= not w21418 and w21425;
w22152 <= not w21427 and w22151;
w22153 <= not w21666 and w22152;
w22154 <= not w21418 and not w21427;
w22155 <= not w21666 and w22154;
w22156 <= not w21425 and not w22155;
w22157 <= not w22153 and not w22156;
w22158 <= w2162 and not w22138;
w22159 <= not w22148 and w22158;
w22160 <= not w22157 and not w22159;
w22161 <= not w22150 and not w22160;
w22162 <= not w1938 and not w22161;
w22163 <= w21437 and not w21439;
w22164 <= not w21430 and w22163;
w22165 <= not w21666 and w22164;
w22166 <= not w21430 and not w21439;
w22167 <= not w21666 and w22166;
w22168 <= not w21437 and not w22167;
w22169 <= not w22165 and not w22168;
w22170 <= w1938 and not w22150;
w22171 <= not w22160 and w22170;
w22172 <= not w22169 and not w22171;
w22173 <= not w22162 and not w22172;
w22174 <= not w1725 and not w22173;
w22175 <= not w21442 and w21449;
w22176 <= not w21451 and w22175;
w22177 <= not w21666 and w22176;
w22178 <= not w21442 and not w21451;
w22179 <= not w21666 and w22178;
w22180 <= not w21449 and not w22179;
w22181 <= not w22177 and not w22180;
w22182 <= w1725 and not w22162;
w22183 <= not w22172 and w22182;
w22184 <= not w22181 and not w22183;
w22185 <= not w22174 and not w22184;
w22186 <= not w1525 and not w22185;
w22187 <= w21461 and not w21463;
w22188 <= not w21454 and w22187;
w22189 <= not w21666 and w22188;
w22190 <= not w21454 and not w21463;
w22191 <= not w21666 and w22190;
w22192 <= not w21461 and not w22191;
w22193 <= not w22189 and not w22192;
w22194 <= w1525 and not w22174;
w22195 <= not w22184 and w22194;
w22196 <= not w22193 and not w22195;
w22197 <= not w22186 and not w22196;
w22198 <= not w1337 and not w22197;
w22199 <= not w21466 and w21473;
w22200 <= not w21475 and w22199;
w22201 <= not w21666 and w22200;
w22202 <= not w21466 and not w21475;
w22203 <= not w21666 and w22202;
w22204 <= not w21473 and not w22203;
w22205 <= not w22201 and not w22204;
w22206 <= w1337 and not w22186;
w22207 <= not w22196 and w22206;
w22208 <= not w22205 and not w22207;
w22209 <= not w22198 and not w22208;
w22210 <= not w1161 and not w22209;
w22211 <= w21485 and not w21487;
w22212 <= not w21478 and w22211;
w22213 <= not w21666 and w22212;
w22214 <= not w21478 and not w21487;
w22215 <= not w21666 and w22214;
w22216 <= not w21485 and not w22215;
w22217 <= not w22213 and not w22216;
w22218 <= w1161 and not w22198;
w22219 <= not w22208 and w22218;
w22220 <= not w22217 and not w22219;
w22221 <= not w22210 and not w22220;
w22222 <= not w997 and not w22221;
w22223 <= not w21490 and w21497;
w22224 <= not w21499 and w22223;
w22225 <= not w21666 and w22224;
w22226 <= not w21490 and not w21499;
w22227 <= not w21666 and w22226;
w22228 <= not w21497 and not w22227;
w22229 <= not w22225 and not w22228;
w22230 <= w997 and not w22210;
w22231 <= not w22220 and w22230;
w22232 <= not w22229 and not w22231;
w22233 <= not w22222 and not w22232;
w22234 <= not w845 and not w22233;
w22235 <= w21509 and not w21511;
w22236 <= not w21502 and w22235;
w22237 <= not w21666 and w22236;
w22238 <= not w21502 and not w21511;
w22239 <= not w21666 and w22238;
w22240 <= not w21509 and not w22239;
w22241 <= not w22237 and not w22240;
w22242 <= w845 and not w22222;
w22243 <= not w22232 and w22242;
w22244 <= not w22241 and not w22243;
w22245 <= not w22234 and not w22244;
w22246 <= not w705 and not w22245;
w22247 <= not w21514 and w21521;
w22248 <= not w21523 and w22247;
w22249 <= not w21666 and w22248;
w22250 <= not w21514 and not w21523;
w22251 <= not w21666 and w22250;
w22252 <= not w21521 and not w22251;
w22253 <= not w22249 and not w22252;
w22254 <= w705 and not w22234;
w22255 <= not w22244 and w22254;
w22256 <= not w22253 and not w22255;
w22257 <= not w22246 and not w22256;
w22258 <= not w577 and not w22257;
w22259 <= w21533 and not w21535;
w22260 <= not w21526 and w22259;
w22261 <= not w21666 and w22260;
w22262 <= not w21526 and not w21535;
w22263 <= not w21666 and w22262;
w22264 <= not w21533 and not w22263;
w22265 <= not w22261 and not w22264;
w22266 <= w577 and not w22246;
w22267 <= not w22256 and w22266;
w22268 <= not w22265 and not w22267;
w22269 <= not w22258 and not w22268;
w22270 <= not w460 and not w22269;
w22271 <= not w21538 and w21545;
w22272 <= not w21547 and w22271;
w22273 <= not w21666 and w22272;
w22274 <= not w21538 and not w21547;
w22275 <= not w21666 and w22274;
w22276 <= not w21545 and not w22275;
w22277 <= not w22273 and not w22276;
w22278 <= w460 and not w22258;
w22279 <= not w22268 and w22278;
w22280 <= not w22277 and not w22279;
w22281 <= not w22270 and not w22280;
w22282 <= not w356 and not w22281;
w22283 <= w21557 and not w21559;
w22284 <= not w21550 and w22283;
w22285 <= not w21666 and w22284;
w22286 <= not w21550 and not w21559;
w22287 <= not w21666 and w22286;
w22288 <= not w21557 and not w22287;
w22289 <= not w22285 and not w22288;
w22290 <= w356 and not w22270;
w22291 <= not w22280 and w22290;
w22292 <= not w22289 and not w22291;
w22293 <= not w22282 and not w22292;
w22294 <= not w264 and not w22293;
w22295 <= not w21562 and w21569;
w22296 <= not w21571 and w22295;
w22297 <= not w21666 and w22296;
w22298 <= not w21562 and not w21571;
w22299 <= not w21666 and w22298;
w22300 <= not w21569 and not w22299;
w22301 <= not w22297 and not w22300;
w22302 <= w264 and not w22282;
w22303 <= not w22292 and w22302;
w22304 <= not w22301 and not w22303;
w22305 <= not w22294 and not w22304;
w22306 <= not w184 and not w22305;
w22307 <= w21581 and not w21583;
w22308 <= not w21574 and w22307;
w22309 <= not w21666 and w22308;
w22310 <= not w21574 and not w21583;
w22311 <= not w21666 and w22310;
w22312 <= not w21581 and not w22311;
w22313 <= not w22309 and not w22312;
w22314 <= w184 and not w22294;
w22315 <= not w22304 and w22314;
w22316 <= not w22313 and not w22315;
w22317 <= not w22306 and not w22316;
w22318 <= not w115 and not w22317;
w22319 <= not w21586 and w21593;
w22320 <= not w21595 and w22319;
w22321 <= not w21666 and w22320;
w22322 <= not w21586 and not w21595;
w22323 <= not w21666 and w22322;
w22324 <= not w21593 and not w22323;
w22325 <= not w22321 and not w22324;
w22326 <= w115 and not w22306;
w22327 <= not w22316 and w22326;
w22328 <= not w22325 and not w22327;
w22329 <= not w22318 and not w22328;
w22330 <= not w60 and not w22329;
w22331 <= w21605 and not w21607;
w22332 <= not w21598 and w22331;
w22333 <= not w21666 and w22332;
w22334 <= not w21598 and not w21607;
w22335 <= not w21666 and w22334;
w22336 <= not w21605 and not w22335;
w22337 <= not w22333 and not w22336;
w22338 <= w60 and not w22318;
w22339 <= not w22328 and w22338;
w22340 <= not w22337 and not w22339;
w22341 <= not w22330 and not w22340;
w22342 <= not w22 and not w22341;
w22343 <= w22 and not w22330;
w22344 <= not w22340 and w22343;
w22345 <= not w21610 and w21619;
w22346 <= not w21612 and w22345;
w22347 <= not w21666 and w22346;
w22348 <= not w21610 and not w21612;
w22349 <= not w21666 and w22348;
w22350 <= not w21619 and not w22349;
w22351 <= not w22347 and not w22350;
w22352 <= not w22344 and not w22351;
w22353 <= not w22342 and not w22352;
w22354 <= not w5 and not w22353;
w22355 <= w21629 and not w21631;
w22356 <= not w21622 and w22355;
w22357 <= not w21666 and w22356;
w22358 <= not w21622 and not w21631;
w22359 <= not w21666 and w22358;
w22360 <= not w21629 and not w22359;
w22361 <= not w22357 and not w22360;
w22362 <= w5 and not w22342;
w22363 <= not w22352 and w22362;
w22364 <= not w22361 and not w22363;
w22365 <= not w22354 and not w22364;
w22366 <= not w21634 and w21641;
w22367 <= not w21643 and w22366;
w22368 <= not w21666 and w22367;
w22369 <= not w21634 and not w21643;
w22370 <= not w21666 and w22369;
w22371 <= not w21641 and not w22370;
w22372 <= not w22368 and not w22371;
w22373 <= not w21645 and not w21652;
w22374 <= not w21666 and w22373;
w22375 <= not w21660 and not w22374;
w22376 <= not w22372 and w22375;
w22377 <= not w22365 and w22376;
w22378 <= w0 and not w22377;
w22379 <= not w22354 and w22372;
w22380 <= not w22364 and w22379;
w22381 <= not w21652 and not w21666;
w22382 <= w21645 and not w22381;
w22383 <= not w0 and not w22373;
w22384 <= not w22382 and w22383;
w22385 <= not w22380 and not w22384;
w22386 <= not w22378 and w22385;
w22387 <= a(6) and not w22386;
w22388 <= not a(4) and not a(5);
w22389 <= not a(6) and w22388;
w22390 <= not w22387 and not w22389;
w22391 <= not w21666 and not w22390;
w22392 <= not w21664 and not w22389;
w22393 <= not w21660 and w22392;
w22394 <= not w21658 and w22393;
w22395 <= not w22387 and w22394;
w22396 <= not a(6) and not w22386;
w22397 <= a(7) and not w22396;
w22398 <= w21668 and not w22386;
w22399 <= not w22397 and not w22398;
w22400 <= not w22395 and w22399;
w22401 <= not w22391 and not w22400;
w22402 <= not w20957 and not w22401;
w22403 <= w20957 and not w22391;
w22404 <= not w22400 and w22403;
w22405 <= not w21666 and not w22384;
w22406 <= not w22380 and w22405;
w22407 <= not w22378 and w22406;
w22408 <= not w22398 and not w22407;
w22409 <= a(8) and not w22408;
w22410 <= not a(8) and not w22407;
w22411 <= not w22398 and w22410;
w22412 <= not w22409 and not w22411;
w22413 <= not w22404 and not w22412;
w22414 <= not w22402 and not w22413;
w22415 <= not w20259 and not w22414;
w22416 <= not w21671 and not w21675;
w22417 <= not w21679 and w22416;
w22418 <= not w22386 and w22417;
w22419 <= not w22386 and w22416;
w22420 <= w21679 and not w22419;
w22421 <= not w22418 and not w22420;
w22422 <= w20259 and not w22402;
w22423 <= not w22413 and w22422;
w22424 <= not w22421 and not w22423;
w22425 <= not w22415 and not w22424;
w22426 <= not w19567 and not w22425;
w22427 <= not w21684 and w21692;
w22428 <= not w21682 and w22427;
w22429 <= not w22386 and w22428;
w22430 <= not w21682 and not w21684;
w22431 <= not w22386 and w22430;
w22432 <= not w21692 and not w22431;
w22433 <= not w22429 and not w22432;
w22434 <= w19567 and not w22415;
w22435 <= not w22424 and w22434;
w22436 <= not w22433 and not w22435;
w22437 <= not w22426 and not w22436;
w22438 <= not w18887 and not w22437;
w22439 <= not w21695 and w21701;
w22440 <= not w21703 and w22439;
w22441 <= not w22386 and w22440;
w22442 <= not w21695 and not w21703;
w22443 <= not w22386 and w22442;
w22444 <= not w21701 and not w22443;
w22445 <= not w22441 and not w22444;
w22446 <= w18887 and not w22426;
w22447 <= not w22436 and w22446;
w22448 <= not w22445 and not w22447;
w22449 <= not w22438 and not w22448;
w22450 <= not w18219 and not w22449;
w22451 <= w21713 and not w21715;
w22452 <= not w21706 and w22451;
w22453 <= not w22386 and w22452;
w22454 <= not w21706 and not w21715;
w22455 <= not w22386 and w22454;
w22456 <= not w21713 and not w22455;
w22457 <= not w22453 and not w22456;
w22458 <= w18219 and not w22438;
w22459 <= not w22448 and w22458;
w22460 <= not w22457 and not w22459;
w22461 <= not w22450 and not w22460;
w22462 <= not w17563 and not w22461;
w22463 <= not w21718 and w21725;
w22464 <= not w21727 and w22463;
w22465 <= not w22386 and w22464;
w22466 <= not w21718 and not w21727;
w22467 <= not w22386 and w22466;
w22468 <= not w21725 and not w22467;
w22469 <= not w22465 and not w22468;
w22470 <= w17563 and not w22450;
w22471 <= not w22460 and w22470;
w22472 <= not w22469 and not w22471;
w22473 <= not w22462 and not w22472;
w22474 <= not w16919 and not w22473;
w22475 <= w21737 and not w21739;
w22476 <= not w21730 and w22475;
w22477 <= not w22386 and w22476;
w22478 <= not w21730 and not w21739;
w22479 <= not w22386 and w22478;
w22480 <= not w21737 and not w22479;
w22481 <= not w22477 and not w22480;
w22482 <= w16919 and not w22462;
w22483 <= not w22472 and w22482;
w22484 <= not w22481 and not w22483;
w22485 <= not w22474 and not w22484;
w22486 <= not w16287 and not w22485;
w22487 <= not w21742 and w21749;
w22488 <= not w21751 and w22487;
w22489 <= not w22386 and w22488;
w22490 <= not w21742 and not w21751;
w22491 <= not w22386 and w22490;
w22492 <= not w21749 and not w22491;
w22493 <= not w22489 and not w22492;
w22494 <= w16287 and not w22474;
w22495 <= not w22484 and w22494;
w22496 <= not w22493 and not w22495;
w22497 <= not w22486 and not w22496;
w22498 <= not w15667 and not w22497;
w22499 <= w21761 and not w21763;
w22500 <= not w21754 and w22499;
w22501 <= not w22386 and w22500;
w22502 <= not w21754 and not w21763;
w22503 <= not w22386 and w22502;
w22504 <= not w21761 and not w22503;
w22505 <= not w22501 and not w22504;
w22506 <= w15667 and not w22486;
w22507 <= not w22496 and w22506;
w22508 <= not w22505 and not w22507;
w22509 <= not w22498 and not w22508;
w22510 <= not w15059 and not w22509;
w22511 <= not w21766 and w21773;
w22512 <= not w21775 and w22511;
w22513 <= not w22386 and w22512;
w22514 <= not w21766 and not w21775;
w22515 <= not w22386 and w22514;
w22516 <= not w21773 and not w22515;
w22517 <= not w22513 and not w22516;
w22518 <= w15059 and not w22498;
w22519 <= not w22508 and w22518;
w22520 <= not w22517 and not w22519;
w22521 <= not w22510 and not w22520;
w22522 <= not w14463 and not w22521;
w22523 <= w21785 and not w21787;
w22524 <= not w21778 and w22523;
w22525 <= not w22386 and w22524;
w22526 <= not w21778 and not w21787;
w22527 <= not w22386 and w22526;
w22528 <= not w21785 and not w22527;
w22529 <= not w22525 and not w22528;
w22530 <= w14463 and not w22510;
w22531 <= not w22520 and w22530;
w22532 <= not w22529 and not w22531;
w22533 <= not w22522 and not w22532;
w22534 <= not w13879 and not w22533;
w22535 <= not w21790 and w21797;
w22536 <= not w21799 and w22535;
w22537 <= not w22386 and w22536;
w22538 <= not w21790 and not w21799;
w22539 <= not w22386 and w22538;
w22540 <= not w21797 and not w22539;
w22541 <= not w22537 and not w22540;
w22542 <= w13879 and not w22522;
w22543 <= not w22532 and w22542;
w22544 <= not w22541 and not w22543;
w22545 <= not w22534 and not w22544;
w22546 <= not w13307 and not w22545;
w22547 <= w21809 and not w21811;
w22548 <= not w21802 and w22547;
w22549 <= not w22386 and w22548;
w22550 <= not w21802 and not w21811;
w22551 <= not w22386 and w22550;
w22552 <= not w21809 and not w22551;
w22553 <= not w22549 and not w22552;
w22554 <= w13307 and not w22534;
w22555 <= not w22544 and w22554;
w22556 <= not w22553 and not w22555;
w22557 <= not w22546 and not w22556;
w22558 <= not w12747 and not w22557;
w22559 <= not w21814 and w21821;
w22560 <= not w21823 and w22559;
w22561 <= not w22386 and w22560;
w22562 <= not w21814 and not w21823;
w22563 <= not w22386 and w22562;
w22564 <= not w21821 and not w22563;
w22565 <= not w22561 and not w22564;
w22566 <= w12747 and not w22546;
w22567 <= not w22556 and w22566;
w22568 <= not w22565 and not w22567;
w22569 <= not w22558 and not w22568;
w22570 <= not w12199 and not w22569;
w22571 <= w21833 and not w21835;
w22572 <= not w21826 and w22571;
w22573 <= not w22386 and w22572;
w22574 <= not w21826 and not w21835;
w22575 <= not w22386 and w22574;
w22576 <= not w21833 and not w22575;
w22577 <= not w22573 and not w22576;
w22578 <= w12199 and not w22558;
w22579 <= not w22568 and w22578;
w22580 <= not w22577 and not w22579;
w22581 <= not w22570 and not w22580;
w22582 <= not w11663 and not w22581;
w22583 <= not w21838 and w21845;
w22584 <= not w21847 and w22583;
w22585 <= not w22386 and w22584;
w22586 <= not w21838 and not w21847;
w22587 <= not w22386 and w22586;
w22588 <= not w21845 and not w22587;
w22589 <= not w22585 and not w22588;
w22590 <= w11663 and not w22570;
w22591 <= not w22580 and w22590;
w22592 <= not w22589 and not w22591;
w22593 <= not w22582 and not w22592;
w22594 <= not w11139 and not w22593;
w22595 <= w21857 and not w21859;
w22596 <= not w21850 and w22595;
w22597 <= not w22386 and w22596;
w22598 <= not w21850 and not w21859;
w22599 <= not w22386 and w22598;
w22600 <= not w21857 and not w22599;
w22601 <= not w22597 and not w22600;
w22602 <= w11139 and not w22582;
w22603 <= not w22592 and w22602;
w22604 <= not w22601 and not w22603;
w22605 <= not w22594 and not w22604;
w22606 <= not w10627 and not w22605;
w22607 <= not w21862 and w21869;
w22608 <= not w21871 and w22607;
w22609 <= not w22386 and w22608;
w22610 <= not w21862 and not w21871;
w22611 <= not w22386 and w22610;
w22612 <= not w21869 and not w22611;
w22613 <= not w22609 and not w22612;
w22614 <= w10627 and not w22594;
w22615 <= not w22604 and w22614;
w22616 <= not w22613 and not w22615;
w22617 <= not w22606 and not w22616;
w22618 <= not w10127 and not w22617;
w22619 <= w21881 and not w21883;
w22620 <= not w21874 and w22619;
w22621 <= not w22386 and w22620;
w22622 <= not w21874 and not w21883;
w22623 <= not w22386 and w22622;
w22624 <= not w21881 and not w22623;
w22625 <= not w22621 and not w22624;
w22626 <= w10127 and not w22606;
w22627 <= not w22616 and w22626;
w22628 <= not w22625 and not w22627;
w22629 <= not w22618 and not w22628;
w22630 <= not w9639 and not w22629;
w22631 <= not w21886 and w21893;
w22632 <= not w21895 and w22631;
w22633 <= not w22386 and w22632;
w22634 <= not w21886 and not w21895;
w22635 <= not w22386 and w22634;
w22636 <= not w21893 and not w22635;
w22637 <= not w22633 and not w22636;
w22638 <= w9639 and not w22618;
w22639 <= not w22628 and w22638;
w22640 <= not w22637 and not w22639;
w22641 <= not w22630 and not w22640;
w22642 <= not w9163 and not w22641;
w22643 <= w21905 and not w21907;
w22644 <= not w21898 and w22643;
w22645 <= not w22386 and w22644;
w22646 <= not w21898 and not w21907;
w22647 <= not w22386 and w22646;
w22648 <= not w21905 and not w22647;
w22649 <= not w22645 and not w22648;
w22650 <= w9163 and not w22630;
w22651 <= not w22640 and w22650;
w22652 <= not w22649 and not w22651;
w22653 <= not w22642 and not w22652;
w22654 <= not w8699 and not w22653;
w22655 <= not w21910 and w21917;
w22656 <= not w21919 and w22655;
w22657 <= not w22386 and w22656;
w22658 <= not w21910 and not w21919;
w22659 <= not w22386 and w22658;
w22660 <= not w21917 and not w22659;
w22661 <= not w22657 and not w22660;
w22662 <= w8699 and not w22642;
w22663 <= not w22652 and w22662;
w22664 <= not w22661 and not w22663;
w22665 <= not w22654 and not w22664;
w22666 <= not w8247 and not w22665;
w22667 <= w21929 and not w21931;
w22668 <= not w21922 and w22667;
w22669 <= not w22386 and w22668;
w22670 <= not w21922 and not w21931;
w22671 <= not w22386 and w22670;
w22672 <= not w21929 and not w22671;
w22673 <= not w22669 and not w22672;
w22674 <= w8247 and not w22654;
w22675 <= not w22664 and w22674;
w22676 <= not w22673 and not w22675;
w22677 <= not w22666 and not w22676;
w22678 <= not w7807 and not w22677;
w22679 <= not w21934 and w21941;
w22680 <= not w21943 and w22679;
w22681 <= not w22386 and w22680;
w22682 <= not w21934 and not w21943;
w22683 <= not w22386 and w22682;
w22684 <= not w21941 and not w22683;
w22685 <= not w22681 and not w22684;
w22686 <= w7807 and not w22666;
w22687 <= not w22676 and w22686;
w22688 <= not w22685 and not w22687;
w22689 <= not w22678 and not w22688;
w22690 <= not w7379 and not w22689;
w22691 <= w21953 and not w21955;
w22692 <= not w21946 and w22691;
w22693 <= not w22386 and w22692;
w22694 <= not w21946 and not w21955;
w22695 <= not w22386 and w22694;
w22696 <= not w21953 and not w22695;
w22697 <= not w22693 and not w22696;
w22698 <= w7379 and not w22678;
w22699 <= not w22688 and w22698;
w22700 <= not w22697 and not w22699;
w22701 <= not w22690 and not w22700;
w22702 <= not w6963 and not w22701;
w22703 <= not w21958 and w21965;
w22704 <= not w21967 and w22703;
w22705 <= not w22386 and w22704;
w22706 <= not w21958 and not w21967;
w22707 <= not w22386 and w22706;
w22708 <= not w21965 and not w22707;
w22709 <= not w22705 and not w22708;
w22710 <= w6963 and not w22690;
w22711 <= not w22700 and w22710;
w22712 <= not w22709 and not w22711;
w22713 <= not w22702 and not w22712;
w22714 <= not w6558 and not w22713;
w22715 <= w21977 and not w21979;
w22716 <= not w21970 and w22715;
w22717 <= not w22386 and w22716;
w22718 <= not w21970 and not w21979;
w22719 <= not w22386 and w22718;
w22720 <= not w21977 and not w22719;
w22721 <= not w22717 and not w22720;
w22722 <= w6558 and not w22702;
w22723 <= not w22712 and w22722;
w22724 <= not w22721 and not w22723;
w22725 <= not w22714 and not w22724;
w22726 <= not w6166 and not w22725;
w22727 <= not w21982 and w21989;
w22728 <= not w21991 and w22727;
w22729 <= not w22386 and w22728;
w22730 <= not w21982 and not w21991;
w22731 <= not w22386 and w22730;
w22732 <= not w21989 and not w22731;
w22733 <= not w22729 and not w22732;
w22734 <= w6166 and not w22714;
w22735 <= not w22724 and w22734;
w22736 <= not w22733 and not w22735;
w22737 <= not w22726 and not w22736;
w22738 <= not w5786 and not w22737;
w22739 <= w22001 and not w22003;
w22740 <= not w21994 and w22739;
w22741 <= not w22386 and w22740;
w22742 <= not w21994 and not w22003;
w22743 <= not w22386 and w22742;
w22744 <= not w22001 and not w22743;
w22745 <= not w22741 and not w22744;
w22746 <= w5786 and not w22726;
w22747 <= not w22736 and w22746;
w22748 <= not w22745 and not w22747;
w22749 <= not w22738 and not w22748;
w22750 <= not w5418 and not w22749;
w22751 <= not w22006 and w22013;
w22752 <= not w22015 and w22751;
w22753 <= not w22386 and w22752;
w22754 <= not w22006 and not w22015;
w22755 <= not w22386 and w22754;
w22756 <= not w22013 and not w22755;
w22757 <= not w22753 and not w22756;
w22758 <= w5418 and not w22738;
w22759 <= not w22748 and w22758;
w22760 <= not w22757 and not w22759;
w22761 <= not w22750 and not w22760;
w22762 <= not w5062 and not w22761;
w22763 <= w22025 and not w22027;
w22764 <= not w22018 and w22763;
w22765 <= not w22386 and w22764;
w22766 <= not w22018 and not w22027;
w22767 <= not w22386 and w22766;
w22768 <= not w22025 and not w22767;
w22769 <= not w22765 and not w22768;
w22770 <= w5062 and not w22750;
w22771 <= not w22760 and w22770;
w22772 <= not w22769 and not w22771;
w22773 <= not w22762 and not w22772;
w22774 <= not w4718 and not w22773;
w22775 <= not w22030 and w22037;
w22776 <= not w22039 and w22775;
w22777 <= not w22386 and w22776;
w22778 <= not w22030 and not w22039;
w22779 <= not w22386 and w22778;
w22780 <= not w22037 and not w22779;
w22781 <= not w22777 and not w22780;
w22782 <= w4718 and not w22762;
w22783 <= not w22772 and w22782;
w22784 <= not w22781 and not w22783;
w22785 <= not w22774 and not w22784;
w22786 <= not w4386 and not w22785;
w22787 <= w22049 and not w22051;
w22788 <= not w22042 and w22787;
w22789 <= not w22386 and w22788;
w22790 <= not w22042 and not w22051;
w22791 <= not w22386 and w22790;
w22792 <= not w22049 and not w22791;
w22793 <= not w22789 and not w22792;
w22794 <= w4386 and not w22774;
w22795 <= not w22784 and w22794;
w22796 <= not w22793 and not w22795;
w22797 <= not w22786 and not w22796;
w22798 <= not w4066 and not w22797;
w22799 <= not w22054 and w22061;
w22800 <= not w22063 and w22799;
w22801 <= not w22386 and w22800;
w22802 <= not w22054 and not w22063;
w22803 <= not w22386 and w22802;
w22804 <= not w22061 and not w22803;
w22805 <= not w22801 and not w22804;
w22806 <= w4066 and not w22786;
w22807 <= not w22796 and w22806;
w22808 <= not w22805 and not w22807;
w22809 <= not w22798 and not w22808;
w22810 <= not w3758 and not w22809;
w22811 <= w22073 and not w22075;
w22812 <= not w22066 and w22811;
w22813 <= not w22386 and w22812;
w22814 <= not w22066 and not w22075;
w22815 <= not w22386 and w22814;
w22816 <= not w22073 and not w22815;
w22817 <= not w22813 and not w22816;
w22818 <= w3758 and not w22798;
w22819 <= not w22808 and w22818;
w22820 <= not w22817 and not w22819;
w22821 <= not w22810 and not w22820;
w22822 <= not w3462 and not w22821;
w22823 <= not w22078 and w22085;
w22824 <= not w22087 and w22823;
w22825 <= not w22386 and w22824;
w22826 <= not w22078 and not w22087;
w22827 <= not w22386 and w22826;
w22828 <= not w22085 and not w22827;
w22829 <= not w22825 and not w22828;
w22830 <= w3462 and not w22810;
w22831 <= not w22820 and w22830;
w22832 <= not w22829 and not w22831;
w22833 <= not w22822 and not w22832;
w22834 <= not w3178 and not w22833;
w22835 <= w22097 and not w22099;
w22836 <= not w22090 and w22835;
w22837 <= not w22386 and w22836;
w22838 <= not w22090 and not w22099;
w22839 <= not w22386 and w22838;
w22840 <= not w22097 and not w22839;
w22841 <= not w22837 and not w22840;
w22842 <= w3178 and not w22822;
w22843 <= not w22832 and w22842;
w22844 <= not w22841 and not w22843;
w22845 <= not w22834 and not w22844;
w22846 <= not w2906 and not w22845;
w22847 <= not w22102 and w22109;
w22848 <= not w22111 and w22847;
w22849 <= not w22386 and w22848;
w22850 <= not w22102 and not w22111;
w22851 <= not w22386 and w22850;
w22852 <= not w22109 and not w22851;
w22853 <= not w22849 and not w22852;
w22854 <= w2906 and not w22834;
w22855 <= not w22844 and w22854;
w22856 <= not w22853 and not w22855;
w22857 <= not w22846 and not w22856;
w22858 <= not w2646 and not w22857;
w22859 <= w22121 and not w22123;
w22860 <= not w22114 and w22859;
w22861 <= not w22386 and w22860;
w22862 <= not w22114 and not w22123;
w22863 <= not w22386 and w22862;
w22864 <= not w22121 and not w22863;
w22865 <= not w22861 and not w22864;
w22866 <= w2646 and not w22846;
w22867 <= not w22856 and w22866;
w22868 <= not w22865 and not w22867;
w22869 <= not w22858 and not w22868;
w22870 <= not w2398 and not w22869;
w22871 <= not w22126 and w22133;
w22872 <= not w22135 and w22871;
w22873 <= not w22386 and w22872;
w22874 <= not w22126 and not w22135;
w22875 <= not w22386 and w22874;
w22876 <= not w22133 and not w22875;
w22877 <= not w22873 and not w22876;
w22878 <= w2398 and not w22858;
w22879 <= not w22868 and w22878;
w22880 <= not w22877 and not w22879;
w22881 <= not w22870 and not w22880;
w22882 <= not w2162 and not w22881;
w22883 <= w22145 and not w22147;
w22884 <= not w22138 and w22883;
w22885 <= not w22386 and w22884;
w22886 <= not w22138 and not w22147;
w22887 <= not w22386 and w22886;
w22888 <= not w22145 and not w22887;
w22889 <= not w22885 and not w22888;
w22890 <= w2162 and not w22870;
w22891 <= not w22880 and w22890;
w22892 <= not w22889 and not w22891;
w22893 <= not w22882 and not w22892;
w22894 <= not w1938 and not w22893;
w22895 <= not w22150 and w22157;
w22896 <= not w22159 and w22895;
w22897 <= not w22386 and w22896;
w22898 <= not w22150 and not w22159;
w22899 <= not w22386 and w22898;
w22900 <= not w22157 and not w22899;
w22901 <= not w22897 and not w22900;
w22902 <= w1938 and not w22882;
w22903 <= not w22892 and w22902;
w22904 <= not w22901 and not w22903;
w22905 <= not w22894 and not w22904;
w22906 <= not w1725 and not w22905;
w22907 <= w22169 and not w22171;
w22908 <= not w22162 and w22907;
w22909 <= not w22386 and w22908;
w22910 <= not w22162 and not w22171;
w22911 <= not w22386 and w22910;
w22912 <= not w22169 and not w22911;
w22913 <= not w22909 and not w22912;
w22914 <= w1725 and not w22894;
w22915 <= not w22904 and w22914;
w22916 <= not w22913 and not w22915;
w22917 <= not w22906 and not w22916;
w22918 <= not w1525 and not w22917;
w22919 <= not w22174 and w22181;
w22920 <= not w22183 and w22919;
w22921 <= not w22386 and w22920;
w22922 <= not w22174 and not w22183;
w22923 <= not w22386 and w22922;
w22924 <= not w22181 and not w22923;
w22925 <= not w22921 and not w22924;
w22926 <= w1525 and not w22906;
w22927 <= not w22916 and w22926;
w22928 <= not w22925 and not w22927;
w22929 <= not w22918 and not w22928;
w22930 <= not w1337 and not w22929;
w22931 <= w22193 and not w22195;
w22932 <= not w22186 and w22931;
w22933 <= not w22386 and w22932;
w22934 <= not w22186 and not w22195;
w22935 <= not w22386 and w22934;
w22936 <= not w22193 and not w22935;
w22937 <= not w22933 and not w22936;
w22938 <= w1337 and not w22918;
w22939 <= not w22928 and w22938;
w22940 <= not w22937 and not w22939;
w22941 <= not w22930 and not w22940;
w22942 <= not w1161 and not w22941;
w22943 <= not w22198 and w22205;
w22944 <= not w22207 and w22943;
w22945 <= not w22386 and w22944;
w22946 <= not w22198 and not w22207;
w22947 <= not w22386 and w22946;
w22948 <= not w22205 and not w22947;
w22949 <= not w22945 and not w22948;
w22950 <= w1161 and not w22930;
w22951 <= not w22940 and w22950;
w22952 <= not w22949 and not w22951;
w22953 <= not w22942 and not w22952;
w22954 <= not w997 and not w22953;
w22955 <= w22217 and not w22219;
w22956 <= not w22210 and w22955;
w22957 <= not w22386 and w22956;
w22958 <= not w22210 and not w22219;
w22959 <= not w22386 and w22958;
w22960 <= not w22217 and not w22959;
w22961 <= not w22957 and not w22960;
w22962 <= w997 and not w22942;
w22963 <= not w22952 and w22962;
w22964 <= not w22961 and not w22963;
w22965 <= not w22954 and not w22964;
w22966 <= not w845 and not w22965;
w22967 <= not w22222 and w22229;
w22968 <= not w22231 and w22967;
w22969 <= not w22386 and w22968;
w22970 <= not w22222 and not w22231;
w22971 <= not w22386 and w22970;
w22972 <= not w22229 and not w22971;
w22973 <= not w22969 and not w22972;
w22974 <= w845 and not w22954;
w22975 <= not w22964 and w22974;
w22976 <= not w22973 and not w22975;
w22977 <= not w22966 and not w22976;
w22978 <= not w705 and not w22977;
w22979 <= w22241 and not w22243;
w22980 <= not w22234 and w22979;
w22981 <= not w22386 and w22980;
w22982 <= not w22234 and not w22243;
w22983 <= not w22386 and w22982;
w22984 <= not w22241 and not w22983;
w22985 <= not w22981 and not w22984;
w22986 <= w705 and not w22966;
w22987 <= not w22976 and w22986;
w22988 <= not w22985 and not w22987;
w22989 <= not w22978 and not w22988;
w22990 <= not w577 and not w22989;
w22991 <= not w22246 and w22253;
w22992 <= not w22255 and w22991;
w22993 <= not w22386 and w22992;
w22994 <= not w22246 and not w22255;
w22995 <= not w22386 and w22994;
w22996 <= not w22253 and not w22995;
w22997 <= not w22993 and not w22996;
w22998 <= w577 and not w22978;
w22999 <= not w22988 and w22998;
w23000 <= not w22997 and not w22999;
w23001 <= not w22990 and not w23000;
w23002 <= not w460 and not w23001;
w23003 <= w22265 and not w22267;
w23004 <= not w22258 and w23003;
w23005 <= not w22386 and w23004;
w23006 <= not w22258 and not w22267;
w23007 <= not w22386 and w23006;
w23008 <= not w22265 and not w23007;
w23009 <= not w23005 and not w23008;
w23010 <= w460 and not w22990;
w23011 <= not w23000 and w23010;
w23012 <= not w23009 and not w23011;
w23013 <= not w23002 and not w23012;
w23014 <= not w356 and not w23013;
w23015 <= not w22270 and w22277;
w23016 <= not w22279 and w23015;
w23017 <= not w22386 and w23016;
w23018 <= not w22270 and not w22279;
w23019 <= not w22386 and w23018;
w23020 <= not w22277 and not w23019;
w23021 <= not w23017 and not w23020;
w23022 <= w356 and not w23002;
w23023 <= not w23012 and w23022;
w23024 <= not w23021 and not w23023;
w23025 <= not w23014 and not w23024;
w23026 <= not w264 and not w23025;
w23027 <= w22289 and not w22291;
w23028 <= not w22282 and w23027;
w23029 <= not w22386 and w23028;
w23030 <= not w22282 and not w22291;
w23031 <= not w22386 and w23030;
w23032 <= not w22289 and not w23031;
w23033 <= not w23029 and not w23032;
w23034 <= w264 and not w23014;
w23035 <= not w23024 and w23034;
w23036 <= not w23033 and not w23035;
w23037 <= not w23026 and not w23036;
w23038 <= not w184 and not w23037;
w23039 <= not w22294 and w22301;
w23040 <= not w22303 and w23039;
w23041 <= not w22386 and w23040;
w23042 <= not w22294 and not w22303;
w23043 <= not w22386 and w23042;
w23044 <= not w22301 and not w23043;
w23045 <= not w23041 and not w23044;
w23046 <= w184 and not w23026;
w23047 <= not w23036 and w23046;
w23048 <= not w23045 and not w23047;
w23049 <= not w23038 and not w23048;
w23050 <= not w115 and not w23049;
w23051 <= w22313 and not w22315;
w23052 <= not w22306 and w23051;
w23053 <= not w22386 and w23052;
w23054 <= not w22306 and not w22315;
w23055 <= not w22386 and w23054;
w23056 <= not w22313 and not w23055;
w23057 <= not w23053 and not w23056;
w23058 <= w115 and not w23038;
w23059 <= not w23048 and w23058;
w23060 <= not w23057 and not w23059;
w23061 <= not w23050 and not w23060;
w23062 <= not w60 and not w23061;
w23063 <= not w22318 and w22325;
w23064 <= not w22327 and w23063;
w23065 <= not w22386 and w23064;
w23066 <= not w22318 and not w22327;
w23067 <= not w22386 and w23066;
w23068 <= not w22325 and not w23067;
w23069 <= not w23065 and not w23068;
w23070 <= w60 and not w23050;
w23071 <= not w23060 and w23070;
w23072 <= not w23069 and not w23071;
w23073 <= not w23062 and not w23072;
w23074 <= not w22 and not w23073;
w23075 <= w22337 and not w22339;
w23076 <= not w22330 and w23075;
w23077 <= not w22386 and w23076;
w23078 <= not w22330 and not w22339;
w23079 <= not w22386 and w23078;
w23080 <= not w22337 and not w23079;
w23081 <= not w23077 and not w23080;
w23082 <= w22 and not w23062;
w23083 <= not w23072 and w23082;
w23084 <= not w23081 and not w23083;
w23085 <= not w23074 and not w23084;
w23086 <= not w5 and not w23085;
w23087 <= w5 and not w23074;
w23088 <= not w23084 and w23087;
w23089 <= not w22342 and w22351;
w23090 <= not w22344 and w23089;
w23091 <= not w22386 and w23090;
w23092 <= not w22342 and not w22344;
w23093 <= not w22386 and w23092;
w23094 <= not w22351 and not w23093;
w23095 <= not w23091 and not w23094;
w23096 <= not w23088 and not w23095;
w23097 <= not w23086 and not w23096;
w23098 <= w22361 and not w22363;
w23099 <= not w22354 and w23098;
w23100 <= not w22386 and w23099;
w23101 <= not w22354 and not w22363;
w23102 <= not w22386 and w23101;
w23103 <= not w22361 and not w23102;
w23104 <= not w23100 and not w23103;
w23105 <= not w22365 and not w22372;
w23106 <= not w22386 and w23105;
w23107 <= not w22380 and not w23106;
w23108 <= not w23104 and w23107;
w23109 <= not w23097 and w23108;
w23110 <= w0 and not w23109;
w23111 <= not w23086 and w23104;
w23112 <= not w23096 and w23111;
w23113 <= not w22372 and not w22386;
w23114 <= w22365 and not w23113;
w23115 <= not w0 and not w23105;
w23116 <= not w23114 and w23115;
w23117 <= not w23112 and not w23116;
w23118 <= not w23110 and w23117;
w23119 <= not w23062 and w23069;
w23120 <= not w23071 and w23119;
w23121 <= not w23118 and w23120;
w23122 <= not w23062 and not w23071;
w23123 <= not w23118 and w23122;
w23124 <= not w23069 and not w23123;
w23125 <= not w23121 and not w23124;
w23126 <= a(4) and not w23118;
w23127 <= not a(2) and not a(3);
w23128 <= not a(4) and w23127;
w23129 <= not w23126 and not w23128;
w23130 <= not w22386 and not w23129;
w23131 <= not w22384 and not w23128;
w23132 <= not w22380 and w23131;
w23133 <= not w22378 and w23132;
w23134 <= not w23126 and w23133;
w23135 <= not a(4) and not w23118;
w23136 <= a(5) and not w23135;
w23137 <= w22388 and not w23118;
w23138 <= not w23136 and not w23137;
w23139 <= not w23134 and w23138;
w23140 <= not w23130 and not w23139;
w23141 <= not w21666 and not w23140;
w23142 <= w21666 and not w23130;
w23143 <= not w23139 and w23142;
w23144 <= not w22386 and not w23116;
w23145 <= not w23112 and w23144;
w23146 <= not w23110 and w23145;
w23147 <= not w23137 and not w23146;
w23148 <= a(6) and not w23147;
w23149 <= not a(6) and not w23146;
w23150 <= not w23137 and w23149;
w23151 <= not w23148 and not w23150;
w23152 <= not w23143 and not w23151;
w23153 <= not w23141 and not w23152;
w23154 <= not w20957 and not w23153;
w23155 <= not w22391 and not w22395;
w23156 <= not w22399 and w23155;
w23157 <= not w23118 and w23156;
w23158 <= not w23118 and w23155;
w23159 <= w22399 and not w23158;
w23160 <= not w23157 and not w23159;
w23161 <= w20957 and not w23141;
w23162 <= not w23152 and w23161;
w23163 <= not w23160 and not w23162;
w23164 <= not w23154 and not w23163;
w23165 <= not w20259 and not w23164;
w23166 <= not w22404 and w22412;
w23167 <= not w22402 and w23166;
w23168 <= not w23118 and w23167;
w23169 <= not w22402 and not w22404;
w23170 <= not w23118 and w23169;
w23171 <= not w22412 and not w23170;
w23172 <= not w23168 and not w23171;
w23173 <= w20259 and not w23154;
w23174 <= not w23163 and w23173;
w23175 <= not w23172 and not w23174;
w23176 <= not w23165 and not w23175;
w23177 <= not w19567 and not w23176;
w23178 <= not w22415 and w22421;
w23179 <= not w22423 and w23178;
w23180 <= not w23118 and w23179;
w23181 <= not w22415 and not w22423;
w23182 <= not w23118 and w23181;
w23183 <= not w22421 and not w23182;
w23184 <= not w23180 and not w23183;
w23185 <= w19567 and not w23165;
w23186 <= not w23175 and w23185;
w23187 <= not w23184 and not w23186;
w23188 <= not w23177 and not w23187;
w23189 <= not w18887 and not w23188;
w23190 <= w22433 and not w22435;
w23191 <= not w22426 and w23190;
w23192 <= not w23118 and w23191;
w23193 <= not w22426 and not w22435;
w23194 <= not w23118 and w23193;
w23195 <= not w22433 and not w23194;
w23196 <= not w23192 and not w23195;
w23197 <= w18887 and not w23177;
w23198 <= not w23187 and w23197;
w23199 <= not w23196 and not w23198;
w23200 <= not w23189 and not w23199;
w23201 <= not w18219 and not w23200;
w23202 <= not w22438 and w22445;
w23203 <= not w22447 and w23202;
w23204 <= not w23118 and w23203;
w23205 <= not w22438 and not w22447;
w23206 <= not w23118 and w23205;
w23207 <= not w22445 and not w23206;
w23208 <= not w23204 and not w23207;
w23209 <= w18219 and not w23189;
w23210 <= not w23199 and w23209;
w23211 <= not w23208 and not w23210;
w23212 <= not w23201 and not w23211;
w23213 <= not w17563 and not w23212;
w23214 <= w22457 and not w22459;
w23215 <= not w22450 and w23214;
w23216 <= not w23118 and w23215;
w23217 <= not w22450 and not w22459;
w23218 <= not w23118 and w23217;
w23219 <= not w22457 and not w23218;
w23220 <= not w23216 and not w23219;
w23221 <= w17563 and not w23201;
w23222 <= not w23211 and w23221;
w23223 <= not w23220 and not w23222;
w23224 <= not w23213 and not w23223;
w23225 <= not w16919 and not w23224;
w23226 <= not w22462 and w22469;
w23227 <= not w22471 and w23226;
w23228 <= not w23118 and w23227;
w23229 <= not w22462 and not w22471;
w23230 <= not w23118 and w23229;
w23231 <= not w22469 and not w23230;
w23232 <= not w23228 and not w23231;
w23233 <= w16919 and not w23213;
w23234 <= not w23223 and w23233;
w23235 <= not w23232 and not w23234;
w23236 <= not w23225 and not w23235;
w23237 <= not w16287 and not w23236;
w23238 <= w22481 and not w22483;
w23239 <= not w22474 and w23238;
w23240 <= not w23118 and w23239;
w23241 <= not w22474 and not w22483;
w23242 <= not w23118 and w23241;
w23243 <= not w22481 and not w23242;
w23244 <= not w23240 and not w23243;
w23245 <= w16287 and not w23225;
w23246 <= not w23235 and w23245;
w23247 <= not w23244 and not w23246;
w23248 <= not w23237 and not w23247;
w23249 <= not w15667 and not w23248;
w23250 <= not w22486 and w22493;
w23251 <= not w22495 and w23250;
w23252 <= not w23118 and w23251;
w23253 <= not w22486 and not w22495;
w23254 <= not w23118 and w23253;
w23255 <= not w22493 and not w23254;
w23256 <= not w23252 and not w23255;
w23257 <= w15667 and not w23237;
w23258 <= not w23247 and w23257;
w23259 <= not w23256 and not w23258;
w23260 <= not w23249 and not w23259;
w23261 <= not w15059 and not w23260;
w23262 <= w22505 and not w22507;
w23263 <= not w22498 and w23262;
w23264 <= not w23118 and w23263;
w23265 <= not w22498 and not w22507;
w23266 <= not w23118 and w23265;
w23267 <= not w22505 and not w23266;
w23268 <= not w23264 and not w23267;
w23269 <= w15059 and not w23249;
w23270 <= not w23259 and w23269;
w23271 <= not w23268 and not w23270;
w23272 <= not w23261 and not w23271;
w23273 <= not w14463 and not w23272;
w23274 <= not w22510 and w22517;
w23275 <= not w22519 and w23274;
w23276 <= not w23118 and w23275;
w23277 <= not w22510 and not w22519;
w23278 <= not w23118 and w23277;
w23279 <= not w22517 and not w23278;
w23280 <= not w23276 and not w23279;
w23281 <= w14463 and not w23261;
w23282 <= not w23271 and w23281;
w23283 <= not w23280 and not w23282;
w23284 <= not w23273 and not w23283;
w23285 <= not w13879 and not w23284;
w23286 <= w22529 and not w22531;
w23287 <= not w22522 and w23286;
w23288 <= not w23118 and w23287;
w23289 <= not w22522 and not w22531;
w23290 <= not w23118 and w23289;
w23291 <= not w22529 and not w23290;
w23292 <= not w23288 and not w23291;
w23293 <= w13879 and not w23273;
w23294 <= not w23283 and w23293;
w23295 <= not w23292 and not w23294;
w23296 <= not w23285 and not w23295;
w23297 <= not w13307 and not w23296;
w23298 <= not w22534 and w22541;
w23299 <= not w22543 and w23298;
w23300 <= not w23118 and w23299;
w23301 <= not w22534 and not w22543;
w23302 <= not w23118 and w23301;
w23303 <= not w22541 and not w23302;
w23304 <= not w23300 and not w23303;
w23305 <= w13307 and not w23285;
w23306 <= not w23295 and w23305;
w23307 <= not w23304 and not w23306;
w23308 <= not w23297 and not w23307;
w23309 <= not w12747 and not w23308;
w23310 <= w22553 and not w22555;
w23311 <= not w22546 and w23310;
w23312 <= not w23118 and w23311;
w23313 <= not w22546 and not w22555;
w23314 <= not w23118 and w23313;
w23315 <= not w22553 and not w23314;
w23316 <= not w23312 and not w23315;
w23317 <= w12747 and not w23297;
w23318 <= not w23307 and w23317;
w23319 <= not w23316 and not w23318;
w23320 <= not w23309 and not w23319;
w23321 <= not w12199 and not w23320;
w23322 <= not w22558 and w22565;
w23323 <= not w22567 and w23322;
w23324 <= not w23118 and w23323;
w23325 <= not w22558 and not w22567;
w23326 <= not w23118 and w23325;
w23327 <= not w22565 and not w23326;
w23328 <= not w23324 and not w23327;
w23329 <= w12199 and not w23309;
w23330 <= not w23319 and w23329;
w23331 <= not w23328 and not w23330;
w23332 <= not w23321 and not w23331;
w23333 <= not w11663 and not w23332;
w23334 <= w22577 and not w22579;
w23335 <= not w22570 and w23334;
w23336 <= not w23118 and w23335;
w23337 <= not w22570 and not w22579;
w23338 <= not w23118 and w23337;
w23339 <= not w22577 and not w23338;
w23340 <= not w23336 and not w23339;
w23341 <= w11663 and not w23321;
w23342 <= not w23331 and w23341;
w23343 <= not w23340 and not w23342;
w23344 <= not w23333 and not w23343;
w23345 <= not w11139 and not w23344;
w23346 <= not w22582 and w22589;
w23347 <= not w22591 and w23346;
w23348 <= not w23118 and w23347;
w23349 <= not w22582 and not w22591;
w23350 <= not w23118 and w23349;
w23351 <= not w22589 and not w23350;
w23352 <= not w23348 and not w23351;
w23353 <= w11139 and not w23333;
w23354 <= not w23343 and w23353;
w23355 <= not w23352 and not w23354;
w23356 <= not w23345 and not w23355;
w23357 <= not w10627 and not w23356;
w23358 <= w22601 and not w22603;
w23359 <= not w22594 and w23358;
w23360 <= not w23118 and w23359;
w23361 <= not w22594 and not w22603;
w23362 <= not w23118 and w23361;
w23363 <= not w22601 and not w23362;
w23364 <= not w23360 and not w23363;
w23365 <= w10627 and not w23345;
w23366 <= not w23355 and w23365;
w23367 <= not w23364 and not w23366;
w23368 <= not w23357 and not w23367;
w23369 <= not w10127 and not w23368;
w23370 <= not w22606 and w22613;
w23371 <= not w22615 and w23370;
w23372 <= not w23118 and w23371;
w23373 <= not w22606 and not w22615;
w23374 <= not w23118 and w23373;
w23375 <= not w22613 and not w23374;
w23376 <= not w23372 and not w23375;
w23377 <= w10127 and not w23357;
w23378 <= not w23367 and w23377;
w23379 <= not w23376 and not w23378;
w23380 <= not w23369 and not w23379;
w23381 <= not w9639 and not w23380;
w23382 <= w22625 and not w22627;
w23383 <= not w22618 and w23382;
w23384 <= not w23118 and w23383;
w23385 <= not w22618 and not w22627;
w23386 <= not w23118 and w23385;
w23387 <= not w22625 and not w23386;
w23388 <= not w23384 and not w23387;
w23389 <= w9639 and not w23369;
w23390 <= not w23379 and w23389;
w23391 <= not w23388 and not w23390;
w23392 <= not w23381 and not w23391;
w23393 <= not w9163 and not w23392;
w23394 <= not w22630 and w22637;
w23395 <= not w22639 and w23394;
w23396 <= not w23118 and w23395;
w23397 <= not w22630 and not w22639;
w23398 <= not w23118 and w23397;
w23399 <= not w22637 and not w23398;
w23400 <= not w23396 and not w23399;
w23401 <= w9163 and not w23381;
w23402 <= not w23391 and w23401;
w23403 <= not w23400 and not w23402;
w23404 <= not w23393 and not w23403;
w23405 <= not w8699 and not w23404;
w23406 <= w22649 and not w22651;
w23407 <= not w22642 and w23406;
w23408 <= not w23118 and w23407;
w23409 <= not w22642 and not w22651;
w23410 <= not w23118 and w23409;
w23411 <= not w22649 and not w23410;
w23412 <= not w23408 and not w23411;
w23413 <= w8699 and not w23393;
w23414 <= not w23403 and w23413;
w23415 <= not w23412 and not w23414;
w23416 <= not w23405 and not w23415;
w23417 <= not w8247 and not w23416;
w23418 <= not w22654 and w22661;
w23419 <= not w22663 and w23418;
w23420 <= not w23118 and w23419;
w23421 <= not w22654 and not w22663;
w23422 <= not w23118 and w23421;
w23423 <= not w22661 and not w23422;
w23424 <= not w23420 and not w23423;
w23425 <= w8247 and not w23405;
w23426 <= not w23415 and w23425;
w23427 <= not w23424 and not w23426;
w23428 <= not w23417 and not w23427;
w23429 <= not w7807 and not w23428;
w23430 <= w22673 and not w22675;
w23431 <= not w22666 and w23430;
w23432 <= not w23118 and w23431;
w23433 <= not w22666 and not w22675;
w23434 <= not w23118 and w23433;
w23435 <= not w22673 and not w23434;
w23436 <= not w23432 and not w23435;
w23437 <= w7807 and not w23417;
w23438 <= not w23427 and w23437;
w23439 <= not w23436 and not w23438;
w23440 <= not w23429 and not w23439;
w23441 <= not w7379 and not w23440;
w23442 <= not w22678 and w22685;
w23443 <= not w22687 and w23442;
w23444 <= not w23118 and w23443;
w23445 <= not w22678 and not w22687;
w23446 <= not w23118 and w23445;
w23447 <= not w22685 and not w23446;
w23448 <= not w23444 and not w23447;
w23449 <= w7379 and not w23429;
w23450 <= not w23439 and w23449;
w23451 <= not w23448 and not w23450;
w23452 <= not w23441 and not w23451;
w23453 <= not w6963 and not w23452;
w23454 <= w22697 and not w22699;
w23455 <= not w22690 and w23454;
w23456 <= not w23118 and w23455;
w23457 <= not w22690 and not w22699;
w23458 <= not w23118 and w23457;
w23459 <= not w22697 and not w23458;
w23460 <= not w23456 and not w23459;
w23461 <= w6963 and not w23441;
w23462 <= not w23451 and w23461;
w23463 <= not w23460 and not w23462;
w23464 <= not w23453 and not w23463;
w23465 <= not w6558 and not w23464;
w23466 <= not w22702 and w22709;
w23467 <= not w22711 and w23466;
w23468 <= not w23118 and w23467;
w23469 <= not w22702 and not w22711;
w23470 <= not w23118 and w23469;
w23471 <= not w22709 and not w23470;
w23472 <= not w23468 and not w23471;
w23473 <= w6558 and not w23453;
w23474 <= not w23463 and w23473;
w23475 <= not w23472 and not w23474;
w23476 <= not w23465 and not w23475;
w23477 <= not w6166 and not w23476;
w23478 <= w22721 and not w22723;
w23479 <= not w22714 and w23478;
w23480 <= not w23118 and w23479;
w23481 <= not w22714 and not w22723;
w23482 <= not w23118 and w23481;
w23483 <= not w22721 and not w23482;
w23484 <= not w23480 and not w23483;
w23485 <= w6166 and not w23465;
w23486 <= not w23475 and w23485;
w23487 <= not w23484 and not w23486;
w23488 <= not w23477 and not w23487;
w23489 <= not w5786 and not w23488;
w23490 <= not w22726 and w22733;
w23491 <= not w22735 and w23490;
w23492 <= not w23118 and w23491;
w23493 <= not w22726 and not w22735;
w23494 <= not w23118 and w23493;
w23495 <= not w22733 and not w23494;
w23496 <= not w23492 and not w23495;
w23497 <= w5786 and not w23477;
w23498 <= not w23487 and w23497;
w23499 <= not w23496 and not w23498;
w23500 <= not w23489 and not w23499;
w23501 <= not w5418 and not w23500;
w23502 <= w22745 and not w22747;
w23503 <= not w22738 and w23502;
w23504 <= not w23118 and w23503;
w23505 <= not w22738 and not w22747;
w23506 <= not w23118 and w23505;
w23507 <= not w22745 and not w23506;
w23508 <= not w23504 and not w23507;
w23509 <= w5418 and not w23489;
w23510 <= not w23499 and w23509;
w23511 <= not w23508 and not w23510;
w23512 <= not w23501 and not w23511;
w23513 <= not w5062 and not w23512;
w23514 <= not w22750 and w22757;
w23515 <= not w22759 and w23514;
w23516 <= not w23118 and w23515;
w23517 <= not w22750 and not w22759;
w23518 <= not w23118 and w23517;
w23519 <= not w22757 and not w23518;
w23520 <= not w23516 and not w23519;
w23521 <= w5062 and not w23501;
w23522 <= not w23511 and w23521;
w23523 <= not w23520 and not w23522;
w23524 <= not w23513 and not w23523;
w23525 <= not w4718 and not w23524;
w23526 <= w22769 and not w22771;
w23527 <= not w22762 and w23526;
w23528 <= not w23118 and w23527;
w23529 <= not w22762 and not w22771;
w23530 <= not w23118 and w23529;
w23531 <= not w22769 and not w23530;
w23532 <= not w23528 and not w23531;
w23533 <= w4718 and not w23513;
w23534 <= not w23523 and w23533;
w23535 <= not w23532 and not w23534;
w23536 <= not w23525 and not w23535;
w23537 <= not w4386 and not w23536;
w23538 <= not w22774 and w22781;
w23539 <= not w22783 and w23538;
w23540 <= not w23118 and w23539;
w23541 <= not w22774 and not w22783;
w23542 <= not w23118 and w23541;
w23543 <= not w22781 and not w23542;
w23544 <= not w23540 and not w23543;
w23545 <= w4386 and not w23525;
w23546 <= not w23535 and w23545;
w23547 <= not w23544 and not w23546;
w23548 <= not w23537 and not w23547;
w23549 <= not w4066 and not w23548;
w23550 <= w22793 and not w22795;
w23551 <= not w22786 and w23550;
w23552 <= not w23118 and w23551;
w23553 <= not w22786 and not w22795;
w23554 <= not w23118 and w23553;
w23555 <= not w22793 and not w23554;
w23556 <= not w23552 and not w23555;
w23557 <= w4066 and not w23537;
w23558 <= not w23547 and w23557;
w23559 <= not w23556 and not w23558;
w23560 <= not w23549 and not w23559;
w23561 <= not w3758 and not w23560;
w23562 <= not w22798 and w22805;
w23563 <= not w22807 and w23562;
w23564 <= not w23118 and w23563;
w23565 <= not w22798 and not w22807;
w23566 <= not w23118 and w23565;
w23567 <= not w22805 and not w23566;
w23568 <= not w23564 and not w23567;
w23569 <= w3758 and not w23549;
w23570 <= not w23559 and w23569;
w23571 <= not w23568 and not w23570;
w23572 <= not w23561 and not w23571;
w23573 <= not w3462 and not w23572;
w23574 <= w22817 and not w22819;
w23575 <= not w22810 and w23574;
w23576 <= not w23118 and w23575;
w23577 <= not w22810 and not w22819;
w23578 <= not w23118 and w23577;
w23579 <= not w22817 and not w23578;
w23580 <= not w23576 and not w23579;
w23581 <= w3462 and not w23561;
w23582 <= not w23571 and w23581;
w23583 <= not w23580 and not w23582;
w23584 <= not w23573 and not w23583;
w23585 <= not w3178 and not w23584;
w23586 <= not w22822 and w22829;
w23587 <= not w22831 and w23586;
w23588 <= not w23118 and w23587;
w23589 <= not w22822 and not w22831;
w23590 <= not w23118 and w23589;
w23591 <= not w22829 and not w23590;
w23592 <= not w23588 and not w23591;
w23593 <= w3178 and not w23573;
w23594 <= not w23583 and w23593;
w23595 <= not w23592 and not w23594;
w23596 <= not w23585 and not w23595;
w23597 <= not w2906 and not w23596;
w23598 <= w22841 and not w22843;
w23599 <= not w22834 and w23598;
w23600 <= not w23118 and w23599;
w23601 <= not w22834 and not w22843;
w23602 <= not w23118 and w23601;
w23603 <= not w22841 and not w23602;
w23604 <= not w23600 and not w23603;
w23605 <= w2906 and not w23585;
w23606 <= not w23595 and w23605;
w23607 <= not w23604 and not w23606;
w23608 <= not w23597 and not w23607;
w23609 <= not w2646 and not w23608;
w23610 <= not w22846 and w22853;
w23611 <= not w22855 and w23610;
w23612 <= not w23118 and w23611;
w23613 <= not w22846 and not w22855;
w23614 <= not w23118 and w23613;
w23615 <= not w22853 and not w23614;
w23616 <= not w23612 and not w23615;
w23617 <= w2646 and not w23597;
w23618 <= not w23607 and w23617;
w23619 <= not w23616 and not w23618;
w23620 <= not w23609 and not w23619;
w23621 <= not w2398 and not w23620;
w23622 <= w22865 and not w22867;
w23623 <= not w22858 and w23622;
w23624 <= not w23118 and w23623;
w23625 <= not w22858 and not w22867;
w23626 <= not w23118 and w23625;
w23627 <= not w22865 and not w23626;
w23628 <= not w23624 and not w23627;
w23629 <= w2398 and not w23609;
w23630 <= not w23619 and w23629;
w23631 <= not w23628 and not w23630;
w23632 <= not w23621 and not w23631;
w23633 <= not w2162 and not w23632;
w23634 <= not w22870 and w22877;
w23635 <= not w22879 and w23634;
w23636 <= not w23118 and w23635;
w23637 <= not w22870 and not w22879;
w23638 <= not w23118 and w23637;
w23639 <= not w22877 and not w23638;
w23640 <= not w23636 and not w23639;
w23641 <= w2162 and not w23621;
w23642 <= not w23631 and w23641;
w23643 <= not w23640 and not w23642;
w23644 <= not w23633 and not w23643;
w23645 <= not w1938 and not w23644;
w23646 <= w22889 and not w22891;
w23647 <= not w22882 and w23646;
w23648 <= not w23118 and w23647;
w23649 <= not w22882 and not w22891;
w23650 <= not w23118 and w23649;
w23651 <= not w22889 and not w23650;
w23652 <= not w23648 and not w23651;
w23653 <= w1938 and not w23633;
w23654 <= not w23643 and w23653;
w23655 <= not w23652 and not w23654;
w23656 <= not w23645 and not w23655;
w23657 <= not w1725 and not w23656;
w23658 <= not w22894 and w22901;
w23659 <= not w22903 and w23658;
w23660 <= not w23118 and w23659;
w23661 <= not w22894 and not w22903;
w23662 <= not w23118 and w23661;
w23663 <= not w22901 and not w23662;
w23664 <= not w23660 and not w23663;
w23665 <= w1725 and not w23645;
w23666 <= not w23655 and w23665;
w23667 <= not w23664 and not w23666;
w23668 <= not w23657 and not w23667;
w23669 <= not w1525 and not w23668;
w23670 <= w22913 and not w22915;
w23671 <= not w22906 and w23670;
w23672 <= not w23118 and w23671;
w23673 <= not w22906 and not w22915;
w23674 <= not w23118 and w23673;
w23675 <= not w22913 and not w23674;
w23676 <= not w23672 and not w23675;
w23677 <= w1525 and not w23657;
w23678 <= not w23667 and w23677;
w23679 <= not w23676 and not w23678;
w23680 <= not w23669 and not w23679;
w23681 <= not w1337 and not w23680;
w23682 <= not w22918 and w22925;
w23683 <= not w22927 and w23682;
w23684 <= not w23118 and w23683;
w23685 <= not w22918 and not w22927;
w23686 <= not w23118 and w23685;
w23687 <= not w22925 and not w23686;
w23688 <= not w23684 and not w23687;
w23689 <= w1337 and not w23669;
w23690 <= not w23679 and w23689;
w23691 <= not w23688 and not w23690;
w23692 <= not w23681 and not w23691;
w23693 <= not w1161 and not w23692;
w23694 <= w22937 and not w22939;
w23695 <= not w22930 and w23694;
w23696 <= not w23118 and w23695;
w23697 <= not w22930 and not w22939;
w23698 <= not w23118 and w23697;
w23699 <= not w22937 and not w23698;
w23700 <= not w23696 and not w23699;
w23701 <= w1161 and not w23681;
w23702 <= not w23691 and w23701;
w23703 <= not w23700 and not w23702;
w23704 <= not w23693 and not w23703;
w23705 <= not w997 and not w23704;
w23706 <= not w22942 and w22949;
w23707 <= not w22951 and w23706;
w23708 <= not w23118 and w23707;
w23709 <= not w22942 and not w22951;
w23710 <= not w23118 and w23709;
w23711 <= not w22949 and not w23710;
w23712 <= not w23708 and not w23711;
w23713 <= w997 and not w23693;
w23714 <= not w23703 and w23713;
w23715 <= not w23712 and not w23714;
w23716 <= not w23705 and not w23715;
w23717 <= not w845 and not w23716;
w23718 <= w22961 and not w22963;
w23719 <= not w22954 and w23718;
w23720 <= not w23118 and w23719;
w23721 <= not w22954 and not w22963;
w23722 <= not w23118 and w23721;
w23723 <= not w22961 and not w23722;
w23724 <= not w23720 and not w23723;
w23725 <= w845 and not w23705;
w23726 <= not w23715 and w23725;
w23727 <= not w23724 and not w23726;
w23728 <= not w23717 and not w23727;
w23729 <= not w705 and not w23728;
w23730 <= not w22966 and w22973;
w23731 <= not w22975 and w23730;
w23732 <= not w23118 and w23731;
w23733 <= not w22966 and not w22975;
w23734 <= not w23118 and w23733;
w23735 <= not w22973 and not w23734;
w23736 <= not w23732 and not w23735;
w23737 <= w705 and not w23717;
w23738 <= not w23727 and w23737;
w23739 <= not w23736 and not w23738;
w23740 <= not w23729 and not w23739;
w23741 <= not w577 and not w23740;
w23742 <= w22985 and not w22987;
w23743 <= not w22978 and w23742;
w23744 <= not w23118 and w23743;
w23745 <= not w22978 and not w22987;
w23746 <= not w23118 and w23745;
w23747 <= not w22985 and not w23746;
w23748 <= not w23744 and not w23747;
w23749 <= w577 and not w23729;
w23750 <= not w23739 and w23749;
w23751 <= not w23748 and not w23750;
w23752 <= not w23741 and not w23751;
w23753 <= not w460 and not w23752;
w23754 <= not w22990 and w22997;
w23755 <= not w22999 and w23754;
w23756 <= not w23118 and w23755;
w23757 <= not w22990 and not w22999;
w23758 <= not w23118 and w23757;
w23759 <= not w22997 and not w23758;
w23760 <= not w23756 and not w23759;
w23761 <= w460 and not w23741;
w23762 <= not w23751 and w23761;
w23763 <= not w23760 and not w23762;
w23764 <= not w23753 and not w23763;
w23765 <= not w356 and not w23764;
w23766 <= w23009 and not w23011;
w23767 <= not w23002 and w23766;
w23768 <= not w23118 and w23767;
w23769 <= not w23002 and not w23011;
w23770 <= not w23118 and w23769;
w23771 <= not w23009 and not w23770;
w23772 <= not w23768 and not w23771;
w23773 <= w356 and not w23753;
w23774 <= not w23763 and w23773;
w23775 <= not w23772 and not w23774;
w23776 <= not w23765 and not w23775;
w23777 <= not w264 and not w23776;
w23778 <= not w23014 and w23021;
w23779 <= not w23023 and w23778;
w23780 <= not w23118 and w23779;
w23781 <= not w23014 and not w23023;
w23782 <= not w23118 and w23781;
w23783 <= not w23021 and not w23782;
w23784 <= not w23780 and not w23783;
w23785 <= w264 and not w23765;
w23786 <= not w23775 and w23785;
w23787 <= not w23784 and not w23786;
w23788 <= not w23777 and not w23787;
w23789 <= not w184 and not w23788;
w23790 <= w23033 and not w23035;
w23791 <= not w23026 and w23790;
w23792 <= not w23118 and w23791;
w23793 <= not w23026 and not w23035;
w23794 <= not w23118 and w23793;
w23795 <= not w23033 and not w23794;
w23796 <= not w23792 and not w23795;
w23797 <= w184 and not w23777;
w23798 <= not w23787 and w23797;
w23799 <= not w23796 and not w23798;
w23800 <= not w23789 and not w23799;
w23801 <= not w115 and not w23800;
w23802 <= not w23038 and w23045;
w23803 <= not w23047 and w23802;
w23804 <= not w23118 and w23803;
w23805 <= not w23038 and not w23047;
w23806 <= not w23118 and w23805;
w23807 <= not w23045 and not w23806;
w23808 <= not w23804 and not w23807;
w23809 <= w115 and not w23789;
w23810 <= not w23799 and w23809;
w23811 <= not w23808 and not w23810;
w23812 <= not w23801 and not w23811;
w23813 <= not w60 and not w23812;
w23814 <= w23057 and not w23059;
w23815 <= not w23050 and w23814;
w23816 <= not w23118 and w23815;
w23817 <= not w23050 and not w23059;
w23818 <= not w23118 and w23817;
w23819 <= not w23057 and not w23818;
w23820 <= not w23816 and not w23819;
w23821 <= w60 and not w23801;
w23822 <= not w23811 and w23821;
w23823 <= not w23820 and not w23822;
w23824 <= not w23813 and not w23823;
w23825 <= not w22 and not w23824;
w23826 <= w22 and not w23813;
w23827 <= not w23823 and w23826;
w23828 <= not w23125 and not w23827;
w23829 <= not w23825 and not w23828;
w23830 <= not w5 and not w23829;
w23831 <= w23081 and not w23083;
w23832 <= not w23074 and w23831;
w23833 <= not w23118 and w23832;
w23834 <= not w23074 and not w23083;
w23835 <= not w23118 and w23834;
w23836 <= not w23081 and not w23835;
w23837 <= not w23833 and not w23836;
w23838 <= w5 and not w23825;
w23839 <= not w23828 and w23838;
w23840 <= not w23837 and not w23839;
w23841 <= not w23830 and not w23840;
w23842 <= not w23086 and w23095;
w23843 <= not w23088 and w23842;
w23844 <= not w23118 and w23843;
w23845 <= not w23086 and not w23088;
w23846 <= not w23118 and w23845;
w23847 <= not w23095 and not w23846;
w23848 <= not w23844 and not w23847;
w23849 <= not w23097 and not w23104;
w23850 <= not w23118 and w23849;
w23851 <= not w23112 and not w23850;
w23852 <= not w23848 and w23851;
w23853 <= not w23841 and w23852;
w23854 <= w0 and not w23853;
w23855 <= not w23830 and w23848;
w23856 <= not w23840 and w23855;
w23857 <= not w23104 and not w23118;
w23858 <= w23097 and not w23857;
w23859 <= not w0 and not w23849;
w23860 <= not w23858 and w23859;
w23861 <= not w23856 and not w23860;
w23862 <= not w23854 and w23861;
w23863 <= not w23825 and not w23827;
w23864 <= not w23862 and w23863;
w23865 <= not w23125 and not w23864;
w23866 <= w23125 and not w23825;
w23867 <= not w23827 and w23866;
w23868 <= not w23862 and w23867;
w23869 <= not w23865 and not w23868;
w23870 <= not w23801 and not w23810;
w23871 <= not w23862 and w23870;
w23872 <= not w23808 and not w23871;
w23873 <= not w23801 and w23808;
w23874 <= not w23810 and w23873;
w23875 <= not w23862 and w23874;
w23876 <= not w23872 and not w23875;
w23877 <= not w23777 and not w23786;
w23878 <= not w23862 and w23877;
w23879 <= not w23784 and not w23878;
w23880 <= not w23777 and w23784;
w23881 <= not w23786 and w23880;
w23882 <= not w23862 and w23881;
w23883 <= not w23879 and not w23882;
w23884 <= not w23753 and not w23762;
w23885 <= not w23862 and w23884;
w23886 <= not w23760 and not w23885;
w23887 <= not w23753 and w23760;
w23888 <= not w23762 and w23887;
w23889 <= not w23862 and w23888;
w23890 <= not w23886 and not w23889;
w23891 <= not w23729 and not w23738;
w23892 <= not w23862 and w23891;
w23893 <= not w23736 and not w23892;
w23894 <= not w23729 and w23736;
w23895 <= not w23738 and w23894;
w23896 <= not w23862 and w23895;
w23897 <= not w23893 and not w23896;
w23898 <= not w23705 and not w23714;
w23899 <= not w23862 and w23898;
w23900 <= not w23712 and not w23899;
w23901 <= not w23705 and w23712;
w23902 <= not w23714 and w23901;
w23903 <= not w23862 and w23902;
w23904 <= not w23900 and not w23903;
w23905 <= not w23681 and not w23690;
w23906 <= not w23862 and w23905;
w23907 <= not w23688 and not w23906;
w23908 <= not w23681 and w23688;
w23909 <= not w23690 and w23908;
w23910 <= not w23862 and w23909;
w23911 <= not w23907 and not w23910;
w23912 <= not w23657 and not w23666;
w23913 <= not w23862 and w23912;
w23914 <= not w23664 and not w23913;
w23915 <= not w23657 and w23664;
w23916 <= not w23666 and w23915;
w23917 <= not w23862 and w23916;
w23918 <= not w23914 and not w23917;
w23919 <= not w23633 and not w23642;
w23920 <= not w23862 and w23919;
w23921 <= not w23640 and not w23920;
w23922 <= not w23633 and w23640;
w23923 <= not w23642 and w23922;
w23924 <= not w23862 and w23923;
w23925 <= not w23921 and not w23924;
w23926 <= not w23609 and not w23618;
w23927 <= not w23862 and w23926;
w23928 <= not w23616 and not w23927;
w23929 <= not w23609 and w23616;
w23930 <= not w23618 and w23929;
w23931 <= not w23862 and w23930;
w23932 <= not w23928 and not w23931;
w23933 <= not w23585 and not w23594;
w23934 <= not w23862 and w23933;
w23935 <= not w23592 and not w23934;
w23936 <= not w23585 and w23592;
w23937 <= not w23594 and w23936;
w23938 <= not w23862 and w23937;
w23939 <= not w23935 and not w23938;
w23940 <= not w23561 and not w23570;
w23941 <= not w23862 and w23940;
w23942 <= not w23568 and not w23941;
w23943 <= not w23561 and w23568;
w23944 <= not w23570 and w23943;
w23945 <= not w23862 and w23944;
w23946 <= not w23942 and not w23945;
w23947 <= not w23537 and not w23546;
w23948 <= not w23862 and w23947;
w23949 <= not w23544 and not w23948;
w23950 <= not w23537 and w23544;
w23951 <= not w23546 and w23950;
w23952 <= not w23862 and w23951;
w23953 <= not w23949 and not w23952;
w23954 <= not w23513 and not w23522;
w23955 <= not w23862 and w23954;
w23956 <= not w23520 and not w23955;
w23957 <= not w23513 and w23520;
w23958 <= not w23522 and w23957;
w23959 <= not w23862 and w23958;
w23960 <= not w23956 and not w23959;
w23961 <= not w23489 and not w23498;
w23962 <= not w23862 and w23961;
w23963 <= not w23496 and not w23962;
w23964 <= not w23489 and w23496;
w23965 <= not w23498 and w23964;
w23966 <= not w23862 and w23965;
w23967 <= not w23963 and not w23966;
w23968 <= not w23465 and not w23474;
w23969 <= not w23862 and w23968;
w23970 <= not w23472 and not w23969;
w23971 <= not w23465 and w23472;
w23972 <= not w23474 and w23971;
w23973 <= not w23862 and w23972;
w23974 <= not w23970 and not w23973;
w23975 <= not w23441 and not w23450;
w23976 <= not w23862 and w23975;
w23977 <= not w23448 and not w23976;
w23978 <= not w23441 and w23448;
w23979 <= not w23450 and w23978;
w23980 <= not w23862 and w23979;
w23981 <= not w23977 and not w23980;
w23982 <= not w23417 and not w23426;
w23983 <= not w23862 and w23982;
w23984 <= not w23424 and not w23983;
w23985 <= not w23417 and w23424;
w23986 <= not w23426 and w23985;
w23987 <= not w23862 and w23986;
w23988 <= not w23984 and not w23987;
w23989 <= not w23393 and not w23402;
w23990 <= not w23862 and w23989;
w23991 <= not w23400 and not w23990;
w23992 <= not w23393 and w23400;
w23993 <= not w23402 and w23992;
w23994 <= not w23862 and w23993;
w23995 <= not w23991 and not w23994;
w23996 <= not w23369 and not w23378;
w23997 <= not w23862 and w23996;
w23998 <= not w23376 and not w23997;
w23999 <= not w23369 and w23376;
w24000 <= not w23378 and w23999;
w24001 <= not w23862 and w24000;
w24002 <= not w23998 and not w24001;
w24003 <= not w23345 and not w23354;
w24004 <= not w23862 and w24003;
w24005 <= not w23352 and not w24004;
w24006 <= not w23345 and w23352;
w24007 <= not w23354 and w24006;
w24008 <= not w23862 and w24007;
w24009 <= not w24005 and not w24008;
w24010 <= not w23321 and not w23330;
w24011 <= not w23862 and w24010;
w24012 <= not w23328 and not w24011;
w24013 <= not w23321 and w23328;
w24014 <= not w23330 and w24013;
w24015 <= not w23862 and w24014;
w24016 <= not w24012 and not w24015;
w24017 <= not w23297 and not w23306;
w24018 <= not w23862 and w24017;
w24019 <= not w23304 and not w24018;
w24020 <= not w23297 and w23304;
w24021 <= not w23306 and w24020;
w24022 <= not w23862 and w24021;
w24023 <= not w24019 and not w24022;
w24024 <= not w23273 and not w23282;
w24025 <= not w23862 and w24024;
w24026 <= not w23280 and not w24025;
w24027 <= not w23273 and w23280;
w24028 <= not w23282 and w24027;
w24029 <= not w23862 and w24028;
w24030 <= not w24026 and not w24029;
w24031 <= not w23249 and not w23258;
w24032 <= not w23862 and w24031;
w24033 <= not w23256 and not w24032;
w24034 <= not w23249 and w23256;
w24035 <= not w23258 and w24034;
w24036 <= not w23862 and w24035;
w24037 <= not w24033 and not w24036;
w24038 <= not w23225 and not w23234;
w24039 <= not w23862 and w24038;
w24040 <= not w23232 and not w24039;
w24041 <= not w23225 and w23232;
w24042 <= not w23234 and w24041;
w24043 <= not w23862 and w24042;
w24044 <= not w24040 and not w24043;
w24045 <= not w23201 and not w23210;
w24046 <= not w23862 and w24045;
w24047 <= not w23208 and not w24046;
w24048 <= not w23201 and w23208;
w24049 <= not w23210 and w24048;
w24050 <= not w23862 and w24049;
w24051 <= not w24047 and not w24050;
w24052 <= not w23177 and not w23186;
w24053 <= not w23862 and w24052;
w24054 <= not w23184 and not w24053;
w24055 <= not w23177 and w23184;
w24056 <= not w23186 and w24055;
w24057 <= not w23862 and w24056;
w24058 <= not w24054 and not w24057;
w24059 <= not w23154 and w23160;
w24060 <= not w23162 and w24059;
w24061 <= not w23862 and w24060;
w24062 <= not w23154 and not w23162;
w24063 <= not w23862 and w24062;
w24064 <= not w23160 and not w24063;
w24065 <= not w24061 and not w24064;
w24066 <= not w23130 and not w23134;
w24067 <= not w23138 and w24066;
w24068 <= not w23862 and w24067;
w24069 <= not w23862 and w24066;
w24070 <= w23138 and not w24069;
w24071 <= not w24068 and not w24070;
w24072 <= w23127 and not w23862;
w24073 <= not w23118 and not w23860;
w24074 <= not w23856 and w24073;
w24075 <= not w23854 and w24074;
w24076 <= not w24072 and not w24075;
w24077 <= a(4) and not w24076;
w24078 <= not a(4) and not w24075;
w24079 <= not w24072 and w24078;
w24080 <= not w24077 and not w24079;
w24081 <= not a(2) and not w23862;
w24082 <= a(3) and not w24081;
w24083 <= not a(0) and not a(1);
w24084 <= not a(2) and not w24083;
w24085 <= a(2) and not w23860;
w24086 <= not w23856 and w24085;
w24087 <= not w23854 and w24086;
w24088 <= not w24084 and not w24087;
w24089 <= not w24072 and w24088;
w24090 <= not w24082 and w24089;
w24091 <= w23118 and not w24090;
w24092 <= not w24072 and not w24082;
w24093 <= not w24088 and not w24092;
w24094 <= not w24091 and not w24093;
w24095 <= not w24080 and w24094;
w24096 <= w22386 and not w24095;
w24097 <= w24080 and not w24094;
w24098 <= not w24096 and not w24097;
w24099 <= w24071 and not w24098;
w24100 <= not w24071 and not w24097;
w24101 <= not w24096 and w24100;
w24102 <= w21666 and not w24101;
w24103 <= not w23141 and not w23143;
w24104 <= not w23862 and w24103;
w24105 <= not w23151 and not w24104;
w24106 <= not w23143 and w23151;
w24107 <= not w23141 and w24106;
w24108 <= not w23862 and w24107;
w24109 <= not w24105 and not w24108;
w24110 <= not w24102 and not w24109;
w24111 <= not w24099 and w24110;
w24112 <= w20957 and not w24111;
w24113 <= not w24099 and not w24102;
w24114 <= w24109 and not w24113;
w24115 <= not w24112 and not w24114;
w24116 <= w24065 and not w24115;
w24117 <= not w24065 and not w24114;
w24118 <= not w24112 and w24117;
w24119 <= w20259 and not w24118;
w24120 <= not w23165 and not w23174;
w24121 <= not w23862 and w24120;
w24122 <= not w23172 and not w24121;
w24123 <= w23172 and not w23174;
w24124 <= not w23165 and w24123;
w24125 <= not w23862 and w24124;
w24126 <= not w24122 and not w24125;
w24127 <= not w24119 and not w24126;
w24128 <= not w24116 and w24127;
w24129 <= w19567 and not w24128;
w24130 <= not w24116 and not w24119;
w24131 <= w24126 and not w24130;
w24132 <= not w24129 and not w24131;
w24133 <= w24058 and not w24132;
w24134 <= not w24058 and not w24131;
w24135 <= not w24129 and w24134;
w24136 <= w18887 and not w24135;
w24137 <= not w23189 and not w23198;
w24138 <= not w23862 and w24137;
w24139 <= not w23196 and not w24138;
w24140 <= w23196 and not w23198;
w24141 <= not w23189 and w24140;
w24142 <= not w23862 and w24141;
w24143 <= not w24139 and not w24142;
w24144 <= not w24136 and not w24143;
w24145 <= not w24133 and w24144;
w24146 <= w18219 and not w24145;
w24147 <= not w24133 and not w24136;
w24148 <= w24143 and not w24147;
w24149 <= not w24146 and not w24148;
w24150 <= w24051 and not w24149;
w24151 <= not w24051 and not w24148;
w24152 <= not w24146 and w24151;
w24153 <= w17563 and not w24152;
w24154 <= not w23213 and not w23222;
w24155 <= not w23862 and w24154;
w24156 <= not w23220 and not w24155;
w24157 <= w23220 and not w23222;
w24158 <= not w23213 and w24157;
w24159 <= not w23862 and w24158;
w24160 <= not w24156 and not w24159;
w24161 <= not w24153 and not w24160;
w24162 <= not w24150 and w24161;
w24163 <= w16919 and not w24162;
w24164 <= not w24150 and not w24153;
w24165 <= w24160 and not w24164;
w24166 <= not w24163 and not w24165;
w24167 <= w24044 and not w24166;
w24168 <= not w24044 and not w24165;
w24169 <= not w24163 and w24168;
w24170 <= w16287 and not w24169;
w24171 <= not w23237 and not w23246;
w24172 <= not w23862 and w24171;
w24173 <= not w23244 and not w24172;
w24174 <= w23244 and not w23246;
w24175 <= not w23237 and w24174;
w24176 <= not w23862 and w24175;
w24177 <= not w24173 and not w24176;
w24178 <= not w24170 and not w24177;
w24179 <= not w24167 and w24178;
w24180 <= w15667 and not w24179;
w24181 <= not w24167 and not w24170;
w24182 <= w24177 and not w24181;
w24183 <= not w24180 and not w24182;
w24184 <= w24037 and not w24183;
w24185 <= not w24037 and not w24182;
w24186 <= not w24180 and w24185;
w24187 <= w15059 and not w24186;
w24188 <= not w23261 and not w23270;
w24189 <= not w23862 and w24188;
w24190 <= not w23268 and not w24189;
w24191 <= w23268 and not w23270;
w24192 <= not w23261 and w24191;
w24193 <= not w23862 and w24192;
w24194 <= not w24190 and not w24193;
w24195 <= not w24187 and not w24194;
w24196 <= not w24184 and w24195;
w24197 <= w14463 and not w24196;
w24198 <= not w24184 and not w24187;
w24199 <= w24194 and not w24198;
w24200 <= not w24197 and not w24199;
w24201 <= w24030 and not w24200;
w24202 <= not w24030 and not w24199;
w24203 <= not w24197 and w24202;
w24204 <= w13879 and not w24203;
w24205 <= not w23285 and not w23294;
w24206 <= not w23862 and w24205;
w24207 <= not w23292 and not w24206;
w24208 <= w23292 and not w23294;
w24209 <= not w23285 and w24208;
w24210 <= not w23862 and w24209;
w24211 <= not w24207 and not w24210;
w24212 <= not w24204 and not w24211;
w24213 <= not w24201 and w24212;
w24214 <= w13307 and not w24213;
w24215 <= not w24201 and not w24204;
w24216 <= w24211 and not w24215;
w24217 <= not w24214 and not w24216;
w24218 <= w24023 and not w24217;
w24219 <= not w24023 and not w24216;
w24220 <= not w24214 and w24219;
w24221 <= w12747 and not w24220;
w24222 <= not w23309 and not w23318;
w24223 <= not w23862 and w24222;
w24224 <= not w23316 and not w24223;
w24225 <= w23316 and not w23318;
w24226 <= not w23309 and w24225;
w24227 <= not w23862 and w24226;
w24228 <= not w24224 and not w24227;
w24229 <= not w24221 and not w24228;
w24230 <= not w24218 and w24229;
w24231 <= w12199 and not w24230;
w24232 <= not w24218 and not w24221;
w24233 <= w24228 and not w24232;
w24234 <= not w24231 and not w24233;
w24235 <= w24016 and not w24234;
w24236 <= not w24016 and not w24233;
w24237 <= not w24231 and w24236;
w24238 <= w11663 and not w24237;
w24239 <= not w23333 and not w23342;
w24240 <= not w23862 and w24239;
w24241 <= not w23340 and not w24240;
w24242 <= w23340 and not w23342;
w24243 <= not w23333 and w24242;
w24244 <= not w23862 and w24243;
w24245 <= not w24241 and not w24244;
w24246 <= not w24238 and not w24245;
w24247 <= not w24235 and w24246;
w24248 <= w11139 and not w24247;
w24249 <= not w24235 and not w24238;
w24250 <= w24245 and not w24249;
w24251 <= not w24248 and not w24250;
w24252 <= w24009 and not w24251;
w24253 <= not w24009 and not w24250;
w24254 <= not w24248 and w24253;
w24255 <= w10627 and not w24254;
w24256 <= not w23357 and not w23366;
w24257 <= not w23862 and w24256;
w24258 <= not w23364 and not w24257;
w24259 <= w23364 and not w23366;
w24260 <= not w23357 and w24259;
w24261 <= not w23862 and w24260;
w24262 <= not w24258 and not w24261;
w24263 <= not w24255 and not w24262;
w24264 <= not w24252 and w24263;
w24265 <= w10127 and not w24264;
w24266 <= not w24252 and not w24255;
w24267 <= w24262 and not w24266;
w24268 <= not w24265 and not w24267;
w24269 <= w24002 and not w24268;
w24270 <= not w24002 and not w24267;
w24271 <= not w24265 and w24270;
w24272 <= w9639 and not w24271;
w24273 <= not w23381 and not w23390;
w24274 <= not w23862 and w24273;
w24275 <= not w23388 and not w24274;
w24276 <= w23388 and not w23390;
w24277 <= not w23381 and w24276;
w24278 <= not w23862 and w24277;
w24279 <= not w24275 and not w24278;
w24280 <= not w24272 and not w24279;
w24281 <= not w24269 and w24280;
w24282 <= w9163 and not w24281;
w24283 <= not w24269 and not w24272;
w24284 <= w24279 and not w24283;
w24285 <= not w24282 and not w24284;
w24286 <= w23995 and not w24285;
w24287 <= not w23995 and not w24284;
w24288 <= not w24282 and w24287;
w24289 <= w8699 and not w24288;
w24290 <= not w23405 and not w23414;
w24291 <= not w23862 and w24290;
w24292 <= not w23412 and not w24291;
w24293 <= w23412 and not w23414;
w24294 <= not w23405 and w24293;
w24295 <= not w23862 and w24294;
w24296 <= not w24292 and not w24295;
w24297 <= not w24289 and not w24296;
w24298 <= not w24286 and w24297;
w24299 <= w8247 and not w24298;
w24300 <= not w24286 and not w24289;
w24301 <= w24296 and not w24300;
w24302 <= not w24299 and not w24301;
w24303 <= w23988 and not w24302;
w24304 <= not w23988 and not w24301;
w24305 <= not w24299 and w24304;
w24306 <= w7807 and not w24305;
w24307 <= not w23429 and not w23438;
w24308 <= not w23862 and w24307;
w24309 <= not w23436 and not w24308;
w24310 <= w23436 and not w23438;
w24311 <= not w23429 and w24310;
w24312 <= not w23862 and w24311;
w24313 <= not w24309 and not w24312;
w24314 <= not w24306 and not w24313;
w24315 <= not w24303 and w24314;
w24316 <= w7379 and not w24315;
w24317 <= not w24303 and not w24306;
w24318 <= w24313 and not w24317;
w24319 <= not w24316 and not w24318;
w24320 <= w23981 and not w24319;
w24321 <= not w23981 and not w24318;
w24322 <= not w24316 and w24321;
w24323 <= w6963 and not w24322;
w24324 <= not w23453 and not w23462;
w24325 <= not w23862 and w24324;
w24326 <= not w23460 and not w24325;
w24327 <= w23460 and not w23462;
w24328 <= not w23453 and w24327;
w24329 <= not w23862 and w24328;
w24330 <= not w24326 and not w24329;
w24331 <= not w24323 and not w24330;
w24332 <= not w24320 and w24331;
w24333 <= w6558 and not w24332;
w24334 <= not w24320 and not w24323;
w24335 <= w24330 and not w24334;
w24336 <= not w24333 and not w24335;
w24337 <= w23974 and not w24336;
w24338 <= not w23974 and not w24335;
w24339 <= not w24333 and w24338;
w24340 <= w6166 and not w24339;
w24341 <= not w23477 and not w23486;
w24342 <= not w23862 and w24341;
w24343 <= not w23484 and not w24342;
w24344 <= w23484 and not w23486;
w24345 <= not w23477 and w24344;
w24346 <= not w23862 and w24345;
w24347 <= not w24343 and not w24346;
w24348 <= not w24340 and not w24347;
w24349 <= not w24337 and w24348;
w24350 <= w5786 and not w24349;
w24351 <= not w24337 and not w24340;
w24352 <= w24347 and not w24351;
w24353 <= not w24350 and not w24352;
w24354 <= w23967 and not w24353;
w24355 <= not w23967 and not w24352;
w24356 <= not w24350 and w24355;
w24357 <= w5418 and not w24356;
w24358 <= not w23501 and not w23510;
w24359 <= not w23862 and w24358;
w24360 <= not w23508 and not w24359;
w24361 <= w23508 and not w23510;
w24362 <= not w23501 and w24361;
w24363 <= not w23862 and w24362;
w24364 <= not w24360 and not w24363;
w24365 <= not w24357 and not w24364;
w24366 <= not w24354 and w24365;
w24367 <= w5062 and not w24366;
w24368 <= not w24354 and not w24357;
w24369 <= w24364 and not w24368;
w24370 <= not w24367 and not w24369;
w24371 <= w23960 and not w24370;
w24372 <= not w23960 and not w24369;
w24373 <= not w24367 and w24372;
w24374 <= w4718 and not w24373;
w24375 <= not w23525 and not w23534;
w24376 <= not w23862 and w24375;
w24377 <= not w23532 and not w24376;
w24378 <= w23532 and not w23534;
w24379 <= not w23525 and w24378;
w24380 <= not w23862 and w24379;
w24381 <= not w24377 and not w24380;
w24382 <= not w24374 and not w24381;
w24383 <= not w24371 and w24382;
w24384 <= w4386 and not w24383;
w24385 <= not w24371 and not w24374;
w24386 <= w24381 and not w24385;
w24387 <= not w24384 and not w24386;
w24388 <= w23953 and not w24387;
w24389 <= not w23953 and not w24386;
w24390 <= not w24384 and w24389;
w24391 <= w4066 and not w24390;
w24392 <= not w23549 and not w23558;
w24393 <= not w23862 and w24392;
w24394 <= not w23556 and not w24393;
w24395 <= w23556 and not w23558;
w24396 <= not w23549 and w24395;
w24397 <= not w23862 and w24396;
w24398 <= not w24394 and not w24397;
w24399 <= not w24391 and not w24398;
w24400 <= not w24388 and w24399;
w24401 <= w3758 and not w24400;
w24402 <= not w24388 and not w24391;
w24403 <= w24398 and not w24402;
w24404 <= not w24401 and not w24403;
w24405 <= w23946 and not w24404;
w24406 <= not w23946 and not w24403;
w24407 <= not w24401 and w24406;
w24408 <= w3462 and not w24407;
w24409 <= not w23573 and not w23582;
w24410 <= not w23862 and w24409;
w24411 <= not w23580 and not w24410;
w24412 <= w23580 and not w23582;
w24413 <= not w23573 and w24412;
w24414 <= not w23862 and w24413;
w24415 <= not w24411 and not w24414;
w24416 <= not w24408 and not w24415;
w24417 <= not w24405 and w24416;
w24418 <= w3178 and not w24417;
w24419 <= not w24405 and not w24408;
w24420 <= w24415 and not w24419;
w24421 <= not w24418 and not w24420;
w24422 <= w23939 and not w24421;
w24423 <= not w23939 and not w24420;
w24424 <= not w24418 and w24423;
w24425 <= w2906 and not w24424;
w24426 <= not w23597 and not w23606;
w24427 <= not w23862 and w24426;
w24428 <= not w23604 and not w24427;
w24429 <= w23604 and not w23606;
w24430 <= not w23597 and w24429;
w24431 <= not w23862 and w24430;
w24432 <= not w24428 and not w24431;
w24433 <= not w24425 and not w24432;
w24434 <= not w24422 and w24433;
w24435 <= w2646 and not w24434;
w24436 <= not w24422 and not w24425;
w24437 <= w24432 and not w24436;
w24438 <= not w24435 and not w24437;
w24439 <= w23932 and not w24438;
w24440 <= not w23932 and not w24437;
w24441 <= not w24435 and w24440;
w24442 <= w2398 and not w24441;
w24443 <= not w23621 and not w23630;
w24444 <= not w23862 and w24443;
w24445 <= not w23628 and not w24444;
w24446 <= w23628 and not w23630;
w24447 <= not w23621 and w24446;
w24448 <= not w23862 and w24447;
w24449 <= not w24445 and not w24448;
w24450 <= not w24442 and not w24449;
w24451 <= not w24439 and w24450;
w24452 <= w2162 and not w24451;
w24453 <= not w24439 and not w24442;
w24454 <= w24449 and not w24453;
w24455 <= not w24452 and not w24454;
w24456 <= w23925 and not w24455;
w24457 <= not w23925 and not w24454;
w24458 <= not w24452 and w24457;
w24459 <= w1938 and not w24458;
w24460 <= not w23645 and not w23654;
w24461 <= not w23862 and w24460;
w24462 <= not w23652 and not w24461;
w24463 <= w23652 and not w23654;
w24464 <= not w23645 and w24463;
w24465 <= not w23862 and w24464;
w24466 <= not w24462 and not w24465;
w24467 <= not w24459 and not w24466;
w24468 <= not w24456 and w24467;
w24469 <= w1725 and not w24468;
w24470 <= not w24456 and not w24459;
w24471 <= w24466 and not w24470;
w24472 <= not w24469 and not w24471;
w24473 <= w23918 and not w24472;
w24474 <= not w23918 and not w24471;
w24475 <= not w24469 and w24474;
w24476 <= w1525 and not w24475;
w24477 <= not w23669 and not w23678;
w24478 <= not w23862 and w24477;
w24479 <= not w23676 and not w24478;
w24480 <= w23676 and not w23678;
w24481 <= not w23669 and w24480;
w24482 <= not w23862 and w24481;
w24483 <= not w24479 and not w24482;
w24484 <= not w24476 and not w24483;
w24485 <= not w24473 and w24484;
w24486 <= w1337 and not w24485;
w24487 <= not w24473 and not w24476;
w24488 <= w24483 and not w24487;
w24489 <= not w24486 and not w24488;
w24490 <= w23911 and not w24489;
w24491 <= not w23911 and not w24488;
w24492 <= not w24486 and w24491;
w24493 <= w1161 and not w24492;
w24494 <= not w23693 and not w23702;
w24495 <= not w23862 and w24494;
w24496 <= not w23700 and not w24495;
w24497 <= w23700 and not w23702;
w24498 <= not w23693 and w24497;
w24499 <= not w23862 and w24498;
w24500 <= not w24496 and not w24499;
w24501 <= not w24493 and not w24500;
w24502 <= not w24490 and w24501;
w24503 <= w997 and not w24502;
w24504 <= not w24490 and not w24493;
w24505 <= w24500 and not w24504;
w24506 <= not w24503 and not w24505;
w24507 <= w23904 and not w24506;
w24508 <= not w23904 and not w24505;
w24509 <= not w24503 and w24508;
w24510 <= w845 and not w24509;
w24511 <= not w23717 and not w23726;
w24512 <= not w23862 and w24511;
w24513 <= not w23724 and not w24512;
w24514 <= w23724 and not w23726;
w24515 <= not w23717 and w24514;
w24516 <= not w23862 and w24515;
w24517 <= not w24513 and not w24516;
w24518 <= not w24510 and not w24517;
w24519 <= not w24507 and w24518;
w24520 <= w705 and not w24519;
w24521 <= not w24507 and not w24510;
w24522 <= w24517 and not w24521;
w24523 <= not w24520 and not w24522;
w24524 <= w23897 and not w24523;
w24525 <= not w23897 and not w24522;
w24526 <= not w24520 and w24525;
w24527 <= w577 and not w24526;
w24528 <= not w23741 and not w23750;
w24529 <= not w23862 and w24528;
w24530 <= not w23748 and not w24529;
w24531 <= w23748 and not w23750;
w24532 <= not w23741 and w24531;
w24533 <= not w23862 and w24532;
w24534 <= not w24530 and not w24533;
w24535 <= not w24527 and not w24534;
w24536 <= not w24524 and w24535;
w24537 <= w460 and not w24536;
w24538 <= not w24524 and not w24527;
w24539 <= w24534 and not w24538;
w24540 <= not w24537 and not w24539;
w24541 <= w23890 and not w24540;
w24542 <= not w23890 and not w24539;
w24543 <= not w24537 and w24542;
w24544 <= w356 and not w24543;
w24545 <= not w23765 and not w23774;
w24546 <= not w23862 and w24545;
w24547 <= not w23772 and not w24546;
w24548 <= w23772 and not w23774;
w24549 <= not w23765 and w24548;
w24550 <= not w23862 and w24549;
w24551 <= not w24547 and not w24550;
w24552 <= not w24544 and not w24551;
w24553 <= not w24541 and w24552;
w24554 <= w264 and not w24553;
w24555 <= not w24541 and not w24544;
w24556 <= w24551 and not w24555;
w24557 <= not w24554 and not w24556;
w24558 <= w23883 and not w24557;
w24559 <= not w23883 and not w24556;
w24560 <= not w24554 and w24559;
w24561 <= w184 and not w24560;
w24562 <= not w23789 and not w23798;
w24563 <= not w23862 and w24562;
w24564 <= not w23796 and not w24563;
w24565 <= w23796 and not w23798;
w24566 <= not w23789 and w24565;
w24567 <= not w23862 and w24566;
w24568 <= not w24564 and not w24567;
w24569 <= not w24561 and not w24568;
w24570 <= not w24558 and w24569;
w24571 <= w115 and not w24570;
w24572 <= not w24558 and not w24561;
w24573 <= w24568 and not w24572;
w24574 <= not w24571 and not w24573;
w24575 <= w23876 and not w24574;
w24576 <= not w23876 and not w24573;
w24577 <= not w24571 and w24576;
w24578 <= w60 and not w24577;
w24579 <= not w23813 and not w23822;
w24580 <= not w23862 and w24579;
w24581 <= not w23820 and not w24580;
w24582 <= w23820 and not w23822;
w24583 <= not w23813 and w24582;
w24584 <= not w23862 and w24583;
w24585 <= not w24581 and not w24584;
w24586 <= not w24578 and not w24585;
w24587 <= not w24575 and w24586;
w24588 <= w22 and not w24587;
w24589 <= not w24575 and not w24578;
w24590 <= w24585 and not w24589;
w24591 <= not w24588 and not w24590;
w24592 <= w23869 and not w24591;
w24593 <= not w23869 and not w24590;
w24594 <= not w24588 and w24593;
w24595 <= w5 and not w24594;
w24596 <= not w23830 and not w23839;
w24597 <= not w23862 and w24596;
w24598 <= not w23837 and not w24597;
w24599 <= w23837 and not w23839;
w24600 <= not w23830 and w24599;
w24601 <= not w23862 and w24600;
w24602 <= not w24598 and not w24601;
w24603 <= not w23841 and not w23848;
w24604 <= not w23862 and w24603;
w24605 <= not w23856 and not w24604;
w24606 <= not w24602 and w24605;
w24607 <= not w24595 and w24606;
w24608 <= not w24592 and w24607;
w24609 <= w0 and not w24608;
w24610 <= not w24592 and not w24595;
w24611 <= w24602 and not w24610;
w24612 <= not w23848 and not w23862;
w24613 <= w23841 and not w24612;
w24614 <= not w0 and not w24603;
w24615 <= not w24613 and w24614;
w24616 <= not w24611 and not w24615;
w24617 <= not w24609 and w24616;
one <= '1';
asqrt(0) <= not w24617;-- level 5058
asqrt(1) <= not w23862;-- level 4900
asqrt(2) <= not w23118;-- level 4745
asqrt(3) <= not w22386;-- level 4592
asqrt(4) <= not w21666;-- level 4442
asqrt(5) <= not w20957;-- level 4294
asqrt(6) <= not w20259;-- level 4149
asqrt(7) <= not w19567;-- level 4006
asqrt(8) <= not w18887;-- level 3866
asqrt(9) <= not w18219;-- level 3728
asqrt(10) <= not w17563;-- level 3593
asqrt(11) <= not w16919;-- level 3460
asqrt(12) <= not w16287;-- level 3330
asqrt(13) <= not w15667;-- level 3202
asqrt(14) <= not w15059;-- level 3077
asqrt(15) <= not w14463;-- level 2954
asqrt(16) <= not w13879;-- level 2834
asqrt(17) <= not w13307;-- level 2716
asqrt(18) <= not w12747;-- level 2601
asqrt(19) <= not w12199;-- level 2488
asqrt(20) <= not w11663;-- level 2378
asqrt(21) <= not w11139;-- level 2270
asqrt(22) <= not w10627;-- level 2165
asqrt(23) <= not w10127;-- level 2062
asqrt(24) <= not w9639;-- level 1962
asqrt(25) <= not w9163;-- level 1864
asqrt(26) <= not w8699;-- level 1769
asqrt(27) <= not w8247;-- level 1676
asqrt(28) <= not w7807;-- level 1586
asqrt(29) <= not w7379;-- level 1498
asqrt(30) <= not w6963;-- level 1413
asqrt(31) <= not w6558;-- level 1330
asqrt(32) <= not w6166;-- level 1250
asqrt(33) <= not w5786;-- level 1172
asqrt(34) <= not w5418;-- level 1097
asqrt(35) <= not w5062;-- level 1024
asqrt(36) <= not w4718;-- level 954
asqrt(37) <= not w4386;-- level 886
asqrt(38) <= not w4066;-- level 821
asqrt(39) <= not w3758;-- level 758
asqrt(40) <= not w3462;-- level 698
asqrt(41) <= not w3178;-- level 640
asqrt(42) <= not w2906;-- level 585
asqrt(43) <= not w2646;-- level 532
asqrt(44) <= not w2398;-- level 482
asqrt(45) <= not w2162;-- level 434
asqrt(46) <= not w1938;-- level 389
asqrt(47) <= not w1725;-- level 346
asqrt(48) <= not w1525;-- level 306
asqrt(49) <= not w1337;-- level 268
asqrt(50) <= not w1161;-- level 233
asqrt(51) <= not w997;-- level 200
asqrt(52) <= not w845;-- level 170
asqrt(53) <= not w705;-- level 142
asqrt(54) <= not w577;-- level 117
asqrt(55) <= not w460;-- level 94
asqrt(56) <= not w356;-- level 74
asqrt(57) <= not w264;-- level 56
asqrt(58) <= not w184;-- level 41
asqrt(59) <= not w115;-- level 28
asqrt(60) <= not w60;-- level 18
asqrt(61) <= not w22;-- level 10
asqrt(62) <= not w5;-- level 4
asqrt(63) <= not w0;-- level 1
end Behavioral;