//-----------------------------------------------------------------------------
//      RapidSilicon
//      Author: Pankil Patel
//      Date:   6/5/2022
//-----------------------------------------------------------------------------

module mode_ctrl (
	input				testmode,
	output				scanmode,
	output				bscanmode,
	output				funcmode
	);
endmodule
