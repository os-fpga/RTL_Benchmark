-- $Id: input.vhdl,v 1.1.1.1 2005-12-06 02:47:46 arif_endro Exp $
-------------------------------------------------------------------------------
-- Title       : Input
-- Project     : Mini AES 128 
-------------------------------------------------------------------------------
-- File        : input.vhdl
-- Author      : "Arif E. Nugroho" <arif_endro@yahoo.com>
-- Created     : 2005/12/03
-- Last update : 
-- Simulators  : ModelSim SE PLUS 6.0
-- Synthesizers: ISE Xilinx 6.3i
-- Target      : 
-------------------------------------------------------------------------------
-- Description : Input stimuli file for test bench.
-------------------------------------------------------------------------------
-- Copyright (C) 2005 Arif E. Nugroho
-- This VHDL design file is an open design; you can redistribute it and/or
-- modify it and/or implement it after contacting the author
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- 
--         THIS SOURCE FILE MAY BE USED AND DISTRIBUTED WITHOUT RESTRICTION
-- PROVIDED THAT THIS COPYRIGHT STATEMENT IS NOT REMOVED FROM THE FILE AND THAT
-- ANY DERIVATIVE WORK CONTAINS THE ORIGINAL COPYRIGHT NOTICE AND THE
-- ASSOCIATED DISCLAIMER.
-- 
-------------------------------------------------------------------------------
-- 
--         THIS SOFTWARE IS PROVIDED BY THE AUTHOR ``AS IS'' AND ANY EXPRESS OR
-- IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF
-- MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.  IN NO
-- EVENT SHALL THE AUTHOR BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
-- SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO,
-- PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
-- OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY,
-- WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR
-- OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_textio.all;
use std.textio.all;

library std_developerskit;
use std_developerskit.std_iopak.all;    -- Function From_HexString

entity input is
  port (
    clock          : out std_logic;
    clear          : out std_logic;
    done           : in  std_logic;
    test_iteration : out integer;
    data_i         : out std_logic_vector (127 downto 000);
    cipher_o       : out std_logic_vector (127 downto 000);
    key_i          : out std_logic_vector (127 downto 000)
    );
end input;

architecture test_bench of input is

--
  file in_file_ptr            : text open read_mode is "../data/ecb_tbl.txt";
--
  signal     clock_int        : std_logic := '0';
--
begin
--
  clock_int          <= not(clock_int) after 1 ns;
  clock              <= clock_int;
--
  process
--
    variable delay            : time      := 1 ns;
    variable in_line          : line;
    variable cipher_text      : string ( 01 to 32 );
    variable plain_text       : string ( 01 to 32 );
    variable key              : string ( 01 to 32 );
    variable test             : integer;
    variable junk_test        : string ( 01 to 02 );
    variable junk_plain_text  : string ( 01 to 03 );
    variable junk_cipher_text : string (01 to 03 );
    variable junk_key         : string ( 01 to 04 );
--
  begin
--
    while not (endfile(in_file_ptr)) loop
--
      readline(in_file_ptr, in_line);   -- blank lines
--
      readline(in_file_ptr, in_line);
      read(in_line, junk_test);
      read(in_line, test);
      readline(in_file_ptr, in_line);
      read(in_line, junk_key);
      read(in_line, key);
      readline(in_file_ptr, in_line);
      read(in_line, junk_plain_text);
      read(in_line, plain_text);
      readline(in_file_ptr, in_line);
      read(in_line, junk_cipher_text);
      read(in_line, cipher_text);
--
      wait until rising_edge(clock_int);
      key_i          <= to_StdLogicVector(From_HexString(key( 01 to 32)));
      data_i         <= to_StdLogicVector(From_HexString(plain_text( 01 to 32 )));
      cipher_o       <= to_StdLogicVector(From_HexString(cipher_text( 01 to 32 )));
      test_iteration <= test;
--
      clear          <= '1';
      wait until rising_edge(clock_int);
      clear          <= '0';
      wait until rising_edge(done);
      wait until rising_edge(clock_int);
--
    end loop;
    wait;
  end process;
--
end test_bench;
